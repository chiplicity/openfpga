VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_core
  CLASS BLOCK ;
  FOREIGN fpga_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2486.000 BY 2546.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END IO_ISOL_N
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2482.000 2386.840 2486.000 2387.440 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END clk
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 2542.000 46.370 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 477.400 2486.000 478.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 795.640 2486.000 796.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 1113.880 2486.000 1114.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 1432.120 2486.000 1432.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 1750.360 2486.000 1750.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 2068.600 2486.000 2069.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2180.490 0.000 2180.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2191.990 0.000 2192.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2203.490 0.000 2203.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2214.990 0.000 2215.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.090 2542.000 138.370 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.490 0.000 2226.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2237.990 0.000 2238.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2249.490 0.000 2249.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2260.990 0.000 2261.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2272.490 0.000 2272.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.990 0.000 1870.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1881.490 0.000 1881.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1892.990 0.000 1893.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1904.490 0.000 1904.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1915.990 0.000 1916.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 230.090 2542.000 230.370 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1927.490 0.000 1927.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1938.990 0.000 1939.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1950.490 0.000 1950.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1961.990 0.000 1962.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1559.030 0.000 1559.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1570.530 0.000 1570.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1582.030 0.000 1582.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1593.530 0.000 1593.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1605.030 0.000 1605.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1616.530 0.000 1616.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 322.090 2542.000 322.370 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1628.030 0.000 1628.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1639.530 0.000 1639.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1651.030 0.000 1651.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1248.530 0.000 1248.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1260.030 0.000 1260.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1271.530 0.000 1271.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1283.030 0.000 1283.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1306.030 0.000 1306.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1317.530 0.000 1317.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 414.090 2542.000 414.370 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1329.030 0.000 1329.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1340.530 0.000 1340.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 937.570 0.000 937.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 949.070 0.000 949.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 960.570 0.000 960.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 972.070 0.000 972.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 983.570 0.000 983.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1006.570 0.000 1006.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1018.070 0.000 1018.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 506.090 2542.000 506.370 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1029.570 0.000 1029.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.070 0.000 627.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 684.570 0.000 684.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 696.070 0.000 696.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 598.090 2542.000 598.370 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 690.550 2542.000 690.830 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 657.600 4.000 658.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 782.550 2542.000 782.830 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1184.600 4.000 1185.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1447.760 4.000 1448.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.920 4.000 1711.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1974.760 4.000 1975.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2237.920 4.000 2238.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 159.160 2486.000 159.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 874.550 2542.000 874.830 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2482.000 583.480 2486.000 584.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2482.000 901.720 2486.000 902.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2482.000 1219.960 2486.000 1220.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2482.000 1538.200 2486.000 1538.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2482.000 1856.440 2486.000 1857.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2482.000 2174.680 2486.000 2175.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2283.990 0.000 2284.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2295.490 0.000 2295.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2306.990 0.000 2307.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2318.490 0.000 2318.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 966.550 2542.000 966.830 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2329.990 0.000 2330.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2341.490 0.000 2341.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2352.990 0.000 2353.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2364.490 0.000 2364.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.990 0.000 2376.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1973.490 0.000 1973.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1984.990 0.000 1985.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1996.490 0.000 1996.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2007.990 0.000 2008.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2019.490 0.000 2019.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1058.550 2542.000 1058.830 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2030.990 0.000 2031.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.490 0.000 2042.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2053.990 0.000 2054.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2065.490 0.000 2065.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1662.530 0.000 1662.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1674.030 0.000 1674.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.530 0.000 1685.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.030 0.000 1697.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1708.530 0.000 1708.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1720.030 0.000 1720.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.550 2542.000 1150.830 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1731.530 0.000 1731.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1743.030 0.000 1743.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1754.530 0.000 1754.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1352.030 0.000 1352.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1363.530 0.000 1363.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1375.030 0.000 1375.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1386.530 0.000 1386.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1398.030 0.000 1398.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1409.530 0.000 1409.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1421.030 0.000 1421.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1242.550 2542.000 1242.830 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1432.530 0.000 1432.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1444.030 0.000 1444.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1041.070 0.000 1041.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1052.570 0.000 1052.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1064.070 0.000 1064.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.070 0.000 1087.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1098.570 0.000 1098.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.070 0.000 1110.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1121.570 0.000 1121.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1335.010 2542.000 1335.290 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1133.070 0.000 1133.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 730.570 0.000 730.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 742.070 0.000 742.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 765.070 0.000 765.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 788.070 0.000 788.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 799.570 0.000 799.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 822.570 0.000 822.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1427.010 2542.000 1427.290 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1519.010 2542.000 1519.290 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.160 4.000 482.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.320 4.000 745.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1611.010 2542.000 1611.290 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.160 4.000 1009.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1272.320 4.000 1272.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1535.480 4.000 1536.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1799.320 4.000 1799.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2062.480 4.000 2063.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2325.640 4.000 2326.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2482.000 265.240 2486.000 265.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1703.010 2542.000 1703.290 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 689.560 2486.000 690.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 1007.800 2486.000 1008.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 1326.040 2486.000 1326.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 1644.280 2486.000 1644.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 1962.520 2486.000 1963.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 2280.760 2486.000 2281.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.490 0.000 2387.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2398.990 0.000 2399.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2410.490 0.000 2410.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2421.990 0.000 2422.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1795.010 2542.000 1795.290 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2433.490 0.000 2433.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2444.990 0.000 2445.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2456.490 0.000 2456.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2467.990 0.000 2468.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2479.490 0.000 2479.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2076.990 0.000 2077.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2088.490 0.000 2088.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2099.990 0.000 2100.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2111.490 0.000 2111.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2122.990 0.000 2123.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.010 2542.000 1887.290 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2134.490 0.000 2134.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2145.990 0.000 2146.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2157.490 0.000 2157.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2168.990 0.000 2169.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1766.030 0.000 1766.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1777.530 0.000 1777.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1789.030 0.000 1789.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1800.530 0.000 1800.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1812.030 0.000 1812.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1823.530 0.000 1823.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1979.470 2542.000 1979.750 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1835.030 0.000 1835.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1846.530 0.000 1846.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1858.030 0.000 1858.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1467.030 0.000 1467.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1478.530 0.000 1478.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1490.030 0.000 1490.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1501.530 0.000 1501.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1513.030 0.000 1513.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1524.530 0.000 1524.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2071.470 2542.000 2071.750 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1536.030 0.000 1536.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1547.530 0.000 1547.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1144.570 0.000 1144.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1167.570 0.000 1167.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1179.070 0.000 1179.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1190.570 0.000 1190.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1202.070 0.000 1202.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1213.570 0.000 1213.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1225.070 0.000 1225.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2163.470 2542.000 2163.750 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 857.070 0.000 857.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 868.570 0.000 868.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.070 0.000 880.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 891.570 0.000 891.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 903.070 0.000 903.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 926.070 0.000 926.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2255.470 2542.000 2255.750 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2347.470 2542.000 2347.750 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2439.470 2542.000 2439.750 2546.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.880 4.000 1097.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1623.200 4.000 1623.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1887.040 4.000 1887.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2150.200 4.000 2150.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2413.360 4.000 2413.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 371.320 2486.000 371.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2482.000 53.080 2486.000 53.680 ;
    END
  END prog_clk
  PIN sc_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2501.080 4.000 2501.680 ;
    END
  END sc_head
  PIN sc_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2482.000 2492.920 2486.000 2493.520 ;
    END
  END sc_tail
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 95.080 2480.320 96.680 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 125.080 2480.320 126.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 40.165 15.385 2436.015 2541.205 ;
      LAYER met1 ;
        RECT 5.590 4.460 2479.790 2541.360 ;
      LAYER met2 ;
        RECT 5.620 2541.720 45.810 2542.000 ;
        RECT 46.650 2541.720 137.810 2542.000 ;
        RECT 138.650 2541.720 229.810 2542.000 ;
        RECT 230.650 2541.720 321.810 2542.000 ;
        RECT 322.650 2541.720 413.810 2542.000 ;
        RECT 414.650 2541.720 505.810 2542.000 ;
        RECT 506.650 2541.720 597.810 2542.000 ;
        RECT 598.650 2541.720 690.270 2542.000 ;
        RECT 691.110 2541.720 782.270 2542.000 ;
        RECT 783.110 2541.720 874.270 2542.000 ;
        RECT 875.110 2541.720 966.270 2542.000 ;
        RECT 967.110 2541.720 1058.270 2542.000 ;
        RECT 1059.110 2541.720 1150.270 2542.000 ;
        RECT 1151.110 2541.720 1242.270 2542.000 ;
        RECT 1243.110 2541.720 1334.730 2542.000 ;
        RECT 1335.570 2541.720 1426.730 2542.000 ;
        RECT 1427.570 2541.720 1518.730 2542.000 ;
        RECT 1519.570 2541.720 1610.730 2542.000 ;
        RECT 1611.570 2541.720 1702.730 2542.000 ;
        RECT 1703.570 2541.720 1794.730 2542.000 ;
        RECT 1795.570 2541.720 1886.730 2542.000 ;
        RECT 1887.570 2541.720 1979.190 2542.000 ;
        RECT 1980.030 2541.720 2071.190 2542.000 ;
        RECT 2072.030 2541.720 2163.190 2542.000 ;
        RECT 2164.030 2541.720 2255.190 2542.000 ;
        RECT 2256.030 2541.720 2347.190 2542.000 ;
        RECT 2348.030 2541.720 2439.190 2542.000 ;
        RECT 2440.030 2541.720 2479.760 2542.000 ;
        RECT 5.620 4.280 2479.760 2541.720 ;
        RECT 6.170 4.000 16.830 4.280 ;
        RECT 17.670 4.000 28.330 4.280 ;
        RECT 29.170 4.000 39.830 4.280 ;
        RECT 40.670 4.000 51.330 4.280 ;
        RECT 52.170 4.000 62.830 4.280 ;
        RECT 63.670 4.000 74.330 4.280 ;
        RECT 75.170 4.000 85.830 4.280 ;
        RECT 86.670 4.000 97.330 4.280 ;
        RECT 98.170 4.000 108.830 4.280 ;
        RECT 109.670 4.000 120.330 4.280 ;
        RECT 121.170 4.000 131.830 4.280 ;
        RECT 132.670 4.000 143.330 4.280 ;
        RECT 144.170 4.000 154.830 4.280 ;
        RECT 155.670 4.000 166.330 4.280 ;
        RECT 167.170 4.000 177.830 4.280 ;
        RECT 178.670 4.000 189.330 4.280 ;
        RECT 190.170 4.000 200.830 4.280 ;
        RECT 201.670 4.000 212.330 4.280 ;
        RECT 213.170 4.000 223.830 4.280 ;
        RECT 224.670 4.000 235.330 4.280 ;
        RECT 236.170 4.000 246.830 4.280 ;
        RECT 247.670 4.000 258.330 4.280 ;
        RECT 259.170 4.000 269.830 4.280 ;
        RECT 270.670 4.000 281.330 4.280 ;
        RECT 282.170 4.000 292.830 4.280 ;
        RECT 293.670 4.000 304.330 4.280 ;
        RECT 305.170 4.000 315.830 4.280 ;
        RECT 316.670 4.000 327.330 4.280 ;
        RECT 328.170 4.000 338.830 4.280 ;
        RECT 339.670 4.000 350.330 4.280 ;
        RECT 351.170 4.000 361.830 4.280 ;
        RECT 362.670 4.000 373.330 4.280 ;
        RECT 374.170 4.000 384.830 4.280 ;
        RECT 385.670 4.000 396.330 4.280 ;
        RECT 397.170 4.000 407.830 4.280 ;
        RECT 408.670 4.000 419.330 4.280 ;
        RECT 420.170 4.000 430.830 4.280 ;
        RECT 431.670 4.000 442.330 4.280 ;
        RECT 443.170 4.000 453.830 4.280 ;
        RECT 454.670 4.000 465.330 4.280 ;
        RECT 466.170 4.000 476.830 4.280 ;
        RECT 477.670 4.000 488.330 4.280 ;
        RECT 489.170 4.000 499.830 4.280 ;
        RECT 500.670 4.000 511.330 4.280 ;
        RECT 512.170 4.000 522.830 4.280 ;
        RECT 523.670 4.000 534.330 4.280 ;
        RECT 535.170 4.000 545.830 4.280 ;
        RECT 546.670 4.000 557.330 4.280 ;
        RECT 558.170 4.000 568.830 4.280 ;
        RECT 569.670 4.000 580.330 4.280 ;
        RECT 581.170 4.000 591.830 4.280 ;
        RECT 592.670 4.000 603.330 4.280 ;
        RECT 604.170 4.000 614.830 4.280 ;
        RECT 615.670 4.000 626.790 4.280 ;
        RECT 627.630 4.000 638.290 4.280 ;
        RECT 639.130 4.000 649.790 4.280 ;
        RECT 650.630 4.000 661.290 4.280 ;
        RECT 662.130 4.000 672.790 4.280 ;
        RECT 673.630 4.000 684.290 4.280 ;
        RECT 685.130 4.000 695.790 4.280 ;
        RECT 696.630 4.000 707.290 4.280 ;
        RECT 708.130 4.000 718.790 4.280 ;
        RECT 719.630 4.000 730.290 4.280 ;
        RECT 731.130 4.000 741.790 4.280 ;
        RECT 742.630 4.000 753.290 4.280 ;
        RECT 754.130 4.000 764.790 4.280 ;
        RECT 765.630 4.000 776.290 4.280 ;
        RECT 777.130 4.000 787.790 4.280 ;
        RECT 788.630 4.000 799.290 4.280 ;
        RECT 800.130 4.000 810.790 4.280 ;
        RECT 811.630 4.000 822.290 4.280 ;
        RECT 823.130 4.000 833.790 4.280 ;
        RECT 834.630 4.000 845.290 4.280 ;
        RECT 846.130 4.000 856.790 4.280 ;
        RECT 857.630 4.000 868.290 4.280 ;
        RECT 869.130 4.000 879.790 4.280 ;
        RECT 880.630 4.000 891.290 4.280 ;
        RECT 892.130 4.000 902.790 4.280 ;
        RECT 903.630 4.000 914.290 4.280 ;
        RECT 915.130 4.000 925.790 4.280 ;
        RECT 926.630 4.000 937.290 4.280 ;
        RECT 938.130 4.000 948.790 4.280 ;
        RECT 949.630 4.000 960.290 4.280 ;
        RECT 961.130 4.000 971.790 4.280 ;
        RECT 972.630 4.000 983.290 4.280 ;
        RECT 984.130 4.000 994.790 4.280 ;
        RECT 995.630 4.000 1006.290 4.280 ;
        RECT 1007.130 4.000 1017.790 4.280 ;
        RECT 1018.630 4.000 1029.290 4.280 ;
        RECT 1030.130 4.000 1040.790 4.280 ;
        RECT 1041.630 4.000 1052.290 4.280 ;
        RECT 1053.130 4.000 1063.790 4.280 ;
        RECT 1064.630 4.000 1075.290 4.280 ;
        RECT 1076.130 4.000 1086.790 4.280 ;
        RECT 1087.630 4.000 1098.290 4.280 ;
        RECT 1099.130 4.000 1109.790 4.280 ;
        RECT 1110.630 4.000 1121.290 4.280 ;
        RECT 1122.130 4.000 1132.790 4.280 ;
        RECT 1133.630 4.000 1144.290 4.280 ;
        RECT 1145.130 4.000 1155.790 4.280 ;
        RECT 1156.630 4.000 1167.290 4.280 ;
        RECT 1168.130 4.000 1178.790 4.280 ;
        RECT 1179.630 4.000 1190.290 4.280 ;
        RECT 1191.130 4.000 1201.790 4.280 ;
        RECT 1202.630 4.000 1213.290 4.280 ;
        RECT 1214.130 4.000 1224.790 4.280 ;
        RECT 1225.630 4.000 1236.290 4.280 ;
        RECT 1237.130 4.000 1248.250 4.280 ;
        RECT 1249.090 4.000 1259.750 4.280 ;
        RECT 1260.590 4.000 1271.250 4.280 ;
        RECT 1272.090 4.000 1282.750 4.280 ;
        RECT 1283.590 4.000 1294.250 4.280 ;
        RECT 1295.090 4.000 1305.750 4.280 ;
        RECT 1306.590 4.000 1317.250 4.280 ;
        RECT 1318.090 4.000 1328.750 4.280 ;
        RECT 1329.590 4.000 1340.250 4.280 ;
        RECT 1341.090 4.000 1351.750 4.280 ;
        RECT 1352.590 4.000 1363.250 4.280 ;
        RECT 1364.090 4.000 1374.750 4.280 ;
        RECT 1375.590 4.000 1386.250 4.280 ;
        RECT 1387.090 4.000 1397.750 4.280 ;
        RECT 1398.590 4.000 1409.250 4.280 ;
        RECT 1410.090 4.000 1420.750 4.280 ;
        RECT 1421.590 4.000 1432.250 4.280 ;
        RECT 1433.090 4.000 1443.750 4.280 ;
        RECT 1444.590 4.000 1455.250 4.280 ;
        RECT 1456.090 4.000 1466.750 4.280 ;
        RECT 1467.590 4.000 1478.250 4.280 ;
        RECT 1479.090 4.000 1489.750 4.280 ;
        RECT 1490.590 4.000 1501.250 4.280 ;
        RECT 1502.090 4.000 1512.750 4.280 ;
        RECT 1513.590 4.000 1524.250 4.280 ;
        RECT 1525.090 4.000 1535.750 4.280 ;
        RECT 1536.590 4.000 1547.250 4.280 ;
        RECT 1548.090 4.000 1558.750 4.280 ;
        RECT 1559.590 4.000 1570.250 4.280 ;
        RECT 1571.090 4.000 1581.750 4.280 ;
        RECT 1582.590 4.000 1593.250 4.280 ;
        RECT 1594.090 4.000 1604.750 4.280 ;
        RECT 1605.590 4.000 1616.250 4.280 ;
        RECT 1617.090 4.000 1627.750 4.280 ;
        RECT 1628.590 4.000 1639.250 4.280 ;
        RECT 1640.090 4.000 1650.750 4.280 ;
        RECT 1651.590 4.000 1662.250 4.280 ;
        RECT 1663.090 4.000 1673.750 4.280 ;
        RECT 1674.590 4.000 1685.250 4.280 ;
        RECT 1686.090 4.000 1696.750 4.280 ;
        RECT 1697.590 4.000 1708.250 4.280 ;
        RECT 1709.090 4.000 1719.750 4.280 ;
        RECT 1720.590 4.000 1731.250 4.280 ;
        RECT 1732.090 4.000 1742.750 4.280 ;
        RECT 1743.590 4.000 1754.250 4.280 ;
        RECT 1755.090 4.000 1765.750 4.280 ;
        RECT 1766.590 4.000 1777.250 4.280 ;
        RECT 1778.090 4.000 1788.750 4.280 ;
        RECT 1789.590 4.000 1800.250 4.280 ;
        RECT 1801.090 4.000 1811.750 4.280 ;
        RECT 1812.590 4.000 1823.250 4.280 ;
        RECT 1824.090 4.000 1834.750 4.280 ;
        RECT 1835.590 4.000 1846.250 4.280 ;
        RECT 1847.090 4.000 1857.750 4.280 ;
        RECT 1858.590 4.000 1869.710 4.280 ;
        RECT 1870.550 4.000 1881.210 4.280 ;
        RECT 1882.050 4.000 1892.710 4.280 ;
        RECT 1893.550 4.000 1904.210 4.280 ;
        RECT 1905.050 4.000 1915.710 4.280 ;
        RECT 1916.550 4.000 1927.210 4.280 ;
        RECT 1928.050 4.000 1938.710 4.280 ;
        RECT 1939.550 4.000 1950.210 4.280 ;
        RECT 1951.050 4.000 1961.710 4.280 ;
        RECT 1962.550 4.000 1973.210 4.280 ;
        RECT 1974.050 4.000 1984.710 4.280 ;
        RECT 1985.550 4.000 1996.210 4.280 ;
        RECT 1997.050 4.000 2007.710 4.280 ;
        RECT 2008.550 4.000 2019.210 4.280 ;
        RECT 2020.050 4.000 2030.710 4.280 ;
        RECT 2031.550 4.000 2042.210 4.280 ;
        RECT 2043.050 4.000 2053.710 4.280 ;
        RECT 2054.550 4.000 2065.210 4.280 ;
        RECT 2066.050 4.000 2076.710 4.280 ;
        RECT 2077.550 4.000 2088.210 4.280 ;
        RECT 2089.050 4.000 2099.710 4.280 ;
        RECT 2100.550 4.000 2111.210 4.280 ;
        RECT 2112.050 4.000 2122.710 4.280 ;
        RECT 2123.550 4.000 2134.210 4.280 ;
        RECT 2135.050 4.000 2145.710 4.280 ;
        RECT 2146.550 4.000 2157.210 4.280 ;
        RECT 2158.050 4.000 2168.710 4.280 ;
        RECT 2169.550 4.000 2180.210 4.280 ;
        RECT 2181.050 4.000 2191.710 4.280 ;
        RECT 2192.550 4.000 2203.210 4.280 ;
        RECT 2204.050 4.000 2214.710 4.280 ;
        RECT 2215.550 4.000 2226.210 4.280 ;
        RECT 2227.050 4.000 2237.710 4.280 ;
        RECT 2238.550 4.000 2249.210 4.280 ;
        RECT 2250.050 4.000 2260.710 4.280 ;
        RECT 2261.550 4.000 2272.210 4.280 ;
        RECT 2273.050 4.000 2283.710 4.280 ;
        RECT 2284.550 4.000 2295.210 4.280 ;
        RECT 2296.050 4.000 2306.710 4.280 ;
        RECT 2307.550 4.000 2318.210 4.280 ;
        RECT 2319.050 4.000 2329.710 4.280 ;
        RECT 2330.550 4.000 2341.210 4.280 ;
        RECT 2342.050 4.000 2352.710 4.280 ;
        RECT 2353.550 4.000 2364.210 4.280 ;
        RECT 2365.050 4.000 2375.710 4.280 ;
        RECT 2376.550 4.000 2387.210 4.280 ;
        RECT 2388.050 4.000 2398.710 4.280 ;
        RECT 2399.550 4.000 2410.210 4.280 ;
        RECT 2411.050 4.000 2421.710 4.280 ;
        RECT 2422.550 4.000 2433.210 4.280 ;
        RECT 2434.050 4.000 2444.710 4.280 ;
        RECT 2445.550 4.000 2456.210 4.280 ;
        RECT 2457.050 4.000 2467.710 4.280 ;
        RECT 2468.550 4.000 2479.210 4.280 ;
      LAYER met3 ;
        RECT 4.000 2502.080 2482.000 2541.285 ;
        RECT 4.400 2500.680 2482.000 2502.080 ;
        RECT 4.000 2493.920 2482.000 2500.680 ;
        RECT 4.000 2492.520 2481.600 2493.920 ;
        RECT 4.000 2414.360 2482.000 2492.520 ;
        RECT 4.400 2412.960 2482.000 2414.360 ;
        RECT 4.000 2387.840 2482.000 2412.960 ;
        RECT 4.000 2386.440 2481.600 2387.840 ;
        RECT 4.000 2326.640 2482.000 2386.440 ;
        RECT 4.400 2325.240 2482.000 2326.640 ;
        RECT 4.000 2281.760 2482.000 2325.240 ;
        RECT 4.000 2280.360 2481.600 2281.760 ;
        RECT 4.000 2238.920 2482.000 2280.360 ;
        RECT 4.400 2237.520 2482.000 2238.920 ;
        RECT 4.000 2175.680 2482.000 2237.520 ;
        RECT 4.000 2174.280 2481.600 2175.680 ;
        RECT 4.000 2151.200 2482.000 2174.280 ;
        RECT 4.400 2149.800 2482.000 2151.200 ;
        RECT 4.000 2069.600 2482.000 2149.800 ;
        RECT 4.000 2068.200 2481.600 2069.600 ;
        RECT 4.000 2063.480 2482.000 2068.200 ;
        RECT 4.400 2062.080 2482.000 2063.480 ;
        RECT 4.000 1975.760 2482.000 2062.080 ;
        RECT 4.400 1974.360 2482.000 1975.760 ;
        RECT 4.000 1963.520 2482.000 1974.360 ;
        RECT 4.000 1962.120 2481.600 1963.520 ;
        RECT 4.000 1888.040 2482.000 1962.120 ;
        RECT 4.400 1886.640 2482.000 1888.040 ;
        RECT 4.000 1857.440 2482.000 1886.640 ;
        RECT 4.000 1856.040 2481.600 1857.440 ;
        RECT 4.000 1800.320 2482.000 1856.040 ;
        RECT 4.400 1798.920 2482.000 1800.320 ;
        RECT 4.000 1751.360 2482.000 1798.920 ;
        RECT 4.000 1749.960 2481.600 1751.360 ;
        RECT 4.000 1711.920 2482.000 1749.960 ;
        RECT 4.400 1710.520 2482.000 1711.920 ;
        RECT 4.000 1645.280 2482.000 1710.520 ;
        RECT 4.000 1643.880 2481.600 1645.280 ;
        RECT 4.000 1624.200 2482.000 1643.880 ;
        RECT 4.400 1622.800 2482.000 1624.200 ;
        RECT 4.000 1539.200 2482.000 1622.800 ;
        RECT 4.000 1537.800 2481.600 1539.200 ;
        RECT 4.000 1536.480 2482.000 1537.800 ;
        RECT 4.400 1535.080 2482.000 1536.480 ;
        RECT 4.000 1448.760 2482.000 1535.080 ;
        RECT 4.400 1447.360 2482.000 1448.760 ;
        RECT 4.000 1433.120 2482.000 1447.360 ;
        RECT 4.000 1431.720 2481.600 1433.120 ;
        RECT 4.000 1361.040 2482.000 1431.720 ;
        RECT 4.400 1359.640 2482.000 1361.040 ;
        RECT 4.000 1327.040 2482.000 1359.640 ;
        RECT 4.000 1325.640 2481.600 1327.040 ;
        RECT 4.000 1273.320 2482.000 1325.640 ;
        RECT 4.400 1271.920 2482.000 1273.320 ;
        RECT 4.000 1220.960 2482.000 1271.920 ;
        RECT 4.000 1219.560 2481.600 1220.960 ;
        RECT 4.000 1185.600 2482.000 1219.560 ;
        RECT 4.400 1184.200 2482.000 1185.600 ;
        RECT 4.000 1114.880 2482.000 1184.200 ;
        RECT 4.000 1113.480 2481.600 1114.880 ;
        RECT 4.000 1097.880 2482.000 1113.480 ;
        RECT 4.400 1096.480 2482.000 1097.880 ;
        RECT 4.000 1010.160 2482.000 1096.480 ;
        RECT 4.400 1008.800 2482.000 1010.160 ;
        RECT 4.400 1008.760 2481.600 1008.800 ;
        RECT 4.000 1007.400 2481.600 1008.760 ;
        RECT 4.000 922.440 2482.000 1007.400 ;
        RECT 4.400 921.040 2482.000 922.440 ;
        RECT 4.000 902.720 2482.000 921.040 ;
        RECT 4.000 901.320 2481.600 902.720 ;
        RECT 4.000 834.040 2482.000 901.320 ;
        RECT 4.400 832.640 2482.000 834.040 ;
        RECT 4.000 796.640 2482.000 832.640 ;
        RECT 4.000 795.240 2481.600 796.640 ;
        RECT 4.000 746.320 2482.000 795.240 ;
        RECT 4.400 744.920 2482.000 746.320 ;
        RECT 4.000 690.560 2482.000 744.920 ;
        RECT 4.000 689.160 2481.600 690.560 ;
        RECT 4.000 658.600 2482.000 689.160 ;
        RECT 4.400 657.200 2482.000 658.600 ;
        RECT 4.000 584.480 2482.000 657.200 ;
        RECT 4.000 583.080 2481.600 584.480 ;
        RECT 4.000 570.880 2482.000 583.080 ;
        RECT 4.400 569.480 2482.000 570.880 ;
        RECT 4.000 483.160 2482.000 569.480 ;
        RECT 4.400 481.760 2482.000 483.160 ;
        RECT 4.000 478.400 2482.000 481.760 ;
        RECT 4.000 477.000 2481.600 478.400 ;
        RECT 4.000 395.440 2482.000 477.000 ;
        RECT 4.400 394.040 2482.000 395.440 ;
        RECT 4.000 372.320 2482.000 394.040 ;
        RECT 4.000 370.920 2481.600 372.320 ;
        RECT 4.000 307.720 2482.000 370.920 ;
        RECT 4.400 306.320 2482.000 307.720 ;
        RECT 4.000 266.240 2482.000 306.320 ;
        RECT 4.000 264.840 2481.600 266.240 ;
        RECT 4.000 220.000 2482.000 264.840 ;
        RECT 4.400 218.600 2482.000 220.000 ;
        RECT 4.000 160.160 2482.000 218.600 ;
        RECT 4.000 158.760 2481.600 160.160 ;
        RECT 4.000 132.280 2482.000 158.760 ;
        RECT 4.400 130.880 2482.000 132.280 ;
        RECT 4.000 54.080 2482.000 130.880 ;
        RECT 4.000 52.680 2481.600 54.080 ;
        RECT 4.000 44.560 2482.000 52.680 ;
        RECT 4.400 43.695 2482.000 44.560 ;
      LAYER met4 ;
        RECT 64.695 76.335 2434.945 2541.360 ;
      LAYER met5 ;
        RECT 5.520 155.080 2480.320 2526.680 ;
  END
END fpga_core
END LIBRARY

