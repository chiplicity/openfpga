VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__2_
  CLASS BLOCK ;
  FOREIGN cbx_1__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 119.130 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 116.730 56.030 119.130 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 116.730 93.750 119.130 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.370 2.400 60.970 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.290 2.400 90.890 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.010 2.400 93.610 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.730 2.400 96.330 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.130 2.400 99.730 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.850 2.400 102.450 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.250 2.400 105.850 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.970 2.400 108.570 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.690 2.400 111.290 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.090 2.400 114.690 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.810 2.400 117.410 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.090 2.400 63.690 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.810 2.400 66.410 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.210 2.400 69.810 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.930 2.400 72.530 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.330 2.400 75.930 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.050 2.400 78.650 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.770 2.400 81.370 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.170 2.400 84.770 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.890 2.400 87.490 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.530 2.400 1.130 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.450 2.400 31.050 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.170 2.400 33.770 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.890 2.400 36.490 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.290 2.400 39.890 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.010 2.400 42.610 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.410 2.400 46.010 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.130 2.400 48.730 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.850 2.400 51.450 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.250 2.400 54.850 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.970 2.400 57.570 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.250 2.400 3.850 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.970 2.400 6.570 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.370 2.400 9.970 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.090 2.400 12.690 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.490 2.400 16.090 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.210 2.400 18.810 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.930 2.400 21.530 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.330 2.400 24.930 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.050 2.400 27.650 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 60.370 150.000 60.970 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 90.290 150.000 90.890 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 93.010 150.000 93.610 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 95.730 150.000 96.330 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 99.130 150.000 99.730 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 101.850 150.000 102.450 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 105.250 150.000 105.850 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 107.970 150.000 108.570 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 110.690 150.000 111.290 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 114.090 150.000 114.690 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 116.810 150.000 117.410 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 63.090 150.000 63.690 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 65.810 150.000 66.410 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 69.210 150.000 69.810 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 71.930 150.000 72.530 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 75.330 150.000 75.930 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 78.050 150.000 78.650 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 80.770 150.000 81.370 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 84.170 150.000 84.770 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 86.890 150.000 87.490 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 0.530 150.000 1.130 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 30.450 150.000 31.050 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 33.170 150.000 33.770 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 35.890 150.000 36.490 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 39.290 150.000 39.890 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 42.010 150.000 42.610 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 45.410 150.000 46.010 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 48.130 150.000 48.730 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 50.850 150.000 51.450 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 54.250 150.000 54.850 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 56.970 150.000 57.570 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 3.250 150.000 3.850 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 5.970 150.000 6.570 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 9.370 150.000 9.970 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 12.090 150.000 12.690 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 15.490 150.000 16.090 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 18.210 150.000 18.810 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 20.930 150.000 21.530 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 24.330 150.000 24.930 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 27.050 150.000 27.650 ;
    END
  END chanx_right_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 116.730 18.770 119.130 ;
    END
  END prog_clk
  PIN top_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 116.730 131.010 119.130 ;
    END
  END top_grid_pin_0_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.720 9.770 31.320 108.170 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 54.720 9.770 56.320 108.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 9.925 144.440 108.015 ;
      LAYER met1 ;
        RECT 5.520 9.770 144.440 108.170 ;
      LAYER met2 ;
        RECT 6.990 116.450 18.210 117.295 ;
        RECT 19.050 116.450 55.470 117.295 ;
        RECT 56.310 116.450 93.190 117.295 ;
        RECT 94.030 116.450 130.450 117.295 ;
        RECT 6.990 0.645 131.260 116.450 ;
      LAYER met3 ;
        RECT 2.800 116.410 147.200 117.275 ;
        RECT 2.400 115.090 147.600 116.410 ;
        RECT 2.800 113.690 147.200 115.090 ;
        RECT 2.400 111.690 147.600 113.690 ;
        RECT 2.800 110.290 147.200 111.690 ;
        RECT 2.400 108.970 147.600 110.290 ;
        RECT 2.800 107.570 147.200 108.970 ;
        RECT 2.400 106.250 147.600 107.570 ;
        RECT 2.800 104.850 147.200 106.250 ;
        RECT 2.400 102.850 147.600 104.850 ;
        RECT 2.800 101.450 147.200 102.850 ;
        RECT 2.400 100.130 147.600 101.450 ;
        RECT 2.800 98.730 147.200 100.130 ;
        RECT 2.400 96.730 147.600 98.730 ;
        RECT 2.800 95.330 147.200 96.730 ;
        RECT 2.400 94.010 147.600 95.330 ;
        RECT 2.800 92.610 147.200 94.010 ;
        RECT 2.400 91.290 147.600 92.610 ;
        RECT 2.800 89.890 147.200 91.290 ;
        RECT 2.400 87.890 147.600 89.890 ;
        RECT 2.800 86.490 147.200 87.890 ;
        RECT 2.400 85.170 147.600 86.490 ;
        RECT 2.800 83.770 147.200 85.170 ;
        RECT 2.400 81.770 147.600 83.770 ;
        RECT 2.800 80.370 147.200 81.770 ;
        RECT 2.400 79.050 147.600 80.370 ;
        RECT 2.800 77.650 147.200 79.050 ;
        RECT 2.400 76.330 147.600 77.650 ;
        RECT 2.800 74.930 147.200 76.330 ;
        RECT 2.400 72.930 147.600 74.930 ;
        RECT 2.800 71.530 147.200 72.930 ;
        RECT 2.400 70.210 147.600 71.530 ;
        RECT 2.800 68.810 147.200 70.210 ;
        RECT 2.400 66.810 147.600 68.810 ;
        RECT 2.800 65.410 147.200 66.810 ;
        RECT 2.400 64.090 147.600 65.410 ;
        RECT 2.800 62.690 147.200 64.090 ;
        RECT 2.400 61.370 147.600 62.690 ;
        RECT 2.800 59.970 147.200 61.370 ;
        RECT 2.400 57.970 147.600 59.970 ;
        RECT 2.800 56.570 147.200 57.970 ;
        RECT 2.400 55.250 147.600 56.570 ;
        RECT 2.800 53.850 147.200 55.250 ;
        RECT 2.400 51.850 147.600 53.850 ;
        RECT 2.800 50.450 147.200 51.850 ;
        RECT 2.400 49.130 147.600 50.450 ;
        RECT 2.800 47.730 147.200 49.130 ;
        RECT 2.400 46.410 147.600 47.730 ;
        RECT 2.800 45.010 147.200 46.410 ;
        RECT 2.400 43.010 147.600 45.010 ;
        RECT 2.800 41.610 147.200 43.010 ;
        RECT 2.400 40.290 147.600 41.610 ;
        RECT 2.800 38.890 147.200 40.290 ;
        RECT 2.400 36.890 147.600 38.890 ;
        RECT 2.800 35.490 147.200 36.890 ;
        RECT 2.400 34.170 147.600 35.490 ;
        RECT 2.800 32.770 147.200 34.170 ;
        RECT 2.400 31.450 147.600 32.770 ;
        RECT 2.800 30.050 147.200 31.450 ;
        RECT 2.400 28.050 147.600 30.050 ;
        RECT 2.800 26.650 147.200 28.050 ;
        RECT 2.400 25.330 147.600 26.650 ;
        RECT 2.800 23.930 147.200 25.330 ;
        RECT 2.400 21.930 147.600 23.930 ;
        RECT 2.800 20.530 147.200 21.930 ;
        RECT 2.400 19.210 147.600 20.530 ;
        RECT 2.800 17.810 147.200 19.210 ;
        RECT 2.400 16.490 147.600 17.810 ;
        RECT 2.800 15.090 147.200 16.490 ;
        RECT 2.400 13.090 147.600 15.090 ;
        RECT 2.800 11.690 147.200 13.090 ;
        RECT 2.400 10.370 147.600 11.690 ;
        RECT 2.800 8.970 147.200 10.370 ;
        RECT 2.400 6.970 147.600 8.970 ;
        RECT 2.800 5.570 147.200 6.970 ;
        RECT 2.400 4.250 147.600 5.570 ;
        RECT 2.800 2.850 147.200 4.250 ;
        RECT 2.400 1.530 147.600 2.850 ;
        RECT 2.800 0.130 147.200 1.530 ;
        RECT 2.400 0.000 147.600 0.130 ;
      LAYER met4 ;
        RECT 79.720 9.770 131.320 108.170 ;
  END
END cbx_1__2_
END LIBRARY

