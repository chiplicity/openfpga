* NGSPICE file created from grid_io_top.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_and4_4 abstract view
.subckt scs8hd_and4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

.subckt grid_io_top address[0] address[1] address[2] address[3] bottom_width_0_height_0__pin_0_
+ bottom_width_0_height_0__pin_10_ bottom_width_0_height_0__pin_11_ bottom_width_0_height_0__pin_12_
+ bottom_width_0_height_0__pin_13_ bottom_width_0_height_0__pin_14_ bottom_width_0_height_0__pin_15_
+ bottom_width_0_height_0__pin_1_ bottom_width_0_height_0__pin_2_ bottom_width_0_height_0__pin_3_
+ bottom_width_0_height_0__pin_4_ bottom_width_0_height_0__pin_5_ bottom_width_0_height_0__pin_6_
+ bottom_width_0_height_0__pin_7_ bottom_width_0_height_0__pin_8_ bottom_width_0_height_0__pin_9_
+ data_in enable gfpga_pad_GPIO_PAD[0] gfpga_pad_GPIO_PAD[1] gfpga_pad_GPIO_PAD[2]
+ gfpga_pad_GPIO_PAD[3] gfpga_pad_GPIO_PAD[4] gfpga_pad_GPIO_PAD[5] gfpga_pad_GPIO_PAD[6]
+ gfpga_pad_GPIO_PAD[7] vpwr vgnd
XFILLER_22_166 vgnd vpwr scs8hd_decap_12
XFILLER_9_159 vgnd vpwr scs8hd_decap_12
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_23_86 vgnd vpwr scs8hd_decap_12
XFILLER_2_154 vgnd vpwr scs8hd_decap_8
XFILLER_2_198 vgnd vpwr scs8hd_decap_8
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XFILLER_29_74 vgnd vpwr scs8hd_decap_12
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_227 vgnd vpwr scs8hd_decap_3
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_15_98 vgnd vpwr scs8hd_decap_12
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_12
XFILLER_22_178 vgnd vpwr scs8hd_decap_12
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_5_196 vpwr vgnd scs8hd_fill_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
XFILLER_23_98 vgnd vpwr scs8hd_decap_12
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XFILLER_2_177 vpwr vgnd scs8hd_fill_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XFILLER_11_232 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _09_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_29_86 vgnd vpwr scs8hd_decap_12
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_4_206 vpwr vgnd scs8hd_fill_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_110 vgnd vpwr scs8hd_decap_12
XFILLER_1_209 vpwr vgnd scs8hd_fill_2
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vgnd vpwr scs8hd_decap_12
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_253 vgnd vpwr scs8hd_decap_12
XFILLER_39_257 vgnd vpwr scs8hd_decap_12
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_135 vgnd vpwr scs8hd_decap_12
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XFILLER_12_190 vgnd vpwr scs8hd_decap_12
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XFILLER_29_98 vgnd vpwr scs8hd_decap_12
XFILLER_28_141 vgnd vpwr scs8hd_decap_12
XFILLER_3_240 vgnd vpwr scs8hd_decap_4
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_16_166 vgnd vpwr scs8hd_decap_12
XANTENNA__04__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_265 vgnd vpwr scs8hd_decap_12
XFILLER_39_269 vgnd vpwr scs8hd_decap_8
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_147 vgnd vpwr scs8hd_decap_12
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_10_117 vgnd vpwr scs8hd_decap_12
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XFILLER_23_220 vgnd vpwr scs8hd_decap_12
XANTENNA__12__A _07_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XANTENNA__07__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XFILLER_4_219 vpwr vgnd scs8hd_fill_2
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XFILLER_0_244 vgnd vpwr scs8hd_fill_1
XFILLER_0_222 vgnd vpwr scs8hd_fill_1
XFILLER_31_159 vgnd vpwr scs8hd_decap_12
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_178 vgnd vpwr scs8hd_decap_12
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_159 vgnd vpwr scs8hd_decap_12
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XFILLER_8_141 vgnd vpwr scs8hd_decap_12
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_232 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch/Q
+ _10_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__12__B _05_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_20_202 vgnd vpwr scs8hd_decap_12
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
XANTENNA__07__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_6_272 vgnd vpwr scs8hd_decap_3
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XFILLER_19_110 vgnd vpwr scs8hd_decap_12
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_25_135 vgnd vpwr scs8hd_decap_12
XFILLER_24_190 vgnd vpwr scs8hd_decap_12
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_105 vgnd vpwr scs8hd_decap_12
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
XFILLER_21_171 vgnd vpwr scs8hd_decap_12
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XANTENNA__12__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
XANTENNA__07__C _07_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_240 vgnd vpwr scs8hd_decap_12
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_3_221 vpwr vgnd scs8hd_fill_2
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_202 vpwr vgnd scs8hd_fill_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_117 vgnd vpwr scs8hd_decap_12
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_190 vpwr vgnd scs8hd_fill_2
XANTENNA__12__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XANTENNA__07__D enable vgnd vpwr scs8hd_diode_2
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_252 vgnd vpwr scs8hd_decap_12
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_28_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_159 vgnd vpwr scs8hd_decap_12
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
X_09_ _07_/C enable address[3] _08_/D _09_/X vgnd vpwr scs8hd_and4_4
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_225 vpwr vgnd scs8hd_fill_2
XFILLER_0_214 vgnd vpwr scs8hd_fill_1
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_129 vgnd vpwr scs8hd_decap_12
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XFILLER_14_202 vgnd vpwr scs8hd_decap_12
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XFILLER_20_227 vgnd vpwr scs8hd_decap_12
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_264 vgnd vpwr scs8hd_decap_8
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_135 vgnd vpwr scs8hd_decap_12
X_08_ address[1] enable address[3] _08_/D _08_/X vgnd vpwr scs8hd_and4_4
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XFILLER_18_190 vgnd vpwr scs8hd_decap_12
XFILLER_16_105 vgnd vpwr scs8hd_decap_12
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_208 vgnd vpwr scs8hd_decap_12
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_171 vgnd vpwr scs8hd_decap_12
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_12_141 vgnd vpwr scs8hd_decap_12
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
XFILLER_4_170 vgnd vpwr scs8hd_fill_1
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XFILLER_1_162 vpwr vgnd scs8hd_fill_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_239 vgnd vpwr scs8hd_decap_12
XFILLER_24_93 vgnd vpwr scs8hd_decap_12
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_147 vgnd vpwr scs8hd_decap_12
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XFILLER_0_249 vpwr vgnd scs8hd_fill_2
X_07_ address[3] address[2] _07_/C enable _07_/X vgnd vpwr scs8hd_and4_4
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_117 vgnd vpwr scs8hd_decap_12
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _10_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XFILLER_19_159 vgnd vpwr scs8hd_decap_12
XFILLER_3_236 vpwr vgnd scs8hd_fill_2
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_206 vgnd vpwr scs8hd_decap_8
X_06_ address[3] address[2] address[1] enable _06_/X vgnd vpwr scs8hd_and4_4
XFILLER_21_62 vgnd vpwr scs8hd_decap_12
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_129 vgnd vpwr scs8hd_decap_12
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XFILLER_21_110 vgnd vpwr scs8hd_decap_12
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
XFILLER_12_154 vgnd vpwr scs8hd_decap_12
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_202 vgnd vpwr scs8hd_decap_12
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_194 vgnd vpwr scs8hd_decap_12
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
Xlogical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch/Q
+ _06_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
XFILLER_27_171 vgnd vpwr scs8hd_decap_12
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_204 vpwr vgnd scs8hd_fill_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
X_05_ enable _05_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_141 vgnd vpwr scs8hd_decap_12
XFILLER_21_74 vgnd vpwr scs8hd_decap_12
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_218 vgnd vpwr scs8hd_decap_4
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XFILLER_12_166 vgnd vpwr scs8hd_decap_12
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
XFILLER_13_86 vgnd vpwr scs8hd_decap_12
XFILLER_9_232 vgnd vpwr scs8hd_decap_12
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
XFILLER_6_224 vpwr vgnd scs8hd_fill_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_12
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_04_ address[2] _08_/D vgnd vpwr scs8hd_inv_8
Xlogical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch/Q
+ _11_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XFILLER_21_86 vgnd vpwr scs8hd_decap_12
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XFILLER_12_178 vgnd vpwr scs8hd_decap_12
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_7_171 vgnd vpwr scs8hd_decap_12
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_74 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XFILLER_22_251 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_98 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_129 vgnd vpwr scs8hd_decap_12
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_217 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_19_86 vgnd vpwr scs8hd_decap_12
X_03_ address[1] _07_/C vgnd vpwr scs8hd_inv_8
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_12
XFILLER_21_98 vgnd vpwr scs8hd_decap_12
XFILLER_15_110 vgnd vpwr scs8hd_decap_12
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_135 vgnd vpwr scs8hd_decap_12
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_190 vgnd vpwr scs8hd_decap_12
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _06_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_86 vgnd vpwr scs8hd_decap_12
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XFILLER_23_208 vgnd vpwr scs8hd_decap_12
XFILLER_22_263 vgnd vpwr scs8hd_decap_12
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XFILLER_39_171 vgnd vpwr scs8hd_decap_12
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_19_98 vgnd vpwr scs8hd_decap_12
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_18_141 vgnd vpwr scs8hd_decap_12
XFILLER_24_166 vgnd vpwr scs8hd_decap_12
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XFILLER_21_147 vgnd vpwr scs8hd_decap_12
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
XFILLER_27_98 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XFILLER_24_178 vgnd vpwr scs8hd_decap_12
XANTENNA__10__A _07_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_21_159 vgnd vpwr scs8hd_decap_12
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XANTENNA__05__A enable vgnd vpwr scs8hd_diode_2
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_166 vgnd vpwr scs8hd_decap_4
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_232 vgnd vpwr scs8hd_decap_12
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_202 vgnd vpwr scs8hd_decap_12
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XANTENNA__13__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_228 vgnd vpwr scs8hd_decap_12
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_27_110 vgnd vpwr scs8hd_decap_12
XANTENNA__08__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
XFILLER_15_135 vgnd vpwr scs8hd_decap_12
XANTENNA__10__B _05_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_14_190 vgnd vpwr scs8hd_decap_12
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XFILLER_11_171 vgnd vpwr scs8hd_decap_12
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_159 vgnd vpwr scs8hd_fill_1
XFILLER_39_196 vgnd vpwr scs8hd_decap_12
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_24_68 vgnd vpwr scs8hd_decap_12
XANTENNA__13__B _05_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XANTENNA__08__B enable vgnd vpwr scs8hd_diode_2
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XFILLER_18_166 vgnd vpwr scs8hd_decap_12
XFILLER_2_210 vgnd vpwr scs8hd_decap_4
XFILLER_2_232 vpwr vgnd scs8hd_fill_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_147 vgnd vpwr scs8hd_decap_12
XANTENNA__10__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
XFILLER_25_220 vgnd vpwr scs8hd_decap_12
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XANTENNA__13__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
XFILLER_5_230 vpwr vgnd scs8hd_fill_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
XANTENNA__08__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XFILLER_18_178 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _11_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_159 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch/Q
+ _07_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__10__D _08_/D vgnd vpwr scs8hd_diode_2
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_129 vgnd vpwr scs8hd_decap_12
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_80 vgnd vpwr scs8hd_decap_12
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XFILLER_25_232 vgnd vpwr scs8hd_decap_12
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_22_202 vgnd vpwr scs8hd_decap_12
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XANTENNA__13__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_5_242 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_27_135 vgnd vpwr scs8hd_decap_12
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XANTENNA__08__D _08_/D vgnd vpwr scs8hd_diode_2
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_190 vgnd vpwr scs8hd_decap_12
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_105 vgnd vpwr scs8hd_decap_12
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
XFILLER_23_171 vgnd vpwr scs8hd_decap_12
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_20_141 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch/Q
+ _12_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XFILLER_28_80 vgnd vpwr scs8hd_decap_12
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_147 vgnd vpwr scs8hd_decap_12
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_117 vgnd vpwr scs8hd_decap_12
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_93 vgnd vpwr scs8hd_decap_12
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_174 vpwr vgnd scs8hd_fill_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_27_159 vgnd vpwr scs8hd_decap_12
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_236 vpwr vgnd scs8hd_fill_2
XFILLER_24_129 vgnd vpwr scs8hd_decap_12
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XFILLER_20_154 vgnd vpwr scs8hd_decap_12
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XFILLER_11_110 vgnd vpwr scs8hd_decap_12
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _07_/X vgnd vpwr scs8hd_diode_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_202 vgnd vpwr scs8hd_decap_12
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XFILLER_0_164 vgnd vpwr scs8hd_decap_8
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_39_135 vgnd vpwr scs8hd_decap_12
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XFILLER_5_234 vgnd vpwr scs8hd_decap_8
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_18_105 vgnd vpwr scs8hd_decap_12
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XFILLER_17_171 vgnd vpwr scs8hd_decap_12
XFILLER_1_270 vgnd vpwr scs8hd_decap_6
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_141 vgnd vpwr scs8hd_decap_12
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_166 vgnd vpwr scs8hd_decap_12
XFILLER_7_159 vgnd vpwr scs8hd_decap_12
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_239 vgnd vpwr scs8hd_decap_12
XFILLER_3_195 vpwr vgnd scs8hd_fill_2
XFILLER_0_198 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_147 vgnd vpwr scs8hd_decap_12
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_5_213 vpwr vgnd scs8hd_fill_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XFILLER_18_117 vgnd vpwr scs8hd_decap_12
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_178 vgnd vpwr scs8hd_decap_12
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_74 vgnd vpwr scs8hd_decap_12
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_3_163 vgnd vpwr scs8hd_fill_1
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XFILLER_12_251 vgnd vpwr scs8hd_decap_12
XFILLER_39_159 vgnd vpwr scs8hd_decap_12
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_2_206 vpwr vgnd scs8hd_fill_2
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_74 vgnd vpwr scs8hd_decap_12
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
XFILLER_23_110 vgnd vpwr scs8hd_decap_12
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
XFILLER_11_98 vgnd vpwr scs8hd_decap_12
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_28_202 vgnd vpwr scs8hd_decap_12
XFILLER_11_135 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_190 vgnd vpwr scs8hd_decap_12
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_86 vgnd vpwr scs8hd_decap_12
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_6
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_171 vgnd vpwr scs8hd_decap_12
XFILLER_5_226 vpwr vgnd scs8hd_fill_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_decap_12
XFILLER_25_86 vgnd vpwr scs8hd_decap_12
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_14_166 vgnd vpwr scs8hd_decap_12
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XFILLER_11_147 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_98 vgnd vpwr scs8hd_decap_12
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch/Q
+ _08_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_98 vgnd vpwr scs8hd_decap_12
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XFILLER_23_123 vgnd vpwr scs8hd_decap_12
XFILLER_14_178 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _12_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XFILLER_9_171 vgnd vpwr scs8hd_decap_12
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XFILLER_11_159 vgnd vpwr scs8hd_decap_12
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_199 vgnd vpwr scs8hd_decap_3
XFILLER_21_232 vgnd vpwr scs8hd_decap_12
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XANTENNA__03__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch/Q
+ _13_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_12
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XFILLER_17_110 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_135 vgnd vpwr scs8hd_decap_12
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XFILLER_22_190 vgnd vpwr scs8hd_decap_12
XFILLER_20_105 vgnd vpwr scs8hd_decap_12
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_22_56 vgnd vpwr scs8hd_decap_12
XANTENNA__11__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XFILLER_25_208 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XANTENNA__06__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XFILLER_4_273 vpwr vgnd scs8hd_fill_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_166 vgnd vpwr scs8hd_decap_12
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XFILLER_1_221 vpwr vgnd scs8hd_fill_2
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_254 vpwr vgnd scs8hd_fill_2
XFILLER_1_276 vgnd vpwr scs8hd_fill_1
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_23_147 vgnd vpwr scs8hd_decap_12
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XANTENNA__09__A _07_/C vgnd vpwr scs8hd_diode_2
XFILLER_20_117 vgnd vpwr scs8hd_decap_12
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_22_68 vgnd vpwr scs8hd_decap_12
XANTENNA__11__B _05_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XANTENNA__06__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XFILLER_21_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_4_241 vgnd vpwr scs8hd_decap_12
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_26_178 vgnd vpwr scs8hd_decap_12
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_23_159 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XANTENNA__09__B enable vgnd vpwr scs8hd_diode_2
XFILLER_20_129 vgnd vpwr scs8hd_decap_12
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
XANTENNA__11__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
X_13_ address[1] _05_/Y address[3] address[2] _13_/Y vgnd vpwr scs8hd_nor4_4
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XANTENNA__06__C address[1] vgnd vpwr scs8hd_diode_2
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _08_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XFILLER_21_257 vgnd vpwr scs8hd_decap_12
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_12_202 vgnd vpwr scs8hd_decap_12
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_110 vgnd vpwr scs8hd_decap_12
XFILLER_5_209 vpwr vgnd scs8hd_fill_2
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XFILLER_20_80 vgnd vpwr scs8hd_decap_12
XFILLER_4_253 vgnd vpwr scs8hd_decap_12
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XPHY_69 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XFILLER_1_201 vpwr vgnd scs8hd_fill_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_17_135 vgnd vpwr scs8hd_decap_12
XFILLER_31_171 vgnd vpwr scs8hd_decap_12
XFILLER_16_190 vgnd vpwr scs8hd_decap_12
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XANTENNA__09__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_13_171 vgnd vpwr scs8hd_decap_12
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_141 vgnd vpwr scs8hd_decap_12
XANTENNA__11__D _08_/D vgnd vpwr scs8hd_diode_2
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
X_12_ _07_/C _05_/Y address[3] address[2] _12_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_159 vgnd vpwr scs8hd_decap_4
XANTENNA__06__D enable vgnd vpwr scs8hd_diode_2
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XFILLER_18_80 vgnd vpwr scs8hd_decap_12
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XFILLER_4_210 vgnd vpwr scs8hd_decap_4
XFILLER_4_265 vgnd vpwr scs8hd_decap_8
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XFILLER_17_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_213 vpwr vgnd scs8hd_fill_2
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
XFILLER_14_117 vgnd vpwr scs8hd_decap_12
XANTENNA__09__D _08_/D vgnd vpwr scs8hd_diode_2
XFILLER_26_80 vgnd vpwr scs8hd_decap_12
XFILLER_9_110 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
X_11_ address[1] _05_/Y address[3] _08_/D _11_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XFILLER_20_93 vgnd vpwr scs8hd_decap_12
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_159 vgnd vpwr scs8hd_decap_12
XFILLER_1_236 vpwr vgnd scs8hd_fill_2
XFILLER_1_258 vgnd vpwr scs8hd_decap_12
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_129 vgnd vpwr scs8hd_decap_12
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_232 vgnd vpwr scs8hd_decap_12
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_10_154 vgnd vpwr scs8hd_decap_12
X_10_ _07_/C _05_/Y address[3] _08_/D _10_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XFILLER_4_223 vpwr vgnd scs8hd_fill_2
XFILLER_28_190 vgnd vpwr scs8hd_decap_12
XFILLER_26_105 vgnd vpwr scs8hd_decap_12
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_171 vgnd vpwr scs8hd_decap_12
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
Xlogical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch/Q
+ _09_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_22_141 vgnd vpwr scs8hd_decap_12
XFILLER_26_93 vgnd vpwr scs8hd_decap_12
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
XFILLER_10_166 vgnd vpwr scs8hd_decap_12
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_2_173 vpwr vgnd scs8hd_fill_2
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_232 vgnd vpwr scs8hd_decap_12
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_29_147 vgnd vpwr scs8hd_decap_12
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_117 vgnd vpwr scs8hd_decap_12
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_1_205 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_39_220 vgnd vpwr scs8hd_decap_12
XFILLER_9_135 vgnd vpwr scs8hd_decap_12
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
XFILLER_27_245 vgnd vpwr scs8hd_decap_12
XFILLER_10_178 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _13_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XFILLER_23_62 vgnd vpwr scs8hd_decap_12
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
XFILLER_20_251 vgnd vpwr scs8hd_decap_12
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_129 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_1_217 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XFILLER_25_184 vgnd vpwr scs8hd_decap_12
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_39_232 vgnd vpwr scs8hd_decap_12
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_154 vgnd vpwr scs8hd_decap_12
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_13_110 vgnd vpwr scs8hd_decap_12
XFILLER_9_147 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XFILLER_18_202 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
XFILLER_23_74 vgnd vpwr scs8hd_decap_12
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_20_263 vgnd vpwr scs8hd_decap_12
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
XFILLER_4_215 vpwr vgnd scs8hd_fill_2
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_25_196 vgnd vpwr scs8hd_decap_12
XFILLER_15_86 vgnd vpwr scs8hd_decap_12
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_141 vgnd vpwr scs8hd_decap_12
XFILLER_0_240 vgnd vpwr scs8hd_decap_4
.ends

