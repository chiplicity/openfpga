magic
tech sky130A
magscale 1 2
timestamp 1604675407
<< locali >>
rect 28785 145215 28819 146881
rect 36145 142087 36179 142597
rect 43965 142087 43999 142529
rect 48197 142087 48231 142529
rect 51693 142087 51727 142257
rect 132101 137429 132285 137463
rect 132101 136987 132135 137429
rect 132377 137191 132411 141849
rect 132101 136953 132285 136987
rect 132561 127399 132595 127569
rect 132561 114955 132595 118253
rect 132653 118151 132687 136953
rect 132745 117947 132779 127365
rect 222721 124815 222755 127501
rect 132561 113731 132595 114921
rect 132653 113799 132687 117709
rect 132745 110263 132779 115057
rect 222813 107951 222847 110229
rect 54821 86123 54855 90237
rect 54821 76467 54855 85953
rect 35961 69259 35995 69497
rect 35961 69225 36053 69259
rect 36145 68647 36179 69225
rect 54821 68647 54855 69361
rect 55189 68851 55223 69293
rect 123821 68579 123855 68749
rect 222537 28187 222571 37741
<< viali >>
rect 28785 146881 28819 146915
rect 28785 145181 28819 145215
rect 36145 142597 36179 142631
rect 36145 142053 36179 142087
rect 43965 142529 43999 142563
rect 43965 142053 43999 142087
rect 48197 142529 48231 142563
rect 48197 142053 48231 142087
rect 51693 142257 51727 142291
rect 51693 142053 51727 142087
rect 132377 141849 132411 141883
rect 132285 137429 132319 137463
rect 132377 137157 132411 137191
rect 132285 136953 132319 136987
rect 132653 136953 132687 136987
rect 132561 127569 132595 127603
rect 132561 127365 132595 127399
rect 132561 118253 132595 118287
rect 222721 127501 222755 127535
rect 132653 118117 132687 118151
rect 132745 127365 132779 127399
rect 222721 124781 222755 124815
rect 132745 117913 132779 117947
rect 132561 114921 132595 114955
rect 132653 117709 132687 117743
rect 132653 113765 132687 113799
rect 132745 115057 132779 115091
rect 132561 113697 132595 113731
rect 132745 110229 132779 110263
rect 222813 110229 222847 110263
rect 222813 107917 222847 107951
rect 54821 90237 54855 90271
rect 54821 86089 54855 86123
rect 54821 85953 54855 85987
rect 54821 76433 54855 76467
rect 35961 69497 35995 69531
rect 54821 69361 54855 69395
rect 36053 69225 36087 69259
rect 36145 69225 36179 69259
rect 36145 68613 36179 68647
rect 55189 69293 55223 69327
rect 55189 68817 55223 68851
rect 54821 68613 54855 68647
rect 123821 68749 123855 68783
rect 123821 68545 123855 68579
rect 222537 37741 222571 37775
rect 222537 28153 222571 28187
<< metal1 >>
rect 23526 244860 23532 244912
rect 23584 244900 23590 244912
rect 70538 244900 70544 244912
rect 23584 244872 70544 244900
rect 23584 244860 23590 244872
rect 70538 244860 70544 244872
rect 70596 244860 70602 244912
rect 105222 244860 105228 244912
rect 105280 244900 105286 244912
rect 149658 244900 149664 244912
rect 105280 244872 149664 244900
rect 105280 244860 105286 244872
rect 149658 244860 149664 244872
rect 149716 244860 149722 244912
rect 50758 244792 50764 244844
rect 50816 244832 50822 244844
rect 142390 244832 142396 244844
rect 50816 244804 142396 244832
rect 50816 244792 50822 244804
rect 142390 244792 142396 244804
rect 142448 244792 142454 244844
rect 157478 244792 157484 244844
rect 157536 244832 157542 244844
rect 159778 244832 159784 244844
rect 157536 244804 159784 244832
rect 157536 244792 157542 244804
rect 159778 244792 159784 244804
rect 159836 244792 159842 244844
rect 85626 242412 85632 242464
rect 85684 242412 85690 242464
rect 85644 242180 85672 242412
rect 132546 242180 132552 242192
rect 85644 242152 132552 242180
rect 132546 242140 132552 242152
rect 132604 242140 132610 242192
rect 165298 242140 165304 242192
rect 165356 242180 165362 242192
rect 214242 242180 214248 242192
rect 165356 242152 214248 242180
rect 165356 242140 165362 242152
rect 214242 242140 214248 242152
rect 214300 242140 214306 242192
rect 93354 242072 93360 242124
rect 93412 242112 93418 242124
rect 187010 242112 187016 242124
rect 93412 242084 187016 242112
rect 93412 242072 93418 242084
rect 187010 242072 187016 242084
rect 187068 242072 187074 242124
rect 167782 229764 167788 229816
rect 167840 229804 167846 229816
rect 168518 229804 168524 229816
rect 167840 229776 168524 229804
rect 167840 229764 167846 229776
rect 168518 229764 168524 229776
rect 168576 229764 168582 229816
rect 207250 223372 207256 223424
rect 207308 223412 207314 223424
rect 223074 223412 223080 223424
rect 207308 223384 223080 223412
rect 207308 223372 207314 223384
rect 223074 223372 223080 223384
rect 223132 223372 223138 223424
rect 170082 222760 170088 222812
rect 170140 222800 170146 222812
rect 207250 222800 207256 222812
rect 170140 222772 207256 222800
rect 170140 222760 170146 222772
rect 207250 222760 207256 222772
rect 207308 222760 207314 222812
rect 71366 217932 71372 217984
rect 71424 217972 71430 217984
rect 71424 217944 98460 217972
rect 71424 217932 71430 217944
rect 98432 217916 98460 217944
rect 143678 217932 143684 217984
rect 143736 217972 143742 217984
rect 170082 217972 170088 217984
rect 143736 217944 170088 217972
rect 143736 217932 143742 217944
rect 170082 217932 170088 217944
rect 170140 217932 170146 217984
rect 46526 217864 46532 217916
rect 46584 217904 46590 217916
rect 98230 217904 98236 217916
rect 46584 217876 98236 217904
rect 46584 217864 46590 217876
rect 98230 217864 98236 217876
rect 98288 217864 98294 217916
rect 98414 217864 98420 217916
rect 98472 217904 98478 217916
rect 109270 217904 109276 217916
rect 98472 217876 109276 217904
rect 98472 217864 98478 217876
rect 109270 217864 109276 217876
rect 109328 217864 109334 217916
rect 118838 217864 118844 217916
rect 118896 217904 118902 217916
rect 169990 217904 169996 217916
rect 118896 217876 169996 217904
rect 118896 217864 118902 217876
rect 169990 217864 169996 217876
rect 170048 217864 170054 217916
rect 109270 217252 109276 217304
rect 109328 217292 109334 217304
rect 143678 217292 143684 217304
rect 109328 217264 143684 217292
rect 109328 217252 109334 217264
rect 143678 217252 143684 217264
rect 143736 217252 143742 217304
rect 37234 217184 37240 217236
rect 37292 217224 37298 217236
rect 71366 217224 71372 217236
rect 37292 217196 71372 217224
rect 37292 217184 37298 217196
rect 71366 217184 71372 217196
rect 71424 217184 71430 217236
rect 79370 217184 79376 217236
rect 79428 217224 79434 217236
rect 127762 217224 127768 217236
rect 79428 217196 127768 217224
rect 79428 217184 79434 217196
rect 127762 217184 127768 217196
rect 127820 217184 127826 217236
rect 81762 216572 81768 216624
rect 81820 216612 81826 216624
rect 93998 216612 94004 216624
rect 81820 216584 94004 216612
rect 81820 216572 81826 216584
rect 93998 216572 94004 216584
rect 94056 216572 94062 216624
rect 158582 216572 158588 216624
rect 158640 216612 158646 216624
rect 167230 216612 167236 216624
rect 158640 216584 167236 216612
rect 158640 216572 158646 216584
rect 167230 216572 167236 216584
rect 167288 216572 167294 216624
rect 91790 216504 91796 216556
rect 91848 216544 91854 216556
rect 102370 216544 102376 216556
rect 91848 216516 102376 216544
rect 91848 216504 91854 216516
rect 102370 216504 102376 216516
rect 102428 216504 102434 216556
rect 164102 216504 164108 216556
rect 164160 216544 164166 216556
rect 174222 216544 174228 216556
rect 164160 216516 174228 216544
rect 164160 216504 164166 216516
rect 174222 216504 174228 216516
rect 174280 216504 174286 216556
rect 86914 216436 86920 216488
rect 86972 216476 86978 216488
rect 98322 216476 98328 216488
rect 86972 216448 98328 216476
rect 86972 216436 86978 216448
rect 98322 216436 98328 216448
rect 98380 216436 98386 216488
rect 154074 216436 154080 216488
rect 154132 216476 154138 216488
rect 166034 216476 166040 216488
rect 154132 216448 166040 216476
rect 154132 216436 154138 216448
rect 166034 216436 166040 216448
rect 166092 216436 166098 216488
rect 62534 215756 62540 215808
rect 62592 215796 62598 215808
rect 71826 215796 71832 215808
rect 62592 215768 71832 215796
rect 62592 215756 62598 215768
rect 71826 215756 71832 215768
rect 71884 215756 71890 215808
rect 135398 215756 135404 215808
rect 135456 215796 135462 215808
rect 143770 215796 143776 215808
rect 135456 215768 143776 215796
rect 135456 215756 135462 215768
rect 143770 215756 143776 215768
rect 143828 215756 143834 215808
rect 100990 214600 100996 214652
rect 101048 214640 101054 214652
rect 102554 214640 102560 214652
rect 101048 214612 102560 214640
rect 101048 214600 101054 214612
rect 102554 214600 102560 214612
rect 102612 214600 102618 214652
rect 135398 214600 135404 214652
rect 135456 214640 135462 214652
rect 136778 214640 136784 214652
rect 135456 214612 136784 214640
rect 135456 214600 135462 214612
rect 136778 214600 136784 214612
rect 136836 214600 136842 214652
rect 62626 214532 62632 214584
rect 62684 214572 62690 214584
rect 65018 214572 65024 214584
rect 62684 214544 65024 214572
rect 62684 214532 62690 214544
rect 65018 214532 65024 214544
rect 65076 214532 65082 214584
rect 172014 213988 172020 214040
rect 172072 214028 172078 214040
rect 174038 214028 174044 214040
rect 172072 214000 174044 214028
rect 172072 213988 172078 214000
rect 174038 213988 174044 214000
rect 174096 213988 174102 214040
rect 135398 213648 135404 213700
rect 135456 213688 135462 213700
rect 136870 213688 136876 213700
rect 135456 213660 136876 213688
rect 135456 213648 135462 213660
rect 136870 213648 136876 213660
rect 136928 213648 136934 213700
rect 100990 213308 100996 213360
rect 101048 213348 101054 213360
rect 103106 213348 103112 213360
rect 101048 213320 103112 213348
rect 101048 213308 101054 213320
rect 103106 213308 103112 213320
rect 103164 213308 103170 213360
rect 62534 213240 62540 213292
rect 62592 213280 62598 213292
rect 65018 213280 65024 213292
rect 62592 213252 65024 213280
rect 62592 213240 62598 213252
rect 65018 213240 65024 213252
rect 65076 213240 65082 213292
rect 135030 213240 135036 213292
rect 135088 213280 135094 213292
rect 137054 213280 137060 213292
rect 135088 213252 137060 213280
rect 135088 213240 135094 213252
rect 137054 213240 137060 213252
rect 137112 213240 137118 213292
rect 102370 213144 102376 213156
rect 102296 213116 102376 213144
rect 63730 213036 63736 213088
rect 63788 213076 63794 213088
rect 66398 213076 66404 213088
rect 63788 213048 66404 213076
rect 63788 213036 63794 213048
rect 66398 213036 66404 213048
rect 66456 213036 66462 213088
rect 100530 213036 100536 213088
rect 100588 213076 100594 213088
rect 102296 213076 102324 213116
rect 102370 213104 102376 213116
rect 102428 213104 102434 213156
rect 174222 213144 174228 213156
rect 172768 213116 174228 213144
rect 100588 213048 102324 213076
rect 100588 213036 100594 213048
rect 172658 213036 172664 213088
rect 172716 213076 172722 213088
rect 172768 213076 172796 213116
rect 174222 213104 174228 213116
rect 174280 213104 174286 213156
rect 172716 213048 172796 213076
rect 172716 213036 172722 213048
rect 172658 212628 172664 212680
rect 172716 212668 172722 212680
rect 174038 212668 174044 212680
rect 172716 212640 174044 212668
rect 172716 212628 172722 212640
rect 174038 212628 174044 212640
rect 174096 212628 174102 212680
rect 135398 212152 135404 212204
rect 135456 212192 135462 212204
rect 136962 212192 136968 212204
rect 135456 212164 136968 212192
rect 135456 212152 135462 212164
rect 136962 212152 136968 212164
rect 137020 212152 137026 212204
rect 100990 211880 100996 211932
rect 101048 211920 101054 211932
rect 102370 211920 102376 211932
rect 101048 211892 102376 211920
rect 101048 211880 101054 211892
rect 102370 211880 102376 211892
rect 102428 211880 102434 211932
rect 135398 211880 135404 211932
rect 135456 211920 135462 211932
rect 136870 211920 136876 211932
rect 135456 211892 136876 211920
rect 135456 211880 135462 211892
rect 136870 211880 136876 211892
rect 136928 211880 136934 211932
rect 62350 211744 62356 211796
rect 62408 211784 62414 211796
rect 64926 211784 64932 211796
rect 62408 211756 64932 211784
rect 62408 211744 62414 211756
rect 64926 211744 64932 211756
rect 64984 211744 64990 211796
rect 62626 211676 62632 211728
rect 62684 211716 62690 211728
rect 65018 211716 65024 211728
rect 62684 211688 65024 211716
rect 62684 211676 62690 211688
rect 65018 211676 65024 211688
rect 65076 211676 65082 211728
rect 102462 211716 102468 211728
rect 102204 211688 102468 211716
rect 100806 211608 100812 211660
rect 100864 211648 100870 211660
rect 102204 211648 102232 211688
rect 102462 211676 102468 211688
rect 102520 211676 102526 211728
rect 172750 211676 172756 211728
rect 172808 211716 172814 211728
rect 174222 211716 174228 211728
rect 172808 211688 174228 211716
rect 172808 211676 172814 211688
rect 174222 211676 174228 211688
rect 174280 211676 174286 211728
rect 100864 211620 102232 211648
rect 100864 211608 100870 211620
rect 172382 211268 172388 211320
rect 172440 211308 172446 211320
rect 174038 211308 174044 211320
rect 172440 211280 174044 211308
rect 172440 211268 172446 211280
rect 174038 211268 174044 211280
rect 174096 211268 174102 211320
rect 62534 210792 62540 210844
rect 62592 210832 62598 210844
rect 65478 210832 65484 210844
rect 62592 210804 65484 210832
rect 62592 210792 62598 210804
rect 65478 210792 65484 210804
rect 65536 210792 65542 210844
rect 100898 210792 100904 210844
rect 100956 210832 100962 210844
rect 103658 210832 103664 210844
rect 100956 210804 103664 210832
rect 100956 210792 100962 210804
rect 103658 210792 103664 210804
rect 103716 210792 103722 210844
rect 172658 210588 172664 210640
rect 172716 210628 172722 210640
rect 174222 210628 174228 210640
rect 172716 210600 174228 210628
rect 172716 210588 172722 210600
rect 174222 210588 174228 210600
rect 174280 210588 174286 210640
rect 100990 210520 100996 210572
rect 101048 210560 101054 210572
rect 102370 210560 102376 210572
rect 101048 210532 102376 210560
rect 101048 210520 101054 210532
rect 102370 210520 102376 210532
rect 102428 210520 102434 210572
rect 134662 210520 134668 210572
rect 134720 210560 134726 210572
rect 136870 210560 136876 210572
rect 134720 210532 136876 210560
rect 134720 210520 134726 210532
rect 136870 210520 136876 210532
rect 136928 210520 136934 210572
rect 62626 210384 62632 210436
rect 62684 210424 62690 210436
rect 65018 210424 65024 210436
rect 62684 210396 65024 210424
rect 62684 210384 62690 210396
rect 65018 210384 65024 210396
rect 65076 210384 65082 210436
rect 207894 210316 207900 210368
rect 207952 210356 207958 210368
rect 223534 210356 223540 210368
rect 207952 210328 223540 210356
rect 207952 210316 207958 210328
rect 223534 210316 223540 210328
rect 223592 210316 223598 210368
rect 172658 210044 172664 210096
rect 172716 210084 172722 210096
rect 174038 210084 174044 210096
rect 172716 210056 174044 210084
rect 172716 210044 172722 210056
rect 174038 210044 174044 210056
rect 174096 210044 174102 210096
rect 62626 209840 62632 209892
rect 62684 209880 62690 209892
rect 66398 209880 66404 209892
rect 62684 209852 66404 209880
rect 62684 209840 62690 209852
rect 66398 209840 66404 209852
rect 66456 209840 66462 209892
rect 171646 209364 171652 209416
rect 171704 209404 171710 209416
rect 174130 209404 174136 209416
rect 171704 209376 174136 209404
rect 171704 209364 171710 209376
rect 174130 209364 174136 209376
rect 174188 209364 174194 209416
rect 62718 209024 62724 209076
rect 62776 209064 62782 209076
rect 65018 209064 65024 209076
rect 62776 209036 65024 209064
rect 62776 209024 62782 209036
rect 65018 209024 65024 209036
rect 65076 209024 65082 209076
rect 135306 209024 135312 209076
rect 135364 209064 135370 209076
rect 137698 209064 137704 209076
rect 135364 209036 137704 209064
rect 135364 209024 135370 209036
rect 137698 209024 137704 209036
rect 137756 209024 137762 209076
rect 174590 208996 174596 209008
rect 172768 208968 174596 208996
rect 172106 208888 172112 208940
rect 172164 208928 172170 208940
rect 172768 208928 172796 208968
rect 174590 208956 174596 208968
rect 174648 208956 174654 209008
rect 172164 208900 172796 208928
rect 172164 208888 172170 208900
rect 62626 208344 62632 208396
rect 62684 208384 62690 208396
rect 66398 208384 66404 208396
rect 62684 208356 66404 208384
rect 62684 208344 62690 208356
rect 66398 208344 66404 208356
rect 66456 208344 66462 208396
rect 135398 207800 135404 207852
rect 135456 207840 135462 207852
rect 136870 207840 136876 207852
rect 135456 207812 136876 207840
rect 135456 207800 135462 207812
rect 136870 207800 136876 207812
rect 136928 207800 136934 207852
rect 63730 207460 63736 207512
rect 63788 207500 63794 207512
rect 65294 207500 65300 207512
rect 63788 207472 65300 207500
rect 63788 207460 63794 207472
rect 65294 207460 65300 207472
rect 65352 207460 65358 207512
rect 171646 206780 171652 206832
rect 171704 206820 171710 206832
rect 174130 206820 174136 206832
rect 171704 206792 174136 206820
rect 171704 206780 171710 206792
rect 174130 206780 174136 206792
rect 174188 206780 174194 206832
rect 62534 206712 62540 206764
rect 62592 206752 62598 206764
rect 65662 206752 65668 206764
rect 62592 206724 65668 206752
rect 62592 206712 62598 206724
rect 65662 206712 65668 206724
rect 65720 206712 65726 206764
rect 135398 206304 135404 206356
rect 135456 206344 135462 206356
rect 136870 206344 136876 206356
rect 135456 206316 136876 206344
rect 135456 206304 135462 206316
rect 136870 206304 136876 206316
rect 136928 206304 136934 206356
rect 62626 206168 62632 206220
rect 62684 206208 62690 206220
rect 64926 206208 64932 206220
rect 62684 206180 64932 206208
rect 62684 206168 62690 206180
rect 64926 206168 64932 206180
rect 64984 206168 64990 206220
rect 171830 205964 171836 206016
rect 171888 206004 171894 206016
rect 174038 206004 174044 206016
rect 171888 205976 174044 206004
rect 171888 205964 171894 205976
rect 174038 205964 174044 205976
rect 174096 205964 174102 206016
rect 62626 205420 62632 205472
rect 62684 205460 62690 205472
rect 66398 205460 66404 205472
rect 62684 205432 66404 205460
rect 62684 205420 62690 205432
rect 66398 205420 66404 205432
rect 66456 205420 66462 205472
rect 62626 204332 62632 204384
rect 62684 204372 62690 204384
rect 65662 204372 65668 204384
rect 62684 204344 65668 204372
rect 62684 204332 62690 204344
rect 65662 204332 65668 204344
rect 65720 204332 65726 204384
rect 62534 204196 62540 204248
rect 62592 204236 62598 204248
rect 65478 204236 65484 204248
rect 62592 204208 65484 204236
rect 62592 204196 62598 204208
rect 65478 204196 65484 204208
rect 65536 204196 65542 204248
rect 100898 200660 100904 200712
rect 100956 200700 100962 200712
rect 102370 200700 102376 200712
rect 100956 200672 102376 200700
rect 100956 200660 100962 200672
rect 102370 200660 102376 200672
rect 102428 200660 102434 200712
rect 135398 200456 135404 200508
rect 135456 200496 135462 200508
rect 136778 200496 136784 200508
rect 135456 200468 136784 200496
rect 135456 200456 135462 200468
rect 136778 200456 136784 200468
rect 136836 200456 136842 200508
rect 172198 199368 172204 199420
rect 172256 199408 172262 199420
rect 175234 199408 175240 199420
rect 172256 199380 175240 199408
rect 172256 199368 172262 199380
rect 175234 199368 175240 199380
rect 175292 199368 175298 199420
rect 100898 199300 100904 199352
rect 100956 199340 100962 199352
rect 102370 199340 102376 199352
rect 100956 199312 102376 199340
rect 100956 199300 100962 199312
rect 102370 199300 102376 199312
rect 102428 199300 102434 199352
rect 62350 199096 62356 199148
rect 62408 199136 62414 199148
rect 65018 199136 65024 199148
rect 62408 199108 65024 199136
rect 62408 199096 62414 199108
rect 65018 199096 65024 199108
rect 65076 199096 65082 199148
rect 134754 199096 134760 199148
rect 134812 199136 134818 199148
rect 136778 199136 136784 199148
rect 134812 199108 136784 199136
rect 134812 199096 134818 199108
rect 136778 199096 136784 199108
rect 136836 199096 136842 199148
rect 172198 198008 172204 198060
rect 172256 198048 172262 198060
rect 174222 198048 174228 198060
rect 172256 198020 174228 198048
rect 172256 198008 172262 198020
rect 174222 198008 174228 198020
rect 174280 198008 174286 198060
rect 100898 197872 100904 197924
rect 100956 197912 100962 197924
rect 102370 197912 102376 197924
rect 100956 197884 102376 197912
rect 100956 197872 100962 197884
rect 102370 197872 102376 197884
rect 102428 197872 102434 197924
rect 62626 197736 62632 197788
rect 62684 197776 62690 197788
rect 65018 197776 65024 197788
rect 62684 197748 65024 197776
rect 62684 197736 62690 197748
rect 65018 197736 65024 197748
rect 65076 197736 65082 197788
rect 135398 197736 135404 197788
rect 135456 197776 135462 197788
rect 136778 197776 136784 197788
rect 135456 197748 136784 197776
rect 135456 197736 135462 197748
rect 136778 197736 136784 197748
rect 136836 197736 136842 197788
rect 172658 196784 172664 196836
rect 172716 196824 172722 196836
rect 174130 196824 174136 196836
rect 172716 196796 174136 196824
rect 172716 196784 172722 196796
rect 174130 196784 174136 196796
rect 174188 196784 174194 196836
rect 100898 196648 100904 196700
rect 100956 196688 100962 196700
rect 102370 196688 102376 196700
rect 100956 196660 102376 196688
rect 100956 196648 100962 196660
rect 102370 196648 102376 196660
rect 102428 196648 102434 196700
rect 172198 196648 172204 196700
rect 172256 196688 172262 196700
rect 174222 196688 174228 196700
rect 172256 196660 174228 196688
rect 172256 196648 172262 196660
rect 174222 196648 174228 196660
rect 174280 196648 174286 196700
rect 63730 196512 63736 196564
rect 63788 196552 63794 196564
rect 66398 196552 66404 196564
rect 63788 196524 66404 196552
rect 63788 196512 63794 196524
rect 66398 196512 66404 196524
rect 66456 196512 66462 196564
rect 100898 196512 100904 196564
rect 100956 196552 100962 196564
rect 102462 196552 102468 196564
rect 100956 196524 102468 196552
rect 100956 196512 100962 196524
rect 102462 196512 102468 196524
rect 102520 196512 102526 196564
rect 62626 196444 62632 196496
rect 62684 196484 62690 196496
rect 65018 196484 65024 196496
rect 62684 196456 65024 196484
rect 62684 196444 62690 196456
rect 65018 196444 65024 196456
rect 65076 196444 65082 196496
rect 135398 196376 135404 196428
rect 135456 196416 135462 196428
rect 136778 196416 136784 196428
rect 135456 196388 136784 196416
rect 135456 196376 135462 196388
rect 136778 196376 136784 196388
rect 136836 196376 136842 196428
rect 134294 196036 134300 196088
rect 134352 196076 134358 196088
rect 136686 196076 136692 196088
rect 134352 196048 136692 196076
rect 134352 196036 134358 196048
rect 136686 196036 136692 196048
rect 136744 196036 136750 196088
rect 171462 195560 171468 195612
rect 171520 195600 171526 195612
rect 174130 195600 174136 195612
rect 171520 195572 174136 195600
rect 171520 195560 171526 195572
rect 174130 195560 174136 195572
rect 174188 195560 174194 195612
rect 100714 195288 100720 195340
rect 100772 195328 100778 195340
rect 102462 195328 102468 195340
rect 100772 195300 102468 195328
rect 100772 195288 100778 195300
rect 102462 195288 102468 195300
rect 102520 195288 102526 195340
rect 66398 195192 66404 195204
rect 63748 195164 66404 195192
rect 62534 195084 62540 195136
rect 62592 195124 62598 195136
rect 63748 195124 63776 195164
rect 66398 195152 66404 195164
rect 66456 195152 66462 195204
rect 100898 195152 100904 195204
rect 100956 195192 100962 195204
rect 102370 195192 102376 195204
rect 100956 195164 102376 195192
rect 100956 195152 100962 195164
rect 102370 195152 102376 195164
rect 102428 195152 102434 195204
rect 136870 195192 136876 195204
rect 136428 195164 136876 195192
rect 62592 195096 63776 195124
rect 62592 195084 62598 195096
rect 135398 195084 135404 195136
rect 135456 195124 135462 195136
rect 136428 195124 136456 195164
rect 136870 195152 136876 195164
rect 136928 195152 136934 195204
rect 172658 195152 172664 195204
rect 172716 195192 172722 195204
rect 174222 195192 174228 195204
rect 172716 195164 174228 195192
rect 172716 195152 172722 195164
rect 174222 195152 174228 195164
rect 174280 195152 174286 195204
rect 135456 195096 136456 195124
rect 135456 195084 135462 195096
rect 62626 194948 62632 195000
rect 62684 194988 62690 195000
rect 65018 194988 65024 195000
rect 62684 194960 65024 194988
rect 62684 194948 62690 194960
rect 65018 194948 65024 194960
rect 65076 194948 65082 195000
rect 135398 194812 135404 194864
rect 135456 194852 135462 194864
rect 136778 194852 136784 194864
rect 135456 194824 136784 194852
rect 135456 194812 135462 194824
rect 136778 194812 136784 194824
rect 136836 194812 136842 194864
rect 100622 194200 100628 194252
rect 100680 194240 100686 194252
rect 102462 194240 102468 194252
rect 100680 194212 102468 194240
rect 100680 194200 100686 194212
rect 102462 194200 102468 194212
rect 102520 194200 102526 194252
rect 171554 194200 171560 194252
rect 171612 194240 171618 194252
rect 174130 194240 174136 194252
rect 171612 194212 174136 194240
rect 171612 194200 171618 194212
rect 174130 194200 174136 194212
rect 174188 194200 174194 194252
rect 100622 193792 100628 193844
rect 100680 193832 100686 193844
rect 102370 193832 102376 193844
rect 100680 193804 102376 193832
rect 100680 193792 100686 193804
rect 102370 193792 102376 193804
rect 102428 193792 102434 193844
rect 172658 193792 172664 193844
rect 172716 193832 172722 193844
rect 174222 193832 174228 193844
rect 172716 193804 174228 193832
rect 172716 193792 172722 193804
rect 174222 193792 174228 193804
rect 174280 193792 174286 193844
rect 135398 193656 135404 193708
rect 135456 193696 135462 193708
rect 136778 193696 136784 193708
rect 135456 193668 136784 193696
rect 135456 193656 135462 193668
rect 136778 193656 136784 193668
rect 136836 193656 136842 193708
rect 135398 193452 135404 193504
rect 135456 193492 135462 193504
rect 136686 193492 136692 193504
rect 135456 193464 136692 193492
rect 135456 193452 135462 193464
rect 136686 193452 136692 193464
rect 136744 193452 136750 193504
rect 62350 193248 62356 193300
rect 62408 193288 62414 193300
rect 65018 193288 65024 193300
rect 62408 193260 65024 193288
rect 62408 193248 62414 193260
rect 65018 193248 65024 193260
rect 65076 193248 65082 193300
rect 171646 192976 171652 193028
rect 171704 193016 171710 193028
rect 174222 193016 174228 193028
rect 171704 192988 174228 193016
rect 171704 192976 171710 192988
rect 174222 192976 174228 192988
rect 174280 192976 174286 193028
rect 99702 192840 99708 192892
rect 99760 192880 99766 192892
rect 102462 192880 102468 192892
rect 99760 192852 102468 192880
rect 99760 192840 99766 192852
rect 102462 192840 102468 192852
rect 102520 192840 102526 192892
rect 172198 192568 172204 192620
rect 172256 192608 172262 192620
rect 174130 192608 174136 192620
rect 172256 192580 174136 192608
rect 172256 192568 172262 192580
rect 174130 192568 174136 192580
rect 174188 192568 174194 192620
rect 100622 192432 100628 192484
rect 100680 192472 100686 192484
rect 102370 192472 102376 192484
rect 100680 192444 102376 192472
rect 100680 192432 100686 192444
rect 102370 192432 102376 192444
rect 102428 192432 102434 192484
rect 135398 192296 135404 192348
rect 135456 192336 135462 192348
rect 136778 192336 136784 192348
rect 135456 192308 136784 192336
rect 135456 192296 135462 192308
rect 136778 192296 136784 192308
rect 136836 192296 136842 192348
rect 62534 192228 62540 192280
rect 62592 192268 62598 192280
rect 64926 192268 64932 192280
rect 62592 192240 64932 192268
rect 62592 192228 62598 192240
rect 64926 192228 64932 192240
rect 64984 192228 64990 192280
rect 134294 192228 134300 192280
rect 134352 192268 134358 192280
rect 136686 192268 136692 192280
rect 134352 192240 136692 192268
rect 134352 192228 134358 192240
rect 136686 192228 136692 192240
rect 136744 192228 136750 192280
rect 99886 191888 99892 191940
rect 99944 191928 99950 191940
rect 102278 191928 102284 191940
rect 99944 191900 102284 191928
rect 99944 191888 99950 191900
rect 102278 191888 102284 191900
rect 102336 191888 102342 191940
rect 62350 191548 62356 191600
rect 62408 191588 62414 191600
rect 65018 191588 65024 191600
rect 62408 191560 65024 191588
rect 62408 191548 62414 191560
rect 65018 191548 65024 191560
rect 65076 191548 65082 191600
rect 172198 191344 172204 191396
rect 172256 191384 172262 191396
rect 174038 191384 174044 191396
rect 172256 191356 174044 191384
rect 172256 191344 172262 191356
rect 174038 191344 174044 191356
rect 174096 191344 174102 191396
rect 172658 191276 172664 191328
rect 172716 191316 172722 191328
rect 173946 191316 173952 191328
rect 172716 191288 173952 191316
rect 172716 191276 172722 191288
rect 173946 191276 173952 191288
rect 174004 191276 174010 191328
rect 100622 191208 100628 191260
rect 100680 191248 100686 191260
rect 102186 191248 102192 191260
rect 100680 191220 102192 191248
rect 100680 191208 100686 191220
rect 102186 191208 102192 191220
rect 102244 191208 102250 191260
rect 66306 191044 66312 191056
rect 63748 191016 66312 191044
rect 62442 190936 62448 190988
rect 62500 190976 62506 190988
rect 63748 190976 63776 191016
rect 66306 191004 66312 191016
rect 66364 191004 66370 191056
rect 100898 191004 100904 191056
rect 100956 191044 100962 191056
rect 102554 191044 102560 191056
rect 100956 191016 102560 191044
rect 100956 191004 100962 191016
rect 102554 191004 102560 191016
rect 102612 191004 102618 191056
rect 134294 191004 134300 191056
rect 134352 191044 134358 191056
rect 136962 191044 136968 191056
rect 134352 191016 136968 191044
rect 134352 191004 134358 191016
rect 136962 191004 136968 191016
rect 137020 191004 137026 191056
rect 172658 191004 172664 191056
rect 172716 191044 172722 191056
rect 174958 191044 174964 191056
rect 172716 191016 174964 191044
rect 172716 191004 172722 191016
rect 174958 191004 174964 191016
rect 175016 191004 175022 191056
rect 62500 190948 63776 190976
rect 62500 190936 62506 190948
rect 135398 190936 135404 190988
rect 135456 190976 135462 190988
rect 136778 190976 136784 190988
rect 135456 190948 136784 190976
rect 135456 190936 135462 190948
rect 136778 190936 136784 190948
rect 136836 190936 136842 190988
rect 62626 190868 62632 190920
rect 62684 190908 62690 190920
rect 65018 190908 65024 190920
rect 62684 190880 65024 190908
rect 62684 190868 62690 190880
rect 65018 190868 65024 190880
rect 65076 190868 65082 190920
rect 134754 190868 134760 190920
rect 134812 190908 134818 190920
rect 136686 190908 136692 190920
rect 134812 190880 136692 190908
rect 134812 190868 134818 190880
rect 136686 190868 136692 190880
rect 136744 190868 136750 190920
rect 172382 190120 172388 190172
rect 172440 190160 172446 190172
rect 174406 190160 174412 190172
rect 172440 190132 174412 190160
rect 172440 190120 172446 190132
rect 174406 190120 174412 190132
rect 174464 190120 174470 190172
rect 100530 190052 100536 190104
rect 100588 190092 100594 190104
rect 102462 190092 102468 190104
rect 100588 190064 102468 190092
rect 100588 190052 100594 190064
rect 102462 190052 102468 190064
rect 102520 190052 102526 190104
rect 99886 189780 99892 189832
rect 99944 189820 99950 189832
rect 102370 189820 102376 189832
rect 99944 189792 102376 189820
rect 99944 189780 99950 189792
rect 102370 189780 102376 189792
rect 102428 189780 102434 189832
rect 172014 189712 172020 189764
rect 172072 189752 172078 189764
rect 175418 189752 175424 189764
rect 172072 189724 175424 189752
rect 172072 189712 172078 189724
rect 175418 189712 175424 189724
rect 175476 189712 175482 189764
rect 63638 189644 63644 189696
rect 63696 189684 63702 189696
rect 66398 189684 66404 189696
rect 63696 189656 66404 189684
rect 63696 189644 63702 189656
rect 66398 189644 66404 189656
rect 66456 189644 66462 189696
rect 62626 189508 62632 189560
rect 62684 189548 62690 189560
rect 65202 189548 65208 189560
rect 62684 189520 65208 189548
rect 62684 189508 62690 189520
rect 65202 189508 65208 189520
rect 65260 189508 65266 189560
rect 134754 189236 134760 189288
rect 134812 189276 134818 189288
rect 136778 189276 136784 189288
rect 134812 189248 136784 189276
rect 134812 189236 134818 189248
rect 136778 189236 136784 189248
rect 136836 189236 136842 189288
rect 62626 189032 62632 189084
rect 62684 189072 62690 189084
rect 65018 189072 65024 189084
rect 62684 189044 65024 189072
rect 62684 189032 62690 189044
rect 65018 189032 65024 189044
rect 65076 189032 65082 189084
rect 135030 188148 135036 188200
rect 135088 188188 135094 188200
rect 137422 188188 137428 188200
rect 135088 188160 137428 188188
rect 135088 188148 135094 188160
rect 137422 188148 137428 188160
rect 137480 188148 137486 188200
rect 116446 187604 116452 187656
rect 116504 187644 116510 187656
rect 117412 187644 117418 187656
rect 116504 187616 117418 187644
rect 116504 187604 116510 187616
rect 117412 187604 117418 187616
rect 117470 187604 117476 187656
rect 132638 186924 132644 186976
rect 132696 186964 132702 186976
rect 144874 186964 144880 186976
rect 132696 186936 144880 186964
rect 132696 186924 132702 186936
rect 144874 186924 144880 186936
rect 144932 186924 144938 186976
rect 121874 186856 121880 186908
rect 121932 186896 121938 186908
rect 125186 186896 125192 186908
rect 121932 186868 125192 186896
rect 121932 186856 121938 186868
rect 125186 186856 125192 186868
rect 125244 186856 125250 186908
rect 132086 186856 132092 186908
rect 132144 186896 132150 186908
rect 164838 186896 164844 186908
rect 132144 186868 164844 186896
rect 132144 186856 132150 186868
rect 164838 186856 164844 186868
rect 164896 186856 164902 186908
rect 35578 185428 35584 185480
rect 35636 185468 35642 185480
rect 37878 185468 37884 185480
rect 35636 185440 37884 185468
rect 35636 185428 35642 185440
rect 37878 185428 37884 185440
rect 37936 185428 37942 185480
rect 41006 185428 41012 185480
rect 41064 185468 41070 185480
rect 43398 185468 43404 185480
rect 41064 185440 43404 185468
rect 41064 185428 41070 185440
rect 43398 185428 43404 185440
rect 43456 185428 43462 185480
rect 43766 185428 43772 185480
rect 43824 185468 43830 185480
rect 44686 185468 44692 185480
rect 43824 185440 44692 185468
rect 43824 185428 43830 185440
rect 44686 185428 44692 185440
rect 44744 185428 44750 185480
rect 49010 185428 49016 185480
rect 49068 185468 49074 185480
rect 50574 185468 50580 185480
rect 49068 185440 50580 185468
rect 49068 185428 49074 185440
rect 50574 185428 50580 185440
rect 50632 185428 50638 185480
rect 50666 185428 50672 185480
rect 50724 185468 50730 185480
rect 53334 185468 53340 185480
rect 50724 185440 53340 185468
rect 50724 185428 50730 185440
rect 53334 185428 53340 185440
rect 53392 185428 53398 185480
rect 53426 185428 53432 185480
rect 53484 185468 53490 185480
rect 58118 185468 58124 185480
rect 53484 185440 58124 185468
rect 53484 185428 53490 185440
rect 58118 185428 58124 185440
rect 58176 185428 58182 185480
rect 110098 185428 110104 185480
rect 110156 185468 110162 185480
rect 111110 185468 111116 185480
rect 110156 185440 111116 185468
rect 110156 185428 110162 185440
rect 111110 185428 111116 185440
rect 111168 185428 111174 185480
rect 125922 185428 125928 185480
rect 125980 185468 125986 185480
rect 128130 185468 128136 185480
rect 125980 185440 128136 185468
rect 125980 185428 125986 185440
rect 128130 185428 128136 185440
rect 128188 185428 128194 185480
rect 182870 185428 182876 185480
rect 182928 185468 182934 185480
rect 183606 185468 183612 185480
rect 182928 185440 183612 185468
rect 182928 185428 182934 185440
rect 183606 185428 183612 185440
rect 183664 185428 183670 185480
rect 190138 185428 190144 185480
rect 190196 185468 190202 185480
rect 191426 185468 191432 185480
rect 190196 185440 191432 185468
rect 190196 185428 190202 185440
rect 191426 185428 191432 185440
rect 191484 185428 191490 185480
rect 197314 185428 197320 185480
rect 197372 185468 197378 185480
rect 201638 185468 201644 185480
rect 197372 185440 201644 185468
rect 197372 185428 197378 185440
rect 201638 185428 201644 185440
rect 201696 185428 201702 185480
rect 40362 185360 40368 185412
rect 40420 185400 40426 185412
rect 43030 185400 43036 185412
rect 40420 185372 43036 185400
rect 40420 185360 40426 185372
rect 43030 185360 43036 185372
rect 43088 185360 43094 185412
rect 43122 185360 43128 185412
rect 43180 185400 43186 185412
rect 44594 185400 44600 185412
rect 43180 185372 44600 185400
rect 43180 185360 43186 185372
rect 44594 185360 44600 185372
rect 44652 185360 44658 185412
rect 50206 185360 50212 185412
rect 50264 185400 50270 185412
rect 52690 185400 52696 185412
rect 50264 185372 52696 185400
rect 50264 185360 50270 185372
rect 52690 185360 52696 185372
rect 52748 185360 52754 185412
rect 110742 185360 110748 185412
rect 110800 185400 110806 185412
rect 111478 185400 111484 185412
rect 110800 185372 111484 185400
rect 110800 185360 110806 185372
rect 111478 185360 111484 185372
rect 111536 185360 111542 185412
rect 127210 185360 127216 185412
rect 127268 185400 127274 185412
rect 129970 185400 129976 185412
rect 127268 185372 129976 185400
rect 127268 185360 127274 185372
rect 129970 185360 129976 185372
rect 130028 185360 130034 185412
rect 190598 185360 190604 185412
rect 190656 185400 190662 185412
rect 192530 185400 192536 185412
rect 190656 185372 192536 185400
rect 190656 185360 190662 185372
rect 192530 185360 192536 185372
rect 192588 185360 192594 185412
rect 192898 185360 192904 185412
rect 192956 185400 192962 185412
rect 195382 185400 195388 185412
rect 192956 185372 195388 185400
rect 192956 185360 192962 185372
rect 195382 185360 195388 185372
rect 195440 185360 195446 185412
rect 195750 185360 195756 185412
rect 195808 185400 195814 185412
rect 199338 185400 199344 185412
rect 195808 185372 199344 185400
rect 195808 185360 195814 185372
rect 199338 185360 199344 185372
rect 199396 185360 199402 185412
rect 36314 185292 36320 185344
rect 36372 185332 36378 185344
rect 40638 185332 40644 185344
rect 36372 185304 40644 185332
rect 36372 185292 36378 185304
rect 40638 185292 40644 185304
rect 40696 185292 40702 185344
rect 41742 185292 41748 185344
rect 41800 185332 41806 185344
rect 43858 185332 43864 185344
rect 41800 185304 43864 185332
rect 41800 185292 41806 185304
rect 43858 185292 43864 185304
rect 43916 185292 43922 185344
rect 52230 185292 52236 185344
rect 52288 185332 52294 185344
rect 56094 185332 56100 185344
rect 52288 185304 56100 185332
rect 52288 185292 52294 185304
rect 56094 185292 56100 185304
rect 56152 185292 56158 185344
rect 125922 185292 125928 185344
rect 125980 185332 125986 185344
rect 127302 185332 127308 185344
rect 125980 185304 127308 185332
rect 125980 185292 125986 185304
rect 127302 185292 127308 185304
rect 127360 185292 127366 185344
rect 193358 185292 193364 185344
rect 193416 185332 193422 185344
rect 195934 185332 195940 185344
rect 193416 185304 195940 185332
rect 193416 185292 193422 185304
rect 195934 185292 195940 185304
rect 195992 185292 195998 185344
rect 196118 185292 196124 185344
rect 196176 185332 196182 185344
rect 199982 185332 199988 185344
rect 196176 185304 199988 185332
rect 196176 185292 196182 185304
rect 199982 185292 199988 185304
rect 200040 185292 200046 185344
rect 39718 185224 39724 185276
rect 39776 185264 39782 185276
rect 42662 185264 42668 185276
rect 39776 185236 42668 185264
rect 39776 185224 39782 185236
rect 42662 185224 42668 185236
rect 42720 185224 42726 185276
rect 49470 185224 49476 185276
rect 49528 185264 49534 185276
rect 51310 185264 51316 185276
rect 49528 185236 51316 185264
rect 49528 185224 49534 185236
rect 51310 185224 51316 185236
rect 51368 185224 51374 185276
rect 53058 185224 53064 185276
rect 53116 185264 53122 185276
rect 57382 185264 57388 185276
rect 53116 185236 57388 185264
rect 53116 185224 53122 185236
rect 57382 185224 57388 185236
rect 57440 185224 57446 185276
rect 105590 185224 105596 185276
rect 105648 185264 105654 185276
rect 109270 185264 109276 185276
rect 105648 185236 109276 185264
rect 105648 185224 105654 185236
rect 109270 185224 109276 185236
rect 109328 185224 109334 185276
rect 124818 185224 124824 185276
rect 124876 185264 124882 185276
rect 126382 185264 126388 185276
rect 124876 185236 126388 185264
rect 124876 185224 124882 185236
rect 126382 185224 126388 185236
rect 126440 185224 126446 185276
rect 192530 185224 192536 185276
rect 192588 185264 192594 185276
rect 194830 185264 194836 185276
rect 192588 185236 194836 185264
rect 192588 185224 192594 185236
rect 194830 185224 194836 185236
rect 194888 185224 194894 185276
rect 195290 185224 195296 185276
rect 195348 185264 195354 185276
rect 198786 185264 198792 185276
rect 195348 185236 198792 185264
rect 195348 185224 195354 185236
rect 198786 185224 198792 185236
rect 198844 185224 198850 185276
rect 37602 185156 37608 185208
rect 37660 185196 37666 185208
rect 41466 185196 41472 185208
rect 37660 185168 41472 185196
rect 37660 185156 37666 185168
rect 41466 185156 41472 185168
rect 41524 185156 41530 185208
rect 51034 185156 51040 185208
rect 51092 185196 51098 185208
rect 53978 185196 53984 185208
rect 51092 185168 53984 185196
rect 51092 185156 51098 185168
rect 53978 185156 53984 185168
rect 54036 185156 54042 185208
rect 194094 185156 194100 185208
rect 194152 185196 194158 185208
rect 197130 185196 197136 185208
rect 194152 185168 197136 185196
rect 194152 185156 194158 185168
rect 197130 185156 197136 185168
rect 197188 185156 197194 185208
rect 38982 185088 38988 185140
rect 39040 185128 39046 185140
rect 42202 185128 42208 185140
rect 39040 185100 42208 185128
rect 39040 185088 39046 185100
rect 42202 185088 42208 185100
rect 42260 185088 42266 185140
rect 42386 185088 42392 185140
rect 42444 185128 42450 185140
rect 44226 185128 44232 185140
rect 42444 185100 44232 185128
rect 42444 185088 42450 185100
rect 44226 185088 44232 185100
rect 44284 185088 44290 185140
rect 49838 185088 49844 185140
rect 49896 185128 49902 185140
rect 51954 185128 51960 185140
rect 49896 185100 51960 185128
rect 49896 185088 49902 185100
rect 51954 185088 51960 185100
rect 52012 185088 52018 185140
rect 52598 185088 52604 185140
rect 52656 185128 52662 185140
rect 56738 185128 56744 185140
rect 52656 185100 56744 185128
rect 52656 185088 52662 185100
rect 56738 185088 56744 185100
rect 56796 185088 56802 185140
rect 190414 185088 190420 185140
rect 190472 185128 190478 185140
rect 191978 185128 191984 185140
rect 190472 185100 191984 185128
rect 190472 185088 190478 185100
rect 191978 185088 191984 185100
rect 192036 185088 192042 185140
rect 194554 185088 194560 185140
rect 194612 185128 194618 185140
rect 197682 185128 197688 185140
rect 194612 185100 197688 185128
rect 194612 185088 194618 185100
rect 197682 185088 197688 185100
rect 197740 185088 197746 185140
rect 38338 185020 38344 185072
rect 38396 185060 38402 185072
rect 41834 185060 41840 185072
rect 38396 185032 41840 185060
rect 38396 185020 38402 185032
rect 41834 185020 41840 185032
rect 41892 185020 41898 185072
rect 48642 185020 48648 185072
rect 48700 185060 48706 185072
rect 49930 185060 49936 185072
rect 48700 185032 49936 185060
rect 48700 185020 48706 185032
rect 49930 185020 49936 185032
rect 49988 185020 49994 185072
rect 51402 185020 51408 185072
rect 51460 185060 51466 185072
rect 54714 185060 54720 185072
rect 51460 185032 54720 185060
rect 51460 185020 51466 185032
rect 54714 185020 54720 185032
rect 54772 185020 54778 185072
rect 127210 185020 127216 185072
rect 127268 185060 127274 185072
rect 130430 185060 130436 185072
rect 127268 185032 130436 185060
rect 127268 185020 127274 185032
rect 130430 185020 130436 185032
rect 130488 185020 130494 185072
rect 194646 185020 194652 185072
rect 194704 185060 194710 185072
rect 198234 185060 198240 185072
rect 194704 185032 198240 185060
rect 194704 185020 194710 185032
rect 198234 185020 198240 185032
rect 198292 185020 198298 185072
rect 51862 184952 51868 185004
rect 51920 184992 51926 185004
rect 55358 184992 55364 185004
rect 51920 184964 55364 184992
rect 51920 184952 51926 184964
rect 55358 184952 55364 184964
rect 55416 184952 55422 185004
rect 177718 184952 177724 185004
rect 177776 184992 177782 185004
rect 181122 184992 181128 185004
rect 177776 184964 181128 184992
rect 177776 184952 177782 184964
rect 181122 184952 181128 184964
rect 181180 184952 181186 185004
rect 181674 184952 181680 185004
rect 181732 184992 181738 185004
rect 183100 184992 183106 185004
rect 181732 184964 183106 184992
rect 181732 184952 181738 184964
rect 183100 184952 183106 184964
rect 183158 184952 183164 185004
rect 189080 184952 189086 185004
rect 189138 184992 189144 185004
rect 190230 184992 190236 185004
rect 189138 184964 190236 184992
rect 189138 184952 189144 184964
rect 190230 184952 190236 184964
rect 190288 184952 190294 185004
rect 191104 184952 191110 185004
rect 191162 184992 191168 185004
rect 193082 184992 193088 185004
rect 191162 184964 193088 184992
rect 191162 184952 191168 184964
rect 193082 184952 193088 184964
rect 193140 184952 193146 185004
rect 193496 184952 193502 185004
rect 193554 184992 193560 185004
rect 196486 184992 196492 185004
rect 193554 184964 196492 184992
rect 193554 184952 193560 184964
rect 196486 184952 196492 184964
rect 196544 184952 196550 185004
rect 197820 184952 197826 185004
rect 197878 184992 197884 185004
rect 202834 184992 202840 185004
rect 197878 184964 202840 184992
rect 197878 184952 197884 184964
rect 202834 184952 202840 184964
rect 202892 184952 202898 185004
rect 36958 184884 36964 184936
rect 37016 184924 37022 184936
rect 41006 184924 41012 184936
rect 37016 184896 41012 184924
rect 37016 184884 37022 184896
rect 41006 184884 41012 184896
rect 41064 184884 41070 184936
rect 127210 184884 127216 184936
rect 127268 184924 127274 184936
rect 129326 184924 129332 184936
rect 127268 184896 129332 184924
rect 127268 184884 127274 184896
rect 129326 184884 129332 184896
rect 129384 184884 129390 184936
rect 182226 184884 182232 184936
rect 182284 184924 182290 184936
rect 183468 184924 183474 184936
rect 182284 184896 183474 184924
rect 182284 184884 182290 184896
rect 183468 184884 183474 184896
rect 183526 184884 183532 184936
rect 189448 184884 189454 184936
rect 189506 184924 189512 184936
rect 190782 184924 190788 184936
rect 189506 184896 190788 184924
rect 189506 184884 189512 184896
rect 190782 184884 190788 184896
rect 190840 184884 190846 184936
rect 191472 184884 191478 184936
rect 191530 184924 191536 184936
rect 193634 184924 193640 184936
rect 191530 184896 193640 184924
rect 191530 184884 191536 184896
rect 193634 184884 193640 184896
rect 193692 184884 193698 184936
rect 196624 184884 196630 184936
rect 196682 184924 196688 184936
rect 201086 184924 201092 184936
rect 196682 184896 201092 184924
rect 196682 184884 196688 184896
rect 201086 184884 201092 184896
rect 201144 184884 201150 184936
rect 191978 184816 191984 184868
rect 192036 184856 192042 184868
rect 194002 184856 194008 184868
rect 192036 184828 194008 184856
rect 192036 184816 192042 184828
rect 194002 184816 194008 184828
rect 194060 184816 194066 184868
rect 196486 184816 196492 184868
rect 196544 184856 196550 184868
rect 200534 184856 200540 184868
rect 196544 184828 200540 184856
rect 196544 184816 196550 184828
rect 200534 184816 200540 184828
rect 200592 184816 200598 184868
rect 127026 184680 127032 184732
rect 127084 184720 127090 184732
rect 128682 184720 128688 184732
rect 127084 184692 128688 184720
rect 127084 184680 127090 184692
rect 128682 184680 128688 184692
rect 128740 184680 128746 184732
rect 53978 184544 53984 184596
rect 54036 184584 54042 184596
rect 58762 184584 58768 184596
rect 54036 184556 58768 184584
rect 54036 184544 54042 184556
rect 58762 184544 58768 184556
rect 58820 184544 58826 184596
rect 127026 184476 127032 184528
rect 127084 184516 127090 184528
rect 127578 184516 127584 184528
rect 127084 184488 127584 184516
rect 127084 184476 127090 184488
rect 127578 184476 127584 184488
rect 127636 184476 127642 184528
rect 39258 184408 39264 184460
rect 39316 184408 39322 184460
rect 54530 184408 54536 184460
rect 54588 184408 54594 184460
rect 34934 184272 34940 184324
rect 34992 184312 34998 184324
rect 37970 184312 37976 184324
rect 34992 184284 37976 184312
rect 34992 184272 34998 184284
rect 37970 184272 37976 184284
rect 38028 184272 38034 184324
rect 34198 184204 34204 184256
rect 34256 184244 34262 184256
rect 39276 184244 39304 184408
rect 34256 184216 39304 184244
rect 54548 184244 54576 184408
rect 59498 184244 59504 184256
rect 54548 184216 59504 184244
rect 34256 184204 34262 184216
rect 59498 184204 59504 184216
rect 59556 184204 59562 184256
rect 106050 184204 106056 184256
rect 106108 184244 106114 184256
rect 107154 184244 107160 184256
rect 106108 184216 107160 184244
rect 106108 184204 106114 184216
rect 107154 184204 107160 184216
rect 107212 184204 107218 184256
rect 177074 184204 177080 184256
rect 177132 184244 177138 184256
rect 179374 184244 179380 184256
rect 177132 184216 179380 184244
rect 177132 184204 177138 184216
rect 179374 184204 179380 184216
rect 179432 184204 179438 184256
rect 177626 184136 177632 184188
rect 177684 184176 177690 184188
rect 178822 184176 178828 184188
rect 177684 184148 178828 184176
rect 177684 184136 177690 184148
rect 178822 184136 178828 184148
rect 178880 184136 178886 184188
rect 33554 184068 33560 184120
rect 33612 184108 33618 184120
rect 38890 184108 38896 184120
rect 33612 184080 38896 184108
rect 33612 184068 33618 184080
rect 38890 184068 38896 184080
rect 38948 184068 38954 184120
rect 105958 184068 105964 184120
rect 106016 184108 106022 184120
rect 106602 184108 106608 184120
rect 106016 184080 106608 184108
rect 106016 184068 106022 184080
rect 106602 184068 106608 184080
rect 106660 184068 106666 184120
rect 108350 184108 108356 184120
rect 106712 184080 108356 184108
rect 106142 184000 106148 184052
rect 106200 184040 106206 184052
rect 106712 184040 106740 184080
rect 108350 184068 108356 184080
rect 108408 184068 108414 184120
rect 177534 184068 177540 184120
rect 177592 184108 177598 184120
rect 178270 184108 178276 184120
rect 177592 184080 178276 184108
rect 177592 184068 177598 184080
rect 178270 184068 178276 184080
rect 178328 184068 178334 184120
rect 180570 184108 180576 184120
rect 178380 184080 180576 184108
rect 106200 184012 106740 184040
rect 106200 184000 106206 184012
rect 177442 184000 177448 184052
rect 177500 184040 177506 184052
rect 178380 184040 178408 184080
rect 180570 184068 180576 184080
rect 180628 184068 180634 184120
rect 177500 184012 178408 184040
rect 177500 184000 177506 184012
rect 176982 182436 176988 182488
rect 177040 182476 177046 182488
rect 180018 182476 180024 182488
rect 177040 182448 180024 182476
rect 177040 182436 177046 182448
rect 180018 182436 180024 182448
rect 180076 182436 180082 182488
rect 105590 182368 105596 182420
rect 105648 182408 105654 182420
rect 107890 182408 107896 182420
rect 105648 182380 107896 182408
rect 105648 182368 105654 182380
rect 107890 182368 107896 182380
rect 107948 182368 107954 182420
rect 105406 180328 105412 180380
rect 105464 180368 105470 180380
rect 108074 180368 108080 180380
rect 105464 180340 108080 180368
rect 105464 180328 105470 180340
rect 108074 180328 108080 180340
rect 108132 180328 108138 180380
rect 106326 178560 106332 178612
rect 106384 178600 106390 178612
rect 107890 178600 107896 178612
rect 106384 178572 107896 178600
rect 106384 178560 106390 178572
rect 107890 178560 107896 178572
rect 107948 178560 107954 178612
rect 32634 177200 32640 177252
rect 32692 177240 32698 177252
rect 37418 177240 37424 177252
rect 32692 177212 37424 177240
rect 32692 177200 32698 177212
rect 37418 177200 37424 177212
rect 37476 177200 37482 177252
rect 57566 177200 57572 177252
rect 57624 177240 57630 177252
rect 59590 177240 59596 177252
rect 57624 177212 59596 177240
rect 57624 177200 57630 177212
rect 59590 177200 59596 177212
rect 59648 177200 59654 177252
rect 106418 175840 106424 175892
rect 106476 175880 106482 175892
rect 107890 175880 107896 175892
rect 106476 175852 107896 175880
rect 106476 175840 106482 175852
rect 107890 175840 107896 175852
rect 107948 175840 107954 175892
rect 177718 175840 177724 175892
rect 177776 175880 177782 175892
rect 179650 175880 179656 175892
rect 177776 175852 179656 175880
rect 177776 175840 177782 175852
rect 179650 175840 179656 175852
rect 179708 175840 179714 175892
rect 106142 174344 106148 174396
rect 106200 174384 106206 174396
rect 108534 174384 108540 174396
rect 106200 174356 108540 174384
rect 106200 174344 106206 174356
rect 108534 174344 108540 174356
rect 108592 174344 108598 174396
rect 177350 174344 177356 174396
rect 177408 174384 177414 174396
rect 180294 174384 180300 174396
rect 177408 174356 180300 174384
rect 177408 174344 177414 174356
rect 180294 174344 180300 174356
rect 180352 174344 180358 174396
rect 176982 174276 176988 174328
rect 177040 174316 177046 174328
rect 179926 174316 179932 174328
rect 177040 174288 179932 174316
rect 177040 174276 177046 174288
rect 179926 174276 179932 174288
rect 179984 174276 179990 174328
rect 106050 173052 106056 173104
rect 106108 173092 106114 173104
rect 108166 173092 108172 173104
rect 106108 173064 108172 173092
rect 106108 173052 106114 173064
rect 108166 173052 108172 173064
rect 108224 173052 108230 173104
rect 177626 173052 177632 173104
rect 177684 173092 177690 173104
rect 179650 173092 179656 173104
rect 177684 173064 179656 173092
rect 177684 173052 177690 173064
rect 179650 173052 179656 173064
rect 179708 173052 179714 173104
rect 177534 172916 177540 172968
rect 177592 172956 177598 172968
rect 179742 172956 179748 172968
rect 177592 172928 179748 172956
rect 177592 172916 177598 172928
rect 179742 172916 179748 172928
rect 179800 172916 179806 172968
rect 105222 171692 105228 171744
rect 105280 171732 105286 171744
rect 107890 171732 107896 171744
rect 105280 171704 107896 171732
rect 105280 171692 105286 171704
rect 107890 171692 107896 171704
rect 107948 171692 107954 171744
rect 178086 171692 178092 171744
rect 178144 171732 178150 171744
rect 179650 171732 179656 171744
rect 178144 171704 179656 171732
rect 178144 171692 178150 171704
rect 179650 171692 179656 171704
rect 179708 171692 179714 171744
rect 222798 169108 222804 169160
rect 222856 169148 222862 169160
rect 223534 169148 223540 169160
rect 222856 169120 223540 169148
rect 222856 169108 222862 169120
rect 223534 169108 223540 169120
rect 223592 169108 223598 169160
rect 105958 168904 105964 168956
rect 106016 168944 106022 168956
rect 107890 168944 107896 168956
rect 106016 168916 107896 168944
rect 106016 168904 106022 168916
rect 107890 168904 107896 168916
rect 107948 168904 107954 168956
rect 177534 168904 177540 168956
rect 177592 168944 177598 168956
rect 179650 168944 179656 168956
rect 177592 168916 179656 168944
rect 177592 168904 177598 168916
rect 179650 168904 179656 168916
rect 179708 168904 179714 168956
rect 106418 166116 106424 166168
rect 106476 166156 106482 166168
rect 107798 166156 107804 166168
rect 106476 166128 107804 166156
rect 106476 166116 106482 166128
rect 107798 166116 107804 166128
rect 107856 166116 107862 166168
rect 177534 166116 177540 166168
rect 177592 166156 177598 166168
rect 179558 166156 179564 166168
rect 177592 166128 179564 166156
rect 177592 166116 177598 166128
rect 179558 166116 179564 166128
rect 179616 166116 179622 166168
rect 201086 166116 201092 166168
rect 201144 166156 201150 166168
rect 204490 166156 204496 166168
rect 201144 166128 204496 166156
rect 201144 166116 201150 166128
rect 204490 166116 204496 166128
rect 204548 166116 204554 166168
rect 28862 164756 28868 164808
rect 28920 164796 28926 164808
rect 37418 164796 37424 164808
rect 28920 164768 37424 164796
rect 28920 164756 28926 164768
rect 37418 164756 37424 164768
rect 37476 164756 37482 164808
rect 54898 164756 54904 164808
rect 54956 164796 54962 164808
rect 59590 164796 59596 164808
rect 54956 164768 59596 164796
rect 54956 164756 54962 164768
rect 59590 164756 59596 164768
rect 59648 164756 59654 164808
rect 106418 163464 106424 163516
rect 106476 163504 106482 163516
rect 107798 163504 107804 163516
rect 106476 163476 107804 163504
rect 106476 163464 106482 163476
rect 107798 163464 107804 163476
rect 107856 163464 107862 163516
rect 177718 163464 177724 163516
rect 177776 163504 177782 163516
rect 179558 163504 179564 163516
rect 177776 163476 179564 163504
rect 177776 163464 177782 163476
rect 179558 163464 179564 163476
rect 179616 163464 179622 163516
rect 106142 162104 106148 162156
rect 106200 162144 106206 162156
rect 108534 162144 108540 162156
rect 106200 162116 108540 162144
rect 106200 162104 106206 162116
rect 108534 162104 108540 162116
rect 108592 162104 108598 162156
rect 176982 162036 176988 162088
rect 177040 162076 177046 162088
rect 179650 162076 179656 162088
rect 177040 162048 179656 162076
rect 177040 162036 177046 162048
rect 179650 162036 179656 162048
rect 179708 162036 179714 162088
rect 176982 160812 176988 160864
rect 177040 160852 177046 160864
rect 179558 160852 179564 160864
rect 177040 160824 179564 160852
rect 177040 160812 177046 160824
rect 179558 160812 179564 160824
rect 179616 160812 179622 160864
rect 105774 160608 105780 160660
rect 105832 160648 105838 160660
rect 107798 160648 107804 160660
rect 105832 160620 107804 160648
rect 105832 160608 105838 160620
rect 107798 160608 107804 160620
rect 107856 160608 107862 160660
rect 106418 159248 106424 159300
rect 106476 159288 106482 159300
rect 107706 159288 107712 159300
rect 106476 159260 107712 159288
rect 106476 159248 106482 159260
rect 107706 159248 107712 159260
rect 107764 159248 107770 159300
rect 177534 159248 177540 159300
rect 177592 159288 177598 159300
rect 179466 159288 179472 159300
rect 177592 159260 179472 159288
rect 177592 159248 177598 159260
rect 179466 159248 179472 159260
rect 179524 159248 179530 159300
rect 105406 158160 105412 158212
rect 105464 158200 105470 158212
rect 107890 158200 107896 158212
rect 105464 158172 107896 158200
rect 105464 158160 105470 158172
rect 107890 158160 107896 158172
rect 107948 158160 107954 158212
rect 177350 157888 177356 157940
rect 177408 157928 177414 157940
rect 179650 157928 179656 157940
rect 177408 157900 179656 157928
rect 177408 157888 177414 157900
rect 179650 157888 179656 157900
rect 179708 157888 179714 157940
rect 105406 156936 105412 156988
rect 105464 156976 105470 156988
rect 107246 156976 107252 156988
rect 105464 156948 107252 156976
rect 105464 156936 105470 156948
rect 107246 156936 107252 156948
rect 107304 156936 107310 156988
rect 222798 156868 222804 156920
rect 222856 156908 222862 156920
rect 223534 156908 223540 156920
rect 222856 156880 223540 156908
rect 222856 156868 222862 156880
rect 223534 156868 223540 156880
rect 223592 156868 223598 156920
rect 177534 156460 177540 156512
rect 177592 156500 177598 156512
rect 180478 156500 180484 156512
rect 177592 156472 180484 156500
rect 177592 156460 177598 156472
rect 180478 156460 180484 156472
rect 180536 156460 180542 156512
rect 105222 155712 105228 155764
rect 105280 155752 105286 155764
rect 107154 155752 107160 155764
rect 105280 155724 107160 155752
rect 105280 155712 105286 155724
rect 107154 155712 107160 155724
rect 107212 155712 107218 155764
rect 177534 155100 177540 155152
rect 177592 155140 177598 155152
rect 180386 155140 180392 155152
rect 177592 155112 180392 155140
rect 177592 155100 177598 155112
rect 180386 155100 180392 155112
rect 180444 155100 180450 155152
rect 105590 153808 105596 153860
rect 105648 153848 105654 153860
rect 107982 153848 107988 153860
rect 105648 153820 107988 153848
rect 105648 153808 105654 153820
rect 107982 153808 107988 153820
rect 108040 153808 108046 153860
rect 177350 153808 177356 153860
rect 177408 153848 177414 153860
rect 180294 153848 180300 153860
rect 177408 153820 180300 153848
rect 177408 153808 177414 153820
rect 180294 153808 180300 153820
rect 180352 153808 180358 153860
rect 105774 153740 105780 153792
rect 105832 153780 105838 153792
rect 108534 153780 108540 153792
rect 105832 153752 108540 153780
rect 105832 153740 105838 153752
rect 108534 153740 108540 153752
rect 108592 153740 108598 153792
rect 178178 153740 178184 153792
rect 178236 153780 178242 153792
rect 179742 153780 179748 153792
rect 178236 153752 179748 153780
rect 178236 153740 178242 153752
rect 179742 153740 179748 153752
rect 179800 153740 179806 153792
rect 57474 151496 57480 151548
rect 57532 151536 57538 151548
rect 59590 151536 59596 151548
rect 57532 151508 59596 151536
rect 57532 151496 57538 151508
rect 59590 151496 59596 151508
rect 59648 151496 59654 151548
rect 200534 151496 200540 151548
rect 200592 151536 200598 151548
rect 207434 151536 207440 151548
rect 200592 151508 207440 151536
rect 200592 151496 200598 151508
rect 207434 151496 207440 151508
rect 207492 151496 207498 151548
rect 28770 146912 28776 146924
rect 28731 146884 28776 146912
rect 28770 146872 28776 146884
rect 28828 146872 28834 146924
rect 178270 146600 178276 146652
rect 178328 146640 178334 146652
rect 179006 146640 179012 146652
rect 178328 146612 179012 146640
rect 178328 146600 178334 146612
rect 179006 146600 179012 146612
rect 179064 146600 179070 146652
rect 105866 145444 105872 145496
rect 105924 145484 105930 145496
rect 105924 145456 107752 145484
rect 105924 145444 105930 145456
rect 107724 145416 107752 145456
rect 109270 145416 109276 145428
rect 107724 145388 109276 145416
rect 109270 145376 109276 145388
rect 109328 145376 109334 145428
rect 178270 145240 178276 145292
rect 178328 145280 178334 145292
rect 181122 145280 181128 145292
rect 178328 145252 181128 145280
rect 178328 145240 178334 145252
rect 181122 145240 181128 145252
rect 181180 145240 181186 145292
rect 22238 145172 22244 145224
rect 22296 145212 22302 145224
rect 28773 145215 28831 145221
rect 28773 145212 28785 145215
rect 22296 145184 28785 145212
rect 22296 145172 22302 145184
rect 28773 145181 28785 145184
rect 28819 145181 28831 145215
rect 28773 145175 28831 145181
rect 177442 145036 177448 145088
rect 177500 145076 177506 145088
rect 180570 145076 180576 145088
rect 177500 145048 180576 145076
rect 177500 145036 177506 145048
rect 180570 145036 180576 145048
rect 180628 145036 180634 145088
rect 191840 144696 191846 144748
rect 191898 144736 191904 144748
rect 194278 144736 194284 144748
rect 191898 144708 194284 144736
rect 191898 144696 191904 144708
rect 194278 144696 194284 144708
rect 194336 144696 194342 144748
rect 191472 144628 191478 144680
rect 191530 144668 191536 144680
rect 193634 144668 193640 144680
rect 191530 144640 193640 144668
rect 191530 144628 191536 144640
rect 193634 144628 193640 144640
rect 193692 144628 193698 144680
rect 197820 144628 197826 144680
rect 197878 144668 197884 144680
rect 202834 144668 202840 144680
rect 197878 144640 202840 144668
rect 197878 144628 197884 144640
rect 202834 144628 202840 144640
rect 202892 144628 202898 144680
rect 52506 144492 52512 144544
rect 52564 144532 52570 144544
rect 55358 144532 55364 144544
rect 52564 144504 55364 144532
rect 52564 144492 52570 144504
rect 55358 144492 55364 144504
rect 55416 144492 55422 144544
rect 54622 144220 54628 144272
rect 54680 144260 54686 144272
rect 60418 144260 60424 144272
rect 54680 144232 60424 144260
rect 54680 144220 54686 144232
rect 60418 144220 60424 144232
rect 60476 144220 60482 144272
rect 125830 144220 125836 144272
rect 125888 144260 125894 144272
rect 131442 144260 131448 144272
rect 125888 144232 131448 144260
rect 125888 144220 125894 144232
rect 131442 144220 131448 144232
rect 131500 144220 131506 144272
rect 190598 144220 190604 144272
rect 190656 144260 190662 144272
rect 192530 144260 192536 144272
rect 190656 144232 192536 144260
rect 190656 144220 190662 144232
rect 192530 144220 192536 144232
rect 192588 144220 192594 144272
rect 198510 144220 198516 144272
rect 198568 144260 198574 144272
rect 203386 144260 203392 144272
rect 198568 144232 203392 144260
rect 198568 144220 198574 144232
rect 203386 144220 203392 144232
rect 203444 144220 203450 144272
rect 40638 144152 40644 144204
rect 40696 144192 40702 144204
rect 43030 144192 43036 144204
rect 40696 144164 43036 144192
rect 40696 144152 40702 144164
rect 43030 144152 43036 144164
rect 43088 144152 43094 144204
rect 54254 144152 54260 144204
rect 54312 144192 54318 144204
rect 59774 144192 59780 144204
rect 54312 144164 59780 144192
rect 54312 144152 54318 144164
rect 59774 144152 59780 144164
rect 59832 144152 59838 144204
rect 106418 144152 106424 144204
rect 106476 144192 106482 144204
rect 108350 144192 108356 144204
rect 106476 144164 108356 144192
rect 106476 144152 106482 144164
rect 108350 144152 108356 144164
rect 108408 144152 108414 144204
rect 120310 144152 120316 144204
rect 120368 144192 120374 144204
rect 122334 144192 122340 144204
rect 120368 144164 122340 144192
rect 120368 144152 120374 144164
rect 122334 144152 122340 144164
rect 122392 144152 122398 144204
rect 126658 144152 126664 144204
rect 126716 144192 126722 144204
rect 132178 144192 132184 144204
rect 126716 144164 132184 144192
rect 126716 144152 126722 144164
rect 132178 144152 132184 144164
rect 132236 144152 132242 144204
rect 198878 144152 198884 144204
rect 198936 144192 198942 144204
rect 203938 144192 203944 144204
rect 198936 144164 203944 144192
rect 198936 144152 198942 144164
rect 203938 144152 203944 144164
rect 203996 144152 204002 144204
rect 41282 144084 41288 144136
rect 41340 144124 41346 144136
rect 43398 144124 43404 144136
rect 41340 144096 43404 144124
rect 41340 144084 41346 144096
rect 43398 144084 43404 144096
rect 43456 144084 43462 144136
rect 55358 144084 55364 144136
rect 55416 144084 55422 144136
rect 56370 144124 56376 144136
rect 55468 144096 56376 144124
rect 55376 144056 55404 144084
rect 55468 144056 55496 144096
rect 56370 144084 56376 144096
rect 56428 144084 56434 144136
rect 106510 144084 106516 144136
rect 106568 144124 106574 144136
rect 107154 144124 107160 144136
rect 106568 144096 107160 144124
rect 106568 144084 106574 144096
rect 107154 144084 107160 144096
rect 107212 144084 107218 144136
rect 118930 144084 118936 144136
rect 118988 144124 118994 144136
rect 120586 144124 120592 144136
rect 118988 144096 120592 144124
rect 118988 144084 118994 144096
rect 120586 144084 120592 144096
rect 120644 144084 120650 144136
rect 126290 144084 126296 144136
rect 126348 144124 126354 144136
rect 131626 144124 131632 144136
rect 126348 144096 131632 144124
rect 126348 144084 126354 144096
rect 131626 144084 131632 144096
rect 131684 144084 131690 144136
rect 55376 144028 55496 144056
rect 34106 142656 34112 142708
rect 34164 142696 34170 142708
rect 39074 142696 39080 142708
rect 34164 142668 39080 142696
rect 34164 142656 34170 142668
rect 39074 142656 39080 142668
rect 39132 142656 39138 142708
rect 39994 142656 40000 142708
rect 40052 142696 40058 142708
rect 42294 142696 42300 142708
rect 40052 142668 42300 142696
rect 40052 142656 40058 142668
rect 42294 142656 42300 142668
rect 42352 142656 42358 142708
rect 42662 142656 42668 142708
rect 42720 142696 42726 142708
rect 44226 142696 44232 142708
rect 42720 142668 44232 142696
rect 42720 142656 42726 142668
rect 44226 142656 44232 142668
rect 44284 142656 44290 142708
rect 47814 142656 47820 142708
rect 47872 142696 47878 142708
rect 48826 142696 48832 142708
rect 47872 142668 48832 142696
rect 47872 142656 47878 142668
rect 48826 142656 48832 142668
rect 48884 142656 48890 142708
rect 49010 142656 49016 142708
rect 49068 142696 49074 142708
rect 50850 142696 50856 142708
rect 49068 142668 50856 142696
rect 49068 142656 49074 142668
rect 50850 142656 50856 142668
rect 50908 142656 50914 142708
rect 51034 142656 51040 142708
rect 51092 142696 51098 142708
rect 54254 142696 54260 142708
rect 51092 142668 54260 142696
rect 51092 142656 51098 142668
rect 54254 142656 54260 142668
rect 54312 142656 54318 142708
rect 62810 142656 62816 142708
rect 62868 142696 62874 142708
rect 62868 142668 65156 142696
rect 62868 142656 62874 142668
rect 16626 142588 16632 142640
rect 16684 142628 16690 142640
rect 31806 142628 31812 142640
rect 16684 142600 31812 142628
rect 16684 142588 16690 142600
rect 31806 142588 31812 142600
rect 31864 142628 31870 142640
rect 36133 142631 36191 142637
rect 36133 142628 36145 142631
rect 31864 142600 36145 142628
rect 31864 142588 31870 142600
rect 36133 142597 36145 142600
rect 36179 142597 36191 142631
rect 36133 142591 36191 142597
rect 34658 142520 34664 142572
rect 34716 142560 34722 142572
rect 39442 142560 39448 142572
rect 34716 142532 39448 142560
rect 34716 142520 34722 142532
rect 39442 142520 39448 142532
rect 39500 142520 39506 142572
rect 42018 142520 42024 142572
rect 42076 142560 42082 142572
rect 43858 142560 43864 142572
rect 42076 142532 43864 142560
rect 42076 142520 42082 142532
rect 43858 142520 43864 142532
rect 43916 142520 43922 142572
rect 43953 142563 44011 142569
rect 43953 142529 43965 142563
rect 43999 142560 44011 142563
rect 48185 142563 48243 142569
rect 48185 142560 48197 142563
rect 43999 142532 48197 142560
rect 43999 142529 44011 142532
rect 43953 142523 44011 142529
rect 48185 142529 48197 142532
rect 48231 142529 48243 142563
rect 48185 142523 48243 142529
rect 48274 142520 48280 142572
rect 48332 142560 48338 142572
rect 49470 142560 49476 142572
rect 48332 142532 49476 142560
rect 48332 142520 48338 142532
rect 49470 142520 49476 142532
rect 49528 142520 49534 142572
rect 50482 142520 50488 142572
rect 50540 142560 50546 142572
rect 52966 142560 52972 142572
rect 50540 142532 52972 142560
rect 50540 142520 50546 142532
rect 52966 142520 52972 142532
rect 53024 142520 53030 142572
rect 65128 142560 65156 142668
rect 66490 142656 66496 142708
rect 66548 142696 66554 142708
rect 67870 142696 67876 142708
rect 66548 142668 67876 142696
rect 66548 142656 66554 142668
rect 67870 142656 67876 142668
rect 67928 142656 67934 142708
rect 72838 142656 72844 142708
rect 72896 142696 72902 142708
rect 74494 142696 74500 142708
rect 72896 142668 74500 142696
rect 72896 142656 72902 142668
rect 74494 142656 74500 142668
rect 74552 142656 74558 142708
rect 74770 142656 74776 142708
rect 74828 142696 74834 142708
rect 75598 142696 75604 142708
rect 74828 142668 75604 142696
rect 74828 142656 74834 142668
rect 75598 142656 75604 142668
rect 75656 142656 75662 142708
rect 80106 142656 80112 142708
rect 80164 142696 80170 142708
rect 81670 142696 81676 142708
rect 80164 142668 81676 142696
rect 80164 142656 80170 142668
rect 81670 142656 81676 142668
rect 81728 142656 81734 142708
rect 85626 142656 85632 142708
rect 85684 142696 85690 142708
rect 90962 142696 90968 142708
rect 85684 142668 90968 142696
rect 85684 142656 85690 142668
rect 90962 142656 90968 142668
rect 91020 142656 91026 142708
rect 95470 142656 95476 142708
rect 95528 142696 95534 142708
rect 96758 142696 96764 142708
rect 95528 142668 96764 142696
rect 95528 142656 95534 142668
rect 96758 142656 96764 142668
rect 96816 142656 96822 142708
rect 117458 142656 117464 142708
rect 117516 142696 117522 142708
rect 118838 142696 118844 142708
rect 117516 142668 118844 142696
rect 117516 142656 117522 142668
rect 118838 142656 118844 142668
rect 118896 142656 118902 142708
rect 120678 142656 120684 142708
rect 120736 142696 120742 142708
rect 123438 142696 123444 142708
rect 120736 142668 123444 142696
rect 120736 142656 120742 142668
rect 123438 142656 123444 142668
rect 123496 142656 123502 142708
rect 125094 142656 125100 142708
rect 125152 142696 125158 142708
rect 129878 142696 129884 142708
rect 125152 142668 129884 142696
rect 125152 142656 125158 142668
rect 129878 142656 129884 142668
rect 129936 142656 129942 142708
rect 142666 142656 142672 142708
rect 142724 142696 142730 142708
rect 145426 142696 145432 142708
rect 142724 142668 145432 142696
rect 142724 142656 142730 142668
rect 145426 142656 145432 142668
rect 145484 142656 145490 142708
rect 146438 142656 146444 142708
rect 146496 142696 146502 142708
rect 147634 142696 147640 142708
rect 146496 142668 147640 142696
rect 146496 142656 146502 142668
rect 147634 142656 147640 142668
rect 147692 142656 147698 142708
rect 154350 142656 154356 142708
rect 154408 142696 154414 142708
rect 157662 142696 157668 142708
rect 154408 142668 157668 142696
rect 154408 142656 154414 142668
rect 157662 142656 157668 142668
rect 157720 142656 157726 142708
rect 165850 142656 165856 142708
rect 165908 142696 165914 142708
rect 166586 142696 166592 142708
rect 165908 142668 166592 142696
rect 165908 142656 165914 142668
rect 166586 142656 166592 142668
rect 166644 142656 166650 142708
rect 182226 142656 182232 142708
rect 182284 142696 182290 142708
rect 183238 142696 183244 142708
rect 182284 142668 183244 142696
rect 182284 142656 182290 142668
rect 183238 142656 183244 142668
rect 183296 142656 183302 142708
rect 189678 142656 189684 142708
rect 189736 142696 189742 142708
rect 190782 142696 190788 142708
rect 189736 142668 190788 142696
rect 189736 142656 189742 142668
rect 190782 142656 190788 142668
rect 190840 142656 190846 142708
rect 191334 142656 191340 142708
rect 191392 142696 191398 142708
rect 193082 142696 193088 142708
rect 191392 142668 193088 142696
rect 191392 142656 191398 142668
rect 193082 142656 193088 142668
rect 193140 142656 193146 142708
rect 194094 142656 194100 142708
rect 194152 142696 194158 142708
rect 197130 142696 197136 142708
rect 194152 142668 197136 142696
rect 194152 142656 194158 142668
rect 197130 142656 197136 142668
rect 197188 142656 197194 142708
rect 200994 142656 201000 142708
rect 201052 142696 201058 142708
rect 215898 142696 215904 142708
rect 201052 142668 215904 142696
rect 201052 142656 201058 142668
rect 215898 142656 215904 142668
rect 215956 142656 215962 142708
rect 81210 142588 81216 142640
rect 81268 142628 81274 142640
rect 83510 142628 83516 142640
rect 81268 142600 83516 142628
rect 81268 142588 81274 142600
rect 83510 142588 83516 142600
rect 83568 142588 83574 142640
rect 86730 142588 86736 142640
rect 86788 142628 86794 142640
rect 92802 142628 92808 142640
rect 86788 142600 92808 142628
rect 86788 142588 86794 142600
rect 92802 142588 92808 142600
rect 92860 142588 92866 142640
rect 118286 142588 118292 142640
rect 118344 142628 118350 142640
rect 119942 142628 119948 142640
rect 118344 142600 119948 142628
rect 118344 142588 118350 142600
rect 119942 142588 119948 142600
rect 120000 142588 120006 142640
rect 125462 142588 125468 142640
rect 125520 142628 125526 142640
rect 130430 142628 130436 142640
rect 125520 142600 130436 142628
rect 125520 142588 125526 142600
rect 130430 142588 130436 142600
rect 130488 142588 130494 142640
rect 165482 142588 165488 142640
rect 165540 142628 165546 142640
rect 169346 142628 169352 142640
rect 165540 142600 169352 142628
rect 165540 142588 165546 142600
rect 169346 142588 169352 142600
rect 169404 142588 169410 142640
rect 189310 142588 189316 142640
rect 189368 142628 189374 142640
rect 190230 142628 190236 142640
rect 189368 142600 190236 142628
rect 189368 142588 189374 142600
rect 190230 142588 190236 142600
rect 190288 142588 190294 142640
rect 196946 142588 196952 142640
rect 197004 142628 197010 142640
rect 201086 142628 201092 142640
rect 197004 142600 201092 142628
rect 197004 142588 197010 142600
rect 201086 142588 201092 142600
rect 201144 142588 201150 142640
rect 71182 142560 71188 142572
rect 65128 142532 71188 142560
rect 71182 142520 71188 142532
rect 71240 142520 71246 142572
rect 121046 142520 121052 142572
rect 121104 142560 121110 142572
rect 124450 142560 124456 142572
rect 121104 142532 124456 142560
rect 121104 142520 121110 142532
rect 124450 142520 124456 142532
rect 124508 142520 124514 142572
rect 124634 142520 124640 142572
rect 124692 142560 124698 142572
rect 129326 142560 129332 142572
rect 124692 142532 129332 142560
rect 124692 142520 124698 142532
rect 129326 142520 129332 142532
rect 129384 142520 129390 142572
rect 134478 142520 134484 142572
rect 134536 142560 134542 142572
rect 143218 142560 143224 142572
rect 134536 142532 143224 142560
rect 134536 142520 134542 142532
rect 143218 142520 143224 142532
rect 143276 142520 143282 142572
rect 197314 142520 197320 142572
rect 197372 142560 197378 142572
rect 201638 142560 201644 142572
rect 197372 142532 201644 142560
rect 197372 142520 197378 142532
rect 201638 142520 201644 142532
rect 201696 142520 201702 142572
rect 27574 142452 27580 142504
rect 27632 142492 27638 142504
rect 27632 142464 48596 142492
rect 27632 142452 27638 142464
rect 37234 142384 37240 142436
rect 37292 142424 37298 142436
rect 41006 142424 41012 142436
rect 37292 142396 41012 142424
rect 37292 142384 37298 142396
rect 41006 142384 41012 142396
rect 41064 142384 41070 142436
rect 39258 142316 39264 142368
rect 39316 142356 39322 142368
rect 42202 142356 42208 142368
rect 39316 142328 42208 142356
rect 39316 142316 39322 142328
rect 42202 142316 42208 142328
rect 42260 142316 42266 142368
rect 48568 142356 48596 142464
rect 48642 142452 48648 142504
rect 48700 142492 48706 142504
rect 50206 142492 50212 142504
rect 48700 142464 50212 142492
rect 48700 142452 48706 142464
rect 50206 142452 50212 142464
rect 50264 142452 50270 142504
rect 50666 142452 50672 142504
rect 50724 142492 50730 142504
rect 53610 142492 53616 142504
rect 50724 142464 53616 142492
rect 50724 142452 50730 142464
rect 53610 142452 53616 142464
rect 53668 142452 53674 142504
rect 87834 142452 87840 142504
rect 87892 142492 87898 142504
rect 94734 142492 94740 142504
rect 87892 142464 94740 142492
rect 87892 142452 87898 142464
rect 94734 142452 94740 142464
rect 94792 142452 94798 142504
rect 102278 142452 102284 142504
rect 102336 142492 102342 142504
rect 174314 142492 174320 142504
rect 102336 142464 174320 142492
rect 102336 142452 102342 142464
rect 174314 142452 174320 142464
rect 174372 142452 174378 142504
rect 190138 142452 190144 142504
rect 190196 142492 190202 142504
rect 191426 142492 191432 142504
rect 190196 142464 191432 142492
rect 190196 142452 190202 142464
rect 191426 142452 191432 142464
rect 191484 142452 191490 142504
rect 194554 142452 194560 142504
rect 194612 142492 194618 142504
rect 197682 142492 197688 142504
rect 194612 142464 197688 142492
rect 194612 142452 194618 142464
rect 197682 142452 197688 142464
rect 197740 142452 197746 142504
rect 51402 142384 51408 142436
rect 51460 142424 51466 142436
rect 54990 142424 54996 142436
rect 51460 142396 54996 142424
rect 51460 142384 51466 142396
rect 54990 142384 54996 142396
rect 55048 142384 55054 142436
rect 69158 142384 69164 142436
rect 69216 142424 69222 142436
rect 72286 142424 72292 142436
rect 69216 142396 72292 142424
rect 69216 142384 69222 142396
rect 72286 142384 72292 142396
rect 72344 142384 72350 142436
rect 101450 142384 101456 142436
rect 101508 142424 101514 142436
rect 173210 142424 173216 142436
rect 101508 142396 173216 142424
rect 101508 142384 101514 142396
rect 173210 142384 173216 142396
rect 173268 142384 173274 142436
rect 192898 142384 192904 142436
rect 192956 142424 192962 142436
rect 195382 142424 195388 142436
rect 192956 142396 195388 142424
rect 192956 142384 192962 142396
rect 195382 142384 195388 142396
rect 195440 142384 195446 142436
rect 195750 142384 195756 142436
rect 195808 142424 195814 142436
rect 199062 142424 199068 142436
rect 195808 142396 199068 142424
rect 195808 142384 195814 142396
rect 199062 142384 199068 142396
rect 199120 142384 199126 142436
rect 54714 142356 54720 142368
rect 48568 142328 54720 142356
rect 54714 142316 54720 142328
rect 54772 142316 54778 142368
rect 83418 142316 83424 142368
rect 83476 142356 83482 142368
rect 87282 142356 87288 142368
rect 83476 142328 87288 142356
rect 83476 142316 83482 142328
rect 87282 142316 87288 142328
rect 87340 142316 87346 142368
rect 98966 142316 98972 142368
rect 99024 142356 99030 142368
rect 102278 142356 102284 142368
rect 99024 142328 102284 142356
rect 99024 142316 99030 142328
rect 102278 142316 102284 142328
rect 102336 142316 102342 142368
rect 119482 142316 119488 142368
rect 119540 142356 119546 142368
rect 121690 142356 121696 142368
rect 119540 142328 121696 142356
rect 119540 142316 119546 142328
rect 121690 142316 121696 142328
rect 121748 142316 121754 142368
rect 123898 142316 123904 142368
rect 123956 142356 123962 142368
rect 128130 142356 128136 142368
rect 123956 142328 128136 142356
rect 123956 142316 123962 142328
rect 128130 142316 128136 142328
rect 128188 142316 128194 142368
rect 160974 142316 160980 142368
rect 161032 142356 161038 142368
rect 168886 142356 168892 142368
rect 161032 142328 168892 142356
rect 161032 142316 161038 142328
rect 168886 142316 168892 142328
rect 168944 142316 168950 142368
rect 181674 142316 181680 142368
rect 181732 142356 181738 142368
rect 182778 142356 182784 142368
rect 181732 142328 182784 142356
rect 181732 142316 181738 142328
rect 182778 142316 182784 142328
rect 182836 142316 182842 142368
rect 192438 142316 192444 142368
rect 192496 142356 192502 142368
rect 194830 142356 194836 142368
rect 192496 142328 194836 142356
rect 192496 142316 192502 142328
rect 194830 142316 194836 142328
rect 194888 142316 194894 142368
rect 196118 142316 196124 142368
rect 196176 142356 196182 142368
rect 199614 142356 199620 142368
rect 196176 142328 199620 142356
rect 196176 142316 196182 142328
rect 199614 142316 199620 142328
rect 199672 142316 199678 142368
rect 36590 142248 36596 142300
rect 36648 142288 36654 142300
rect 40362 142288 40368 142300
rect 36648 142260 40368 142288
rect 36648 142248 36654 142260
rect 40362 142248 40368 142260
rect 40420 142248 40426 142300
rect 43398 142248 43404 142300
rect 43456 142288 43462 142300
rect 44594 142288 44600 142300
rect 43456 142260 44600 142288
rect 43456 142248 43462 142260
rect 44594 142248 44600 142260
rect 44652 142248 44658 142300
rect 45422 142248 45428 142300
rect 45480 142288 45486 142300
rect 45790 142288 45796 142300
rect 45480 142260 45796 142288
rect 45480 142248 45486 142260
rect 45790 142248 45796 142260
rect 45848 142248 45854 142300
rect 49746 142248 49752 142300
rect 49804 142288 49810 142300
rect 51586 142288 51592 142300
rect 49804 142260 51592 142288
rect 49804 142248 49810 142260
rect 51586 142248 51592 142260
rect 51644 142248 51650 142300
rect 51681 142291 51739 142297
rect 51681 142257 51693 142291
rect 51727 142288 51739 142291
rect 51727 142260 54944 142288
rect 51727 142257 51739 142260
rect 51681 142251 51739 142257
rect 38614 142180 38620 142232
rect 38672 142220 38678 142232
rect 41834 142220 41840 142232
rect 38672 142192 41840 142220
rect 38672 142180 38678 142192
rect 41834 142180 41840 142192
rect 41892 142180 41898 142232
rect 54916 142220 54944 142260
rect 93446 142248 93452 142300
rect 93504 142288 93510 142300
rect 98138 142288 98144 142300
rect 93504 142260 98144 142288
rect 93504 142248 93510 142260
rect 98138 142248 98144 142260
rect 98196 142248 98202 142300
rect 123714 142248 123720 142300
rect 123772 142288 123778 142300
rect 127578 142288 127584 142300
rect 123772 142260 127584 142288
rect 123772 142248 123778 142260
rect 127578 142248 127584 142260
rect 127636 142248 127642 142300
rect 159870 142248 159876 142300
rect 159928 142288 159934 142300
rect 167046 142288 167052 142300
rect 159928 142260 167052 142288
rect 159928 142248 159934 142260
rect 167046 142248 167052 142260
rect 167104 142248 167110 142300
rect 172106 142248 172112 142300
rect 172164 142288 172170 142300
rect 174590 142288 174596 142300
rect 172164 142260 174596 142288
rect 172164 142248 172170 142260
rect 174590 142248 174596 142260
rect 174648 142248 174654 142300
rect 194646 142248 194652 142300
rect 194704 142288 194710 142300
rect 198234 142288 198240 142300
rect 194704 142260 198240 142288
rect 194704 142248 194710 142260
rect 198234 142248 198240 142260
rect 198292 142248 198298 142300
rect 57474 142220 57480 142232
rect 54916 142192 57480 142220
rect 57474 142180 57480 142192
rect 57532 142180 57538 142232
rect 92342 142180 92348 142232
rect 92400 142220 92406 142232
rect 97218 142220 97224 142232
rect 92400 142192 97224 142220
rect 92400 142180 92406 142192
rect 97218 142180 97224 142192
rect 97276 142180 97282 142232
rect 121506 142180 121512 142232
rect 121564 142220 121570 142232
rect 124634 142220 124640 142232
rect 121564 142192 124640 142220
rect 121564 142180 121570 142192
rect 124634 142180 124640 142192
rect 124692 142180 124698 142232
rect 168794 142180 168800 142232
rect 168852 142220 168858 142232
rect 172750 142220 172756 142232
rect 168852 142192 172756 142220
rect 168852 142180 168858 142192
rect 172750 142180 172756 142192
rect 172808 142180 172814 142232
rect 195290 142180 195296 142232
rect 195348 142220 195354 142232
rect 198786 142220 198792 142232
rect 195348 142192 198792 142220
rect 195348 142180 195354 142192
rect 198786 142180 198792 142192
rect 198844 142180 198850 142232
rect 37878 142112 37884 142164
rect 37936 142152 37942 142164
rect 41466 142152 41472 142164
rect 37936 142124 41472 142152
rect 37936 142112 37942 142124
rect 41466 142112 41472 142124
rect 41524 142112 41530 142164
rect 49838 142112 49844 142164
rect 49896 142152 49902 142164
rect 52230 142152 52236 142164
rect 49896 142124 52236 142152
rect 49896 142112 49902 142124
rect 52230 142112 52236 142124
rect 52288 142112 52294 142164
rect 52598 142112 52604 142164
rect 52656 142152 52662 142164
rect 57014 142152 57020 142164
rect 52656 142124 57020 142152
rect 52656 142112 52662 142124
rect 57014 142112 57020 142124
rect 57072 142112 57078 142164
rect 62350 142112 62356 142164
rect 62408 142152 62414 142164
rect 63454 142152 63460 142164
rect 62408 142124 63460 142152
rect 62408 142112 62414 142124
rect 63454 142112 63460 142124
rect 63512 142112 63518 142164
rect 117090 142112 117096 142164
rect 117148 142152 117154 142164
rect 118194 142152 118200 142164
rect 117148 142124 118200 142152
rect 117148 142112 117154 142124
rect 118194 142112 118200 142124
rect 118252 142112 118258 142164
rect 123070 142112 123076 142164
rect 123128 142152 123134 142164
rect 126934 142152 126940 142164
rect 123128 142124 126940 142152
rect 123128 142112 123134 142124
rect 126934 142112 126940 142124
rect 126992 142112 126998 142164
rect 158766 142112 158772 142164
rect 158824 142152 158830 142164
rect 165114 142152 165120 142164
rect 158824 142124 165120 142152
rect 158824 142112 158830 142124
rect 165114 142112 165120 142124
rect 165172 142112 165178 142164
rect 190506 142112 190512 142164
rect 190564 142152 190570 142164
rect 191978 142152 191984 142164
rect 190564 142124 191984 142152
rect 190564 142112 190570 142124
rect 191978 142112 191984 142124
rect 192036 142112 192042 142164
rect 193358 142112 193364 142164
rect 193416 142152 193422 142164
rect 195934 142152 195940 142164
rect 193416 142124 195940 142152
rect 193416 142112 193422 142124
rect 195934 142112 195940 142124
rect 195992 142112 195998 142164
rect 196486 142112 196492 142164
rect 196544 142152 196550 142164
rect 200534 142152 200540 142164
rect 196544 142124 200540 142152
rect 196544 142112 196550 142124
rect 200534 142112 200540 142124
rect 200592 142112 200598 142164
rect 36133 142087 36191 142093
rect 36133 142053 36145 142087
rect 36179 142084 36191 142087
rect 43953 142087 44011 142093
rect 43953 142084 43965 142087
rect 36179 142056 43965 142084
rect 36179 142053 36191 142056
rect 36133 142047 36191 142053
rect 43953 142053 43965 142056
rect 43999 142053 44011 142087
rect 43953 142047 44011 142053
rect 48185 142087 48243 142093
rect 48185 142053 48197 142087
rect 48231 142084 48243 142087
rect 51681 142087 51739 142093
rect 51681 142084 51693 142087
rect 48231 142056 51693 142084
rect 48231 142053 48243 142056
rect 48185 142047 48243 142053
rect 51681 142053 51693 142056
rect 51727 142053 51739 142087
rect 51681 142047 51739 142053
rect 51862 142044 51868 142096
rect 51920 142084 51926 142096
rect 55358 142084 55364 142096
rect 51920 142056 55364 142084
rect 51920 142044 51926 142056
rect 55358 142044 55364 142056
rect 55416 142044 55422 142096
rect 182870 142044 182876 142096
rect 182928 142084 182934 142096
rect 183606 142084 183612 142096
rect 182928 142056 183612 142084
rect 182928 142044 182934 142056
rect 183606 142044 183612 142056
rect 183664 142044 183670 142096
rect 222522 142044 222528 142096
rect 222580 142084 222586 142096
rect 222798 142084 222804 142096
rect 222580 142056 222804 142084
rect 222580 142044 222586 142056
rect 222798 142044 222804 142056
rect 222856 142044 222862 142096
rect 53058 141976 53064 142028
rect 53116 142016 53122 142028
rect 57658 142016 57664 142028
rect 53116 141988 57664 142016
rect 53116 141976 53122 141988
rect 57658 141976 57664 141988
rect 57716 141976 57722 142028
rect 63454 141976 63460 142028
rect 63512 142016 63518 142028
rect 64558 142016 64564 142028
rect 63512 141988 64564 142016
rect 63512 141976 63518 141988
rect 64558 141976 64564 141988
rect 64616 141976 64622 142028
rect 88938 141976 88944 142028
rect 88996 142016 89002 142028
rect 96850 142016 96856 142028
rect 88996 141988 96856 142016
rect 88996 141976 89002 141988
rect 96850 141976 96856 141988
rect 96908 141976 96914 142028
rect 110420 141976 110426 142028
rect 110478 142016 110484 142028
rect 111478 142016 111484 142028
rect 110478 141988 111484 142016
rect 110478 141976 110484 141988
rect 111478 141976 111484 141988
rect 111536 141976 111542 142028
rect 113272 141976 113278 142028
rect 113330 142016 113336 142028
rect 113502 142016 113508 142028
rect 113330 141988 113508 142016
rect 113330 141976 113336 141988
rect 113502 141976 113508 141988
rect 113560 141976 113566 142028
rect 116262 141976 116268 142028
rect 116320 142016 116326 142028
rect 117412 142016 117418 142028
rect 116320 141988 117418 142016
rect 116320 141976 116326 141988
rect 117412 141976 117418 141988
rect 117470 141976 117476 142028
rect 117826 141976 117832 142028
rect 117884 142016 117890 142028
rect 119712 142016 119718 142028
rect 117884 141988 119718 142016
rect 117884 141976 117890 141988
rect 119712 141976 119718 141988
rect 119770 141976 119776 142028
rect 120494 141976 120500 142028
rect 120552 142016 120558 142028
rect 123208 142016 123214 142028
rect 120552 141988 123214 142016
rect 120552 141976 120558 141988
rect 123208 141976 123214 141988
rect 123266 141976 123272 142028
rect 124266 141976 124272 142028
rect 124324 142016 124330 142028
rect 129004 142016 129010 142028
rect 124324 141988 129010 142016
rect 124324 141976 124330 141988
rect 129004 141976 129010 141988
rect 129062 141976 129068 142028
rect 164378 141976 164384 142028
rect 164436 142016 164442 142028
rect 169254 142016 169260 142028
rect 164436 141988 169260 142016
rect 164436 141976 164442 141988
rect 169254 141976 169260 141988
rect 169312 141976 169318 142028
rect 193726 141976 193732 142028
rect 193784 142016 193790 142028
rect 196486 142016 196492 142028
rect 193784 141988 196492 142016
rect 193784 141976 193790 141988
rect 196486 141976 196492 141988
rect 196544 141976 196550 142028
rect 207986 141976 207992 142028
rect 208044 142016 208050 142028
rect 221234 142016 221240 142028
rect 208044 141988 221240 142016
rect 208044 141976 208050 141988
rect 221234 141976 221240 141988
rect 221292 141976 221298 142028
rect 109776 141908 109782 141960
rect 109834 141948 109840 141960
rect 111110 141948 111116 141960
rect 109834 141920 111116 141948
rect 109834 141908 109840 141920
rect 111110 141908 111116 141920
rect 111168 141908 111174 141960
rect 116630 141908 116636 141960
rect 116688 141948 116694 141960
rect 117964 141948 117970 141960
rect 116688 141920 117970 141948
rect 116688 141908 116694 141920
rect 117964 141908 117970 141920
rect 118022 141908 118028 141960
rect 119114 141908 119120 141960
rect 119172 141948 119178 141960
rect 121460 141948 121466 141960
rect 119172 141920 121466 141948
rect 119172 141908 119178 141920
rect 121460 141908 121466 141920
rect 121518 141908 121524 141960
rect 121874 141908 121880 141960
rect 121932 141948 121938 141960
rect 125508 141948 125514 141960
rect 121932 141920 125514 141948
rect 121932 141908 121938 141920
rect 125508 141908 125514 141920
rect 125566 141908 125572 141960
rect 153246 141908 153252 141960
rect 153304 141948 153310 141960
rect 155822 141948 155828 141960
rect 153304 141920 155828 141948
rect 153304 141908 153310 141920
rect 155822 141908 155828 141920
rect 155880 141908 155886 141960
rect 207894 141908 207900 141960
rect 207952 141948 207958 141960
rect 210562 141948 210568 141960
rect 207952 141920 210568 141948
rect 207952 141908 207958 141920
rect 210562 141908 210568 141920
rect 210620 141908 210626 141960
rect 222522 141908 222528 141960
rect 222580 141948 222586 141960
rect 223534 141948 223540 141960
rect 222580 141920 223540 141948
rect 222580 141908 222586 141920
rect 223534 141908 223540 141920
rect 223592 141908 223598 141960
rect 70998 141840 71004 141892
rect 71056 141880 71062 141892
rect 73390 141880 73396 141892
rect 71056 141852 73396 141880
rect 71056 141840 71062 141852
rect 73390 141840 73396 141852
rect 73448 141840 73454 141892
rect 84522 141840 84528 141892
rect 84580 141880 84586 141892
rect 89122 141880 89128 141892
rect 84580 141852 89128 141880
rect 84580 141840 84586 141852
rect 89122 141840 89128 141852
rect 89180 141840 89186 141892
rect 132362 141880 132368 141892
rect 132323 141852 132368 141880
rect 132362 141840 132368 141852
rect 132420 141840 132426 141892
rect 35578 141772 35584 141824
rect 35636 141812 35642 141824
rect 39810 141812 39816 141824
rect 35636 141784 39816 141812
rect 35636 141772 35642 141784
rect 39810 141772 39816 141784
rect 39868 141772 39874 141824
rect 122886 141772 122892 141824
rect 122944 141812 122950 141824
rect 126382 141812 126388 141824
rect 122944 141784 126388 141812
rect 122944 141772 122950 141784
rect 126382 141772 126388 141784
rect 126440 141772 126446 141824
rect 152142 141772 152148 141824
rect 152200 141812 152206 141824
rect 153890 141812 153896 141824
rect 152200 141784 153896 141812
rect 152200 141772 152206 141784
rect 153890 141772 153896 141784
rect 153948 141772 153954 141824
rect 197406 141772 197412 141824
rect 197464 141812 197470 141824
rect 201822 141812 201828 141824
rect 197464 141784 201828 141812
rect 197464 141772 197470 141784
rect 201822 141772 201828 141784
rect 201880 141772 201886 141824
rect 58670 141744 58676 141756
rect 57216 141716 58676 141744
rect 35946 141636 35952 141688
rect 36004 141636 36010 141688
rect 40178 141636 40184 141688
rect 40236 141636 40242 141688
rect 53426 141636 53432 141688
rect 53484 141636 53490 141688
rect 53794 141636 53800 141688
rect 53852 141676 53858 141688
rect 57216 141676 57244 141716
rect 58670 141704 58676 141716
rect 58728 141704 58734 141756
rect 122242 141704 122248 141756
rect 122300 141744 122306 141756
rect 125830 141744 125836 141756
rect 122300 141716 125836 141744
rect 122300 141704 122306 141716
rect 125830 141704 125836 141716
rect 125888 141704 125894 141756
rect 53852 141648 57244 141676
rect 53852 141636 53858 141648
rect 58210 141636 58216 141688
rect 58268 141636 58274 141688
rect 100070 141636 100076 141688
rect 100128 141676 100134 141688
rect 103474 141676 103480 141688
rect 100128 141648 103480 141676
rect 100128 141636 100134 141648
rect 103474 141636 103480 141648
rect 103532 141636 103538 141688
rect 132086 141636 132092 141688
rect 132144 141676 132150 141688
rect 132638 141676 132644 141688
rect 132144 141648 132644 141676
rect 132144 141636 132150 141648
rect 132638 141636 132644 141648
rect 132696 141636 132702 141688
rect 140826 141636 140832 141688
rect 140884 141676 140890 141688
rect 144322 141676 144328 141688
rect 140884 141648 144328 141676
rect 140884 141636 140890 141648
rect 144322 141636 144328 141648
rect 144380 141636 144386 141688
rect 35964 141336 35992 141636
rect 40196 141336 40224 141636
rect 35964 141308 40224 141336
rect 53444 141336 53472 141636
rect 58228 141336 58256 141636
rect 144506 141568 144512 141620
rect 144564 141608 144570 141620
rect 146530 141608 146536 141620
rect 144564 141580 146536 141608
rect 144564 141568 144570 141580
rect 146530 141568 146536 141580
rect 146588 141568 146594 141620
rect 151038 141568 151044 141620
rect 151096 141608 151102 141620
rect 152050 141608 152056 141620
rect 151096 141580 152056 141608
rect 151096 141568 151102 141580
rect 152050 141568 152056 141580
rect 152108 141568 152114 141620
rect 157938 141568 157944 141620
rect 157996 141608 158002 141620
rect 163274 141608 163280 141620
rect 157996 141580 163280 141608
rect 157996 141568 158002 141580
rect 163274 141568 163280 141580
rect 163332 141568 163338 141620
rect 82314 141500 82320 141552
rect 82372 141540 82378 141552
rect 85350 141540 85356 141552
rect 82372 141512 85356 141540
rect 82372 141500 82378 141512
rect 85350 141500 85356 141512
rect 85408 141500 85414 141552
rect 156558 141500 156564 141552
rect 156616 141540 156622 141552
rect 161434 141540 161440 141552
rect 156616 141512 161440 141540
rect 156616 141500 156622 141512
rect 161434 141500 161440 141512
rect 161492 141500 161498 141552
rect 135122 141432 135128 141484
rect 135180 141472 135186 141484
rect 137698 141472 137704 141484
rect 135180 141444 137704 141472
rect 135180 141432 135186 141444
rect 137698 141432 137704 141444
rect 137756 141432 137762 141484
rect 155454 141364 155460 141416
rect 155512 141404 155518 141416
rect 159502 141404 159508 141416
rect 155512 141376 159508 141404
rect 155512 141364 155518 141376
rect 159502 141364 159508 141376
rect 159560 141364 159566 141416
rect 169898 141364 169904 141416
rect 169956 141404 169962 141416
rect 169956 141376 172888 141404
rect 169956 141364 169962 141376
rect 53444 141308 58256 141336
rect 97862 141296 97868 141348
rect 97920 141336 97926 141348
rect 97920 141308 100944 141336
rect 97920 141296 97926 141308
rect 62810 141228 62816 141280
rect 62868 141268 62874 141280
rect 69250 141268 69256 141280
rect 62868 141240 69256 141268
rect 62868 141228 62874 141240
rect 69250 141228 69256 141240
rect 69308 141228 69314 141280
rect 62718 141160 62724 141212
rect 62776 141200 62782 141212
rect 68054 141200 68060 141212
rect 62776 141172 68060 141200
rect 62776 141160 62782 141172
rect 68054 141160 68060 141172
rect 68112 141160 68118 141212
rect 100916 141200 100944 141308
rect 134570 141296 134576 141348
rect 134628 141336 134634 141348
rect 136594 141336 136600 141348
rect 134628 141308 136600 141336
rect 134628 141296 134634 141308
rect 136594 141296 136600 141308
rect 136652 141296 136658 141348
rect 171002 141296 171008 141348
rect 171060 141336 171066 141348
rect 171060 141308 172796 141336
rect 171060 141296 171066 141308
rect 102370 141200 102376 141212
rect 100916 141172 102376 141200
rect 102370 141160 102376 141172
rect 102428 141160 102434 141212
rect 172768 141200 172796 141308
rect 172860 141268 172888 141376
rect 174222 141268 174228 141280
rect 172860 141240 174228 141268
rect 174222 141228 174228 141240
rect 174280 141228 174286 141280
rect 174406 141200 174412 141212
rect 172768 141172 174412 141200
rect 174406 141160 174412 141172
rect 174464 141160 174470 141212
rect 135306 141092 135312 141144
rect 135364 141132 135370 141144
rect 141102 141132 141108 141144
rect 135364 141104 141108 141132
rect 135364 141092 135370 141104
rect 141102 141092 141108 141104
rect 141160 141092 141166 141144
rect 135306 140684 135312 140736
rect 135364 140724 135370 140736
rect 141010 140724 141016 140736
rect 135364 140696 141016 140724
rect 135364 140684 135370 140696
rect 141010 140684 141016 140696
rect 141068 140684 141074 140736
rect 62810 139868 62816 139920
rect 62868 139908 62874 139920
rect 66490 139908 66496 139920
rect 62868 139880 66496 139908
rect 62868 139868 62874 139880
rect 66490 139868 66496 139880
rect 66548 139868 66554 139920
rect 95470 139868 95476 139920
rect 95528 139908 95534 139920
rect 102370 139908 102376 139920
rect 95528 139880 102376 139908
rect 95528 139868 95534 139880
rect 102370 139868 102376 139880
rect 102428 139868 102434 139920
rect 172750 139868 172756 139920
rect 172808 139908 172814 139920
rect 174314 139908 174320 139920
rect 172808 139880 174320 139908
rect 172808 139868 172814 139880
rect 174314 139868 174320 139880
rect 174372 139868 174378 139920
rect 95562 139800 95568 139852
rect 95620 139840 95626 139852
rect 102462 139840 102468 139852
rect 95620 139812 102468 139840
rect 95620 139800 95626 139812
rect 102462 139800 102468 139812
rect 102520 139800 102526 139852
rect 135306 139800 135312 139852
rect 135364 139840 135370 139852
rect 139538 139840 139544 139852
rect 135364 139812 139544 139840
rect 135364 139800 135370 139812
rect 139538 139800 139544 139812
rect 139596 139800 139602 139852
rect 167230 139800 167236 139852
rect 167288 139840 167294 139852
rect 174130 139840 174136 139852
rect 167288 139812 174136 139840
rect 167288 139800 167294 139812
rect 174130 139800 174136 139812
rect 174188 139800 174194 139852
rect 94090 139732 94096 139784
rect 94148 139772 94154 139784
rect 102554 139772 102560 139784
rect 94148 139744 102560 139772
rect 94148 139732 94154 139744
rect 102554 139732 102560 139744
rect 102612 139732 102618 139784
rect 165850 139732 165856 139784
rect 165908 139772 165914 139784
rect 174222 139772 174228 139784
rect 165908 139744 174228 139772
rect 165908 139732 165914 139744
rect 174222 139732 174228 139744
rect 174280 139732 174286 139784
rect 62350 139664 62356 139716
rect 62408 139704 62414 139716
rect 66582 139704 66588 139716
rect 62408 139676 66588 139704
rect 62408 139664 62414 139676
rect 66582 139664 66588 139676
rect 66640 139664 66646 139716
rect 135306 139460 135312 139512
rect 135364 139500 135370 139512
rect 138250 139500 138256 139512
rect 135364 139472 138256 139500
rect 135364 139460 135370 139472
rect 138250 139460 138256 139472
rect 138308 139460 138314 139512
rect 62810 139256 62816 139308
rect 62868 139296 62874 139308
rect 65110 139296 65116 139308
rect 62868 139268 65116 139296
rect 62868 139256 62874 139268
rect 65110 139256 65116 139268
rect 65168 139256 65174 139308
rect 62902 138644 62908 138696
rect 62960 138684 62966 138696
rect 66398 138684 66404 138696
rect 62960 138656 66404 138684
rect 62960 138644 62966 138656
rect 66398 138644 66404 138656
rect 66456 138644 66462 138696
rect 135398 138644 135404 138696
rect 135456 138684 135462 138696
rect 136962 138684 136968 138696
rect 135456 138656 136968 138684
rect 135456 138644 135462 138656
rect 136962 138644 136968 138656
rect 137020 138644 137026 138696
rect 62810 138576 62816 138628
rect 62868 138616 62874 138628
rect 66214 138616 66220 138628
rect 62868 138588 66220 138616
rect 62868 138576 62874 138588
rect 66214 138576 66220 138588
rect 66272 138576 66278 138628
rect 135306 138576 135312 138628
rect 135364 138616 135370 138628
rect 136870 138616 136876 138628
rect 135364 138588 136876 138616
rect 135364 138576 135370 138588
rect 136870 138576 136876 138588
rect 136928 138576 136934 138628
rect 98138 138508 98144 138560
rect 98196 138548 98202 138560
rect 102370 138548 102376 138560
rect 98196 138520 102376 138548
rect 98196 138508 98202 138520
rect 102370 138508 102376 138520
rect 102428 138508 102434 138560
rect 169254 138508 169260 138560
rect 169312 138548 169318 138560
rect 174222 138548 174228 138560
rect 169312 138520 174228 138548
rect 169312 138508 169318 138520
rect 174222 138508 174228 138520
rect 174280 138508 174286 138560
rect 97218 138440 97224 138492
rect 97276 138480 97282 138492
rect 102462 138480 102468 138492
rect 97276 138452 102468 138480
rect 97276 138440 97282 138452
rect 102462 138440 102468 138452
rect 102520 138440 102526 138492
rect 169346 138440 169352 138492
rect 169404 138480 169410 138492
rect 174130 138480 174136 138492
rect 169404 138452 174136 138480
rect 169404 138440 169410 138452
rect 174130 138440 174136 138452
rect 174188 138440 174194 138492
rect 135214 137488 135220 137540
rect 135272 137528 135278 137540
rect 136870 137528 136876 137540
rect 135272 137500 136876 137528
rect 135272 137488 135278 137500
rect 136870 137488 136876 137500
rect 136928 137488 136934 137540
rect 100070 137420 100076 137472
rect 100128 137460 100134 137472
rect 102278 137460 102284 137472
rect 100128 137432 102284 137460
rect 100128 137420 100134 137432
rect 102278 137420 102284 137432
rect 102336 137420 102342 137472
rect 132273 137463 132331 137469
rect 132273 137429 132285 137463
rect 132319 137460 132331 137463
rect 132638 137460 132644 137472
rect 132319 137432 132644 137460
rect 132319 137429 132331 137432
rect 132273 137423 132331 137429
rect 132638 137420 132644 137432
rect 132696 137420 132702 137472
rect 62626 137216 62632 137268
rect 62684 137256 62690 137268
rect 66398 137256 66404 137268
rect 62684 137228 66404 137256
rect 62684 137216 62690 137228
rect 66398 137216 66404 137228
rect 66456 137216 66462 137268
rect 99702 137216 99708 137268
rect 99760 137256 99766 137268
rect 102186 137256 102192 137268
rect 99760 137228 102192 137256
rect 99760 137216 99766 137228
rect 102186 137216 102192 137228
rect 102244 137216 102250 137268
rect 135122 137216 135128 137268
rect 135180 137256 135186 137268
rect 136870 137256 136876 137268
rect 135180 137228 136876 137256
rect 135180 137216 135186 137228
rect 136870 137216 136876 137228
rect 136928 137216 136934 137268
rect 172658 137216 172664 137268
rect 172716 137256 172722 137268
rect 174038 137256 174044 137268
rect 172716 137228 174044 137256
rect 172716 137216 172722 137228
rect 174038 137216 174044 137228
rect 174096 137216 174102 137268
rect 62718 137148 62724 137200
rect 62776 137188 62782 137200
rect 66306 137188 66312 137200
rect 62776 137160 66312 137188
rect 62776 137148 62782 137160
rect 66306 137148 66312 137160
rect 66364 137148 66370 137200
rect 101450 137148 101456 137200
rect 101508 137188 101514 137200
rect 101910 137188 101916 137200
rect 101508 137160 101916 137188
rect 101508 137148 101514 137160
rect 101910 137148 101916 137160
rect 101968 137148 101974 137200
rect 132365 137191 132423 137197
rect 132365 137157 132377 137191
rect 132411 137188 132423 137191
rect 132638 137188 132644 137200
rect 132411 137160 132644 137188
rect 132411 137157 132423 137160
rect 132365 137151 132423 137157
rect 132638 137148 132644 137160
rect 132696 137148 132702 137200
rect 172566 137080 172572 137132
rect 172624 137120 172630 137132
rect 174130 137120 174136 137132
rect 172624 137092 174136 137120
rect 172624 137080 172630 137092
rect 174130 137080 174136 137092
rect 174188 137080 174194 137132
rect 100622 137012 100628 137064
rect 100680 137052 100686 137064
rect 102370 137052 102376 137064
rect 100680 137024 102376 137052
rect 100680 137012 100686 137024
rect 102370 137012 102376 137024
rect 102428 137012 102434 137064
rect 172198 137012 172204 137064
rect 172256 137052 172262 137064
rect 174222 137052 174228 137064
rect 172256 137024 174228 137052
rect 172256 137012 172262 137024
rect 174222 137012 174228 137024
rect 174280 137012 174286 137064
rect 132273 136987 132331 136993
rect 132273 136953 132285 136987
rect 132319 136984 132331 136987
rect 132641 136987 132699 136993
rect 132641 136984 132653 136987
rect 132319 136956 132653 136984
rect 132319 136953 132331 136956
rect 132273 136947 132331 136953
rect 132641 136953 132653 136956
rect 132687 136953 132699 136987
rect 132641 136947 132699 136953
rect 100530 136740 100536 136792
rect 100588 136780 100594 136792
rect 102646 136780 102652 136792
rect 100588 136752 102652 136780
rect 100588 136740 100594 136752
rect 102646 136740 102652 136752
rect 102704 136740 102710 136792
rect 172658 135992 172664 136044
rect 172716 136032 172722 136044
rect 173946 136032 173952 136044
rect 172716 136004 173952 136032
rect 172716 135992 172722 136004
rect 173946 135992 173952 136004
rect 174004 135992 174010 136044
rect 62994 135856 63000 135908
rect 63052 135896 63058 135908
rect 65662 135896 65668 135908
rect 63052 135868 65668 135896
rect 63052 135856 63058 135868
rect 65662 135856 65668 135868
rect 65720 135856 65726 135908
rect 100898 135856 100904 135908
rect 100956 135896 100962 135908
rect 102002 135896 102008 135908
rect 100956 135868 102008 135896
rect 100956 135856 100962 135868
rect 102002 135856 102008 135868
rect 102060 135856 102066 135908
rect 134294 135856 134300 135908
rect 134352 135896 134358 135908
rect 136962 135896 136968 135908
rect 134352 135868 136968 135896
rect 134352 135856 134358 135868
rect 136962 135856 136968 135868
rect 137020 135856 137026 135908
rect 172658 135856 172664 135908
rect 172716 135896 172722 135908
rect 173762 135896 173768 135908
rect 172716 135868 173768 135896
rect 172716 135856 172722 135868
rect 173762 135856 173768 135868
rect 173820 135856 173826 135908
rect 62902 135788 62908 135840
rect 62960 135828 62966 135840
rect 66398 135828 66404 135840
rect 62960 135800 66404 135828
rect 62960 135788 62966 135800
rect 66398 135788 66404 135800
rect 66456 135788 66462 135840
rect 100622 135788 100628 135840
rect 100680 135828 100686 135840
rect 100680 135800 101956 135828
rect 100680 135788 100686 135800
rect 101928 135760 101956 135800
rect 135306 135788 135312 135840
rect 135364 135828 135370 135840
rect 136870 135828 136876 135840
rect 135364 135800 136876 135828
rect 135364 135788 135370 135800
rect 136870 135788 136876 135800
rect 136928 135788 136934 135840
rect 172566 135788 172572 135840
rect 172624 135828 172630 135840
rect 172624 135800 172796 135828
rect 172624 135788 172630 135800
rect 102370 135760 102376 135772
rect 101928 135732 102376 135760
rect 102370 135720 102376 135732
rect 102428 135720 102434 135772
rect 172768 135760 172796 135800
rect 174222 135760 174228 135772
rect 172768 135732 174228 135760
rect 174222 135720 174228 135732
rect 174280 135720 174286 135772
rect 62810 135652 62816 135704
rect 62868 135692 62874 135704
rect 65018 135692 65024 135704
rect 62868 135664 65024 135692
rect 62868 135652 62874 135664
rect 65018 135652 65024 135664
rect 65076 135652 65082 135704
rect 172750 135652 172756 135704
rect 172808 135692 172814 135704
rect 174130 135692 174136 135704
rect 172808 135664 174136 135692
rect 172808 135652 172814 135664
rect 174130 135652 174136 135664
rect 174188 135652 174194 135704
rect 135214 135380 135220 135432
rect 135272 135420 135278 135432
rect 136778 135420 136784 135432
rect 135272 135392 136784 135420
rect 135272 135380 135278 135392
rect 136778 135380 136784 135392
rect 136836 135380 136842 135432
rect 99886 134632 99892 134684
rect 99944 134672 99950 134684
rect 102278 134672 102284 134684
rect 99944 134644 102284 134672
rect 99944 134632 99950 134644
rect 102278 134632 102284 134644
rect 102336 134632 102342 134684
rect 100898 134564 100904 134616
rect 100956 134604 100962 134616
rect 102094 134604 102100 134616
rect 100956 134576 102100 134604
rect 100956 134564 100962 134576
rect 102094 134564 102100 134576
rect 102152 134564 102158 134616
rect 62718 134496 62724 134548
rect 62776 134536 62782 134548
rect 66214 134536 66220 134548
rect 62776 134508 66220 134536
rect 62776 134496 62782 134508
rect 66214 134496 66220 134508
rect 66272 134496 66278 134548
rect 135122 134496 135128 134548
rect 135180 134536 135186 134548
rect 136962 134536 136968 134548
rect 135180 134508 136968 134536
rect 135180 134496 135186 134508
rect 136962 134496 136968 134508
rect 137020 134496 137026 134548
rect 172658 134496 172664 134548
rect 172716 134536 172722 134548
rect 174038 134536 174044 134548
rect 172716 134508 174044 134536
rect 172716 134496 172722 134508
rect 174038 134496 174044 134508
rect 174096 134496 174102 134548
rect 62810 134428 62816 134480
rect 62868 134468 62874 134480
rect 65846 134468 65852 134480
rect 62868 134440 65852 134468
rect 62868 134428 62874 134440
rect 65846 134428 65852 134440
rect 65904 134428 65910 134480
rect 135398 134428 135404 134480
rect 135456 134468 135462 134480
rect 136870 134468 136876 134480
rect 135456 134440 136876 134468
rect 135456 134428 135462 134440
rect 136870 134428 136876 134440
rect 136928 134428 136934 134480
rect 172566 134428 172572 134480
rect 172624 134468 172630 134480
rect 173854 134468 173860 134480
rect 172624 134440 173860 134468
rect 172624 134428 172630 134440
rect 173854 134428 173860 134440
rect 173912 134428 173918 134480
rect 100990 134360 100996 134412
rect 101048 134400 101054 134412
rect 102370 134400 102376 134412
rect 101048 134372 102376 134400
rect 101048 134360 101054 134372
rect 102370 134360 102376 134372
rect 102428 134360 102434 134412
rect 204766 134360 204772 134412
rect 204824 134400 204830 134412
rect 204950 134400 204956 134412
rect 204824 134372 204956 134400
rect 204824 134360 204830 134372
rect 204950 134360 204956 134372
rect 205008 134360 205014 134412
rect 100898 133204 100904 133256
rect 100956 133244 100962 133256
rect 102002 133244 102008 133256
rect 100956 133216 102008 133244
rect 100956 133204 100962 133216
rect 102002 133204 102008 133216
rect 102060 133204 102066 133256
rect 100254 133136 100260 133188
rect 100312 133176 100318 133188
rect 102186 133176 102192 133188
rect 100312 133148 102192 133176
rect 100312 133136 100318 133148
rect 102186 133136 102192 133148
rect 102244 133136 102250 133188
rect 63454 133068 63460 133120
rect 63512 133108 63518 133120
rect 65478 133108 65484 133120
rect 63512 133080 65484 133108
rect 63512 133068 63518 133080
rect 65478 133068 65484 133080
rect 65536 133068 65542 133120
rect 135214 133068 135220 133120
rect 135272 133108 135278 133120
rect 136962 133108 136968 133120
rect 135272 133080 136968 133108
rect 135272 133068 135278 133080
rect 136962 133068 136968 133080
rect 137020 133068 137026 133120
rect 171646 133068 171652 133120
rect 171704 133108 171710 133120
rect 173210 133108 173216 133120
rect 171704 133080 173216 133108
rect 171704 133068 171710 133080
rect 173210 133068 173216 133080
rect 173268 133068 173274 133120
rect 63546 133000 63552 133052
rect 63604 133040 63610 133052
rect 66398 133040 66404 133052
rect 63604 133012 66404 133040
rect 63604 133000 63610 133012
rect 66398 133000 66404 133012
rect 66456 133000 66462 133052
rect 135306 133000 135312 133052
rect 135364 133040 135370 133052
rect 136870 133040 136876 133052
rect 135364 133012 136876 133040
rect 135364 133000 135370 133012
rect 136870 133000 136876 133012
rect 136928 133000 136934 133052
rect 63086 131708 63092 131760
rect 63144 131748 63150 131760
rect 65662 131748 65668 131760
rect 63144 131720 65668 131748
rect 63144 131708 63150 131720
rect 65662 131708 65668 131720
rect 65720 131708 65726 131760
rect 100898 131708 100904 131760
rect 100956 131748 100962 131760
rect 102094 131748 102100 131760
rect 100956 131720 102100 131748
rect 100956 131708 100962 131720
rect 102094 131708 102100 131720
rect 102152 131708 102158 131760
rect 135030 131708 135036 131760
rect 135088 131748 135094 131760
rect 136962 131748 136968 131760
rect 135088 131720 136968 131748
rect 135088 131708 135094 131720
rect 136962 131708 136968 131720
rect 137020 131708 137026 131760
rect 172014 131708 172020 131760
rect 172072 131748 172078 131760
rect 172750 131748 172756 131760
rect 172072 131720 172756 131748
rect 172072 131708 172078 131720
rect 172750 131708 172756 131720
rect 172808 131708 172814 131760
rect 63638 131640 63644 131692
rect 63696 131680 63702 131692
rect 66398 131680 66404 131692
rect 63696 131652 66404 131680
rect 63696 131640 63702 131652
rect 66398 131640 66404 131652
rect 66456 131640 66462 131692
rect 100254 131640 100260 131692
rect 100312 131680 100318 131692
rect 102278 131680 102284 131692
rect 100312 131652 102284 131680
rect 100312 131640 100318 131652
rect 102278 131640 102284 131652
rect 102336 131640 102342 131692
rect 135398 131640 135404 131692
rect 135456 131680 135462 131692
rect 136870 131680 136876 131692
rect 135456 131652 136876 131680
rect 135456 131640 135462 131652
rect 136870 131640 136876 131652
rect 136928 131640 136934 131692
rect 171646 131640 171652 131692
rect 171704 131680 171710 131692
rect 173026 131680 173032 131692
rect 171704 131652 173032 131680
rect 171704 131640 171710 131652
rect 173026 131640 173032 131652
rect 173084 131640 173090 131692
rect 173118 131572 173124 131624
rect 173176 131612 173182 131624
rect 174130 131612 174136 131624
rect 173176 131584 174136 131612
rect 173176 131572 173182 131584
rect 174130 131572 174136 131584
rect 174188 131572 174194 131624
rect 172934 131300 172940 131352
rect 172992 131340 172998 131352
rect 175050 131340 175056 131352
rect 172992 131312 175056 131340
rect 172992 131300 172998 131312
rect 175050 131300 175056 131312
rect 175108 131300 175114 131352
rect 172750 131028 172756 131080
rect 172808 131068 172814 131080
rect 174130 131068 174136 131080
rect 172808 131040 174136 131068
rect 172808 131028 172814 131040
rect 174130 131028 174136 131040
rect 174188 131028 174194 131080
rect 62810 130756 62816 130808
rect 62868 130796 62874 130808
rect 65018 130796 65024 130808
rect 62868 130768 65024 130796
rect 62868 130756 62874 130768
rect 65018 130756 65024 130768
rect 65076 130756 65082 130808
rect 134294 130756 134300 130808
rect 134352 130796 134358 130808
rect 136778 130796 136784 130808
rect 134352 130768 136784 130796
rect 134352 130756 134358 130768
rect 136778 130756 136784 130768
rect 136836 130756 136842 130808
rect 172382 130552 172388 130604
rect 172440 130592 172446 130604
rect 174038 130592 174044 130604
rect 172440 130564 174044 130592
rect 172440 130552 172446 130564
rect 174038 130552 174044 130564
rect 174096 130552 174102 130604
rect 100254 130416 100260 130468
rect 100312 130456 100318 130468
rect 102278 130456 102284 130468
rect 100312 130428 102284 130456
rect 100312 130416 100318 130428
rect 102278 130416 102284 130428
rect 102336 130416 102342 130468
rect 62902 130348 62908 130400
rect 62960 130388 62966 130400
rect 66398 130388 66404 130400
rect 62960 130360 66404 130388
rect 62960 130348 62966 130360
rect 66398 130348 66404 130360
rect 66456 130348 66462 130400
rect 100898 130348 100904 130400
rect 100956 130388 100962 130400
rect 102002 130388 102008 130400
rect 100956 130360 102008 130388
rect 100956 130348 100962 130360
rect 102002 130348 102008 130360
rect 102060 130348 102066 130400
rect 135122 130348 135128 130400
rect 135180 130388 135186 130400
rect 136962 130388 136968 130400
rect 135180 130360 136968 130388
rect 135180 130348 135186 130360
rect 136962 130348 136968 130360
rect 137020 130348 137026 130400
rect 62718 130280 62724 130332
rect 62776 130320 62782 130332
rect 66306 130320 66312 130332
rect 62776 130292 66312 130320
rect 62776 130280 62782 130292
rect 66306 130280 66312 130292
rect 66364 130280 66370 130332
rect 135306 130280 135312 130332
rect 135364 130320 135370 130332
rect 136870 130320 136876 130332
rect 135364 130292 136876 130320
rect 135364 130280 135370 130292
rect 136870 130280 136876 130292
rect 136928 130280 136934 130332
rect 100990 130212 100996 130264
rect 101048 130252 101054 130264
rect 102370 130252 102376 130264
rect 101048 130224 102376 130252
rect 101048 130212 101054 130224
rect 102370 130212 102376 130224
rect 102428 130212 102434 130264
rect 173026 130212 173032 130264
rect 173084 130252 173090 130264
rect 174130 130252 174136 130264
rect 173084 130224 174136 130252
rect 173084 130212 173090 130224
rect 174130 130212 174136 130224
rect 174188 130212 174194 130264
rect 172842 130144 172848 130196
rect 172900 130184 172906 130196
rect 174498 130184 174504 130196
rect 172900 130156 174504 130184
rect 172900 130144 172906 130156
rect 174498 130144 174504 130156
rect 174556 130144 174562 130196
rect 172658 129192 172664 129244
rect 172716 129232 172722 129244
rect 173946 129232 173952 129244
rect 172716 129204 173952 129232
rect 172716 129192 172722 129204
rect 173946 129192 173952 129204
rect 174004 129192 174010 129244
rect 62626 128988 62632 129040
rect 62684 129028 62690 129040
rect 66398 129028 66404 129040
rect 62684 129000 66404 129028
rect 62684 128988 62690 129000
rect 66398 128988 66404 129000
rect 66456 128988 66462 129040
rect 100254 128988 100260 129040
rect 100312 129028 100318 129040
rect 102094 129028 102100 129040
rect 100312 129000 102100 129028
rect 100312 128988 100318 129000
rect 102094 128988 102100 129000
rect 102152 128988 102158 129040
rect 134294 128988 134300 129040
rect 134352 129028 134358 129040
rect 136962 129028 136968 129040
rect 134352 129000 136968 129028
rect 134352 128988 134358 129000
rect 136962 128988 136968 129000
rect 137020 128988 137026 129040
rect 62810 128920 62816 128972
rect 62868 128960 62874 128972
rect 65478 128960 65484 128972
rect 62868 128932 65484 128960
rect 62868 128920 62874 128932
rect 65478 128920 65484 128932
rect 65536 128920 65542 128972
rect 100898 128920 100904 128972
rect 100956 128960 100962 128972
rect 102186 128960 102192 128972
rect 100956 128932 102192 128960
rect 100956 128920 100962 128932
rect 102186 128920 102192 128932
rect 102244 128920 102250 128972
rect 135214 128920 135220 128972
rect 135272 128960 135278 128972
rect 136870 128960 136876 128972
rect 135272 128932 136876 128960
rect 135272 128920 135278 128932
rect 136870 128920 136876 128932
rect 136928 128920 136934 128972
rect 172658 128920 172664 128972
rect 172716 128960 172722 128972
rect 173854 128960 173860 128972
rect 172716 128932 173860 128960
rect 172716 128920 172722 128932
rect 173854 128920 173860 128932
rect 173912 128920 173918 128972
rect 172750 128852 172756 128904
rect 172808 128892 172814 128904
rect 174130 128892 174136 128904
rect 172808 128864 174136 128892
rect 172808 128852 172814 128864
rect 174130 128852 174136 128864
rect 174188 128852 174194 128904
rect 100070 127832 100076 127884
rect 100128 127872 100134 127884
rect 102278 127872 102284 127884
rect 100128 127844 102284 127872
rect 100128 127832 100134 127844
rect 102278 127832 102284 127844
rect 102336 127832 102342 127884
rect 100806 127560 100812 127612
rect 100864 127600 100870 127612
rect 102002 127600 102008 127612
rect 100864 127572 102008 127600
rect 100864 127560 100870 127572
rect 102002 127560 102008 127572
rect 102060 127560 102066 127612
rect 132549 127603 132607 127609
rect 132549 127569 132561 127603
rect 132595 127600 132607 127603
rect 132638 127600 132644 127612
rect 132595 127572 132644 127600
rect 132595 127569 132607 127572
rect 132549 127563 132607 127569
rect 132638 127560 132644 127572
rect 132696 127560 132702 127612
rect 135122 127560 135128 127612
rect 135180 127600 135186 127612
rect 136870 127600 136876 127612
rect 135180 127572 136876 127600
rect 135180 127560 135186 127572
rect 136870 127560 136876 127572
rect 136928 127560 136934 127612
rect 62902 127492 62908 127544
rect 62960 127532 62966 127544
rect 66398 127532 66404 127544
rect 62960 127504 66404 127532
rect 62960 127492 62966 127504
rect 66398 127492 66404 127504
rect 66456 127492 66462 127544
rect 171646 127492 171652 127544
rect 171704 127532 171710 127544
rect 222709 127535 222767 127541
rect 171704 127504 172796 127532
rect 171704 127492 171710 127504
rect 172768 127464 172796 127504
rect 222709 127501 222721 127535
rect 222755 127532 222767 127535
rect 222798 127532 222804 127544
rect 222755 127504 222804 127532
rect 222755 127501 222767 127504
rect 222709 127495 222767 127501
rect 222798 127492 222804 127504
rect 222856 127492 222862 127544
rect 174222 127464 174228 127476
rect 172768 127436 174228 127464
rect 174222 127424 174228 127436
rect 174280 127424 174286 127476
rect 132549 127399 132607 127405
rect 132549 127365 132561 127399
rect 132595 127396 132607 127399
rect 132638 127396 132644 127408
rect 132595 127368 132644 127396
rect 132595 127365 132607 127368
rect 132549 127359 132607 127365
rect 132638 127356 132644 127368
rect 132696 127356 132702 127408
rect 132730 127356 132736 127408
rect 132788 127396 132794 127408
rect 132788 127368 132833 127396
rect 132788 127356 132794 127368
rect 134662 127152 134668 127204
rect 134720 127192 134726 127204
rect 136778 127192 136784 127204
rect 134720 127164 136784 127192
rect 134720 127152 134726 127164
rect 136778 127152 136784 127164
rect 136836 127152 136842 127204
rect 62810 126880 62816 126932
rect 62868 126920 62874 126932
rect 65018 126920 65024 126932
rect 62868 126892 65024 126920
rect 62868 126880 62874 126892
rect 65018 126880 65024 126892
rect 65076 126880 65082 126932
rect 172382 126336 172388 126388
rect 172440 126376 172446 126388
rect 174038 126376 174044 126388
rect 172440 126348 174044 126376
rect 172440 126336 172446 126348
rect 174038 126336 174044 126348
rect 174096 126336 174102 126388
rect 62718 126200 62724 126252
rect 62776 126240 62782 126252
rect 66306 126240 66312 126252
rect 62776 126212 66312 126240
rect 62776 126200 62782 126212
rect 66306 126200 66312 126212
rect 66364 126200 66370 126252
rect 100622 126200 100628 126252
rect 100680 126240 100686 126252
rect 102278 126240 102284 126252
rect 100680 126212 102284 126240
rect 100680 126200 100686 126212
rect 102278 126200 102284 126212
rect 102336 126200 102342 126252
rect 135398 126200 135404 126252
rect 135456 126240 135462 126252
rect 136962 126240 136968 126252
rect 135456 126212 136968 126240
rect 135456 126200 135462 126212
rect 136962 126200 136968 126212
rect 137020 126200 137026 126252
rect 172658 126200 172664 126252
rect 172716 126240 172722 126252
rect 173854 126240 173860 126252
rect 172716 126212 173860 126240
rect 172716 126200 172722 126212
rect 173854 126200 173860 126212
rect 173912 126200 173918 126252
rect 62626 126132 62632 126184
rect 62684 126172 62690 126184
rect 66398 126172 66404 126184
rect 62684 126144 66404 126172
rect 62684 126132 62690 126144
rect 66398 126132 66404 126144
rect 66456 126132 66462 126184
rect 100530 126132 100536 126184
rect 100588 126172 100594 126184
rect 100588 126144 101036 126172
rect 100588 126132 100594 126144
rect 101008 126104 101036 126144
rect 135306 126132 135312 126184
rect 135364 126172 135370 126184
rect 136870 126172 136876 126184
rect 135364 126144 136876 126172
rect 135364 126132 135370 126144
rect 136870 126132 136876 126144
rect 136928 126132 136934 126184
rect 172014 126132 172020 126184
rect 172072 126172 172078 126184
rect 172072 126144 173532 126172
rect 172072 126132 172078 126144
rect 102370 126104 102376 126116
rect 101008 126076 102376 126104
rect 102370 126064 102376 126076
rect 102428 126064 102434 126116
rect 134846 126064 134852 126116
rect 134904 126104 134910 126116
rect 136778 126104 136784 126116
rect 134904 126076 136784 126104
rect 134904 126064 134910 126076
rect 136778 126064 136784 126076
rect 136836 126064 136842 126116
rect 173504 126104 173532 126144
rect 174130 126104 174136 126116
rect 173504 126076 174136 126104
rect 174130 126064 174136 126076
rect 174188 126064 174194 126116
rect 172750 125996 172756 126048
rect 172808 126036 172814 126048
rect 174222 126036 174228 126048
rect 172808 126008 174228 126036
rect 172808 125996 172814 126008
rect 174222 125996 174228 126008
rect 174280 125996 174286 126048
rect 62810 125520 62816 125572
rect 62868 125560 62874 125572
rect 65018 125560 65024 125572
rect 62868 125532 65024 125560
rect 62868 125520 62874 125532
rect 65018 125520 65024 125532
rect 65076 125520 65082 125572
rect 100622 125112 100628 125164
rect 100680 125152 100686 125164
rect 102094 125152 102100 125164
rect 100680 125124 102100 125152
rect 100680 125112 100686 125124
rect 102094 125112 102100 125124
rect 102152 125112 102158 125164
rect 100622 124840 100628 124892
rect 100680 124880 100686 124892
rect 102002 124880 102008 124892
rect 100680 124852 102008 124880
rect 100680 124840 100686 124852
rect 102002 124840 102008 124852
rect 102060 124840 102066 124892
rect 172658 124840 172664 124892
rect 172716 124880 172722 124892
rect 173946 124880 173952 124892
rect 172716 124852 173952 124880
rect 172716 124840 172722 124852
rect 173946 124840 173952 124852
rect 174004 124840 174010 124892
rect 62902 124772 62908 124824
rect 62960 124812 62966 124824
rect 65846 124812 65852 124824
rect 62960 124784 65852 124812
rect 62960 124772 62966 124784
rect 65846 124772 65852 124784
rect 65904 124772 65910 124824
rect 135122 124772 135128 124824
rect 135180 124812 135186 124824
rect 136870 124812 136876 124824
rect 135180 124784 136876 124812
rect 135180 124772 135186 124784
rect 136870 124772 136876 124784
rect 136928 124772 136934 124824
rect 172014 124772 172020 124824
rect 172072 124812 172078 124824
rect 222706 124812 222712 124824
rect 172072 124784 172796 124812
rect 222667 124784 222712 124812
rect 172072 124772 172078 124784
rect 100990 124704 100996 124756
rect 101048 124744 101054 124756
rect 102370 124744 102376 124756
rect 101048 124716 102376 124744
rect 101048 124704 101054 124716
rect 102370 124704 102376 124716
rect 102428 124704 102434 124756
rect 172768 124744 172796 124784
rect 222706 124772 222712 124784
rect 222764 124772 222770 124824
rect 174222 124744 174228 124756
rect 172768 124716 174228 124744
rect 174222 124704 174228 124716
rect 174280 124704 174286 124756
rect 135214 124364 135220 124416
rect 135272 124404 135278 124416
rect 136778 124404 136784 124416
rect 135272 124376 136784 124404
rect 135272 124364 135278 124376
rect 136778 124364 136784 124376
rect 136836 124364 136842 124416
rect 62810 124092 62816 124144
rect 62868 124132 62874 124144
rect 65018 124132 65024 124144
rect 62868 124104 65024 124132
rect 62868 124092 62874 124104
rect 65018 124092 65024 124104
rect 65076 124092 65082 124144
rect 100622 123616 100628 123668
rect 100680 123656 100686 123668
rect 102278 123656 102284 123668
rect 100680 123628 102284 123656
rect 100680 123616 100686 123628
rect 102278 123616 102284 123628
rect 102336 123616 102342 123668
rect 63546 123344 63552 123396
rect 63604 123384 63610 123396
rect 66398 123384 66404 123396
rect 63604 123356 66404 123384
rect 63604 123344 63610 123356
rect 66398 123344 66404 123356
rect 66456 123344 66462 123396
rect 99886 123344 99892 123396
rect 99944 123384 99950 123396
rect 102186 123384 102192 123396
rect 99944 123356 102192 123384
rect 99944 123344 99950 123356
rect 102186 123344 102192 123356
rect 102244 123344 102250 123396
rect 135398 123344 135404 123396
rect 135456 123384 135462 123396
rect 136870 123384 136876 123396
rect 135456 123356 136876 123384
rect 135456 123344 135462 123356
rect 136870 123344 136876 123356
rect 136928 123344 136934 123396
rect 172382 123344 172388 123396
rect 172440 123384 172446 123396
rect 174038 123384 174044 123396
rect 172440 123356 174044 123384
rect 172440 123344 172446 123356
rect 174038 123344 174044 123356
rect 174096 123344 174102 123396
rect 135306 122868 135312 122920
rect 135364 122908 135370 122920
rect 136778 122908 136784 122920
rect 135364 122880 136784 122908
rect 135364 122868 135370 122880
rect 136778 122868 136784 122880
rect 136836 122868 136842 122920
rect 62810 122596 62816 122648
rect 62868 122636 62874 122648
rect 65018 122636 65024 122648
rect 62868 122608 65024 122636
rect 62868 122596 62874 122608
rect 65018 122596 65024 122608
rect 65076 122596 65082 122648
rect 100162 122188 100168 122240
rect 100220 122228 100226 122240
rect 102278 122228 102284 122240
rect 100220 122200 102284 122228
rect 100220 122188 100226 122200
rect 102278 122188 102284 122200
rect 102336 122188 102342 122240
rect 135122 122120 135128 122172
rect 135180 122160 135186 122172
rect 137054 122160 137060 122172
rect 135180 122132 137060 122160
rect 135180 122120 135186 122132
rect 137054 122120 137060 122132
rect 137112 122120 137118 122172
rect 63454 122052 63460 122104
rect 63512 122092 63518 122104
rect 66306 122092 66312 122104
rect 63512 122064 66312 122092
rect 63512 122052 63518 122064
rect 66306 122052 66312 122064
rect 66364 122052 66370 122104
rect 100898 122052 100904 122104
rect 100956 122092 100962 122104
rect 102094 122092 102100 122104
rect 100956 122064 102100 122092
rect 100956 122052 100962 122064
rect 102094 122052 102100 122064
rect 102152 122052 102158 122104
rect 135214 122052 135220 122104
rect 135272 122092 135278 122104
rect 136962 122092 136968 122104
rect 135272 122064 136968 122092
rect 135272 122052 135278 122064
rect 136962 122052 136968 122064
rect 137020 122052 137026 122104
rect 63638 121984 63644 122036
rect 63696 122024 63702 122036
rect 66398 122024 66404 122036
rect 63696 121996 66404 122024
rect 63696 121984 63702 121996
rect 66398 121984 66404 121996
rect 66456 121984 66462 122036
rect 136870 122024 136876 122036
rect 135508 121996 136876 122024
rect 135306 121916 135312 121968
rect 135364 121956 135370 121968
rect 135508 121956 135536 121996
rect 136870 121984 136876 121996
rect 136928 121984 136934 122036
rect 171554 121984 171560 122036
rect 171612 122024 171618 122036
rect 171612 121996 172796 122024
rect 171612 121984 171618 121996
rect 135364 121928 135536 121956
rect 172768 121956 172796 121996
rect 174130 121956 174136 121968
rect 172768 121928 174136 121956
rect 135364 121916 135370 121928
rect 174130 121916 174136 121928
rect 174188 121916 174194 121968
rect 172842 121780 172848 121832
rect 172900 121820 172906 121832
rect 174314 121820 174320 121832
rect 172900 121792 174320 121820
rect 172900 121780 172906 121792
rect 174314 121780 174320 121792
rect 174372 121780 174378 121832
rect 62810 121440 62816 121492
rect 62868 121480 62874 121492
rect 65018 121480 65024 121492
rect 62868 121452 65024 121480
rect 62868 121440 62874 121452
rect 65018 121440 65024 121452
rect 65076 121440 65082 121492
rect 100622 120896 100628 120948
rect 100680 120936 100686 120948
rect 102278 120936 102284 120948
rect 100680 120908 102284 120936
rect 100680 120896 100686 120908
rect 102278 120896 102284 120908
rect 102336 120896 102342 120948
rect 171738 120896 171744 120948
rect 171796 120936 171802 120948
rect 174038 120936 174044 120948
rect 171796 120908 174044 120936
rect 171796 120896 171802 120908
rect 174038 120896 174044 120908
rect 174096 120896 174102 120948
rect 100622 120624 100628 120676
rect 100680 120664 100686 120676
rect 102186 120664 102192 120676
rect 100680 120636 102192 120664
rect 100680 120624 100686 120636
rect 102186 120624 102192 120636
rect 102244 120624 102250 120676
rect 172658 120624 172664 120676
rect 172716 120664 172722 120676
rect 173946 120664 173952 120676
rect 172716 120636 173952 120664
rect 172716 120624 172722 120636
rect 173946 120624 173952 120636
rect 174004 120624 174010 120676
rect 100990 120556 100996 120608
rect 101048 120596 101054 120608
rect 102370 120596 102376 120608
rect 101048 120568 102376 120596
rect 101048 120556 101054 120568
rect 102370 120556 102376 120568
rect 102428 120556 102434 120608
rect 172934 120556 172940 120608
rect 172992 120596 172998 120608
rect 174130 120596 174136 120608
rect 172992 120568 174136 120596
rect 172992 120556 172998 120568
rect 174130 120556 174136 120568
rect 174188 120556 174194 120608
rect 172750 120488 172756 120540
rect 172808 120528 172814 120540
rect 174314 120528 174320 120540
rect 172808 120500 174320 120528
rect 172808 120488 172814 120500
rect 174314 120488 174320 120500
rect 174372 120488 174378 120540
rect 134846 120216 134852 120268
rect 134904 120256 134910 120268
rect 136778 120256 136784 120268
rect 134904 120228 136784 120256
rect 134904 120216 134910 120228
rect 136778 120216 136784 120228
rect 136836 120216 136842 120268
rect 62810 119944 62816 119996
rect 62868 119984 62874 119996
rect 65018 119984 65024 119996
rect 62868 119956 65024 119984
rect 62868 119944 62874 119956
rect 65018 119944 65024 119956
rect 65076 119944 65082 119996
rect 172658 119536 172664 119588
rect 172716 119576 172722 119588
rect 174038 119576 174044 119588
rect 172716 119548 174044 119576
rect 172716 119536 172722 119548
rect 174038 119536 174044 119548
rect 174096 119536 174102 119588
rect 100622 119400 100628 119452
rect 100680 119440 100686 119452
rect 102278 119440 102284 119452
rect 100680 119412 102284 119440
rect 100680 119400 100686 119412
rect 102278 119400 102284 119412
rect 102336 119400 102342 119452
rect 62902 119264 62908 119316
rect 62960 119304 62966 119316
rect 66398 119304 66404 119316
rect 62960 119276 66404 119304
rect 62960 119264 62966 119276
rect 66398 119264 66404 119276
rect 66456 119264 66462 119316
rect 135214 119264 135220 119316
rect 135272 119304 135278 119316
rect 136962 119304 136968 119316
rect 135272 119276 136968 119304
rect 135272 119264 135278 119276
rect 136962 119264 136968 119276
rect 137020 119264 137026 119316
rect 62718 119128 62724 119180
rect 62776 119168 62782 119180
rect 66214 119168 66220 119180
rect 62776 119140 66220 119168
rect 62776 119128 62782 119140
rect 66214 119128 66220 119140
rect 66272 119128 66278 119180
rect 135306 119060 135312 119112
rect 135364 119100 135370 119112
rect 136870 119100 136876 119112
rect 135364 119072 136876 119100
rect 135364 119060 135370 119072
rect 136870 119060 136876 119072
rect 136928 119060 136934 119112
rect 62810 118720 62816 118772
rect 62868 118760 62874 118772
rect 65018 118760 65024 118772
rect 62868 118732 65024 118760
rect 62868 118720 62874 118732
rect 65018 118720 65024 118732
rect 65076 118720 65082 118772
rect 135030 118652 135036 118704
rect 135088 118692 135094 118704
rect 136778 118692 136784 118704
rect 135088 118664 136784 118692
rect 135088 118652 135094 118664
rect 136778 118652 136784 118664
rect 136836 118652 136842 118704
rect 100622 118312 100628 118364
rect 100680 118352 100686 118364
rect 102186 118352 102192 118364
rect 100680 118324 102192 118352
rect 100680 118312 100686 118324
rect 102186 118312 102192 118324
rect 102244 118312 102250 118364
rect 132549 118287 132607 118293
rect 132549 118253 132561 118287
rect 132595 118284 132607 118287
rect 132638 118284 132644 118296
rect 132595 118256 132644 118284
rect 132595 118253 132607 118256
rect 132549 118247 132607 118253
rect 132638 118244 132644 118256
rect 132696 118244 132702 118296
rect 132641 118151 132699 118157
rect 132641 118117 132653 118151
rect 132687 118148 132699 118151
rect 132730 118148 132736 118160
rect 132687 118120 132736 118148
rect 132687 118117 132699 118120
rect 132641 118111 132699 118117
rect 132730 118108 132736 118120
rect 132788 118108 132794 118160
rect 172658 118040 172664 118092
rect 172716 118080 172722 118092
rect 173946 118080 173952 118092
rect 172716 118052 173952 118080
rect 172716 118040 172722 118052
rect 173946 118040 173952 118052
rect 174004 118040 174010 118092
rect 100622 117904 100628 117956
rect 100680 117944 100686 117956
rect 102278 117944 102284 117956
rect 100680 117916 102284 117944
rect 100680 117904 100686 117916
rect 102278 117904 102284 117916
rect 102336 117904 102342 117956
rect 132730 117904 132736 117956
rect 132788 117944 132794 117956
rect 132788 117916 132833 117944
rect 132788 117904 132794 117916
rect 135306 117904 135312 117956
rect 135364 117944 135370 117956
rect 136870 117944 136876 117956
rect 135364 117916 136876 117944
rect 135364 117904 135370 117916
rect 136870 117904 136876 117916
rect 136928 117904 136934 117956
rect 62718 117836 62724 117888
rect 62776 117876 62782 117888
rect 66398 117876 66404 117888
rect 62776 117848 66404 117876
rect 62776 117836 62782 117848
rect 66398 117836 66404 117848
rect 66456 117836 66462 117888
rect 136962 117876 136968 117888
rect 135508 117848 136968 117876
rect 100990 117768 100996 117820
rect 101048 117808 101054 117820
rect 102370 117808 102376 117820
rect 101048 117780 102376 117808
rect 101048 117768 101054 117780
rect 102370 117768 102376 117780
rect 102428 117768 102434 117820
rect 134110 117768 134116 117820
rect 134168 117808 134174 117820
rect 135508 117808 135536 117848
rect 136962 117836 136968 117848
rect 137020 117836 137026 117888
rect 172014 117836 172020 117888
rect 172072 117876 172078 117888
rect 174038 117876 174044 117888
rect 172072 117848 174044 117876
rect 172072 117836 172078 117848
rect 174038 117836 174044 117848
rect 174096 117836 174102 117888
rect 134168 117780 135536 117808
rect 134168 117768 134174 117780
rect 172750 117768 172756 117820
rect 172808 117808 172814 117820
rect 174130 117808 174136 117820
rect 172808 117780 174136 117808
rect 172808 117768 172814 117780
rect 174130 117768 174136 117780
rect 174188 117768 174194 117820
rect 132638 117740 132644 117752
rect 132599 117712 132644 117740
rect 132638 117700 132644 117712
rect 132696 117700 132702 117752
rect 62810 117292 62816 117344
rect 62868 117332 62874 117344
rect 65018 117332 65024 117344
rect 62868 117304 65024 117332
rect 62868 117292 62874 117304
rect 65018 117292 65024 117304
rect 65076 117292 65082 117344
rect 62810 117156 62816 117208
rect 62868 117196 62874 117208
rect 64926 117196 64932 117208
rect 62868 117168 64932 117196
rect 62868 117156 62874 117168
rect 64926 117156 64932 117168
rect 64984 117156 64990 117208
rect 134662 117156 134668 117208
rect 134720 117196 134726 117208
rect 136778 117196 136784 117208
rect 134720 117168 136784 117196
rect 134720 117156 134726 117168
rect 136778 117156 136784 117168
rect 136836 117156 136842 117208
rect 100622 116612 100628 116664
rect 100680 116652 100686 116664
rect 102186 116652 102192 116664
rect 100680 116624 102192 116652
rect 100680 116612 100686 116624
rect 102186 116612 102192 116624
rect 102244 116612 102250 116664
rect 172566 116544 172572 116596
rect 172624 116584 172630 116596
rect 173854 116584 173860 116596
rect 172624 116556 173860 116584
rect 172624 116544 172630 116556
rect 173854 116544 173860 116556
rect 173912 116544 173918 116596
rect 100530 116476 100536 116528
rect 100588 116516 100594 116528
rect 100588 116488 101036 116516
rect 100588 116476 100594 116488
rect 101008 116448 101036 116488
rect 172658 116476 172664 116528
rect 172716 116516 172722 116528
rect 172716 116488 172796 116516
rect 172716 116476 172722 116488
rect 102370 116448 102376 116460
rect 101008 116420 102376 116448
rect 102370 116408 102376 116420
rect 102428 116408 102434 116460
rect 172768 116448 172796 116488
rect 174222 116448 174228 116460
rect 172768 116420 174228 116448
rect 174222 116408 174228 116420
rect 174280 116408 174286 116460
rect 100714 116340 100720 116392
rect 100772 116380 100778 116392
rect 102462 116380 102468 116392
rect 100772 116352 102468 116380
rect 100772 116340 100778 116352
rect 102462 116340 102468 116352
rect 102520 116340 102526 116392
rect 172474 116340 172480 116392
rect 172532 116380 172538 116392
rect 174130 116380 174136 116392
rect 172532 116352 174136 116380
rect 172532 116340 172538 116352
rect 174130 116340 174136 116352
rect 174188 116340 174194 116392
rect 62810 115728 62816 115780
rect 62868 115768 62874 115780
rect 65018 115768 65024 115780
rect 62868 115740 65024 115768
rect 62868 115728 62874 115740
rect 65018 115728 65024 115740
rect 65076 115728 65082 115780
rect 134478 115728 134484 115780
rect 134536 115768 134542 115780
rect 136778 115768 136784 115780
rect 134536 115740 136784 115768
rect 134536 115728 134542 115740
rect 136778 115728 136784 115740
rect 136836 115728 136842 115780
rect 172658 115592 172664 115644
rect 172716 115632 172722 115644
rect 174038 115632 174044 115644
rect 172716 115604 174044 115632
rect 172716 115592 172722 115604
rect 174038 115592 174044 115604
rect 174096 115592 174102 115644
rect 100622 115184 100628 115236
rect 100680 115224 100686 115236
rect 102278 115224 102284 115236
rect 100680 115196 102284 115224
rect 100680 115184 100686 115196
rect 102278 115184 102284 115196
rect 102336 115184 102342 115236
rect 144874 115116 144880 115168
rect 144932 115156 144938 115168
rect 204766 115156 204772 115168
rect 144932 115128 204772 115156
rect 144932 115116 144938 115128
rect 204766 115116 204772 115128
rect 204824 115116 204830 115168
rect 132638 115048 132644 115100
rect 132696 115088 132702 115100
rect 132733 115091 132791 115097
rect 132733 115088 132745 115091
rect 132696 115060 132745 115088
rect 132696 115048 132702 115060
rect 132733 115057 132745 115060
rect 132779 115057 132791 115091
rect 132733 115051 132791 115057
rect 222614 115048 222620 115100
rect 222672 115088 222678 115100
rect 222982 115088 222988 115100
rect 222672 115060 222988 115088
rect 222672 115048 222678 115060
rect 222982 115048 222988 115060
rect 223040 115048 223046 115100
rect 135306 114980 135312 115032
rect 135364 115020 135370 115032
rect 136870 115020 136876 115032
rect 135364 114992 136876 115020
rect 135364 114980 135370 114992
rect 136870 114980 136876 114992
rect 136928 114980 136934 115032
rect 132549 114955 132607 114961
rect 132549 114921 132561 114955
rect 132595 114952 132607 114955
rect 144874 114952 144880 114964
rect 132595 114924 144880 114952
rect 132595 114921 132607 114924
rect 132549 114915 132607 114921
rect 144874 114912 144880 114924
rect 144932 114912 144938 114964
rect 62810 114844 62816 114896
rect 62868 114884 62874 114896
rect 66398 114884 66404 114896
rect 62868 114856 66404 114884
rect 62868 114844 62874 114856
rect 66398 114844 66404 114856
rect 66456 114844 66462 114896
rect 62810 114572 62816 114624
rect 62868 114612 62874 114624
rect 65018 114612 65024 114624
rect 62868 114584 65024 114612
rect 62868 114572 62874 114584
rect 65018 114572 65024 114584
rect 65076 114572 65082 114624
rect 134846 114436 134852 114488
rect 134904 114476 134910 114488
rect 136778 114476 136784 114488
rect 134904 114448 136784 114476
rect 134904 114436 134910 114448
rect 136778 114436 136784 114448
rect 136836 114436 136842 114488
rect 30426 114300 30432 114352
rect 30484 114340 30490 114352
rect 92710 114340 92716 114352
rect 30484 114312 92716 114340
rect 30484 114300 30490 114312
rect 92710 114300 92716 114312
rect 92768 114300 92774 114352
rect 132086 113756 132092 113808
rect 132144 113796 132150 113808
rect 132641 113799 132699 113805
rect 132641 113796 132653 113799
rect 132144 113768 132653 113796
rect 132144 113756 132150 113768
rect 132641 113765 132653 113768
rect 132687 113765 132699 113799
rect 132641 113759 132699 113765
rect 132454 113688 132460 113740
rect 132512 113728 132518 113740
rect 132549 113731 132607 113737
rect 132549 113728 132561 113731
rect 132512 113700 132561 113728
rect 132512 113688 132518 113700
rect 132549 113697 132561 113700
rect 132595 113697 132607 113731
rect 132549 113691 132607 113697
rect 73206 113620 73212 113672
rect 73264 113660 73270 113672
rect 109454 113660 109460 113672
rect 73264 113632 109460 113660
rect 73264 113620 73270 113632
rect 109454 113620 109460 113632
rect 109512 113620 109518 113672
rect 113502 113620 113508 113672
rect 113560 113660 113566 113672
rect 114376 113660 114382 113672
rect 113560 113632 114382 113660
rect 113560 113620 113566 113632
rect 114376 113620 114382 113632
rect 114434 113620 114440 113672
rect 114514 113620 114520 113672
rect 114572 113660 114578 113672
rect 115480 113660 115486 113672
rect 114572 113632 115486 113660
rect 114572 113620 114578 113632
rect 115480 113620 115486 113632
rect 115538 113620 115544 113672
rect 116630 113620 116636 113672
rect 116688 113660 116694 113672
rect 118792 113660 118798 113672
rect 116688 113632 118798 113660
rect 116688 113620 116694 113632
rect 118792 113620 118798 113632
rect 118850 113620 118856 113672
rect 120126 113620 120132 113672
rect 120184 113660 120190 113672
rect 123116 113660 123122 113672
rect 120184 113632 123122 113660
rect 120184 113620 120190 113632
rect 123116 113620 123122 113632
rect 123174 113620 123180 113672
rect 126290 113620 126296 113672
rect 126348 113660 126354 113672
rect 131948 113660 131954 113672
rect 126348 113632 131954 113660
rect 126348 113620 126354 113632
rect 131948 113620 131954 113632
rect 132006 113620 132012 113672
rect 154810 113620 154816 113672
rect 154868 113660 154874 113672
rect 205042 113660 205048 113672
rect 154868 113632 205048 113660
rect 154868 113620 154874 113632
rect 205042 113620 205048 113632
rect 205100 113620 205106 113672
rect 122702 113552 122708 113604
rect 122760 113592 122766 113604
rect 127026 113592 127032 113604
rect 122760 113564 127032 113592
rect 122760 113552 122766 113564
rect 127026 113552 127032 113564
rect 127084 113552 127090 113604
rect 123070 113416 123076 113468
rect 123128 113456 123134 113468
rect 127486 113456 127492 113468
rect 123128 113428 127492 113456
rect 123128 113416 123134 113428
rect 127486 113416 127492 113428
rect 127544 113416 127550 113468
rect 123898 113348 123904 113400
rect 123956 113388 123962 113400
rect 128590 113388 128596 113400
rect 123956 113360 128596 113388
rect 123956 113348 123962 113360
rect 128590 113348 128596 113360
rect 128648 113348 128654 113400
rect 124634 113280 124640 113332
rect 124692 113320 124698 113332
rect 129694 113320 129700 113332
rect 124692 113292 129700 113320
rect 124692 113280 124698 113292
rect 129694 113280 129700 113292
rect 129752 113280 129758 113332
rect 122242 113212 122248 113264
rect 122300 113252 122306 113264
rect 126382 113252 126388 113264
rect 122300 113224 126388 113252
rect 122300 113212 122306 113224
rect 126382 113212 126388 113224
rect 126440 113212 126446 113264
rect 81670 113144 81676 113196
rect 81728 113184 81734 113196
rect 82498 113184 82504 113196
rect 81728 113156 82504 113184
rect 81728 113144 81734 113156
rect 82498 113144 82504 113156
rect 82556 113144 82562 113196
rect 116262 113144 116268 113196
rect 116320 113184 116326 113196
rect 118194 113184 118200 113196
rect 116320 113156 118200 113184
rect 116320 113144 116326 113156
rect 118194 113144 118200 113156
rect 118252 113144 118258 113196
rect 125462 113144 125468 113196
rect 125520 113184 125526 113196
rect 130798 113184 130804 113196
rect 125520 113156 130804 113184
rect 125520 113144 125526 113156
rect 130798 113144 130804 113156
rect 130856 113144 130862 113196
rect 188942 113144 188948 113196
rect 189000 113184 189006 113196
rect 189678 113184 189684 113196
rect 189000 113156 189684 113184
rect 189000 113144 189006 113156
rect 189678 113144 189684 113156
rect 189736 113144 189742 113196
rect 113870 113076 113876 113128
rect 113928 113116 113934 113128
rect 114882 113116 114888 113128
rect 113928 113088 114888 113116
rect 113928 113076 113934 113088
rect 114882 113076 114888 113088
rect 114940 113076 114946 113128
rect 115066 113076 115072 113128
rect 115124 113116 115130 113128
rect 116538 113116 116544 113128
rect 115124 113088 116544 113116
rect 115124 113076 115130 113088
rect 116538 113076 116544 113088
rect 116596 113076 116602 113128
rect 121874 113076 121880 113128
rect 121932 113116 121938 113128
rect 125830 113116 125836 113128
rect 121932 113088 125836 113116
rect 121932 113076 121938 113088
rect 125830 113076 125836 113088
rect 125888 113076 125894 113128
rect 183974 113076 183980 113128
rect 184032 113116 184038 113128
rect 184434 113116 184440 113128
rect 184032 113088 184440 113116
rect 184032 113076 184038 113088
rect 184434 113076 184440 113088
rect 184492 113076 184498 113128
rect 188482 113076 188488 113128
rect 188540 113116 188546 113128
rect 189126 113116 189132 113128
rect 188540 113088 189132 113116
rect 188540 113076 188546 113088
rect 189126 113076 189132 113088
rect 189184 113076 189190 113128
rect 195750 113076 195756 113128
rect 195808 113116 195814 113128
rect 199338 113116 199344 113128
rect 195808 113088 199344 113116
rect 195808 113076 195814 113088
rect 199338 113076 199344 113088
rect 199396 113076 199402 113128
rect 115434 113008 115440 113060
rect 115492 113048 115498 113060
rect 117090 113048 117096 113060
rect 115492 113020 117096 113048
rect 115492 113008 115498 113020
rect 117090 113008 117096 113020
rect 117148 113008 117154 113060
rect 125094 113008 125100 113060
rect 125152 113048 125158 113060
rect 130246 113048 130252 113060
rect 125152 113020 130252 113048
rect 125152 113008 125158 113020
rect 130246 113008 130252 113020
rect 130304 113008 130310 113060
rect 193726 113008 193732 113060
rect 193784 113048 193790 113060
rect 196486 113048 196492 113060
rect 193784 113020 196492 113048
rect 193784 113008 193790 113020
rect 196486 113008 196492 113020
rect 196544 113008 196550 113060
rect 125830 112940 125836 112992
rect 125888 112980 125894 112992
rect 131350 112980 131356 112992
rect 125888 112952 131356 112980
rect 125888 112940 125894 112952
rect 131350 112940 131356 112952
rect 131408 112940 131414 112992
rect 196118 112940 196124 112992
rect 196176 112980 196182 112992
rect 199982 112980 199988 112992
rect 196176 112952 199988 112980
rect 196176 112940 196182 112952
rect 199982 112940 199988 112952
rect 200040 112940 200046 112992
rect 114698 112872 114704 112924
rect 114756 112912 114762 112924
rect 115986 112912 115992 112924
rect 114756 112884 115992 112912
rect 114756 112872 114762 112884
rect 115986 112872 115992 112884
rect 116044 112872 116050 112924
rect 124266 112872 124272 112924
rect 124324 112912 124330 112924
rect 129142 112912 129148 112924
rect 124324 112884 129148 112912
rect 124324 112872 124330 112884
rect 129142 112872 129148 112884
rect 129200 112872 129206 112924
rect 191334 112872 191340 112924
rect 191392 112912 191398 112924
rect 193082 112912 193088 112924
rect 191392 112884 193088 112912
rect 191392 112872 191398 112884
rect 193082 112872 193088 112884
rect 193140 112872 193146 112924
rect 123438 112804 123444 112856
rect 123496 112844 123502 112856
rect 128038 112844 128044 112856
rect 123496 112816 128044 112844
rect 123496 112804 123502 112816
rect 128038 112804 128044 112816
rect 128096 112804 128102 112856
rect 117826 112736 117832 112788
rect 117884 112776 117890 112788
rect 120218 112776 120224 112788
rect 117884 112748 120224 112776
rect 117884 112736 117890 112748
rect 120218 112736 120224 112748
rect 120276 112736 120282 112788
rect 126658 112736 126664 112788
rect 126716 112776 126722 112788
rect 132546 112776 132552 112788
rect 126716 112748 132552 112776
rect 126716 112736 126722 112748
rect 132546 112736 132552 112748
rect 132604 112736 132610 112788
rect 188022 112736 188028 112788
rect 188080 112776 188086 112788
rect 188574 112776 188580 112788
rect 188080 112748 188580 112776
rect 188080 112736 188086 112748
rect 188574 112736 188580 112748
rect 188632 112736 188638 112788
rect 192898 112736 192904 112788
rect 192956 112776 192962 112788
rect 195382 112776 195388 112788
rect 192956 112748 195388 112776
rect 192956 112736 192962 112748
rect 195382 112736 195388 112748
rect 195440 112736 195446 112788
rect 196486 112736 196492 112788
rect 196544 112776 196550 112788
rect 200534 112776 200540 112788
rect 196544 112748 200540 112776
rect 196544 112736 196550 112748
rect 200534 112736 200540 112748
rect 200592 112736 200598 112788
rect 197314 112668 197320 112720
rect 197372 112708 197378 112720
rect 201638 112708 201644 112720
rect 197372 112680 201644 112708
rect 197372 112668 197378 112680
rect 201638 112668 201644 112680
rect 201696 112668 201702 112720
rect 189218 112600 189224 112652
rect 189276 112640 189282 112652
rect 190230 112640 190236 112652
rect 189276 112612 190236 112640
rect 189276 112600 189282 112612
rect 190230 112600 190236 112612
rect 190288 112600 190294 112652
rect 192530 112600 192536 112652
rect 192588 112640 192594 112652
rect 194738 112640 194744 112652
rect 192588 112612 194744 112640
rect 192588 112600 192594 112612
rect 194738 112600 194744 112612
rect 194796 112600 194802 112652
rect 196946 112600 196952 112652
rect 197004 112640 197010 112652
rect 201086 112640 201092 112652
rect 197004 112612 201092 112640
rect 197004 112600 197010 112612
rect 201086 112600 201092 112612
rect 201144 112600 201150 112652
rect 121506 112532 121512 112584
rect 121564 112572 121570 112584
rect 125278 112572 125284 112584
rect 121564 112544 125284 112572
rect 121564 112532 121570 112544
rect 125278 112532 125284 112544
rect 125336 112532 125342 112584
rect 197406 112532 197412 112584
rect 197464 112572 197470 112584
rect 202190 112572 202196 112584
rect 197464 112544 202196 112572
rect 197464 112532 197470 112544
rect 202190 112532 202196 112544
rect 202248 112532 202254 112584
rect 121046 112464 121052 112516
rect 121104 112504 121110 112516
rect 124726 112504 124732 112516
rect 121104 112476 124732 112504
rect 121104 112464 121110 112476
rect 124726 112464 124732 112476
rect 124784 112464 124790 112516
rect 189586 112464 189592 112516
rect 189644 112504 189650 112516
rect 190782 112504 190788 112516
rect 189644 112476 190788 112504
rect 189644 112464 189650 112476
rect 190782 112464 190788 112476
rect 190840 112464 190846 112516
rect 198142 112464 198148 112516
rect 198200 112504 198206 112516
rect 202834 112504 202840 112516
rect 198200 112476 202840 112504
rect 198200 112464 198206 112476
rect 202834 112464 202840 112476
rect 202892 112464 202898 112516
rect 120310 112396 120316 112448
rect 120368 112436 120374 112448
rect 120368 112408 122104 112436
rect 120368 112396 120374 112408
rect 113042 112328 113048 112380
rect 113100 112368 113106 112380
rect 113778 112368 113784 112380
rect 113100 112340 113784 112368
rect 113100 112328 113106 112340
rect 113778 112328 113784 112340
rect 113836 112328 113842 112380
rect 119114 112328 119120 112380
rect 119172 112368 119178 112380
rect 119172 112340 121552 112368
rect 119172 112328 119178 112340
rect 81670 112260 81676 112312
rect 81728 112300 81734 112312
rect 110466 112300 110472 112312
rect 81728 112272 110472 112300
rect 81728 112260 81734 112272
rect 110466 112260 110472 112272
rect 110524 112260 110530 112312
rect 121524 112300 121552 112340
rect 121966 112300 121972 112312
rect 121524 112272 121972 112300
rect 121966 112260 121972 112272
rect 122024 112260 122030 112312
rect 122076 112300 122104 112408
rect 190506 112396 190512 112448
rect 190564 112436 190570 112448
rect 191978 112436 191984 112448
rect 190564 112408 191984 112436
rect 190564 112396 190570 112408
rect 191978 112396 191984 112408
rect 192036 112396 192042 112448
rect 194554 112396 194560 112448
rect 194612 112436 194618 112448
rect 197682 112436 197688 112448
rect 194612 112408 197688 112436
rect 194612 112396 194618 112408
rect 197682 112396 197688 112408
rect 197740 112396 197746 112448
rect 198878 112396 198884 112448
rect 198936 112436 198942 112448
rect 198936 112408 201868 112436
rect 198936 112396 198942 112408
rect 190138 112328 190144 112380
rect 190196 112368 190202 112380
rect 191426 112368 191432 112380
rect 190196 112340 191432 112368
rect 190196 112328 190202 112340
rect 191426 112328 191432 112340
rect 191484 112328 191490 112380
rect 191702 112328 191708 112380
rect 191760 112368 191766 112380
rect 191760 112340 192116 112368
rect 191760 112328 191766 112340
rect 123622 112300 123628 112312
rect 122076 112272 123628 112300
rect 123622 112260 123628 112272
rect 123680 112260 123686 112312
rect 192088 112300 192116 112340
rect 193174 112328 193180 112380
rect 193232 112368 193238 112380
rect 193232 112340 194692 112368
rect 193232 112328 193238 112340
rect 193634 112300 193640 112312
rect 192088 112272 193640 112300
rect 193634 112260 193640 112272
rect 193692 112260 193698 112312
rect 194664 112300 194692 112340
rect 194738 112328 194744 112380
rect 194796 112368 194802 112380
rect 198234 112368 198240 112380
rect 194796 112340 198240 112368
rect 194796 112328 194802 112340
rect 198234 112328 198240 112340
rect 198292 112328 198298 112380
rect 198510 112328 198516 112380
rect 198568 112368 198574 112380
rect 201840 112368 201868 112408
rect 198568 112340 201776 112368
rect 201840 112340 203524 112368
rect 198568 112328 198574 112340
rect 195934 112300 195940 112312
rect 194664 112272 195940 112300
rect 195934 112260 195940 112272
rect 195992 112260 195998 112312
rect 201748 112300 201776 112340
rect 203386 112300 203392 112312
rect 201748 112272 203392 112300
rect 203386 112260 203392 112272
rect 203444 112260 203450 112312
rect 203496 112300 203524 112340
rect 203938 112300 203944 112312
rect 203496 112272 203944 112300
rect 203938 112260 203944 112272
rect 203996 112260 204002 112312
rect 109454 112192 109460 112244
rect 109512 112232 109518 112244
rect 132454 112232 132460 112244
rect 109512 112204 132460 112232
rect 109512 112192 109518 112204
rect 132454 112192 132460 112204
rect 132512 112192 132518 112244
rect 34474 112124 34480 112176
rect 34532 112164 34538 112176
rect 39442 112164 39448 112176
rect 34532 112136 39448 112164
rect 34532 112124 34538 112136
rect 39442 112124 39448 112136
rect 39500 112124 39506 112176
rect 52598 112124 52604 112176
rect 52656 112164 52662 112176
rect 57014 112164 57020 112176
rect 52656 112136 57020 112164
rect 52656 112124 52662 112136
rect 57014 112124 57020 112136
rect 57072 112124 57078 112176
rect 110006 112124 110012 112176
rect 110064 112164 110070 112176
rect 164470 112164 164476 112176
rect 110064 112136 164476 112164
rect 110064 112124 110070 112136
rect 164470 112124 164476 112136
rect 164528 112124 164534 112176
rect 51034 112056 51040 112108
rect 51092 112096 51098 112108
rect 54254 112096 54260 112108
rect 51092 112068 54260 112096
rect 51092 112056 51098 112068
rect 54254 112056 54260 112068
rect 54312 112056 54318 112108
rect 116170 112056 116176 112108
rect 116228 112096 116234 112108
rect 117642 112096 117648 112108
rect 116228 112068 117648 112096
rect 116228 112056 116234 112068
rect 117642 112056 117648 112068
rect 117700 112056 117706 112108
rect 120954 112056 120960 112108
rect 121012 112096 121018 112108
rect 124174 112096 124180 112108
rect 121012 112068 124180 112096
rect 121012 112056 121018 112068
rect 124174 112056 124180 112068
rect 124232 112056 124238 112108
rect 190598 112056 190604 112108
rect 190656 112096 190662 112108
rect 192438 112096 192444 112108
rect 190656 112068 192444 112096
rect 190656 112056 190662 112068
rect 192438 112056 192444 112068
rect 192496 112056 192502 112108
rect 53058 111988 53064 112040
rect 53116 112028 53122 112040
rect 57658 112028 57664 112040
rect 53116 112000 57664 112028
rect 53116 111988 53122 112000
rect 57658 111988 57664 112000
rect 57716 111988 57722 112040
rect 51862 111920 51868 111972
rect 51920 111960 51926 111972
rect 55634 111960 55640 111972
rect 51920 111932 55640 111960
rect 51920 111920 51926 111932
rect 55634 111920 55640 111932
rect 55692 111920 55698 111972
rect 35210 111852 35216 111904
rect 35268 111892 35274 111904
rect 39810 111892 39816 111904
rect 35268 111864 39816 111892
rect 35268 111852 35274 111864
rect 39810 111852 39816 111864
rect 39868 111852 39874 111904
rect 52506 111852 52512 111904
rect 52564 111892 52570 111904
rect 56370 111892 56376 111904
rect 52564 111864 56376 111892
rect 52564 111852 52570 111864
rect 56370 111852 56376 111864
rect 56428 111852 56434 111904
rect 53794 111784 53800 111836
rect 53852 111824 53858 111836
rect 59038 111824 59044 111836
rect 53852 111796 59044 111824
rect 53852 111784 53858 111796
rect 59038 111784 59044 111796
rect 59096 111784 59102 111836
rect 54254 111716 54260 111768
rect 54312 111756 54318 111768
rect 59774 111756 59780 111768
rect 54312 111728 59780 111756
rect 54312 111716 54318 111728
rect 59774 111716 59780 111728
rect 59832 111716 59838 111768
rect 35854 111648 35860 111700
rect 35912 111688 35918 111700
rect 40270 111688 40276 111700
rect 35912 111660 40276 111688
rect 35912 111648 35918 111660
rect 40270 111648 40276 111660
rect 40328 111648 40334 111700
rect 53426 111648 53432 111700
rect 53484 111688 53490 111700
rect 58394 111688 58400 111700
rect 53484 111660 58400 111688
rect 53484 111648 53490 111660
rect 58394 111648 58400 111660
rect 58452 111648 58458 111700
rect 33830 111580 33836 111632
rect 33888 111620 33894 111632
rect 39074 111620 39080 111632
rect 33888 111592 39080 111620
rect 33888 111580 33894 111592
rect 39074 111580 39080 111592
rect 39132 111580 39138 111632
rect 54622 111580 54628 111632
rect 54680 111620 54686 111632
rect 60418 111620 60424 111632
rect 54680 111592 60424 111620
rect 54680 111580 54686 111592
rect 60418 111580 60424 111592
rect 60476 111580 60482 111632
rect 37878 111512 37884 111564
rect 37936 111552 37942 111564
rect 41466 111552 41472 111564
rect 37936 111524 41472 111552
rect 37936 111512 37942 111524
rect 41466 111512 41472 111524
rect 41524 111512 41530 111564
rect 39258 111444 39264 111496
rect 39316 111484 39322 111496
rect 42202 111484 42208 111496
rect 39316 111456 42208 111484
rect 39316 111444 39322 111456
rect 42202 111444 42208 111456
rect 42260 111444 42266 111496
rect 118838 111444 118844 111496
rect 118896 111484 118902 111496
rect 121414 111484 121420 111496
rect 118896 111456 121420 111484
rect 118896 111444 118902 111456
rect 121414 111444 121420 111456
rect 121472 111444 121478 111496
rect 39994 111376 40000 111428
rect 40052 111416 40058 111428
rect 42294 111416 42300 111428
rect 40052 111388 42300 111416
rect 40052 111376 40058 111388
rect 42294 111376 42300 111388
rect 42352 111376 42358 111428
rect 48274 111376 48280 111428
rect 48332 111416 48338 111428
rect 49470 111416 49476 111428
rect 48332 111388 49476 111416
rect 48332 111376 48338 111388
rect 49470 111376 49476 111388
rect 49528 111376 49534 111428
rect 50666 111376 50672 111428
rect 50724 111416 50730 111428
rect 53610 111416 53616 111428
rect 50724 111388 53616 111416
rect 50724 111376 50730 111388
rect 53610 111376 53616 111388
rect 53668 111376 53674 111428
rect 117458 111376 117464 111428
rect 117516 111416 117522 111428
rect 119758 111416 119764 111428
rect 117516 111388 119764 111416
rect 117516 111376 117522 111388
rect 119758 111376 119764 111388
rect 119816 111376 119822 111428
rect 182226 111376 182232 111428
rect 182284 111416 182290 111428
rect 183238 111416 183244 111428
rect 182284 111388 183244 111416
rect 182284 111376 182290 111388
rect 183238 111376 183244 111388
rect 183296 111376 183302 111428
rect 194094 111376 194100 111428
rect 194152 111416 194158 111428
rect 197130 111416 197136 111428
rect 194152 111388 197136 111416
rect 194152 111376 194158 111388
rect 197130 111376 197136 111388
rect 197188 111376 197194 111428
rect 40638 111308 40644 111360
rect 40696 111348 40702 111360
rect 43030 111348 43036 111360
rect 40696 111320 43036 111348
rect 40696 111308 40702 111320
rect 43030 111308 43036 111320
rect 43088 111308 43094 111360
rect 43398 111308 43404 111360
rect 43456 111348 43462 111360
rect 44594 111348 44600 111360
rect 43456 111320 44600 111348
rect 43456 111308 43462 111320
rect 44594 111308 44600 111320
rect 44652 111308 44658 111360
rect 47814 111308 47820 111360
rect 47872 111348 47878 111360
rect 48826 111348 48832 111360
rect 47872 111320 48832 111348
rect 47872 111308 47878 111320
rect 48826 111308 48832 111320
rect 48884 111308 48890 111360
rect 49838 111308 49844 111360
rect 49896 111348 49902 111360
rect 52230 111348 52236 111360
rect 49896 111320 52236 111348
rect 49896 111308 49902 111320
rect 52230 111308 52236 111320
rect 52288 111308 52294 111360
rect 117366 111308 117372 111360
rect 117424 111348 117430 111360
rect 119206 111348 119212 111360
rect 117424 111320 119212 111348
rect 117424 111308 117430 111320
rect 119206 111308 119212 111320
rect 119264 111308 119270 111360
rect 182870 111308 182876 111360
rect 182928 111348 182934 111360
rect 183790 111348 183796 111360
rect 182928 111320 183796 111348
rect 182928 111308 182934 111320
rect 183790 111308 183796 111320
rect 183848 111308 183854 111360
rect 191978 111308 191984 111360
rect 192036 111348 192042 111360
rect 194278 111348 194284 111360
rect 192036 111320 194284 111348
rect 192036 111308 192042 111320
rect 194278 111308 194284 111320
rect 194336 111308 194342 111360
rect 195290 111308 195296 111360
rect 195348 111348 195354 111360
rect 198786 111348 198792 111360
rect 195348 111320 198792 111348
rect 195348 111308 195354 111320
rect 198786 111308 198792 111320
rect 198844 111308 198850 111360
rect 37234 111240 37240 111292
rect 37292 111280 37298 111292
rect 41006 111280 41012 111292
rect 37292 111252 41012 111280
rect 37292 111240 37298 111252
rect 41006 111240 41012 111252
rect 41064 111240 41070 111292
rect 48642 111240 48648 111292
rect 48700 111280 48706 111292
rect 50206 111280 50212 111292
rect 48700 111252 50212 111280
rect 48700 111240 48706 111252
rect 50206 111240 50212 111252
rect 50264 111240 50270 111292
rect 51402 111240 51408 111292
rect 51460 111280 51466 111292
rect 54990 111280 54996 111292
rect 51460 111252 54996 111280
rect 51460 111240 51466 111252
rect 54990 111240 54996 111252
rect 55048 111240 55054 111292
rect 118562 111240 118568 111292
rect 118620 111280 118626 111292
rect 120862 111280 120868 111292
rect 118620 111252 120868 111280
rect 118620 111240 118626 111252
rect 120862 111240 120868 111252
rect 120920 111240 120926 111292
rect 36590 111172 36596 111224
rect 36648 111212 36654 111224
rect 40638 111212 40644 111224
rect 36648 111184 40644 111212
rect 36648 111172 36654 111184
rect 40638 111172 40644 111184
rect 40696 111172 40702 111224
rect 41282 111172 41288 111224
rect 41340 111212 41346 111224
rect 43398 111212 43404 111224
rect 41340 111184 43404 111212
rect 41340 111172 41346 111184
rect 43398 111172 43404 111184
rect 43456 111172 43462 111224
rect 44318 111172 44324 111224
rect 44376 111212 44382 111224
rect 45054 111212 45060 111224
rect 44376 111184 45060 111212
rect 44376 111172 44382 111184
rect 45054 111172 45060 111184
rect 45112 111172 45118 111224
rect 49470 111172 49476 111224
rect 49528 111212 49534 111224
rect 51586 111212 51592 111224
rect 49528 111184 51592 111212
rect 49528 111172 49534 111184
rect 51586 111172 51592 111184
rect 51644 111172 51650 111224
rect 105222 111172 105228 111224
rect 105280 111212 105286 111224
rect 106602 111212 106608 111224
rect 105280 111184 106608 111212
rect 105280 111172 105286 111184
rect 106602 111172 106608 111184
rect 106660 111172 106666 111224
rect 119758 111172 119764 111224
rect 119816 111212 119822 111224
rect 122518 111212 122524 111224
rect 119816 111184 122524 111212
rect 119816 111172 119822 111184
rect 122518 111172 122524 111184
rect 122576 111172 122582 111224
rect 177258 111172 177264 111224
rect 177316 111212 177322 111224
rect 178270 111212 178276 111224
rect 177316 111184 178276 111212
rect 177316 111172 177322 111184
rect 178270 111172 178276 111184
rect 178328 111172 178334 111224
rect 42018 111104 42024 111156
rect 42076 111144 42082 111156
rect 43858 111144 43864 111156
rect 42076 111116 43864 111144
rect 42076 111104 42082 111116
rect 43858 111104 43864 111116
rect 43916 111104 43922 111156
rect 50206 111104 50212 111156
rect 50264 111144 50270 111156
rect 52966 111144 52972 111156
rect 50264 111116 52972 111144
rect 50264 111104 50270 111116
rect 52966 111104 52972 111116
rect 53024 111104 53030 111156
rect 105498 111104 105504 111156
rect 105556 111144 105562 111156
rect 107154 111144 107160 111156
rect 105556 111116 107160 111144
rect 105556 111104 105562 111116
rect 107154 111104 107160 111116
rect 107212 111104 107218 111156
rect 177074 111104 177080 111156
rect 177132 111144 177138 111156
rect 178822 111144 178828 111156
rect 177132 111116 178828 111144
rect 177132 111104 177138 111116
rect 178822 111104 178828 111116
rect 178880 111104 178886 111156
rect 38614 111036 38620 111088
rect 38672 111076 38678 111088
rect 41834 111076 41840 111088
rect 38672 111048 41840 111076
rect 38672 111036 38678 111048
rect 41834 111036 41840 111048
rect 41892 111036 41898 111088
rect 49010 111036 49016 111088
rect 49068 111076 49074 111088
rect 50850 111076 50856 111088
rect 49068 111048 50856 111076
rect 49068 111036 49074 111048
rect 50850 111036 50856 111048
rect 50908 111036 50914 111088
rect 105682 111036 105688 111088
rect 105740 111076 105746 111088
rect 107706 111076 107712 111088
rect 105740 111048 107712 111076
rect 105740 111036 105746 111048
rect 107706 111036 107712 111048
rect 107764 111036 107770 111088
rect 176890 111036 176896 111088
rect 176948 111076 176954 111088
rect 179374 111076 179380 111088
rect 176948 111048 179380 111076
rect 176948 111036 176954 111048
rect 179374 111036 179380 111048
rect 179432 111036 179438 111088
rect 42662 110968 42668 111020
rect 42720 111008 42726 111020
rect 44226 111008 44232 111020
rect 42720 110980 44232 111008
rect 42720 110968 42726 110980
rect 44226 110968 44232 110980
rect 44284 110968 44290 111020
rect 108810 111008 108816 111020
rect 106528 110980 108816 111008
rect 105958 110900 105964 110952
rect 106016 110940 106022 110952
rect 106528 110940 106556 110980
rect 108810 110968 108816 110980
rect 108868 110968 108874 111020
rect 176982 110968 176988 111020
rect 177040 111008 177046 111020
rect 180018 111008 180024 111020
rect 177040 110980 180024 111008
rect 177040 110968 177046 110980
rect 180018 110968 180024 110980
rect 180076 110968 180082 111020
rect 181674 110968 181680 111020
rect 181732 111008 181738 111020
rect 183100 111008 183106 111020
rect 181732 110980 183106 111008
rect 181732 110968 181738 110980
rect 183100 110968 183106 110980
rect 183158 110968 183164 111020
rect 183422 110968 183428 111020
rect 183480 111008 183486 111020
rect 184296 111008 184302 111020
rect 183480 110980 184302 111008
rect 183480 110968 183486 110980
rect 184296 110968 184302 110980
rect 184354 110968 184360 111020
rect 106016 110912 106556 110940
rect 106016 110900 106022 110912
rect 177718 110900 177724 110952
rect 177776 110940 177782 110952
rect 181122 110940 181128 110952
rect 177776 110912 181128 110940
rect 177776 110900 177782 110912
rect 181122 110900 181128 110912
rect 181180 110900 181186 110952
rect 132546 110220 132552 110272
rect 132604 110260 132610 110272
rect 132733 110263 132791 110269
rect 132733 110260 132745 110263
rect 132604 110232 132745 110260
rect 132604 110220 132610 110232
rect 132733 110229 132745 110232
rect 132779 110229 132791 110263
rect 132733 110223 132791 110229
rect 222706 110220 222712 110272
rect 222764 110260 222770 110272
rect 222801 110263 222859 110269
rect 222801 110260 222813 110263
rect 222764 110232 222813 110260
rect 222764 110220 222770 110232
rect 222801 110229 222813 110232
rect 222847 110229 222859 110263
rect 222801 110223 222859 110229
rect 105774 109472 105780 109524
rect 105832 109512 105838 109524
rect 108258 109512 108264 109524
rect 105832 109484 108264 109512
rect 105832 109472 105838 109484
rect 108258 109472 108264 109484
rect 108316 109472 108322 109524
rect 177350 108996 177356 109048
rect 177408 109036 177414 109048
rect 180570 109036 180576 109048
rect 177408 109008 180576 109036
rect 177408 108996 177414 109008
rect 180570 108996 180576 109008
rect 180628 108996 180634 109048
rect 222798 107948 222804 107960
rect 222759 107920 222804 107948
rect 222798 107908 222804 107920
rect 222856 107908 222862 107960
rect 32634 104032 32640 104084
rect 32692 104072 32698 104084
rect 37418 104072 37424 104084
rect 32692 104044 37424 104072
rect 32692 104032 32698 104044
rect 37418 104032 37424 104044
rect 37476 104032 37482 104084
rect 105682 104032 105688 104084
rect 105740 104072 105746 104084
rect 107890 104072 107896 104084
rect 105740 104044 107896 104072
rect 105740 104032 105746 104044
rect 107890 104032 107896 104044
rect 107948 104032 107954 104084
rect 178178 104032 178184 104084
rect 178236 104072 178242 104084
rect 179650 104072 179656 104084
rect 178236 104044 179656 104072
rect 178236 104032 178242 104044
rect 179650 104032 179656 104044
rect 179708 104032 179714 104084
rect 106326 101312 106332 101364
rect 106384 101352 106390 101364
rect 107890 101352 107896 101364
rect 106384 101324 107896 101352
rect 106384 101312 106390 101324
rect 107890 101312 107896 101324
rect 107948 101312 107954 101364
rect 177626 101312 177632 101364
rect 177684 101352 177690 101364
rect 179650 101352 179656 101364
rect 177684 101324 179656 101352
rect 177684 101312 177690 101324
rect 179650 101312 179656 101324
rect 179708 101312 179714 101364
rect 57566 100972 57572 101024
rect 57624 101012 57630 101024
rect 60510 101012 60516 101024
rect 57624 100984 60516 101012
rect 57624 100972 57630 100984
rect 60510 100972 60516 100984
rect 60568 100972 60574 101024
rect 105958 100768 105964 100820
rect 106016 100808 106022 100820
rect 108626 100808 108632 100820
rect 106016 100780 108632 100808
rect 106016 100768 106022 100780
rect 108626 100768 108632 100780
rect 108684 100768 108690 100820
rect 176982 100768 176988 100820
rect 177040 100808 177046 100820
rect 180294 100808 180300 100820
rect 177040 100780 180300 100808
rect 177040 100768 177046 100780
rect 180294 100768 180300 100780
rect 180352 100768 180358 100820
rect 106418 99884 106424 99936
rect 106476 99924 106482 99936
rect 107890 99924 107896 99936
rect 106476 99896 107896 99924
rect 106476 99884 106482 99896
rect 107890 99884 107896 99896
rect 107948 99884 107954 99936
rect 177718 99884 177724 99936
rect 177776 99924 177782 99936
rect 179650 99924 179656 99936
rect 177776 99896 179656 99924
rect 177776 99884 177782 99896
rect 179650 99884 179656 99896
rect 179708 99884 179714 99936
rect 105590 99408 105596 99460
rect 105648 99448 105654 99460
rect 108534 99448 108540 99460
rect 105648 99420 108540 99448
rect 105648 99408 105654 99420
rect 108534 99408 108540 99420
rect 108592 99408 108598 99460
rect 177350 99272 177356 99324
rect 177408 99312 177414 99324
rect 180386 99312 180392 99324
rect 177408 99284 180392 99312
rect 177408 99272 177414 99284
rect 180386 99272 180392 99284
rect 180444 99272 180450 99324
rect 105774 97164 105780 97216
rect 105832 97204 105838 97216
rect 107890 97204 107896 97216
rect 105832 97176 107896 97204
rect 105832 97164 105838 97176
rect 107890 97164 107896 97176
rect 107948 97164 107954 97216
rect 177534 97164 177540 97216
rect 177592 97204 177598 97216
rect 179650 97204 179656 97216
rect 177592 97176 179656 97204
rect 177592 97164 177598 97176
rect 179650 97164 179656 97176
rect 179708 97164 179714 97216
rect 222982 97096 222988 97148
rect 223040 97136 223046 97148
rect 223534 97136 223540 97148
rect 223040 97108 223540 97136
rect 223040 97096 223046 97108
rect 223534 97096 223540 97108
rect 223592 97096 223598 97148
rect 105774 94308 105780 94360
rect 105832 94348 105838 94360
rect 107798 94348 107804 94360
rect 105832 94320 107804 94348
rect 105832 94308 105838 94320
rect 107798 94308 107804 94320
rect 107856 94308 107862 94360
rect 177350 93900 177356 93952
rect 177408 93940 177414 93952
rect 179558 93940 179564 93952
rect 177408 93912 179564 93940
rect 177408 93900 177414 93912
rect 179558 93900 179564 93912
rect 179616 93900 179622 93952
rect 222798 92540 222804 92592
rect 222856 92580 222862 92592
rect 223534 92580 223540 92592
rect 222856 92552 223540 92580
rect 222856 92540 222862 92552
rect 223534 92540 223540 92552
rect 223592 92540 223598 92592
rect 105222 92064 105228 92116
rect 105280 92104 105286 92116
rect 107798 92104 107804 92116
rect 105280 92076 107804 92104
rect 105280 92064 105286 92076
rect 107798 92064 107804 92076
rect 107856 92064 107862 92116
rect 176982 91996 176988 92048
rect 177040 92036 177046 92048
rect 179558 92036 179564 92048
rect 177040 92008 179564 92036
rect 177040 91996 177046 92008
rect 179558 91996 179564 92008
rect 179616 91996 179622 92048
rect 201086 91588 201092 91640
rect 201144 91628 201150 91640
rect 204490 91628 204496 91640
rect 201144 91600 204496 91628
rect 201144 91588 201150 91600
rect 204490 91588 204496 91600
rect 204548 91588 204554 91640
rect 28862 90228 28868 90280
rect 28920 90268 28926 90280
rect 36406 90268 36412 90280
rect 28920 90240 36412 90268
rect 28920 90228 28926 90240
rect 36406 90228 36412 90240
rect 36464 90228 36470 90280
rect 54809 90271 54867 90277
rect 54809 90237 54821 90271
rect 54855 90268 54867 90271
rect 59590 90268 59596 90280
rect 54855 90240 59596 90268
rect 54855 90237 54867 90240
rect 54809 90231 54867 90237
rect 59590 90228 59596 90240
rect 59648 90228 59654 90280
rect 105774 89208 105780 89260
rect 105832 89248 105838 89260
rect 107798 89248 107804 89260
rect 105832 89220 107804 89248
rect 105832 89208 105838 89220
rect 107798 89208 107804 89220
rect 107856 89208 107862 89260
rect 132362 88868 132368 88920
rect 132420 88868 132426 88920
rect 132380 88840 132408 88868
rect 132546 88840 132552 88852
rect 132380 88812 132552 88840
rect 132546 88800 132552 88812
rect 132604 88800 132610 88852
rect 105406 87848 105412 87900
rect 105464 87888 105470 87900
rect 107890 87888 107896 87900
rect 105464 87860 107896 87888
rect 105464 87848 105470 87860
rect 107890 87848 107896 87860
rect 107948 87848 107954 87900
rect 177350 87508 177356 87560
rect 177408 87548 177414 87560
rect 179650 87548 179656 87560
rect 177408 87520 179656 87548
rect 177408 87508 177414 87520
rect 179650 87508 179656 87520
rect 179708 87508 179714 87560
rect 106418 86352 106424 86404
rect 106476 86392 106482 86404
rect 107982 86392 107988 86404
rect 106476 86364 107988 86392
rect 106476 86352 106482 86364
rect 107982 86352 107988 86364
rect 108040 86352 108046 86404
rect 54806 86120 54812 86132
rect 54767 86092 54812 86120
rect 54806 86080 54812 86092
rect 54864 86080 54870 86132
rect 177534 86080 177540 86132
rect 177592 86120 177598 86132
rect 179742 86120 179748 86132
rect 177592 86092 179748 86120
rect 177592 86080 177598 86092
rect 179742 86080 179748 86092
rect 179800 86080 179806 86132
rect 54806 85984 54812 85996
rect 54767 85956 54812 85984
rect 54806 85944 54812 85956
rect 54864 85944 54870 85996
rect 105130 84788 105136 84840
rect 105188 84828 105194 84840
rect 107798 84828 107804 84840
rect 105188 84800 107804 84828
rect 105188 84788 105194 84800
rect 107798 84788 107804 84800
rect 107856 84788 107862 84840
rect 176982 84788 176988 84840
rect 177040 84828 177046 84840
rect 179558 84828 179564 84840
rect 177040 84800 179564 84828
rect 177040 84788 177046 84800
rect 179558 84788 179564 84800
rect 179616 84788 179622 84840
rect 222798 84788 222804 84840
rect 222856 84828 222862 84840
rect 223534 84828 223540 84840
rect 222856 84800 223540 84828
rect 222856 84788 222862 84800
rect 223534 84788 223540 84800
rect 223592 84788 223598 84840
rect 105682 84720 105688 84772
rect 105740 84760 105746 84772
rect 107614 84760 107620 84772
rect 105740 84732 107620 84760
rect 105740 84720 105746 84732
rect 107614 84720 107620 84732
rect 107672 84720 107678 84772
rect 178178 84720 178184 84772
rect 178236 84760 178242 84772
rect 179650 84760 179656 84772
rect 178236 84732 179656 84760
rect 178236 84720 178242 84732
rect 179650 84720 179656 84732
rect 179708 84720 179714 84772
rect 178086 83428 178092 83480
rect 178144 83468 178150 83480
rect 179466 83468 179472 83480
rect 178144 83440 179472 83468
rect 178144 83428 178150 83440
rect 179466 83428 179472 83440
rect 179524 83428 179530 83480
rect 105222 83360 105228 83412
rect 105280 83400 105286 83412
rect 107706 83400 107712 83412
rect 105280 83372 107712 83400
rect 105280 83360 105286 83372
rect 107706 83360 107712 83372
rect 107764 83360 107770 83412
rect 177718 82272 177724 82324
rect 177776 82312 177782 82324
rect 179742 82312 179748 82324
rect 177776 82284 179748 82312
rect 177776 82272 177782 82284
rect 179742 82272 179748 82284
rect 179800 82272 179806 82324
rect 106418 82136 106424 82188
rect 106476 82176 106482 82188
rect 107890 82176 107896 82188
rect 106476 82148 107896 82176
rect 106476 82136 106482 82148
rect 107890 82136 107896 82148
rect 107948 82136 107954 82188
rect 105958 80776 105964 80828
rect 106016 80816 106022 80828
rect 108534 80816 108540 80828
rect 106016 80788 108540 80816
rect 106016 80776 106022 80788
rect 108534 80776 108540 80788
rect 108592 80776 108598 80828
rect 178086 80572 178092 80624
rect 178144 80612 178150 80624
rect 180294 80612 180300 80624
rect 178144 80584 180300 80612
rect 178144 80572 178150 80584
rect 180294 80572 180300 80584
rect 180352 80572 180358 80624
rect 132546 79280 132552 79332
rect 132604 79280 132610 79332
rect 105406 79212 105412 79264
rect 105464 79252 105470 79264
rect 108074 79252 108080 79264
rect 105464 79224 108080 79252
rect 105464 79212 105470 79224
rect 108074 79212 108080 79224
rect 108132 79212 108138 79264
rect 132564 79196 132592 79280
rect 177626 79212 177632 79264
rect 177684 79252 177690 79264
rect 180018 79252 180024 79264
rect 177684 79224 180024 79252
rect 177684 79212 177690 79224
rect 180018 79212 180024 79224
rect 180076 79212 180082 79264
rect 132546 79144 132552 79196
rect 132604 79144 132610 79196
rect 105222 77852 105228 77904
rect 105280 77892 105286 77904
rect 107522 77892 107528 77904
rect 105280 77864 107528 77892
rect 105280 77852 105286 77864
rect 107522 77852 107528 77864
rect 107580 77852 107586 77904
rect 176982 77852 176988 77904
rect 177040 77892 177046 77904
rect 179374 77892 179380 77904
rect 177040 77864 179380 77892
rect 177040 77852 177046 77864
rect 179374 77852 179380 77864
rect 179432 77852 179438 77904
rect 30518 77784 30524 77836
rect 30576 77824 30582 77836
rect 37418 77824 37424 77836
rect 30576 77796 37424 77824
rect 30576 77784 30582 77796
rect 37418 77784 37424 77796
rect 37476 77784 37482 77836
rect 57474 77580 57480 77632
rect 57532 77620 57538 77632
rect 59590 77620 59596 77632
rect 57532 77592 59596 77620
rect 57532 77580 57538 77592
rect 59590 77580 59596 77592
rect 59648 77580 59654 77632
rect 54809 76467 54867 76473
rect 54809 76433 54821 76467
rect 54855 76464 54867 76467
rect 54990 76464 54996 76476
rect 54855 76436 54996 76464
rect 54855 76433 54867 76436
rect 54809 76427 54867 76433
rect 54990 76424 54996 76436
rect 55048 76424 55054 76476
rect 222982 75064 222988 75116
rect 223040 75104 223046 75116
rect 223534 75104 223540 75116
rect 223040 75076 223540 75104
rect 223040 75064 223046 75076
rect 223534 75064 223540 75076
rect 223592 75064 223598 75116
rect 222798 73568 222804 73620
rect 222856 73608 222862 73620
rect 223074 73608 223080 73620
rect 222856 73580 223080 73608
rect 222856 73568 222862 73580
rect 223074 73568 223080 73580
rect 223132 73568 223138 73620
rect 105866 72412 105872 72464
rect 105924 72452 105930 72464
rect 109178 72452 109184 72464
rect 105924 72424 109184 72452
rect 105924 72412 105930 72424
rect 109178 72412 109184 72424
rect 109236 72412 109242 72464
rect 177626 72344 177632 72396
rect 177684 72384 177690 72396
rect 180938 72384 180944 72396
rect 177684 72356 180944 72384
rect 177684 72344 177690 72356
rect 180938 72344 180944 72356
rect 180996 72344 181002 72396
rect 177350 70916 177356 70968
rect 177408 70956 177414 70968
rect 177408 70928 178316 70956
rect 177408 70916 177414 70928
rect 178288 70888 178316 70928
rect 180570 70888 180576 70900
rect 178288 70860 180576 70888
rect 180570 70848 180576 70860
rect 180628 70848 180634 70900
rect 189816 70712 189822 70764
rect 189874 70752 189880 70764
rect 191426 70752 191432 70764
rect 189874 70724 191432 70752
rect 189874 70712 189880 70724
rect 191426 70712 191432 70724
rect 191484 70712 191490 70764
rect 182870 70644 182876 70696
rect 182928 70684 182934 70696
rect 183836 70684 183842 70696
rect 182928 70656 183842 70684
rect 182928 70644 182934 70656
rect 183836 70644 183842 70656
rect 183894 70644 183900 70696
rect 189448 70644 189454 70696
rect 189506 70684 189512 70696
rect 190782 70684 190788 70696
rect 189506 70656 190788 70684
rect 189506 70644 189512 70656
rect 190782 70644 190788 70656
rect 190840 70644 190846 70696
rect 191840 70644 191846 70696
rect 191898 70684 191904 70696
rect 194278 70684 194284 70696
rect 191898 70656 194284 70684
rect 191898 70644 191904 70656
rect 194278 70644 194284 70656
rect 194336 70644 194342 70696
rect 106510 70304 106516 70356
rect 106568 70344 106574 70356
rect 108350 70344 108356 70356
rect 106568 70316 108356 70344
rect 106568 70304 106574 70316
rect 108350 70304 108356 70316
rect 108408 70304 108414 70356
rect 49470 69760 49476 69812
rect 49528 69800 49534 69812
rect 51586 69800 51592 69812
rect 49528 69772 51592 69800
rect 49528 69760 49534 69772
rect 51586 69760 51592 69772
rect 51644 69760 51650 69812
rect 119850 69760 119856 69812
rect 119908 69800 119914 69812
rect 122334 69800 122340 69812
rect 119908 69772 122340 69800
rect 119908 69760 119914 69772
rect 122334 69760 122340 69772
rect 122392 69760 122398 69812
rect 48642 69692 48648 69744
rect 48700 69732 48706 69744
rect 50206 69732 50212 69744
rect 48700 69704 50212 69732
rect 48700 69692 48706 69704
rect 50206 69692 50212 69704
rect 50264 69692 50270 69744
rect 119482 69692 119488 69744
rect 119540 69732 119546 69744
rect 121690 69732 121696 69744
rect 119540 69704 121696 69732
rect 119540 69692 119546 69704
rect 121690 69692 121696 69704
rect 121748 69692 121754 69744
rect 48274 69624 48280 69676
rect 48332 69664 48338 69676
rect 49470 69664 49476 69676
rect 48332 69636 49476 69664
rect 48332 69624 48338 69636
rect 49470 69624 49476 69636
rect 49528 69624 49534 69676
rect 49838 69624 49844 69676
rect 49896 69664 49902 69676
rect 52230 69664 52236 69676
rect 49896 69636 52236 69664
rect 49896 69624 49902 69636
rect 52230 69624 52236 69636
rect 52288 69624 52294 69676
rect 117090 69624 117096 69676
rect 117148 69664 117154 69676
rect 118194 69664 118200 69676
rect 117148 69636 118200 69664
rect 117148 69624 117154 69636
rect 118194 69624 118200 69636
rect 118252 69624 118258 69676
rect 118654 69624 118660 69676
rect 118712 69664 118718 69676
rect 120586 69664 120592 69676
rect 118712 69636 120592 69664
rect 118712 69624 118718 69636
rect 120586 69624 120592 69636
rect 120644 69624 120650 69676
rect 191702 69624 191708 69676
rect 191760 69664 191766 69676
rect 193634 69664 193640 69676
rect 191760 69636 193640 69664
rect 191760 69624 191766 69636
rect 193634 69624 193640 69636
rect 193692 69624 193698 69676
rect 39258 69556 39264 69608
rect 39316 69596 39322 69608
rect 39316 69568 40408 69596
rect 39316 69556 39322 69568
rect 22238 69488 22244 69540
rect 22296 69528 22302 69540
rect 28678 69528 28684 69540
rect 22296 69500 28684 69528
rect 22296 69488 22302 69500
rect 28678 69488 28684 69500
rect 28736 69488 28742 69540
rect 35949 69531 36007 69537
rect 35949 69528 35961 69531
rect 35228 69500 35961 69528
rect 16626 69420 16632 69472
rect 16684 69460 16690 69472
rect 31898 69460 31904 69472
rect 16684 69432 31904 69460
rect 16684 69420 16690 69432
rect 31898 69420 31904 69432
rect 31956 69460 31962 69472
rect 35228 69460 35256 69500
rect 35949 69497 35961 69500
rect 35995 69497 36007 69531
rect 35949 69491 36007 69497
rect 36038 69488 36044 69540
rect 36096 69528 36102 69540
rect 40270 69528 40276 69540
rect 36096 69500 40276 69528
rect 36096 69488 36102 69500
rect 40270 69488 40276 69500
rect 40328 69488 40334 69540
rect 40380 69528 40408 69568
rect 47814 69556 47820 69608
rect 47872 69596 47878 69608
rect 48826 69596 48832 69608
rect 47872 69568 48832 69596
rect 47872 69556 47878 69568
rect 48826 69556 48832 69568
rect 48884 69556 48890 69608
rect 49010 69556 49016 69608
rect 49068 69596 49074 69608
rect 50850 69596 50856 69608
rect 49068 69568 50856 69596
rect 49068 69556 49074 69568
rect 50850 69556 50856 69568
rect 50908 69556 50914 69608
rect 54990 69596 54996 69608
rect 51788 69568 54996 69596
rect 42202 69528 42208 69540
rect 40380 69500 42208 69528
rect 42202 69488 42208 69500
rect 42260 69488 42266 69540
rect 31956 69432 35256 69460
rect 31956 69420 31962 69432
rect 35578 69420 35584 69472
rect 35636 69460 35642 69472
rect 39810 69460 39816 69472
rect 35636 69432 39816 69460
rect 35636 69420 35642 69432
rect 39810 69420 39816 69432
rect 39868 69420 39874 69472
rect 34658 69352 34664 69404
rect 34716 69392 34722 69404
rect 39442 69392 39448 69404
rect 34716 69364 39448 69392
rect 34716 69352 34722 69364
rect 39442 69352 39448 69364
rect 39500 69352 39506 69404
rect 27574 69284 27580 69336
rect 27632 69324 27638 69336
rect 51788 69324 51816 69568
rect 54990 69556 54996 69568
rect 55048 69556 55054 69608
rect 59038 69596 59044 69608
rect 57216 69568 59044 69596
rect 53794 69488 53800 69540
rect 53852 69528 53858 69540
rect 57216 69528 57244 69568
rect 59038 69556 59044 69568
rect 59096 69556 59102 69608
rect 116630 69556 116636 69608
rect 116688 69596 116694 69608
rect 117642 69596 117648 69608
rect 116688 69568 117648 69596
rect 116688 69556 116694 69568
rect 117642 69556 117648 69568
rect 117700 69556 117706 69608
rect 118286 69556 118292 69608
rect 118344 69596 118350 69608
rect 120310 69596 120316 69608
rect 118344 69568 120316 69596
rect 118344 69556 118350 69568
rect 120310 69556 120316 69568
rect 120368 69556 120374 69608
rect 131626 69596 131632 69608
rect 131276 69568 131632 69596
rect 53852 69500 57244 69528
rect 53852 69488 53858 69500
rect 126290 69488 126296 69540
rect 126348 69528 126354 69540
rect 131276 69528 131304 69568
rect 131626 69556 131632 69568
rect 131684 69556 131690 69608
rect 190414 69556 190420 69608
rect 190472 69596 190478 69608
rect 191978 69596 191984 69608
rect 190472 69568 191984 69596
rect 190472 69556 190478 69568
rect 191978 69556 191984 69568
rect 192036 69556 192042 69608
rect 203938 69596 203944 69608
rect 200920 69568 203944 69596
rect 126348 69500 131304 69528
rect 126348 69488 126354 69500
rect 198878 69488 198884 69540
rect 198936 69528 198942 69540
rect 200920 69528 200948 69568
rect 203938 69556 203944 69568
rect 203996 69556 204002 69608
rect 198936 69500 200948 69528
rect 198936 69488 198942 69500
rect 200994 69488 201000 69540
rect 201052 69528 201058 69540
rect 215898 69528 215904 69540
rect 201052 69500 215904 69528
rect 201052 69488 201058 69500
rect 215898 69488 215904 69500
rect 215956 69488 215962 69540
rect 53426 69420 53432 69472
rect 53484 69460 53490 69472
rect 58118 69460 58124 69472
rect 53484 69432 58124 69460
rect 53484 69420 53490 69432
rect 58118 69420 58124 69432
rect 58176 69420 58182 69472
rect 123438 69420 123444 69472
rect 123496 69460 123502 69472
rect 127578 69460 127584 69472
rect 123496 69432 127584 69460
rect 123496 69420 123502 69432
rect 127578 69420 127584 69432
rect 127636 69420 127642 69472
rect 198510 69420 198516 69472
rect 198568 69460 198574 69472
rect 203018 69460 203024 69472
rect 198568 69432 203024 69460
rect 198568 69420 198574 69432
rect 203018 69420 203024 69432
rect 203076 69420 203082 69472
rect 54809 69395 54867 69401
rect 54809 69361 54821 69395
rect 54855 69392 54867 69395
rect 57474 69392 57480 69404
rect 54855 69364 57480 69392
rect 54855 69361 54867 69364
rect 54809 69355 54867 69361
rect 57474 69352 57480 69364
rect 57532 69352 57538 69404
rect 124634 69352 124640 69404
rect 124692 69392 124698 69404
rect 129326 69392 129332 69404
rect 124692 69364 129332 69392
rect 124692 69352 124698 69364
rect 129326 69352 129332 69364
rect 129384 69352 129390 69404
rect 196118 69352 196124 69404
rect 196176 69392 196182 69404
rect 199982 69392 199988 69404
rect 196176 69364 199988 69392
rect 196176 69352 196182 69364
rect 199982 69352 199988 69364
rect 200040 69352 200046 69404
rect 27632 69296 51816 69324
rect 27632 69284 27638 69296
rect 51862 69284 51868 69336
rect 51920 69324 51926 69336
rect 55177 69327 55235 69333
rect 55177 69324 55189 69327
rect 51920 69296 55189 69324
rect 51920 69284 51926 69296
rect 55177 69293 55189 69296
rect 55223 69293 55235 69327
rect 55177 69287 55235 69293
rect 91238 69284 91244 69336
rect 91296 69324 91302 69336
rect 132086 69324 132092 69336
rect 91296 69296 132092 69324
rect 91296 69284 91302 69296
rect 132086 69284 132092 69296
rect 132144 69284 132150 69336
rect 194554 69284 194560 69336
rect 194612 69324 194618 69336
rect 197682 69324 197688 69336
rect 194612 69296 197688 69324
rect 194612 69284 194618 69296
rect 197682 69284 197688 69296
rect 197740 69284 197746 69336
rect 201086 69284 201092 69336
rect 201144 69324 201150 69336
rect 210562 69324 210568 69336
rect 201144 69296 210568 69324
rect 201144 69284 201150 69296
rect 210562 69284 210568 69296
rect 210620 69284 210626 69336
rect 36041 69259 36099 69265
rect 36041 69225 36053 69259
rect 36087 69256 36099 69259
rect 36133 69259 36191 69265
rect 36133 69256 36145 69259
rect 36087 69228 36145 69256
rect 36087 69225 36099 69228
rect 36041 69219 36099 69225
rect 36133 69225 36145 69228
rect 36179 69225 36191 69259
rect 36133 69219 36191 69225
rect 121874 69216 121880 69268
rect 121932 69256 121938 69268
rect 125186 69256 125192 69268
rect 121932 69228 125192 69256
rect 121932 69216 121938 69228
rect 125186 69216 125192 69228
rect 125244 69216 125250 69268
rect 125462 69216 125468 69268
rect 125520 69256 125526 69268
rect 130430 69256 130436 69268
rect 125520 69228 130436 69256
rect 125520 69216 125526 69228
rect 130430 69216 130436 69228
rect 130488 69216 130494 69268
rect 196486 69216 196492 69268
rect 196544 69256 196550 69268
rect 200534 69256 200540 69268
rect 196544 69228 200540 69256
rect 196544 69216 196550 69228
rect 200534 69216 200540 69228
rect 200592 69216 200598 69268
rect 40178 69148 40184 69200
rect 40236 69188 40242 69200
rect 42662 69188 42668 69200
rect 40236 69160 42668 69188
rect 40236 69148 40242 69160
rect 42662 69148 42668 69160
rect 42720 69148 42726 69200
rect 54622 69148 54628 69200
rect 54680 69188 54686 69200
rect 60142 69188 60148 69200
rect 54680 69160 60148 69188
rect 54680 69148 54686 69160
rect 60142 69148 60148 69160
rect 60200 69148 60206 69200
rect 92342 69148 92348 69200
rect 92400 69188 92406 69200
rect 97494 69188 97500 69200
rect 92400 69160 97500 69188
rect 92400 69148 92406 69160
rect 97494 69148 97500 69160
rect 97552 69148 97558 69200
rect 122242 69148 122248 69200
rect 122300 69188 122306 69200
rect 122300 69160 124588 69188
rect 122300 69148 122306 69160
rect 34106 69080 34112 69132
rect 34164 69120 34170 69132
rect 39074 69120 39080 69132
rect 34164 69092 39080 69120
rect 34164 69080 34170 69092
rect 39074 69080 39080 69092
rect 39132 69080 39138 69132
rect 40638 69080 40644 69132
rect 40696 69120 40702 69132
rect 43030 69120 43036 69132
rect 40696 69092 43036 69120
rect 40696 69080 40702 69092
rect 43030 69080 43036 69092
rect 43088 69080 43094 69132
rect 52598 69080 52604 69132
rect 52656 69120 52662 69132
rect 56738 69120 56744 69132
rect 52656 69092 56744 69120
rect 52656 69080 52662 69092
rect 56738 69080 56744 69092
rect 56796 69080 56802 69132
rect 110558 69080 110564 69132
rect 110616 69120 110622 69132
rect 111478 69120 111484 69132
rect 110616 69092 111484 69120
rect 110616 69080 110622 69092
rect 111478 69080 111484 69092
rect 111536 69080 111542 69132
rect 121046 69080 121052 69132
rect 121104 69120 121110 69132
rect 124450 69120 124456 69132
rect 121104 69092 124456 69120
rect 121104 69080 121110 69092
rect 124450 69080 124456 69092
rect 124508 69080 124514 69132
rect 124560 69120 124588 69160
rect 125830 69148 125836 69200
rect 125888 69188 125894 69200
rect 131258 69188 131264 69200
rect 125888 69160 131264 69188
rect 125888 69148 125894 69160
rect 131258 69148 131264 69160
rect 131316 69148 131322 69200
rect 168886 69188 168892 69200
rect 161728 69160 168892 69188
rect 125922 69120 125928 69132
rect 124560 69092 125928 69120
rect 125922 69080 125928 69092
rect 125980 69080 125986 69132
rect 126658 69080 126664 69132
rect 126716 69120 126722 69132
rect 132178 69120 132184 69132
rect 126716 69092 132184 69120
rect 126716 69080 126722 69092
rect 132178 69080 132184 69092
rect 132236 69080 132242 69132
rect 36590 69012 36596 69064
rect 36648 69052 36654 69064
rect 40362 69052 40368 69064
rect 36648 69024 40368 69052
rect 36648 69012 36654 69024
rect 40362 69012 40368 69024
rect 40420 69012 40426 69064
rect 42018 69012 42024 69064
rect 42076 69052 42082 69064
rect 43858 69052 43864 69064
rect 42076 69024 43864 69052
rect 42076 69012 42082 69024
rect 43858 69012 43864 69024
rect 43916 69012 43922 69064
rect 53058 69012 53064 69064
rect 53116 69052 53122 69064
rect 57658 69052 57664 69064
rect 53116 69024 57664 69052
rect 53116 69012 53122 69024
rect 57658 69012 57664 69024
rect 57716 69012 57722 69064
rect 125094 69012 125100 69064
rect 125152 69052 125158 69064
rect 129878 69052 129884 69064
rect 125152 69024 129884 69052
rect 125152 69012 125158 69024
rect 129878 69012 129884 69024
rect 129936 69012 129942 69064
rect 37234 68944 37240 68996
rect 37292 68984 37298 68996
rect 41006 68984 41012 68996
rect 37292 68956 41012 68984
rect 37292 68944 37298 68956
rect 41006 68944 41012 68956
rect 41064 68944 41070 68996
rect 42662 68944 42668 68996
rect 42720 68984 42726 68996
rect 44226 68984 44232 68996
rect 42720 68956 44232 68984
rect 42720 68944 42726 68956
rect 44226 68944 44232 68956
rect 44284 68944 44290 68996
rect 52506 68944 52512 68996
rect 52564 68984 52570 68996
rect 52564 68956 54208 68984
rect 52564 68944 52570 68956
rect 41282 68876 41288 68928
rect 41340 68916 41346 68928
rect 43398 68916 43404 68928
rect 41340 68888 43404 68916
rect 41340 68876 41346 68888
rect 43398 68876 43404 68888
rect 43456 68876 43462 68928
rect 50666 68876 50672 68928
rect 50724 68916 50730 68928
rect 53610 68916 53616 68928
rect 50724 68888 53616 68916
rect 50724 68876 50730 68888
rect 53610 68876 53616 68888
rect 53668 68876 53674 68928
rect 54180 68916 54208 68956
rect 54254 68944 54260 68996
rect 54312 68984 54318 68996
rect 59498 68984 59504 68996
rect 54312 68956 59504 68984
rect 54312 68944 54318 68956
rect 59498 68944 59504 68956
rect 59556 68944 59562 68996
rect 62902 68944 62908 68996
rect 62960 68984 62966 68996
rect 67870 68984 67876 68996
rect 62960 68956 67876 68984
rect 62960 68944 62966 68956
rect 67870 68944 67876 68956
rect 67928 68944 67934 68996
rect 88938 68944 88944 68996
rect 88996 68984 89002 68996
rect 96850 68984 96856 68996
rect 88996 68956 96856 68984
rect 88996 68944 89002 68956
rect 96850 68944 96856 68956
rect 96908 68944 96914 68996
rect 122702 68944 122708 68996
rect 122760 68984 122766 68996
rect 126382 68984 126388 68996
rect 122760 68956 126388 68984
rect 122760 68944 122766 68956
rect 126382 68944 126388 68956
rect 126440 68944 126446 68996
rect 160974 68944 160980 68996
rect 161032 68984 161038 68996
rect 161728 68984 161756 69160
rect 168886 69148 168892 69160
rect 168944 69148 168950 69200
rect 192530 69148 192536 69200
rect 192588 69188 192594 69200
rect 194830 69188 194836 69200
rect 192588 69160 194836 69188
rect 192588 69148 192594 69160
rect 194830 69148 194836 69160
rect 194888 69148 194894 69200
rect 196946 69148 196952 69200
rect 197004 69188 197010 69200
rect 201086 69188 201092 69200
rect 197004 69160 201092 69188
rect 197004 69148 197010 69160
rect 201086 69148 201092 69160
rect 201144 69148 201150 69200
rect 192898 69080 192904 69132
rect 192956 69120 192962 69132
rect 195382 69120 195388 69132
rect 192956 69092 195388 69120
rect 192956 69080 192962 69092
rect 195382 69080 195388 69092
rect 195440 69080 195446 69132
rect 197406 69080 197412 69132
rect 197464 69120 197470 69132
rect 201822 69120 201828 69132
rect 197464 69092 201828 69120
rect 197464 69080 197470 69092
rect 201822 69080 201828 69092
rect 201880 69080 201886 69132
rect 167690 69012 167696 69064
rect 167748 69052 167754 69064
rect 174130 69052 174136 69064
rect 167748 69024 174136 69052
rect 167748 69012 167754 69024
rect 174130 69012 174136 69024
rect 174188 69012 174194 69064
rect 194094 69012 194100 69064
rect 194152 69052 194158 69064
rect 197130 69052 197136 69064
rect 194152 69024 197136 69052
rect 194152 69012 194158 69024
rect 197130 69012 197136 69024
rect 197188 69012 197194 69064
rect 197314 69012 197320 69064
rect 197372 69052 197378 69064
rect 201638 69052 201644 69064
rect 197372 69024 201644 69052
rect 197372 69012 197378 69024
rect 201638 69012 201644 69024
rect 201696 69012 201702 69064
rect 161032 68956 161756 68984
rect 161032 68944 161038 68956
rect 166586 68944 166592 68996
rect 166644 68984 166650 68996
rect 174222 68984 174228 68996
rect 166644 68956 174228 68984
rect 166644 68944 166650 68956
rect 174222 68944 174228 68956
rect 174280 68944 174286 68996
rect 181674 68944 181680 68996
rect 181732 68984 181738 68996
rect 182778 68984 182784 68996
rect 181732 68956 182784 68984
rect 181732 68944 181738 68956
rect 182778 68944 182784 68956
rect 182836 68944 182842 68996
rect 193358 68944 193364 68996
rect 193416 68984 193422 68996
rect 195934 68984 195940 68996
rect 193416 68956 195940 68984
rect 193416 68944 193422 68956
rect 195934 68944 195940 68956
rect 195992 68944 195998 68996
rect 198142 68944 198148 68996
rect 198200 68984 198206 68996
rect 202834 68984 202840 68996
rect 198200 68956 202840 68984
rect 198200 68944 198206 68956
rect 202834 68944 202840 68956
rect 202892 68944 202898 68996
rect 54180 68888 55128 68916
rect 38614 68808 38620 68860
rect 38672 68848 38678 68860
rect 41834 68848 41840 68860
rect 38672 68820 41840 68848
rect 38672 68808 38678 68820
rect 41834 68808 41840 68820
rect 41892 68808 41898 68860
rect 51034 68808 51040 68860
rect 51092 68848 51098 68860
rect 54254 68848 54260 68860
rect 51092 68820 54260 68848
rect 51092 68808 51098 68820
rect 54254 68808 54260 68820
rect 54312 68808 54318 68860
rect 37878 68740 37884 68792
rect 37936 68780 37942 68792
rect 41466 68780 41472 68792
rect 37936 68752 41472 68780
rect 37936 68740 37942 68752
rect 41466 68740 41472 68752
rect 41524 68740 41530 68792
rect 51402 68740 51408 68792
rect 51460 68780 51466 68792
rect 54990 68780 54996 68792
rect 51460 68752 54996 68780
rect 51460 68740 51466 68752
rect 54990 68740 54996 68752
rect 55048 68740 55054 68792
rect 55100 68780 55128 68888
rect 83418 68876 83424 68928
rect 83476 68916 83482 68928
rect 87190 68916 87196 68928
rect 83476 68888 87196 68916
rect 83476 68876 83482 68888
rect 87190 68876 87196 68888
rect 87248 68876 87254 68928
rect 87834 68876 87840 68928
rect 87892 68916 87898 68928
rect 94734 68916 94740 68928
rect 87892 68888 94740 68916
rect 87892 68876 87898 68888
rect 94734 68876 94740 68888
rect 94792 68876 94798 68928
rect 120494 68876 120500 68928
rect 120552 68916 120558 68928
rect 123070 68916 123076 68928
rect 120552 68888 123076 68916
rect 120552 68876 120558 68888
rect 123070 68876 123076 68888
rect 123128 68876 123134 68928
rect 124266 68876 124272 68928
rect 124324 68916 124330 68928
rect 128682 68916 128688 68928
rect 124324 68888 128688 68916
rect 124324 68876 124330 68888
rect 128682 68876 128688 68888
rect 128740 68876 128746 68928
rect 151038 68876 151044 68928
rect 151096 68916 151102 68928
rect 152050 68916 152056 68928
rect 151096 68888 152056 68916
rect 151096 68876 151102 68888
rect 152050 68876 152056 68888
rect 152108 68876 152114 68928
rect 159870 68876 159876 68928
rect 159928 68916 159934 68928
rect 159928 68888 165252 68916
rect 159928 68876 159934 68888
rect 55177 68851 55235 68857
rect 55177 68817 55189 68851
rect 55223 68848 55235 68851
rect 55634 68848 55640 68860
rect 55223 68820 55640 68848
rect 55223 68817 55235 68820
rect 55177 68811 55235 68817
rect 55634 68808 55640 68820
rect 55692 68808 55698 68860
rect 62718 68808 62724 68860
rect 62776 68848 62782 68860
rect 68974 68848 68980 68860
rect 62776 68820 68980 68848
rect 62776 68808 62782 68820
rect 68974 68808 68980 68820
rect 69032 68808 69038 68860
rect 82314 68808 82320 68860
rect 82372 68848 82378 68860
rect 85350 68848 85356 68860
rect 82372 68820 85356 68848
rect 82372 68808 82378 68820
rect 85350 68808 85356 68820
rect 85408 68808 85414 68860
rect 93446 68808 93452 68860
rect 93504 68848 93510 68860
rect 102554 68848 102560 68860
rect 93504 68820 102560 68848
rect 93504 68808 93510 68820
rect 102554 68808 102560 68820
rect 102612 68808 102618 68860
rect 110098 68808 110104 68860
rect 110156 68848 110162 68860
rect 111110 68848 111116 68860
rect 110156 68820 111116 68848
rect 110156 68808 110162 68820
rect 111110 68808 111116 68820
rect 111168 68808 111174 68860
rect 116262 68808 116268 68860
rect 116320 68848 116326 68860
rect 117090 68848 117096 68860
rect 116320 68820 117096 68848
rect 116320 68808 116326 68820
rect 117090 68808 117096 68820
rect 117148 68808 117154 68860
rect 117458 68808 117464 68860
rect 117516 68848 117522 68860
rect 118930 68848 118936 68860
rect 117516 68820 118936 68848
rect 117516 68808 117522 68820
rect 118930 68808 118936 68820
rect 118988 68808 118994 68860
rect 123346 68808 123352 68860
rect 123404 68848 123410 68860
rect 127302 68848 127308 68860
rect 123404 68820 127308 68848
rect 123404 68808 123410 68820
rect 127302 68808 127308 68820
rect 127360 68808 127366 68860
rect 140826 68808 140832 68860
rect 140884 68848 140890 68860
rect 144322 68848 144328 68860
rect 140884 68820 144328 68848
rect 140884 68808 140890 68820
rect 144322 68808 144328 68820
rect 144380 68808 144386 68860
rect 158766 68808 158772 68860
rect 158824 68848 158830 68860
rect 165114 68848 165120 68860
rect 158824 68820 165120 68848
rect 158824 68808 158830 68820
rect 165114 68808 165120 68820
rect 165172 68808 165178 68860
rect 165224 68848 165252 68888
rect 168794 68876 168800 68928
rect 168852 68916 168858 68928
rect 173854 68916 173860 68928
rect 168852 68888 173860 68916
rect 168852 68876 168858 68888
rect 173854 68876 173860 68888
rect 173912 68876 173918 68928
rect 193726 68876 193732 68928
rect 193784 68916 193790 68928
rect 196486 68916 196492 68928
rect 193784 68888 196492 68916
rect 193784 68876 193790 68888
rect 196486 68876 196492 68888
rect 196544 68876 196550 68928
rect 167046 68848 167052 68860
rect 165224 68820 167052 68848
rect 167046 68808 167052 68820
rect 167104 68808 167110 68860
rect 169898 68808 169904 68860
rect 169956 68848 169962 68860
rect 173946 68848 173952 68860
rect 169956 68820 173952 68848
rect 169956 68808 169962 68820
rect 173946 68808 173952 68820
rect 174004 68808 174010 68860
rect 195750 68808 195756 68860
rect 195808 68848 195814 68860
rect 199338 68848 199344 68860
rect 195808 68820 199344 68848
rect 195808 68808 195814 68820
rect 199338 68808 199344 68820
rect 199396 68808 199402 68860
rect 205134 68808 205140 68860
rect 205192 68848 205198 68860
rect 221234 68848 221240 68860
rect 205192 68820 221240 68848
rect 205192 68808 205198 68820
rect 221234 68808 221240 68820
rect 221292 68808 221298 68860
rect 56370 68780 56376 68792
rect 55100 68752 56376 68780
rect 56370 68740 56376 68752
rect 56428 68740 56434 68792
rect 120678 68740 120684 68792
rect 120736 68780 120742 68792
rect 123438 68780 123444 68792
rect 120736 68752 123444 68780
rect 120736 68740 120742 68752
rect 123438 68740 123444 68752
rect 123496 68740 123502 68792
rect 123809 68783 123867 68789
rect 123809 68749 123821 68783
rect 123855 68780 123867 68783
rect 132546 68780 132552 68792
rect 123855 68752 132552 68780
rect 123855 68749 123867 68752
rect 123809 68743 123867 68749
rect 132546 68740 132552 68752
rect 132604 68740 132610 68792
rect 165482 68740 165488 68792
rect 165540 68780 165546 68792
rect 174406 68780 174412 68792
rect 165540 68752 174412 68780
rect 165540 68740 165546 68752
rect 174406 68740 174412 68752
rect 174464 68740 174470 68792
rect 190598 68740 190604 68792
rect 190656 68780 190662 68792
rect 192530 68780 192536 68792
rect 190656 68752 192536 68780
rect 190656 68740 190662 68752
rect 192530 68740 192536 68752
rect 192588 68740 192594 68792
rect 195290 68740 195296 68792
rect 195348 68780 195354 68792
rect 198786 68780 198792 68792
rect 195348 68752 198792 68780
rect 195348 68740 195354 68752
rect 198786 68740 198792 68752
rect 198844 68740 198850 68792
rect 43398 68672 43404 68724
rect 43456 68712 43462 68724
rect 44594 68712 44600 68724
rect 43456 68684 44600 68712
rect 43456 68672 43462 68684
rect 44594 68672 44600 68684
rect 44652 68672 44658 68724
rect 50482 68672 50488 68724
rect 50540 68712 50546 68724
rect 52966 68712 52972 68724
rect 50540 68684 52972 68712
rect 50540 68672 50546 68684
rect 52966 68672 52972 68684
rect 53024 68672 53030 68724
rect 102278 68672 102284 68724
rect 102336 68712 102342 68724
rect 174314 68712 174320 68724
rect 102336 68684 174320 68712
rect 102336 68672 102342 68684
rect 174314 68672 174320 68684
rect 174372 68672 174378 68724
rect 36133 68647 36191 68653
rect 36133 68613 36145 68647
rect 36179 68644 36191 68647
rect 54809 68647 54867 68653
rect 54809 68644 54821 68647
rect 36179 68616 54821 68644
rect 36179 68613 36191 68616
rect 36133 68607 36191 68613
rect 54809 68613 54821 68616
rect 54855 68613 54867 68647
rect 54809 68607 54867 68613
rect 101174 68604 101180 68656
rect 101232 68644 101238 68656
rect 173210 68644 173216 68656
rect 101232 68616 173216 68644
rect 101232 68604 101238 68616
rect 173210 68604 173216 68616
rect 173268 68604 173274 68656
rect 194646 68604 194652 68656
rect 194704 68644 194710 68656
rect 198234 68644 198240 68656
rect 194704 68616 198240 68644
rect 194704 68604 194710 68616
rect 198234 68604 198240 68616
rect 198292 68604 198298 68656
rect 90134 68536 90140 68588
rect 90192 68576 90198 68588
rect 123809 68579 123867 68585
rect 123809 68576 123821 68579
rect 90192 68548 123821 68576
rect 90192 68536 90198 68548
rect 123809 68545 123821 68548
rect 123855 68545 123867 68579
rect 123809 68539 123867 68545
rect 123898 68536 123904 68588
rect 123956 68576 123962 68588
rect 128130 68576 128136 68588
rect 123956 68548 128136 68576
rect 123956 68536 123962 68548
rect 128130 68536 128136 68548
rect 128188 68536 128194 68588
rect 182226 68536 182232 68588
rect 182284 68576 182290 68588
rect 183238 68576 183244 68588
rect 182284 68548 183244 68576
rect 182284 68536 182290 68548
rect 183238 68536 183244 68548
rect 183296 68536 183302 68588
rect 97862 68468 97868 68520
rect 97920 68508 97926 68520
rect 102370 68508 102376 68520
rect 97920 68480 102376 68508
rect 97920 68468 97926 68480
rect 102370 68468 102376 68480
rect 102428 68468 102434 68520
rect 121506 68468 121512 68520
rect 121564 68508 121570 68520
rect 124634 68508 124640 68520
rect 121564 68480 124640 68508
rect 121564 68468 121570 68480
rect 124634 68468 124640 68480
rect 124692 68468 124698 68520
rect 74586 68400 74592 68452
rect 74644 68440 74650 68452
rect 75598 68440 75604 68452
rect 74644 68412 75604 68440
rect 74644 68400 74650 68412
rect 75598 68400 75604 68412
rect 75656 68400 75662 68452
rect 94550 68400 94556 68452
rect 94608 68440 94614 68452
rect 102646 68440 102652 68452
rect 94608 68412 102652 68440
rect 94608 68400 94614 68412
rect 102646 68400 102652 68412
rect 102704 68400 102710 68452
rect 86730 68332 86736 68384
rect 86788 68372 86794 68384
rect 92802 68372 92808 68384
rect 86788 68344 92808 68372
rect 86788 68332 86794 68344
rect 92802 68332 92808 68344
rect 92860 68332 92866 68384
rect 95654 68332 95660 68384
rect 95712 68372 95718 68384
rect 102738 68372 102744 68384
rect 95712 68344 102744 68372
rect 95712 68332 95718 68344
rect 102738 68332 102744 68344
rect 102796 68332 102802 68384
rect 155454 68332 155460 68384
rect 155512 68372 155518 68384
rect 159502 68372 159508 68384
rect 155512 68344 159508 68372
rect 155512 68332 155518 68344
rect 159502 68332 159508 68344
rect 159560 68332 159566 68384
rect 62994 68264 63000 68316
rect 63052 68304 63058 68316
rect 64558 68304 64564 68316
rect 63052 68276 64564 68304
rect 63052 68264 63058 68276
rect 64558 68264 64564 68276
rect 64616 68264 64622 68316
rect 70998 68264 71004 68316
rect 71056 68304 71062 68316
rect 73390 68304 73396 68316
rect 71056 68276 73396 68304
rect 71056 68264 71062 68276
rect 73390 68264 73396 68276
rect 73448 68264 73454 68316
rect 81210 68264 81216 68316
rect 81268 68304 81274 68316
rect 83510 68304 83516 68316
rect 81268 68276 83516 68304
rect 81268 68264 81274 68276
rect 83510 68264 83516 68276
rect 83568 68264 83574 68316
rect 85626 68264 85632 68316
rect 85684 68304 85690 68316
rect 90962 68304 90968 68316
rect 85684 68276 90968 68304
rect 85684 68264 85690 68276
rect 90962 68264 90968 68276
rect 91020 68264 91026 68316
rect 96758 68264 96764 68316
rect 96816 68304 96822 68316
rect 102462 68304 102468 68316
rect 96816 68276 102468 68304
rect 96816 68264 96822 68276
rect 102462 68264 102468 68276
rect 102520 68264 102526 68316
rect 144506 68264 144512 68316
rect 144564 68304 144570 68316
rect 146530 68304 146536 68316
rect 144564 68276 146536 68304
rect 144564 68264 144570 68276
rect 146530 68264 146536 68276
rect 146588 68264 146594 68316
rect 153246 68264 153252 68316
rect 153304 68304 153310 68316
rect 155822 68304 155828 68316
rect 153304 68276 155828 68304
rect 153304 68264 153310 68276
rect 155822 68264 155828 68276
rect 155880 68264 155886 68316
rect 156558 68264 156564 68316
rect 156616 68304 156622 68316
rect 161434 68304 161440 68316
rect 156616 68276 161440 68304
rect 156616 68264 156622 68276
rect 161434 68264 161440 68276
rect 161492 68264 161498 68316
rect 163274 68304 163280 68316
rect 161636 68276 163280 68304
rect 62350 68196 62356 68248
rect 62408 68236 62414 68248
rect 63454 68236 63460 68248
rect 62408 68208 63460 68236
rect 62408 68196 62414 68208
rect 63454 68196 63460 68208
rect 63512 68196 63518 68248
rect 69158 68196 69164 68248
rect 69216 68236 69222 68248
rect 72286 68236 72292 68248
rect 69216 68208 72292 68236
rect 69216 68196 69222 68208
rect 72286 68196 72292 68208
rect 72344 68196 72350 68248
rect 72838 68196 72844 68248
rect 72896 68236 72902 68248
rect 74494 68236 74500 68248
rect 72896 68208 74500 68236
rect 72896 68196 72902 68208
rect 74494 68196 74500 68208
rect 74552 68196 74558 68248
rect 80106 68196 80112 68248
rect 80164 68236 80170 68248
rect 81670 68236 81676 68248
rect 80164 68208 81676 68236
rect 80164 68196 80170 68208
rect 81670 68196 81676 68208
rect 81728 68196 81734 68248
rect 84522 68196 84528 68248
rect 84580 68236 84586 68248
rect 89122 68236 89128 68248
rect 84580 68208 89128 68236
rect 84580 68196 84586 68208
rect 89122 68196 89128 68208
rect 89180 68196 89186 68248
rect 98966 68196 98972 68248
rect 99024 68236 99030 68248
rect 99024 68208 100944 68236
rect 99024 68196 99030 68208
rect 63362 68128 63368 68180
rect 63420 68168 63426 68180
rect 71182 68168 71188 68180
rect 63420 68140 71188 68168
rect 63420 68128 63426 68140
rect 71182 68128 71188 68140
rect 71240 68128 71246 68180
rect 100916 68168 100944 68208
rect 134478 68196 134484 68248
rect 134536 68236 134542 68248
rect 136594 68236 136600 68248
rect 134536 68208 136600 68236
rect 134536 68196 134542 68208
rect 136594 68196 136600 68208
rect 136652 68196 136658 68248
rect 142666 68196 142672 68248
rect 142724 68236 142730 68248
rect 145426 68236 145432 68248
rect 142724 68208 145432 68236
rect 142724 68196 142730 68208
rect 145426 68196 145432 68208
rect 145484 68196 145490 68248
rect 146438 68196 146444 68248
rect 146496 68236 146502 68248
rect 147634 68236 147640 68248
rect 146496 68208 147640 68236
rect 146496 68196 146502 68208
rect 147634 68196 147640 68208
rect 147692 68196 147698 68248
rect 152142 68196 152148 68248
rect 152200 68236 152206 68248
rect 153890 68236 153896 68248
rect 152200 68208 153896 68236
rect 152200 68196 152206 68208
rect 153890 68196 153896 68208
rect 153948 68196 153954 68248
rect 154350 68196 154356 68248
rect 154408 68236 154414 68248
rect 157662 68236 157668 68248
rect 154408 68208 157668 68236
rect 154408 68196 154414 68208
rect 157662 68196 157668 68208
rect 157720 68196 157726 68248
rect 157938 68196 157944 68248
rect 157996 68236 158002 68248
rect 161636 68236 161664 68276
rect 163274 68264 163280 68276
rect 163332 68264 163338 68316
rect 171002 68264 171008 68316
rect 171060 68304 171066 68316
rect 174038 68304 174044 68316
rect 171060 68276 174044 68304
rect 171060 68264 171066 68276
rect 174038 68264 174044 68276
rect 174096 68264 174102 68316
rect 157996 68208 161664 68236
rect 157996 68196 158002 68208
rect 164378 68196 164384 68248
rect 164436 68236 164442 68248
rect 169438 68236 169444 68248
rect 164436 68208 169444 68236
rect 164436 68196 164442 68208
rect 169438 68196 169444 68208
rect 169496 68196 169502 68248
rect 172106 68196 172112 68248
rect 172164 68236 172170 68248
rect 172164 68208 174084 68236
rect 172164 68196 172170 68208
rect 102922 68168 102928 68180
rect 100916 68140 102928 68168
rect 102922 68128 102928 68140
rect 102980 68128 102986 68180
rect 135306 68128 135312 68180
rect 135364 68168 135370 68180
rect 143218 68168 143224 68180
rect 135364 68140 143224 68168
rect 135364 68128 135370 68140
rect 143218 68128 143224 68140
rect 143276 68128 143282 68180
rect 174056 68168 174084 68208
rect 175050 68168 175056 68180
rect 174056 68140 175056 68168
rect 175050 68128 175056 68140
rect 175108 68128 175114 68180
rect 135030 68060 135036 68112
rect 135088 68100 135094 68112
rect 142114 68100 142120 68112
rect 135088 68072 142120 68100
rect 135088 68060 135094 68072
rect 142114 68060 142120 68072
rect 142172 68060 142178 68112
rect 100070 67652 100076 67704
rect 100128 67692 100134 67704
rect 103474 67692 103480 67704
rect 100128 67664 103480 67692
rect 100128 67652 100134 67664
rect 103474 67652 103480 67664
rect 103532 67652 103538 67704
rect 62810 66700 62816 66752
rect 62868 66740 62874 66752
rect 70078 66740 70084 66752
rect 62868 66712 70084 66740
rect 62868 66700 62874 66712
rect 70078 66700 70084 66712
rect 70136 66700 70142 66752
rect 134662 66700 134668 66752
rect 134720 66740 134726 66752
rect 139906 66740 139912 66752
rect 134720 66712 139912 66740
rect 134720 66700 134726 66712
rect 139906 66700 139912 66712
rect 139964 66700 139970 66752
rect 135306 66428 135312 66480
rect 135364 66468 135370 66480
rect 141010 66468 141016 66480
rect 135364 66440 141016 66468
rect 135364 66428 135370 66440
rect 141010 66428 141016 66440
rect 141068 66428 141074 66480
rect 63362 65544 63368 65596
rect 63420 65584 63426 65596
rect 66398 65584 66404 65596
rect 63420 65556 66404 65584
rect 63420 65544 63426 65556
rect 66398 65544 66404 65556
rect 66456 65544 66462 65596
rect 172658 65544 172664 65596
rect 172716 65584 172722 65596
rect 175326 65584 175332 65596
rect 172716 65556 175332 65584
rect 172716 65544 172722 65556
rect 175326 65544 175332 65556
rect 175384 65544 175390 65596
rect 100898 65408 100904 65460
rect 100956 65448 100962 65460
rect 102370 65448 102376 65460
rect 100956 65420 102376 65448
rect 100956 65408 100962 65420
rect 102370 65408 102376 65420
rect 102428 65408 102434 65460
rect 134662 65408 134668 65460
rect 134720 65448 134726 65460
rect 136870 65448 136876 65460
rect 134720 65420 136876 65448
rect 134720 65408 134726 65420
rect 136870 65408 136876 65420
rect 136928 65408 136934 65460
rect 62810 65340 62816 65392
rect 62868 65380 62874 65392
rect 66306 65380 66312 65392
rect 62868 65352 66312 65380
rect 62868 65340 62874 65352
rect 66306 65340 66312 65352
rect 66364 65340 66370 65392
rect 134846 65340 134852 65392
rect 134904 65380 134910 65392
rect 137698 65380 137704 65392
rect 134904 65352 137704 65380
rect 134904 65340 134910 65352
rect 137698 65340 137704 65352
rect 137756 65340 137762 65392
rect 62718 65272 62724 65324
rect 62776 65312 62782 65324
rect 65662 65312 65668 65324
rect 62776 65284 65668 65312
rect 62776 65272 62782 65284
rect 65662 65272 65668 65284
rect 65720 65272 65726 65324
rect 135306 65204 135312 65256
rect 135364 65244 135370 65256
rect 138158 65244 138164 65256
rect 135364 65216 138164 65244
rect 135364 65204 135370 65216
rect 138158 65204 138164 65216
rect 138216 65204 138222 65256
rect 100622 64456 100628 64508
rect 100680 64496 100686 64508
rect 102738 64496 102744 64508
rect 100680 64468 102744 64496
rect 100680 64456 100686 64468
rect 102738 64456 102744 64468
rect 102796 64456 102802 64508
rect 63546 64320 63552 64372
rect 63604 64360 63610 64372
rect 66398 64360 66404 64372
rect 63604 64332 66404 64360
rect 63604 64320 63610 64332
rect 66398 64320 66404 64332
rect 66456 64320 66462 64372
rect 172658 64320 172664 64372
rect 172716 64360 172722 64372
rect 174222 64360 174228 64372
rect 172716 64332 174228 64360
rect 172716 64320 172722 64332
rect 174222 64320 174228 64332
rect 174280 64320 174286 64372
rect 63454 64184 63460 64236
rect 63512 64224 63518 64236
rect 65662 64224 65668 64236
rect 63512 64196 65668 64224
rect 63512 64184 63518 64196
rect 65662 64184 65668 64196
rect 65720 64184 65726 64236
rect 135306 64116 135312 64168
rect 135364 64156 135370 64168
rect 136962 64156 136968 64168
rect 135364 64128 136968 64156
rect 135364 64116 135370 64128
rect 136962 64116 136968 64128
rect 137020 64116 137026 64168
rect 100898 64048 100904 64100
rect 100956 64088 100962 64100
rect 102462 64088 102468 64100
rect 100956 64060 102468 64088
rect 100956 64048 100962 64060
rect 102462 64048 102468 64060
rect 102520 64048 102526 64100
rect 134846 64048 134852 64100
rect 134904 64088 134910 64100
rect 136870 64088 136876 64100
rect 134904 64060 136876 64088
rect 134904 64048 134910 64060
rect 136870 64048 136876 64060
rect 136928 64048 136934 64100
rect 171830 64048 171836 64100
rect 171888 64088 171894 64100
rect 175234 64088 175240 64100
rect 171888 64060 175240 64088
rect 171888 64048 171894 64060
rect 175234 64048 175240 64060
rect 175292 64048 175298 64100
rect 169438 63980 169444 64032
rect 169496 64020 169502 64032
rect 174130 64020 174136 64032
rect 169496 63992 174136 64020
rect 169496 63980 169502 63992
rect 174130 63980 174136 63992
rect 174188 63980 174194 64032
rect 97494 63776 97500 63828
rect 97552 63816 97558 63828
rect 102554 63816 102560 63828
rect 97552 63788 102560 63816
rect 97552 63776 97558 63788
rect 102554 63776 102560 63788
rect 102612 63776 102618 63828
rect 172658 62960 172664 63012
rect 172716 63000 172722 63012
rect 174130 63000 174136 63012
rect 172716 62972 174136 63000
rect 172716 62960 172722 62972
rect 174130 62960 174136 62972
rect 174188 62960 174194 63012
rect 100622 62824 100628 62876
rect 100680 62864 100686 62876
rect 102370 62864 102376 62876
rect 100680 62836 102376 62864
rect 100680 62824 100686 62836
rect 102370 62824 102376 62836
rect 102428 62824 102434 62876
rect 62718 62688 62724 62740
rect 62776 62728 62782 62740
rect 65662 62728 65668 62740
rect 62776 62700 65668 62728
rect 62776 62688 62782 62700
rect 65662 62688 65668 62700
rect 65720 62688 65726 62740
rect 100622 62688 100628 62740
rect 100680 62728 100686 62740
rect 102554 62728 102560 62740
rect 100680 62700 102560 62728
rect 100680 62688 100686 62700
rect 102554 62688 102560 62700
rect 102612 62688 102618 62740
rect 134478 62688 134484 62740
rect 134536 62728 134542 62740
rect 136962 62728 136968 62740
rect 134536 62700 136968 62728
rect 134536 62688 134542 62700
rect 136962 62688 136968 62700
rect 137020 62688 137026 62740
rect 172658 62688 172664 62740
rect 172716 62728 172722 62740
rect 174314 62728 174320 62740
rect 172716 62700 174320 62728
rect 172716 62688 172722 62700
rect 174314 62688 174320 62700
rect 174372 62688 174378 62740
rect 13314 62620 13320 62672
rect 13372 62660 13378 62672
rect 29230 62660 29236 62672
rect 13372 62632 29236 62660
rect 13372 62620 13378 62632
rect 29230 62620 29236 62632
rect 29288 62620 29294 62672
rect 62810 62620 62816 62672
rect 62868 62660 62874 62672
rect 66398 62660 66404 62672
rect 62868 62632 66404 62660
rect 62868 62620 62874 62632
rect 66398 62620 66404 62632
rect 66456 62620 66462 62672
rect 135398 62620 135404 62672
rect 135456 62660 135462 62672
rect 136870 62660 136876 62672
rect 135456 62632 136876 62660
rect 135456 62620 135462 62632
rect 136870 62620 136876 62632
rect 136928 62620 136934 62672
rect 62902 61464 62908 61516
rect 62960 61504 62966 61516
rect 65662 61504 65668 61516
rect 62960 61476 65668 61504
rect 62960 61464 62966 61476
rect 65662 61464 65668 61476
rect 65720 61464 65726 61516
rect 172658 61464 172664 61516
rect 172716 61504 172722 61516
rect 174222 61504 174228 61516
rect 172716 61476 174228 61504
rect 172716 61464 172722 61476
rect 174222 61464 174228 61476
rect 174280 61464 174286 61516
rect 100622 61328 100628 61380
rect 100680 61368 100686 61380
rect 102462 61368 102468 61380
rect 100680 61340 102468 61368
rect 100680 61328 100686 61340
rect 102462 61328 102468 61340
rect 102520 61328 102526 61380
rect 63730 61260 63736 61312
rect 63788 61300 63794 61312
rect 66398 61300 66404 61312
rect 63788 61272 66404 61300
rect 63788 61260 63794 61272
rect 66398 61260 66404 61272
rect 66456 61260 66462 61312
rect 100530 61260 100536 61312
rect 100588 61300 100594 61312
rect 102738 61300 102744 61312
rect 100588 61272 102744 61300
rect 100588 61260 100594 61272
rect 102738 61260 102744 61272
rect 102796 61260 102802 61312
rect 135306 61260 135312 61312
rect 135364 61300 135370 61312
rect 136870 61300 136876 61312
rect 135364 61272 136876 61300
rect 135364 61260 135370 61272
rect 136870 61260 136876 61272
rect 136928 61260 136934 61312
rect 171830 61260 171836 61312
rect 171888 61300 171894 61312
rect 174406 61300 174412 61312
rect 171888 61272 174412 61300
rect 171888 61260 171894 61272
rect 174406 61260 174412 61272
rect 174464 61260 174470 61312
rect 135030 60920 135036 60972
rect 135088 60960 135094 60972
rect 136778 60960 136784 60972
rect 135088 60932 136784 60960
rect 135088 60920 135094 60932
rect 136778 60920 136784 60932
rect 136836 60920 136842 60972
rect 63822 60580 63828 60632
rect 63880 60620 63886 60632
rect 65478 60620 65484 60632
rect 63880 60592 65484 60620
rect 63880 60580 63886 60592
rect 65478 60580 65484 60592
rect 65536 60580 65542 60632
rect 100622 60376 100628 60428
rect 100680 60416 100686 60428
rect 102646 60416 102652 60428
rect 100680 60388 102652 60416
rect 100680 60376 100686 60388
rect 102646 60376 102652 60388
rect 102704 60376 102710 60428
rect 100622 60240 100628 60292
rect 100680 60280 100686 60292
rect 102370 60280 102376 60292
rect 100680 60252 102376 60280
rect 100680 60240 100686 60252
rect 102370 60240 102376 60252
rect 102428 60240 102434 60292
rect 172658 60240 172664 60292
rect 172716 60280 172722 60292
rect 174314 60280 174320 60292
rect 172716 60252 174320 60280
rect 172716 60240 172722 60252
rect 174314 60240 174320 60252
rect 174372 60240 174378 60292
rect 62626 60104 62632 60156
rect 62684 60144 62690 60156
rect 66398 60144 66404 60156
rect 62684 60116 66404 60144
rect 62684 60104 62690 60116
rect 66398 60104 66404 60116
rect 66456 60104 66462 60156
rect 172198 60104 172204 60156
rect 172256 60144 172262 60156
rect 174130 60144 174136 60156
rect 172256 60116 174136 60144
rect 172256 60104 172262 60116
rect 174130 60104 174136 60116
rect 174188 60104 174194 60156
rect 134478 60036 134484 60088
rect 134536 60076 134542 60088
rect 136962 60076 136968 60088
rect 134536 60048 136968 60076
rect 134536 60036 134542 60048
rect 136962 60036 136968 60048
rect 137020 60036 137026 60088
rect 100622 59968 100628 60020
rect 100680 60008 100686 60020
rect 102554 60008 102560 60020
rect 100680 59980 102560 60008
rect 100680 59968 100686 59980
rect 102554 59968 102560 59980
rect 102612 59968 102618 60020
rect 172658 59968 172664 60020
rect 172716 60008 172722 60020
rect 174498 60008 174504 60020
rect 172716 59980 174504 60008
rect 172716 59968 172722 59980
rect 174498 59968 174504 59980
rect 174556 59968 174562 60020
rect 62718 59900 62724 59952
rect 62776 59940 62782 59952
rect 66306 59940 66312 59952
rect 62776 59912 66312 59940
rect 62776 59900 62782 59912
rect 66306 59900 66312 59912
rect 66364 59900 66370 59952
rect 135398 59900 135404 59952
rect 135456 59940 135462 59952
rect 136870 59940 136876 59952
rect 135456 59912 136876 59940
rect 135456 59900 135462 59912
rect 136870 59900 136876 59912
rect 136928 59900 136934 59952
rect 135030 59832 135036 59884
rect 135088 59872 135094 59884
rect 136778 59872 136784 59884
rect 135088 59844 136784 59872
rect 135088 59832 135094 59844
rect 136778 59832 136784 59844
rect 136836 59832 136842 59884
rect 172198 58880 172204 58932
rect 172256 58920 172262 58932
rect 174590 58920 174596 58932
rect 172256 58892 174596 58920
rect 172256 58880 172262 58892
rect 174590 58880 174596 58892
rect 174648 58880 174654 58932
rect 100622 58744 100628 58796
rect 100680 58784 100686 58796
rect 102462 58784 102468 58796
rect 100680 58756 102468 58784
rect 100680 58744 100686 58756
rect 102462 58744 102468 58756
rect 102520 58744 102526 58796
rect 171830 58744 171836 58796
rect 171888 58784 171894 58796
rect 174222 58784 174228 58796
rect 171888 58756 174228 58784
rect 171888 58744 171894 58756
rect 174222 58744 174228 58756
rect 174280 58744 174286 58796
rect 62810 58608 62816 58660
rect 62868 58648 62874 58660
rect 66306 58648 66312 58660
rect 62868 58620 66312 58648
rect 62868 58608 62874 58620
rect 66306 58608 66312 58620
rect 66364 58608 66370 58660
rect 100622 58608 100628 58660
rect 100680 58648 100686 58660
rect 102646 58648 102652 58660
rect 100680 58620 102652 58648
rect 100680 58608 100686 58620
rect 102646 58608 102652 58620
rect 102704 58608 102710 58660
rect 62902 58540 62908 58592
rect 62960 58580 62966 58592
rect 66398 58580 66404 58592
rect 62960 58552 66404 58580
rect 62960 58540 62966 58552
rect 66398 58540 66404 58552
rect 66456 58540 66462 58592
rect 135306 58540 135312 58592
rect 135364 58580 135370 58592
rect 136870 58580 136876 58592
rect 135364 58552 136876 58580
rect 135364 58540 135370 58552
rect 136870 58540 136876 58552
rect 136928 58540 136934 58592
rect 135030 58404 135036 58456
rect 135088 58444 135094 58456
rect 136778 58444 136784 58456
rect 135088 58416 136784 58444
rect 135088 58404 135094 58416
rect 136778 58404 136784 58416
rect 136836 58404 136842 58456
rect 62718 57384 62724 57436
rect 62776 57424 62782 57436
rect 66398 57424 66404 57436
rect 62776 57396 66404 57424
rect 62776 57384 62782 57396
rect 66398 57384 66404 57396
rect 66456 57384 66462 57436
rect 100622 57384 100628 57436
rect 100680 57424 100686 57436
rect 102370 57424 102376 57436
rect 100680 57396 102376 57424
rect 100680 57384 100686 57396
rect 102370 57384 102376 57396
rect 102428 57384 102434 57436
rect 172658 57384 172664 57436
rect 172716 57424 172722 57436
rect 174314 57424 174320 57436
rect 172716 57396 174320 57424
rect 172716 57384 172722 57396
rect 174314 57384 174320 57396
rect 174372 57384 174378 57436
rect 172658 57248 172664 57300
rect 172716 57288 172722 57300
rect 174406 57288 174412 57300
rect 172716 57260 174412 57288
rect 172716 57248 172722 57260
rect 174406 57248 174412 57260
rect 174464 57248 174470 57300
rect 100622 57180 100628 57232
rect 100680 57220 100686 57232
rect 102462 57220 102468 57232
rect 100680 57192 102468 57220
rect 100680 57180 100686 57192
rect 102462 57180 102468 57192
rect 102520 57180 102526 57232
rect 135398 57180 135404 57232
rect 135456 57220 135462 57232
rect 136962 57220 136968 57232
rect 135456 57192 136968 57220
rect 135456 57180 135462 57192
rect 136962 57180 136968 57192
rect 137020 57180 137026 57232
rect 62626 57112 62632 57164
rect 62684 57152 62690 57164
rect 66398 57152 66404 57164
rect 62684 57124 66404 57152
rect 62684 57112 62690 57124
rect 66398 57112 66404 57124
rect 66456 57112 66462 57164
rect 100530 57112 100536 57164
rect 100588 57152 100594 57164
rect 102554 57152 102560 57164
rect 100588 57124 102560 57152
rect 100588 57112 100594 57124
rect 102554 57112 102560 57124
rect 102612 57112 102618 57164
rect 134754 57112 134760 57164
rect 134812 57152 134818 57164
rect 136870 57152 136876 57164
rect 134812 57124 136876 57152
rect 134812 57112 134818 57124
rect 136870 57112 136876 57124
rect 136928 57112 136934 57164
rect 172014 57112 172020 57164
rect 172072 57152 172078 57164
rect 174130 57152 174136 57164
rect 172072 57124 174136 57152
rect 172072 57112 172078 57124
rect 174130 57112 174136 57124
rect 174188 57112 174194 57164
rect 135030 57044 135036 57096
rect 135088 57084 135094 57096
rect 136778 57084 136784 57096
rect 135088 57056 136784 57084
rect 135088 57044 135094 57056
rect 136778 57044 136784 57056
rect 136836 57044 136842 57096
rect 62534 56976 62540 57028
rect 62592 57016 62598 57028
rect 65018 57016 65024 57028
rect 62592 56988 65024 57016
rect 62592 56976 62598 56988
rect 65018 56976 65024 56988
rect 65076 56976 65082 57028
rect 63638 56296 63644 56348
rect 63696 56336 63702 56348
rect 66398 56336 66404 56348
rect 63696 56308 66404 56336
rect 63696 56296 63702 56308
rect 66398 56296 66404 56308
rect 66456 56296 66462 56348
rect 172658 56024 172664 56076
rect 172716 56064 172722 56076
rect 174222 56064 174228 56076
rect 172716 56036 174228 56064
rect 172716 56024 172722 56036
rect 174222 56024 174228 56036
rect 174280 56024 174286 56076
rect 63270 55888 63276 55940
rect 63328 55928 63334 55940
rect 66398 55928 66404 55940
rect 63328 55900 66404 55928
rect 63328 55888 63334 55900
rect 66398 55888 66404 55900
rect 66456 55888 66462 55940
rect 100622 55888 100628 55940
rect 100680 55928 100686 55940
rect 102370 55928 102376 55940
rect 100680 55900 102376 55928
rect 100680 55888 100686 55900
rect 102370 55888 102376 55900
rect 102428 55888 102434 55940
rect 100898 55752 100904 55804
rect 100956 55792 100962 55804
rect 102646 55792 102652 55804
rect 100956 55764 102652 55792
rect 100956 55752 100962 55764
rect 102646 55752 102652 55764
rect 102704 55752 102710 55804
rect 134202 55752 134208 55804
rect 134260 55792 134266 55804
rect 136870 55792 136876 55804
rect 134260 55764 136876 55792
rect 134260 55752 134266 55764
rect 136870 55752 136876 55764
rect 136928 55752 136934 55804
rect 172658 55752 172664 55804
rect 172716 55792 172722 55804
rect 174958 55792 174964 55804
rect 172716 55764 174964 55792
rect 172716 55752 172722 55764
rect 174958 55752 174964 55764
rect 175016 55752 175022 55804
rect 135030 55412 135036 55464
rect 135088 55452 135094 55464
rect 136778 55452 136784 55464
rect 135088 55424 136784 55452
rect 135088 55412 135094 55424
rect 136778 55412 136784 55424
rect 136836 55412 136842 55464
rect 100622 54800 100628 54852
rect 100680 54840 100686 54852
rect 102462 54840 102468 54852
rect 100680 54812 102468 54840
rect 100680 54800 100686 54812
rect 102462 54800 102468 54812
rect 102520 54800 102526 54852
rect 63362 54664 63368 54716
rect 63420 54704 63426 54716
rect 66398 54704 66404 54716
rect 63420 54676 66404 54704
rect 63420 54664 63426 54676
rect 66398 54664 66404 54676
rect 66456 54664 66462 54716
rect 100806 54528 100812 54580
rect 100864 54568 100870 54580
rect 102554 54568 102560 54580
rect 100864 54540 102560 54568
rect 100864 54528 100870 54540
rect 102554 54528 102560 54540
rect 102612 54528 102618 54580
rect 134294 54528 134300 54580
rect 134352 54568 134358 54580
rect 137146 54568 137152 54580
rect 134352 54540 137152 54568
rect 134352 54528 134358 54540
rect 137146 54528 137152 54540
rect 137204 54528 137210 54580
rect 172106 54528 172112 54580
rect 172164 54568 172170 54580
rect 174774 54568 174780 54580
rect 172164 54540 174780 54568
rect 172164 54528 172170 54540
rect 174774 54528 174780 54540
rect 174832 54528 174838 54580
rect 172658 54460 172664 54512
rect 172716 54500 172722 54512
rect 175326 54500 175332 54512
rect 172716 54472 175332 54500
rect 172716 54460 172722 54472
rect 175326 54460 175332 54472
rect 175384 54460 175390 54512
rect 63546 54392 63552 54444
rect 63604 54432 63610 54444
rect 66306 54432 66312 54444
rect 63604 54404 66312 54432
rect 63604 54392 63610 54404
rect 66306 54392 66312 54404
rect 66364 54392 66370 54444
rect 135122 53916 135128 53968
rect 135180 53956 135186 53968
rect 136778 53956 136784 53968
rect 135180 53928 136784 53956
rect 135180 53916 135186 53928
rect 136778 53916 136784 53928
rect 136836 53916 136842 53968
rect 62810 53304 62816 53356
rect 62868 53344 62874 53356
rect 65294 53344 65300 53356
rect 62868 53316 65300 53344
rect 62868 53304 62874 53316
rect 65294 53304 65300 53316
rect 65352 53304 65358 53356
rect 100622 53236 100628 53288
rect 100680 53276 100686 53288
rect 102738 53276 102744 53288
rect 100680 53248 102744 53276
rect 100680 53236 100686 53248
rect 102738 53236 102744 53248
rect 102796 53236 102802 53288
rect 171646 53168 171652 53220
rect 171704 53208 171710 53220
rect 174130 53208 174136 53220
rect 171704 53180 174136 53208
rect 171704 53168 171710 53180
rect 174130 53168 174136 53180
rect 174188 53168 174194 53220
rect 100622 53032 100628 53084
rect 100680 53072 100686 53084
rect 102370 53072 102376 53084
rect 100680 53044 102376 53072
rect 100680 53032 100686 53044
rect 102370 53032 102376 53044
rect 102428 53032 102434 53084
rect 172658 53032 172664 53084
rect 172716 53072 172722 53084
rect 174498 53072 174504 53084
rect 172716 53044 174504 53072
rect 172716 53032 172722 53044
rect 174498 53032 174504 53044
rect 174556 53032 174562 53084
rect 63730 52964 63736 53016
rect 63788 53004 63794 53016
rect 66398 53004 66404 53016
rect 63788 52976 66404 53004
rect 63788 52964 63794 52976
rect 66398 52964 66404 52976
rect 66456 52964 66462 53016
rect 135398 52964 135404 53016
rect 135456 53004 135462 53016
rect 136870 53004 136876 53016
rect 135456 52976 136876 53004
rect 135456 52964 135462 52976
rect 136870 52964 136876 52976
rect 136928 52964 136934 53016
rect 135122 52556 135128 52608
rect 135180 52596 135186 52608
rect 136778 52596 136784 52608
rect 135180 52568 136784 52596
rect 135180 52556 135186 52568
rect 136778 52556 136784 52568
rect 136836 52556 136842 52608
rect 100622 52216 100628 52268
rect 100680 52256 100686 52268
rect 102646 52256 102652 52268
rect 100680 52228 102652 52256
rect 100680 52216 100686 52228
rect 102646 52216 102652 52228
rect 102704 52216 102710 52268
rect 63362 52080 63368 52132
rect 63420 52120 63426 52132
rect 65294 52120 65300 52132
rect 63420 52092 65300 52120
rect 63420 52080 63426 52092
rect 65294 52080 65300 52092
rect 65352 52080 65358 52132
rect 172566 51944 172572 51996
rect 172624 51984 172630 51996
rect 174314 51984 174320 51996
rect 172624 51956 174320 51984
rect 172624 51944 172630 51956
rect 174314 51944 174320 51956
rect 174372 51944 174378 51996
rect 172658 51808 172664 51860
rect 172716 51848 172722 51860
rect 174406 51848 174412 51860
rect 172716 51820 174412 51848
rect 172716 51808 172722 51820
rect 174406 51808 174412 51820
rect 174464 51808 174470 51860
rect 62718 51672 62724 51724
rect 62776 51712 62782 51724
rect 65662 51712 65668 51724
rect 62776 51684 65668 51712
rect 62776 51672 62782 51684
rect 65662 51672 65668 51684
rect 65720 51672 65726 51724
rect 100622 51672 100628 51724
rect 100680 51712 100686 51724
rect 102462 51712 102468 51724
rect 100680 51684 102468 51712
rect 100680 51672 100686 51684
rect 102462 51672 102468 51684
rect 102520 51672 102526 51724
rect 63730 51604 63736 51656
rect 63788 51644 63794 51656
rect 66306 51644 66312 51656
rect 63788 51616 66312 51644
rect 63788 51604 63794 51616
rect 66306 51604 66312 51616
rect 66364 51604 66370 51656
rect 100530 51604 100536 51656
rect 100588 51644 100594 51656
rect 102554 51644 102560 51656
rect 100588 51616 102560 51644
rect 100588 51604 100594 51616
rect 102554 51604 102560 51616
rect 102612 51604 102618 51656
rect 135306 51604 135312 51656
rect 135364 51644 135370 51656
rect 136870 51644 136876 51656
rect 135364 51616 136876 51644
rect 135364 51604 135370 51616
rect 136870 51604 136876 51616
rect 136928 51604 136934 51656
rect 172014 51604 172020 51656
rect 172072 51644 172078 51656
rect 174222 51644 174228 51656
rect 172072 51616 174228 51644
rect 172072 51604 172078 51616
rect 174222 51604 174228 51616
rect 174280 51604 174286 51656
rect 135030 51332 135036 51384
rect 135088 51372 135094 51384
rect 136778 51372 136784 51384
rect 135088 51344 136784 51372
rect 135088 51332 135094 51344
rect 136778 51332 136784 51344
rect 136836 51332 136842 51384
rect 135398 51060 135404 51112
rect 135456 51100 135462 51112
rect 136686 51100 136692 51112
rect 135456 51072 136692 51100
rect 135456 51060 135462 51072
rect 136686 51060 136692 51072
rect 136744 51060 136750 51112
rect 63822 50584 63828 50636
rect 63880 50624 63886 50636
rect 66398 50624 66404 50636
rect 63880 50596 66404 50624
rect 63880 50584 63886 50596
rect 66398 50584 66404 50596
rect 66456 50584 66462 50636
rect 62810 50448 62816 50500
rect 62868 50488 62874 50500
rect 65662 50488 65668 50500
rect 62868 50460 65668 50488
rect 62868 50448 62874 50460
rect 65662 50448 65668 50460
rect 65720 50448 65726 50500
rect 100622 50448 100628 50500
rect 100680 50488 100686 50500
rect 102646 50488 102652 50500
rect 100680 50460 102652 50488
rect 100680 50448 100686 50460
rect 102646 50448 102652 50460
rect 102704 50448 102710 50500
rect 100622 50312 100628 50364
rect 100680 50352 100686 50364
rect 102370 50352 102376 50364
rect 100680 50324 102376 50352
rect 100680 50312 100686 50324
rect 102370 50312 102376 50324
rect 102428 50312 102434 50364
rect 172198 50312 172204 50364
rect 172256 50352 172262 50364
rect 174130 50352 174136 50364
rect 172256 50324 174136 50352
rect 172256 50312 172262 50324
rect 174130 50312 174136 50324
rect 174188 50312 174194 50364
rect 135398 50244 135404 50296
rect 135456 50284 135462 50296
rect 136870 50284 136876 50296
rect 135456 50256 136876 50284
rect 135456 50244 135462 50256
rect 136870 50244 136876 50256
rect 136928 50244 136934 50296
rect 172658 50244 172664 50296
rect 172716 50284 172722 50296
rect 174314 50284 174320 50296
rect 172716 50256 174320 50284
rect 172716 50244 172722 50256
rect 174314 50244 174320 50256
rect 174372 50244 174378 50296
rect 134846 50176 134852 50228
rect 134904 50216 134910 50228
rect 136778 50216 136784 50228
rect 134904 50188 136784 50216
rect 134904 50176 134910 50188
rect 136778 50176 136784 50188
rect 136836 50176 136842 50228
rect 100622 49224 100628 49276
rect 100680 49264 100686 49276
rect 102462 49264 102468 49276
rect 100680 49236 102468 49264
rect 100680 49224 100686 49236
rect 102462 49224 102468 49236
rect 102520 49224 102526 49276
rect 172658 49224 172664 49276
rect 172716 49264 172722 49276
rect 174222 49264 174228 49276
rect 172716 49236 174228 49264
rect 172716 49224 172722 49236
rect 174222 49224 174228 49236
rect 174280 49224 174286 49276
rect 171830 49088 171836 49140
rect 171888 49128 171894 49140
rect 174406 49128 174412 49140
rect 171888 49100 174412 49128
rect 171888 49088 171894 49100
rect 174406 49088 174412 49100
rect 174464 49088 174470 49140
rect 63730 48952 63736 49004
rect 63788 48992 63794 49004
rect 65478 48992 65484 49004
rect 63788 48964 65484 48992
rect 63788 48952 63794 48964
rect 65478 48952 65484 48964
rect 65536 48952 65542 49004
rect 100622 48952 100628 49004
rect 100680 48992 100686 49004
rect 102554 48992 102560 49004
rect 100680 48964 102560 48992
rect 100680 48952 100686 48964
rect 102554 48952 102560 48964
rect 102612 48952 102618 49004
rect 63362 48884 63368 48936
rect 63420 48924 63426 48936
rect 66398 48924 66404 48936
rect 63420 48896 66404 48924
rect 63420 48884 63426 48896
rect 66398 48884 66404 48896
rect 66456 48884 66462 48936
rect 136870 48924 136876 48936
rect 135508 48896 136876 48924
rect 135306 48816 135312 48868
rect 135364 48856 135370 48868
rect 135508 48856 135536 48896
rect 136870 48884 136876 48896
rect 136928 48884 136934 48936
rect 135364 48828 135536 48856
rect 135364 48816 135370 48828
rect 134754 48408 134760 48460
rect 134812 48448 134818 48460
rect 136778 48448 136784 48460
rect 134812 48420 136784 48448
rect 134812 48408 134818 48420
rect 136778 48408 136784 48420
rect 136836 48408 136842 48460
rect 100622 47864 100628 47916
rect 100680 47904 100686 47916
rect 102646 47904 102652 47916
rect 100680 47876 102652 47904
rect 100680 47864 100686 47876
rect 102646 47864 102652 47876
rect 102704 47864 102710 47916
rect 172566 47864 172572 47916
rect 172624 47904 172630 47916
rect 174222 47904 174228 47916
rect 172624 47876 174228 47904
rect 172624 47864 172630 47876
rect 174222 47864 174228 47876
rect 174280 47864 174286 47916
rect 172658 47728 172664 47780
rect 172716 47768 172722 47780
rect 174130 47768 174136 47780
rect 172716 47740 174136 47768
rect 172716 47728 172722 47740
rect 174130 47728 174136 47740
rect 174188 47728 174194 47780
rect 100622 47592 100628 47644
rect 100680 47632 100686 47644
rect 102370 47632 102376 47644
rect 100680 47604 102376 47632
rect 100680 47592 100686 47604
rect 102370 47592 102376 47604
rect 102428 47592 102434 47644
rect 172658 47592 172664 47644
rect 172716 47632 172722 47644
rect 174314 47632 174320 47644
rect 172716 47604 174320 47632
rect 172716 47592 172722 47604
rect 174314 47592 174320 47604
rect 174372 47592 174378 47644
rect 62810 47456 62816 47508
rect 62868 47496 62874 47508
rect 65662 47496 65668 47508
rect 62868 47468 65668 47496
rect 62868 47456 62874 47468
rect 65662 47456 65668 47468
rect 65720 47456 65726 47508
rect 100622 47456 100628 47508
rect 100680 47496 100686 47508
rect 102462 47496 102468 47508
rect 100680 47468 102468 47496
rect 100680 47456 100686 47468
rect 102462 47456 102468 47468
rect 102520 47456 102526 47508
rect 135398 47456 135404 47508
rect 135456 47496 135462 47508
rect 136870 47496 136876 47508
rect 135456 47468 136876 47496
rect 135456 47456 135462 47468
rect 136870 47456 136876 47468
rect 136928 47456 136934 47508
rect 62902 47388 62908 47440
rect 62960 47428 62966 47440
rect 64926 47428 64932 47440
rect 62960 47400 64932 47428
rect 62960 47388 62966 47400
rect 64926 47388 64932 47400
rect 64984 47388 64990 47440
rect 134846 47320 134852 47372
rect 134904 47360 134910 47372
rect 136778 47360 136784 47372
rect 134904 47332 136784 47360
rect 134904 47320 134910 47332
rect 136778 47320 136784 47332
rect 136836 47320 136842 47372
rect 135306 47116 135312 47168
rect 135364 47156 135370 47168
rect 136686 47156 136692 47168
rect 135364 47128 136692 47156
rect 135364 47116 135370 47128
rect 136686 47116 136692 47128
rect 136744 47116 136750 47168
rect 62718 46912 62724 46964
rect 62776 46952 62782 46964
rect 65018 46952 65024 46964
rect 62776 46924 65024 46952
rect 62776 46912 62782 46924
rect 65018 46912 65024 46924
rect 65076 46912 65082 46964
rect 172658 46504 172664 46556
rect 172716 46544 172722 46556
rect 174222 46544 174228 46556
rect 172716 46516 174228 46544
rect 172716 46504 172722 46516
rect 174222 46504 174228 46516
rect 174280 46504 174286 46556
rect 63730 46368 63736 46420
rect 63788 46408 63794 46420
rect 66398 46408 66404 46420
rect 63788 46380 66404 46408
rect 63788 46368 63794 46380
rect 66398 46368 66404 46380
rect 66456 46368 66462 46420
rect 100622 46232 100628 46284
rect 100680 46272 100686 46284
rect 102554 46272 102560 46284
rect 100680 46244 102560 46272
rect 100680 46232 100686 46244
rect 102554 46232 102560 46244
rect 102612 46232 102618 46284
rect 100898 46096 100904 46148
rect 100956 46136 100962 46148
rect 102370 46136 102376 46148
rect 100956 46108 102376 46136
rect 100956 46096 100962 46108
rect 102370 46096 102376 46108
rect 102428 46096 102434 46148
rect 172658 46096 172664 46148
rect 172716 46136 172722 46148
rect 175326 46136 175332 46148
rect 172716 46108 175332 46136
rect 172716 46096 172722 46108
rect 175326 46096 175332 46108
rect 175384 46096 175390 46148
rect 134662 46028 134668 46080
rect 134720 46068 134726 46080
rect 136778 46068 136784 46080
rect 134720 46040 136784 46068
rect 134720 46028 134726 46040
rect 136778 46028 136784 46040
rect 136836 46028 136842 46080
rect 100530 45212 100536 45264
rect 100588 45252 100594 45264
rect 102462 45252 102468 45264
rect 100588 45224 102468 45252
rect 100588 45212 100594 45224
rect 102462 45212 102468 45224
rect 102520 45212 102526 45264
rect 99978 44940 99984 44992
rect 100036 44980 100042 44992
rect 102554 44980 102560 44992
rect 100036 44952 102560 44980
rect 100036 44940 100042 44952
rect 102554 44940 102560 44952
rect 102612 44940 102618 44992
rect 171646 44940 171652 44992
rect 171704 44980 171710 44992
rect 175418 44980 175424 44992
rect 171704 44952 175424 44980
rect 171704 44940 171710 44952
rect 175418 44940 175424 44952
rect 175476 44940 175482 44992
rect 63730 44804 63736 44856
rect 63788 44844 63794 44856
rect 66306 44844 66312 44856
rect 63788 44816 66312 44844
rect 63788 44804 63794 44816
rect 66306 44804 66312 44816
rect 66364 44804 66370 44856
rect 63638 44736 63644 44788
rect 63696 44776 63702 44788
rect 66398 44776 66404 44788
rect 63696 44748 66404 44776
rect 63696 44736 63702 44748
rect 66398 44736 66404 44748
rect 66456 44736 66462 44788
rect 171830 44736 171836 44788
rect 171888 44776 171894 44788
rect 174774 44776 174780 44788
rect 171888 44748 174780 44776
rect 171888 44736 171894 44748
rect 174774 44736 174780 44748
rect 174832 44736 174838 44788
rect 62810 44668 62816 44720
rect 62868 44708 62874 44720
rect 65202 44708 65208 44720
rect 62868 44680 65208 44708
rect 62868 44668 62874 44680
rect 65202 44668 65208 44680
rect 65260 44668 65266 44720
rect 135030 44668 135036 44720
rect 135088 44708 135094 44720
rect 137514 44708 137520 44720
rect 135088 44680 137520 44708
rect 135088 44668 135094 44680
rect 137514 44668 137520 44680
rect 137572 44668 137578 44720
rect 135398 44396 135404 44448
rect 135456 44436 135462 44448
rect 136686 44436 136692 44448
rect 135456 44408 136692 44436
rect 135456 44396 135462 44408
rect 136686 44396 136692 44408
rect 136744 44396 136750 44448
rect 135030 44260 135036 44312
rect 135088 44300 135094 44312
rect 136778 44300 136784 44312
rect 135088 44272 136784 44300
rect 135088 44260 135094 44272
rect 136778 44260 136784 44272
rect 136836 44260 136842 44312
rect 99886 44056 99892 44108
rect 99944 44096 99950 44108
rect 102278 44096 102284 44108
rect 99944 44068 102284 44096
rect 99944 44056 99950 44068
rect 102278 44056 102284 44068
rect 102336 44056 102342 44108
rect 172658 43580 172664 43632
rect 172716 43620 172722 43632
rect 174038 43620 174044 43632
rect 172716 43592 174044 43620
rect 172716 43580 172722 43592
rect 174038 43580 174044 43592
rect 174096 43580 174102 43632
rect 63730 43512 63736 43564
rect 63788 43552 63794 43564
rect 66214 43552 66220 43564
rect 63788 43524 66220 43552
rect 63788 43512 63794 43524
rect 66214 43512 66220 43524
rect 66272 43512 66278 43564
rect 63822 43308 63828 43360
rect 63880 43348 63886 43360
rect 66398 43348 66404 43360
rect 63880 43320 66404 43348
rect 63880 43308 63886 43320
rect 66398 43308 66404 43320
rect 66456 43308 66462 43360
rect 100622 43308 100628 43360
rect 100680 43348 100686 43360
rect 136870 43348 136876 43360
rect 100680 43320 101036 43348
rect 100680 43308 100686 43320
rect 101008 43280 101036 43320
rect 135508 43320 136876 43348
rect 102370 43280 102376 43292
rect 101008 43252 102376 43280
rect 102370 43240 102376 43252
rect 102428 43240 102434 43292
rect 134938 43240 134944 43292
rect 134996 43280 135002 43292
rect 135508 43280 135536 43320
rect 136870 43308 136876 43320
rect 136928 43308 136934 43360
rect 172566 43308 172572 43360
rect 172624 43348 172630 43360
rect 172624 43320 172796 43348
rect 172624 43308 172630 43320
rect 134996 43252 135536 43280
rect 172768 43280 172796 43320
rect 174130 43280 174136 43292
rect 172768 43252 174136 43280
rect 134996 43240 135002 43252
rect 174130 43240 174136 43252
rect 174188 43240 174194 43292
rect 135398 43036 135404 43088
rect 135456 43076 135462 43088
rect 136778 43076 136784 43088
rect 135456 43048 136784 43076
rect 135456 43036 135462 43048
rect 136778 43036 136784 43048
rect 136836 43036 136842 43088
rect 100622 42628 100628 42680
rect 100680 42668 100686 42680
rect 102554 42668 102560 42680
rect 100680 42640 102560 42668
rect 100680 42628 100686 42640
rect 102554 42628 102560 42640
rect 102612 42628 102618 42680
rect 63822 42288 63828 42340
rect 63880 42328 63886 42340
rect 66398 42328 66404 42340
rect 63880 42300 66404 42328
rect 63880 42288 63886 42300
rect 66398 42288 66404 42300
rect 66456 42288 66462 42340
rect 172198 42288 172204 42340
rect 172256 42328 172262 42340
rect 174222 42328 174228 42340
rect 172256 42300 174228 42328
rect 172256 42288 172262 42300
rect 174222 42288 174228 42300
rect 174280 42288 174286 42340
rect 100622 42152 100628 42204
rect 100680 42192 100686 42204
rect 102462 42192 102468 42204
rect 100680 42164 102468 42192
rect 100680 42152 100686 42164
rect 102462 42152 102468 42164
rect 102520 42152 102526 42204
rect 172658 42152 172664 42204
rect 172716 42192 172722 42204
rect 174314 42192 174320 42204
rect 172716 42164 174320 42192
rect 172716 42152 172722 42164
rect 174314 42152 174320 42164
rect 174372 42152 174378 42204
rect 100622 42016 100628 42068
rect 100680 42056 100686 42068
rect 102370 42056 102376 42068
rect 100680 42028 102376 42056
rect 100680 42016 100686 42028
rect 102370 42016 102376 42028
rect 102428 42016 102434 42068
rect 172658 42016 172664 42068
rect 172716 42056 172722 42068
rect 174130 42056 174136 42068
rect 172716 42028 174136 42056
rect 172716 42016 172722 42028
rect 174130 42016 174136 42028
rect 174188 42016 174194 42068
rect 63730 41948 63736 42000
rect 63788 41988 63794 42000
rect 66306 41988 66312 42000
rect 63788 41960 66312 41988
rect 63788 41948 63794 41960
rect 66306 41948 66312 41960
rect 66364 41948 66370 42000
rect 136870 41988 136876 42000
rect 135508 41960 136876 41988
rect 135398 41880 135404 41932
rect 135456 41920 135462 41932
rect 135508 41920 135536 41960
rect 136870 41948 136876 41960
rect 136928 41948 136934 42000
rect 135456 41892 135536 41920
rect 135456 41880 135462 41892
rect 135306 41812 135312 41864
rect 135364 41852 135370 41864
rect 136686 41852 136692 41864
rect 135364 41824 136692 41852
rect 135364 41812 135370 41824
rect 136686 41812 136692 41824
rect 136744 41812 136750 41864
rect 134846 41472 134852 41524
rect 134904 41512 134910 41524
rect 136778 41512 136784 41524
rect 134904 41484 136784 41512
rect 134904 41472 134910 41484
rect 136778 41472 136784 41484
rect 136836 41472 136842 41524
rect 63178 40520 63184 40572
rect 63236 40560 63242 40572
rect 66398 40560 66404 40572
rect 63236 40532 66404 40560
rect 63236 40520 63242 40532
rect 66398 40520 66404 40532
rect 66456 40520 66462 40572
rect 71918 39908 71924 39960
rect 71976 39948 71982 39960
rect 82498 39948 82504 39960
rect 71976 39920 82504 39948
rect 71976 39908 71982 39920
rect 82498 39908 82504 39920
rect 82556 39908 82562 39960
rect 143586 39908 143592 39960
rect 143644 39948 143650 39960
rect 154810 39948 154816 39960
rect 143644 39920 154816 39948
rect 143644 39908 143650 39920
rect 154810 39908 154816 39920
rect 154868 39908 154874 39960
rect 66306 39840 66312 39892
rect 66364 39880 66370 39892
rect 86270 39880 86276 39892
rect 66364 39852 86276 39880
rect 66364 39840 66370 39852
rect 86270 39840 86276 39852
rect 86328 39840 86334 39892
rect 138066 39840 138072 39892
rect 138124 39880 138130 39892
rect 158582 39880 158588 39892
rect 138124 39852 158588 39880
rect 138124 39840 138130 39852
rect 158582 39840 158588 39852
rect 158640 39840 158646 39892
rect 62810 39160 62816 39212
rect 62868 39200 62874 39212
rect 72562 39200 72568 39212
rect 62868 39172 72568 39200
rect 62868 39160 62874 39172
rect 72562 39160 72568 39172
rect 72620 39160 72626 39212
rect 93170 39160 93176 39212
rect 93228 39200 93234 39212
rect 102370 39200 102376 39212
rect 93228 39172 102376 39200
rect 93228 39160 93234 39172
rect 102370 39160 102376 39172
rect 102428 39160 102434 39212
rect 134478 39160 134484 39212
rect 134536 39200 134542 39212
rect 144874 39200 144880 39212
rect 134536 39172 144880 39200
rect 134536 39160 134542 39172
rect 144874 39160 144880 39172
rect 144932 39160 144938 39212
rect 164838 39160 164844 39212
rect 164896 39200 164902 39212
rect 174130 39200 174136 39212
rect 164896 39172 174136 39200
rect 164896 39160 164902 39172
rect 174130 39160 174136 39172
rect 174188 39160 174194 39212
rect 79370 37732 79376 37784
rect 79428 37772 79434 37784
rect 127762 37772 127768 37784
rect 79428 37744 127768 37772
rect 79428 37732 79434 37744
rect 127762 37732 127768 37744
rect 127820 37732 127826 37784
rect 151038 37732 151044 37784
rect 151096 37772 151102 37784
rect 200074 37772 200080 37784
rect 151096 37744 200080 37772
rect 151096 37732 151102 37744
rect 200074 37732 200080 37744
rect 200132 37732 200138 37784
rect 222522 37772 222528 37784
rect 222483 37744 222528 37772
rect 222522 37732 222528 37744
rect 222580 37732 222586 37784
rect 190782 37664 190788 37716
rect 190840 37704 190846 37716
rect 205134 37704 205140 37716
rect 190840 37676 205140 37704
rect 190840 37664 190846 37676
rect 205134 37664 205140 37676
rect 205192 37664 205198 37716
rect 30518 33584 30524 33636
rect 30576 33624 30582 33636
rect 66214 33624 66220 33636
rect 30576 33596 66220 33624
rect 30576 33584 30582 33596
rect 66214 33584 66220 33596
rect 66272 33584 66278 33636
rect 118838 33584 118844 33636
rect 118896 33624 118902 33636
rect 136870 33624 136876 33636
rect 118896 33596 136876 33624
rect 118896 33584 118902 33596
rect 136870 33584 136876 33596
rect 136928 33584 136934 33636
rect 222525 28187 222583 28193
rect 222525 28153 222537 28187
rect 222571 28184 222583 28187
rect 222706 28184 222712 28196
rect 222571 28156 222712 28184
rect 222571 28153 222583 28156
rect 222525 28147 222583 28153
rect 222706 28144 222712 28156
rect 222764 28144 222770 28196
rect 77990 12572 77996 12624
rect 78048 12612 78054 12624
rect 79048 12612 79054 12624
rect 78048 12584 79054 12612
rect 78048 12572 78054 12584
rect 79048 12572 79054 12584
rect 79106 12572 79112 12624
rect 86914 11688 86920 11740
rect 86972 11728 86978 11740
rect 132546 11728 132552 11740
rect 86972 11700 132552 11728
rect 86972 11688 86978 11700
rect 132546 11688 132552 11700
rect 132604 11688 132610 11740
rect 166034 11688 166040 11740
rect 166092 11728 166098 11740
rect 214242 11728 214248 11740
rect 166092 11700 214248 11728
rect 166092 11688 166098 11700
rect 214242 11688 214248 11700
rect 214300 11688 214306 11740
rect 93998 11620 94004 11672
rect 94056 11660 94062 11672
rect 187010 11660 187016 11672
rect 94056 11632 187016 11660
rect 94056 11620 94062 11632
rect 187010 11620 187016 11632
rect 187068 11620 187074 11672
rect 23526 10940 23532 10992
rect 23584 10980 23590 10992
rect 71274 10980 71280 10992
rect 23584 10952 71280 10980
rect 23584 10940 23590 10952
rect 71274 10940 71280 10952
rect 71332 10940 71338 10992
rect 105222 10940 105228 10992
rect 105280 10980 105286 10992
rect 151038 10980 151044 10992
rect 105280 10952 151044 10980
rect 105280 10940 105286 10952
rect 151038 10940 151044 10952
rect 151096 10940 151102 10992
rect 50758 10872 50764 10924
rect 50816 10912 50822 10924
rect 143586 10912 143592 10924
rect 50816 10884 143592 10912
rect 50816 10872 50822 10884
rect 143586 10872 143592 10884
rect 143644 10872 143650 10924
rect 158582 10396 158588 10448
rect 158640 10436 158646 10448
rect 159778 10436 159784 10448
rect 158640 10408 159784 10436
rect 158640 10396 158646 10408
rect 159778 10396 159784 10408
rect 159836 10396 159842 10448
<< via1 >>
rect 23532 244860 23584 244912
rect 70544 244860 70596 244912
rect 105228 244860 105280 244912
rect 149664 244860 149716 244912
rect 50764 244792 50816 244844
rect 142396 244792 142448 244844
rect 157484 244792 157536 244844
rect 159784 244792 159836 244844
rect 85632 242412 85684 242464
rect 132552 242140 132604 242192
rect 165304 242140 165356 242192
rect 214248 242140 214300 242192
rect 93360 242072 93412 242124
rect 187016 242072 187068 242124
rect 167788 229764 167840 229816
rect 168524 229764 168576 229816
rect 207256 223372 207308 223424
rect 223080 223372 223132 223424
rect 170088 222760 170140 222812
rect 207256 222760 207308 222812
rect 71372 217932 71424 217984
rect 143684 217932 143736 217984
rect 170088 217932 170140 217984
rect 46532 217864 46584 217916
rect 98236 217864 98288 217916
rect 98420 217864 98472 217916
rect 109276 217864 109328 217916
rect 118844 217864 118896 217916
rect 169996 217864 170048 217916
rect 109276 217252 109328 217304
rect 143684 217252 143736 217304
rect 37240 217184 37292 217236
rect 71372 217184 71424 217236
rect 79376 217184 79428 217236
rect 127768 217184 127820 217236
rect 81768 216572 81820 216624
rect 94004 216572 94056 216624
rect 158588 216572 158640 216624
rect 167236 216572 167288 216624
rect 91796 216504 91848 216556
rect 102376 216504 102428 216556
rect 164108 216504 164160 216556
rect 174228 216504 174280 216556
rect 86920 216436 86972 216488
rect 98328 216436 98380 216488
rect 154080 216436 154132 216488
rect 166040 216436 166092 216488
rect 62540 215756 62592 215808
rect 71832 215756 71884 215808
rect 135404 215756 135456 215808
rect 143776 215756 143828 215808
rect 100996 214600 101048 214652
rect 102560 214600 102612 214652
rect 135404 214600 135456 214652
rect 136784 214600 136836 214652
rect 62632 214532 62684 214584
rect 65024 214532 65076 214584
rect 172020 213988 172072 214040
rect 174044 213988 174096 214040
rect 135404 213648 135456 213700
rect 136876 213648 136928 213700
rect 100996 213308 101048 213360
rect 103112 213308 103164 213360
rect 62540 213240 62592 213292
rect 65024 213240 65076 213292
rect 135036 213240 135088 213292
rect 137060 213240 137112 213292
rect 63736 213036 63788 213088
rect 66404 213036 66456 213088
rect 100536 213036 100588 213088
rect 102376 213104 102428 213156
rect 172664 213036 172716 213088
rect 174228 213104 174280 213156
rect 172664 212628 172716 212680
rect 174044 212628 174096 212680
rect 135404 212152 135456 212204
rect 136968 212152 137020 212204
rect 100996 211880 101048 211932
rect 102376 211880 102428 211932
rect 135404 211880 135456 211932
rect 136876 211880 136928 211932
rect 62356 211744 62408 211796
rect 64932 211744 64984 211796
rect 62632 211676 62684 211728
rect 65024 211676 65076 211728
rect 100812 211608 100864 211660
rect 102468 211676 102520 211728
rect 172756 211676 172808 211728
rect 174228 211676 174280 211728
rect 172388 211268 172440 211320
rect 174044 211268 174096 211320
rect 62540 210792 62592 210844
rect 65484 210792 65536 210844
rect 100904 210792 100956 210844
rect 103664 210792 103716 210844
rect 172664 210588 172716 210640
rect 174228 210588 174280 210640
rect 100996 210520 101048 210572
rect 102376 210520 102428 210572
rect 134668 210520 134720 210572
rect 136876 210520 136928 210572
rect 62632 210384 62684 210436
rect 65024 210384 65076 210436
rect 207900 210316 207952 210368
rect 223540 210316 223592 210368
rect 172664 210044 172716 210096
rect 174044 210044 174096 210096
rect 62632 209840 62684 209892
rect 66404 209840 66456 209892
rect 171652 209364 171704 209416
rect 174136 209364 174188 209416
rect 62724 209024 62776 209076
rect 65024 209024 65076 209076
rect 135312 209024 135364 209076
rect 137704 209024 137756 209076
rect 172112 208888 172164 208940
rect 174596 208956 174648 209008
rect 62632 208344 62684 208396
rect 66404 208344 66456 208396
rect 135404 207800 135456 207852
rect 136876 207800 136928 207852
rect 63736 207460 63788 207512
rect 65300 207460 65352 207512
rect 171652 206780 171704 206832
rect 174136 206780 174188 206832
rect 62540 206712 62592 206764
rect 65668 206712 65720 206764
rect 135404 206304 135456 206356
rect 136876 206304 136928 206356
rect 62632 206168 62684 206220
rect 64932 206168 64984 206220
rect 171836 205964 171888 206016
rect 174044 205964 174096 206016
rect 62632 205420 62684 205472
rect 66404 205420 66456 205472
rect 62632 204332 62684 204384
rect 65668 204332 65720 204384
rect 62540 204196 62592 204248
rect 65484 204196 65536 204248
rect 100904 200660 100956 200712
rect 102376 200660 102428 200712
rect 135404 200456 135456 200508
rect 136784 200456 136836 200508
rect 172204 199368 172256 199420
rect 175240 199368 175292 199420
rect 100904 199300 100956 199352
rect 102376 199300 102428 199352
rect 62356 199096 62408 199148
rect 65024 199096 65076 199148
rect 134760 199096 134812 199148
rect 136784 199096 136836 199148
rect 172204 198008 172256 198060
rect 174228 198008 174280 198060
rect 100904 197872 100956 197924
rect 102376 197872 102428 197924
rect 62632 197736 62684 197788
rect 65024 197736 65076 197788
rect 135404 197736 135456 197788
rect 136784 197736 136836 197788
rect 172664 196784 172716 196836
rect 174136 196784 174188 196836
rect 100904 196648 100956 196700
rect 102376 196648 102428 196700
rect 172204 196648 172256 196700
rect 174228 196648 174280 196700
rect 63736 196512 63788 196564
rect 66404 196512 66456 196564
rect 100904 196512 100956 196564
rect 102468 196512 102520 196564
rect 62632 196444 62684 196496
rect 65024 196444 65076 196496
rect 135404 196376 135456 196428
rect 136784 196376 136836 196428
rect 134300 196036 134352 196088
rect 136692 196036 136744 196088
rect 171468 195560 171520 195612
rect 174136 195560 174188 195612
rect 100720 195288 100772 195340
rect 102468 195288 102520 195340
rect 62540 195084 62592 195136
rect 66404 195152 66456 195204
rect 100904 195152 100956 195204
rect 102376 195152 102428 195204
rect 135404 195084 135456 195136
rect 136876 195152 136928 195204
rect 172664 195152 172716 195204
rect 174228 195152 174280 195204
rect 62632 194948 62684 195000
rect 65024 194948 65076 195000
rect 135404 194812 135456 194864
rect 136784 194812 136836 194864
rect 100628 194200 100680 194252
rect 102468 194200 102520 194252
rect 171560 194200 171612 194252
rect 174136 194200 174188 194252
rect 100628 193792 100680 193844
rect 102376 193792 102428 193844
rect 172664 193792 172716 193844
rect 174228 193792 174280 193844
rect 135404 193656 135456 193708
rect 136784 193656 136836 193708
rect 135404 193452 135456 193504
rect 136692 193452 136744 193504
rect 62356 193248 62408 193300
rect 65024 193248 65076 193300
rect 171652 192976 171704 193028
rect 174228 192976 174280 193028
rect 99708 192840 99760 192892
rect 102468 192840 102520 192892
rect 172204 192568 172256 192620
rect 174136 192568 174188 192620
rect 100628 192432 100680 192484
rect 102376 192432 102428 192484
rect 135404 192296 135456 192348
rect 136784 192296 136836 192348
rect 62540 192228 62592 192280
rect 64932 192228 64984 192280
rect 134300 192228 134352 192280
rect 136692 192228 136744 192280
rect 99892 191888 99944 191940
rect 102284 191888 102336 191940
rect 62356 191548 62408 191600
rect 65024 191548 65076 191600
rect 172204 191344 172256 191396
rect 174044 191344 174096 191396
rect 172664 191276 172716 191328
rect 173952 191276 174004 191328
rect 100628 191208 100680 191260
rect 102192 191208 102244 191260
rect 62448 190936 62500 190988
rect 66312 191004 66364 191056
rect 100904 191004 100956 191056
rect 102560 191004 102612 191056
rect 134300 191004 134352 191056
rect 136968 191004 137020 191056
rect 172664 191004 172716 191056
rect 174964 191004 175016 191056
rect 135404 190936 135456 190988
rect 136784 190936 136836 190988
rect 62632 190868 62684 190920
rect 65024 190868 65076 190920
rect 134760 190868 134812 190920
rect 136692 190868 136744 190920
rect 172388 190120 172440 190172
rect 174412 190120 174464 190172
rect 100536 190052 100588 190104
rect 102468 190052 102520 190104
rect 99892 189780 99944 189832
rect 102376 189780 102428 189832
rect 172020 189712 172072 189764
rect 175424 189712 175476 189764
rect 63644 189644 63696 189696
rect 66404 189644 66456 189696
rect 62632 189508 62684 189560
rect 65208 189508 65260 189560
rect 134760 189236 134812 189288
rect 136784 189236 136836 189288
rect 62632 189032 62684 189084
rect 65024 189032 65076 189084
rect 135036 188148 135088 188200
rect 137428 188148 137480 188200
rect 116452 187604 116504 187656
rect 117418 187604 117470 187656
rect 132644 186924 132696 186976
rect 144880 186924 144932 186976
rect 121880 186856 121932 186908
rect 125192 186856 125244 186908
rect 132092 186856 132144 186908
rect 164844 186856 164896 186908
rect 35584 185428 35636 185480
rect 37884 185428 37936 185480
rect 41012 185428 41064 185480
rect 43404 185428 43456 185480
rect 43772 185428 43824 185480
rect 44692 185428 44744 185480
rect 49016 185428 49068 185480
rect 50580 185428 50632 185480
rect 50672 185428 50724 185480
rect 53340 185428 53392 185480
rect 53432 185428 53484 185480
rect 58124 185428 58176 185480
rect 110104 185428 110156 185480
rect 111116 185428 111168 185480
rect 125928 185428 125980 185480
rect 128136 185428 128188 185480
rect 182876 185428 182928 185480
rect 183612 185428 183664 185480
rect 190144 185428 190196 185480
rect 191432 185428 191484 185480
rect 197320 185428 197372 185480
rect 201644 185428 201696 185480
rect 40368 185360 40420 185412
rect 43036 185360 43088 185412
rect 43128 185360 43180 185412
rect 44600 185360 44652 185412
rect 50212 185360 50264 185412
rect 52696 185360 52748 185412
rect 110748 185360 110800 185412
rect 111484 185360 111536 185412
rect 127216 185360 127268 185412
rect 129976 185360 130028 185412
rect 190604 185360 190656 185412
rect 192536 185360 192588 185412
rect 192904 185360 192956 185412
rect 195388 185360 195440 185412
rect 195756 185360 195808 185412
rect 199344 185360 199396 185412
rect 36320 185292 36372 185344
rect 40644 185292 40696 185344
rect 41748 185292 41800 185344
rect 43864 185292 43916 185344
rect 52236 185292 52288 185344
rect 56100 185292 56152 185344
rect 125928 185292 125980 185344
rect 127308 185292 127360 185344
rect 193364 185292 193416 185344
rect 195940 185292 195992 185344
rect 196124 185292 196176 185344
rect 199988 185292 200040 185344
rect 39724 185224 39776 185276
rect 42668 185224 42720 185276
rect 49476 185224 49528 185276
rect 51316 185224 51368 185276
rect 53064 185224 53116 185276
rect 57388 185224 57440 185276
rect 105596 185224 105648 185276
rect 109276 185224 109328 185276
rect 124824 185224 124876 185276
rect 126388 185224 126440 185276
rect 192536 185224 192588 185276
rect 194836 185224 194888 185276
rect 195296 185224 195348 185276
rect 198792 185224 198844 185276
rect 37608 185156 37660 185208
rect 41472 185156 41524 185208
rect 51040 185156 51092 185208
rect 53984 185156 54036 185208
rect 194100 185156 194152 185208
rect 197136 185156 197188 185208
rect 38988 185088 39040 185140
rect 42208 185088 42260 185140
rect 42392 185088 42444 185140
rect 44232 185088 44284 185140
rect 49844 185088 49896 185140
rect 51960 185088 52012 185140
rect 52604 185088 52656 185140
rect 56744 185088 56796 185140
rect 190420 185088 190472 185140
rect 191984 185088 192036 185140
rect 194560 185088 194612 185140
rect 197688 185088 197740 185140
rect 38344 185020 38396 185072
rect 41840 185020 41892 185072
rect 48648 185020 48700 185072
rect 49936 185020 49988 185072
rect 51408 185020 51460 185072
rect 54720 185020 54772 185072
rect 127216 185020 127268 185072
rect 130436 185020 130488 185072
rect 194652 185020 194704 185072
rect 198240 185020 198292 185072
rect 51868 184952 51920 185004
rect 55364 184952 55416 185004
rect 177724 184952 177776 185004
rect 181128 184952 181180 185004
rect 181680 184952 181732 185004
rect 183106 184952 183158 185004
rect 189086 184952 189138 185004
rect 190236 184952 190288 185004
rect 191110 184952 191162 185004
rect 193088 184952 193140 185004
rect 193502 184952 193554 185004
rect 196492 184952 196544 185004
rect 197826 184952 197878 185004
rect 202840 184952 202892 185004
rect 36964 184884 37016 184936
rect 41012 184884 41064 184936
rect 127216 184884 127268 184936
rect 129332 184884 129384 184936
rect 182232 184884 182284 184936
rect 183474 184884 183526 184936
rect 189454 184884 189506 184936
rect 190788 184884 190840 184936
rect 191478 184884 191530 184936
rect 193640 184884 193692 184936
rect 196630 184884 196682 184936
rect 201092 184884 201144 184936
rect 191984 184816 192036 184868
rect 194008 184816 194060 184868
rect 196492 184816 196544 184868
rect 200540 184816 200592 184868
rect 127032 184680 127084 184732
rect 128688 184680 128740 184732
rect 53984 184544 54036 184596
rect 58768 184544 58820 184596
rect 127032 184476 127084 184528
rect 127584 184476 127636 184528
rect 39264 184408 39316 184460
rect 54536 184408 54588 184460
rect 34940 184272 34992 184324
rect 37976 184272 38028 184324
rect 34204 184204 34256 184256
rect 59504 184204 59556 184256
rect 106056 184204 106108 184256
rect 107160 184204 107212 184256
rect 177080 184204 177132 184256
rect 179380 184204 179432 184256
rect 177632 184136 177684 184188
rect 178828 184136 178880 184188
rect 33560 184068 33612 184120
rect 38896 184068 38948 184120
rect 105964 184068 106016 184120
rect 106608 184068 106660 184120
rect 106148 184000 106200 184052
rect 108356 184068 108408 184120
rect 177540 184068 177592 184120
rect 178276 184068 178328 184120
rect 177448 184000 177500 184052
rect 180576 184068 180628 184120
rect 176988 182436 177040 182488
rect 180024 182436 180076 182488
rect 105596 182368 105648 182420
rect 107896 182368 107948 182420
rect 105412 180328 105464 180380
rect 108080 180328 108132 180380
rect 106332 178560 106384 178612
rect 107896 178560 107948 178612
rect 32640 177200 32692 177252
rect 37424 177200 37476 177252
rect 57572 177200 57624 177252
rect 59596 177200 59648 177252
rect 106424 175840 106476 175892
rect 107896 175840 107948 175892
rect 177724 175840 177776 175892
rect 179656 175840 179708 175892
rect 106148 174344 106200 174396
rect 108540 174344 108592 174396
rect 177356 174344 177408 174396
rect 180300 174344 180352 174396
rect 176988 174276 177040 174328
rect 179932 174276 179984 174328
rect 106056 173052 106108 173104
rect 108172 173052 108224 173104
rect 177632 173052 177684 173104
rect 179656 173052 179708 173104
rect 177540 172916 177592 172968
rect 179748 172916 179800 172968
rect 105228 171692 105280 171744
rect 107896 171692 107948 171744
rect 178092 171692 178144 171744
rect 179656 171692 179708 171744
rect 222804 169108 222856 169160
rect 223540 169108 223592 169160
rect 105964 168904 106016 168956
rect 107896 168904 107948 168956
rect 177540 168904 177592 168956
rect 179656 168904 179708 168956
rect 106424 166116 106476 166168
rect 107804 166116 107856 166168
rect 177540 166116 177592 166168
rect 179564 166116 179616 166168
rect 201092 166116 201144 166168
rect 204496 166116 204548 166168
rect 28868 164756 28920 164808
rect 37424 164756 37476 164808
rect 54904 164756 54956 164808
rect 59596 164756 59648 164808
rect 106424 163464 106476 163516
rect 107804 163464 107856 163516
rect 177724 163464 177776 163516
rect 179564 163464 179616 163516
rect 106148 162104 106200 162156
rect 108540 162104 108592 162156
rect 176988 162036 177040 162088
rect 179656 162036 179708 162088
rect 176988 160812 177040 160864
rect 179564 160812 179616 160864
rect 105780 160608 105832 160660
rect 107804 160608 107856 160660
rect 106424 159248 106476 159300
rect 107712 159248 107764 159300
rect 177540 159248 177592 159300
rect 179472 159248 179524 159300
rect 105412 158160 105464 158212
rect 107896 158160 107948 158212
rect 177356 157888 177408 157940
rect 179656 157888 179708 157940
rect 105412 156936 105464 156988
rect 107252 156936 107304 156988
rect 222804 156868 222856 156920
rect 223540 156868 223592 156920
rect 177540 156460 177592 156512
rect 180484 156460 180536 156512
rect 105228 155712 105280 155764
rect 107160 155712 107212 155764
rect 177540 155100 177592 155152
rect 180392 155100 180444 155152
rect 105596 153808 105648 153860
rect 107988 153808 108040 153860
rect 177356 153808 177408 153860
rect 180300 153808 180352 153860
rect 105780 153740 105832 153792
rect 108540 153740 108592 153792
rect 178184 153740 178236 153792
rect 179748 153740 179800 153792
rect 57480 151496 57532 151548
rect 59596 151496 59648 151548
rect 200540 151496 200592 151548
rect 207440 151496 207492 151548
rect 28776 146915 28828 146924
rect 28776 146881 28785 146915
rect 28785 146881 28819 146915
rect 28819 146881 28828 146915
rect 28776 146872 28828 146881
rect 178276 146600 178328 146652
rect 179012 146600 179064 146652
rect 105872 145444 105924 145496
rect 109276 145376 109328 145428
rect 178276 145240 178328 145292
rect 181128 145240 181180 145292
rect 22244 145172 22296 145224
rect 177448 145036 177500 145088
rect 180576 145036 180628 145088
rect 191846 144696 191898 144748
rect 194284 144696 194336 144748
rect 191478 144628 191530 144680
rect 193640 144628 193692 144680
rect 197826 144628 197878 144680
rect 202840 144628 202892 144680
rect 52512 144492 52564 144544
rect 55364 144492 55416 144544
rect 54628 144220 54680 144272
rect 60424 144220 60476 144272
rect 125836 144220 125888 144272
rect 131448 144220 131500 144272
rect 190604 144220 190656 144272
rect 192536 144220 192588 144272
rect 198516 144220 198568 144272
rect 203392 144220 203444 144272
rect 40644 144152 40696 144204
rect 43036 144152 43088 144204
rect 54260 144152 54312 144204
rect 59780 144152 59832 144204
rect 106424 144152 106476 144204
rect 108356 144152 108408 144204
rect 120316 144152 120368 144204
rect 122340 144152 122392 144204
rect 126664 144152 126716 144204
rect 132184 144152 132236 144204
rect 198884 144152 198936 144204
rect 203944 144152 203996 144204
rect 41288 144084 41340 144136
rect 43404 144084 43456 144136
rect 55364 144084 55416 144136
rect 56376 144084 56428 144136
rect 106516 144084 106568 144136
rect 107160 144084 107212 144136
rect 118936 144084 118988 144136
rect 120592 144084 120644 144136
rect 126296 144084 126348 144136
rect 131632 144084 131684 144136
rect 34112 142656 34164 142708
rect 39080 142656 39132 142708
rect 40000 142656 40052 142708
rect 42300 142656 42352 142708
rect 42668 142656 42720 142708
rect 44232 142656 44284 142708
rect 47820 142656 47872 142708
rect 48832 142656 48884 142708
rect 49016 142656 49068 142708
rect 50856 142656 50908 142708
rect 51040 142656 51092 142708
rect 54260 142656 54312 142708
rect 62816 142656 62868 142708
rect 16632 142588 16684 142640
rect 31812 142588 31864 142640
rect 34664 142520 34716 142572
rect 39448 142520 39500 142572
rect 42024 142520 42076 142572
rect 43864 142520 43916 142572
rect 48280 142520 48332 142572
rect 49476 142520 49528 142572
rect 50488 142520 50540 142572
rect 52972 142520 53024 142572
rect 66496 142656 66548 142708
rect 67876 142656 67928 142708
rect 72844 142656 72896 142708
rect 74500 142656 74552 142708
rect 74776 142656 74828 142708
rect 75604 142656 75656 142708
rect 80112 142656 80164 142708
rect 81676 142656 81728 142708
rect 85632 142656 85684 142708
rect 90968 142656 91020 142708
rect 95476 142656 95528 142708
rect 96764 142656 96816 142708
rect 117464 142656 117516 142708
rect 118844 142656 118896 142708
rect 120684 142656 120736 142708
rect 123444 142656 123496 142708
rect 125100 142656 125152 142708
rect 129884 142656 129936 142708
rect 142672 142656 142724 142708
rect 145432 142656 145484 142708
rect 146444 142656 146496 142708
rect 147640 142656 147692 142708
rect 154356 142656 154408 142708
rect 157668 142656 157720 142708
rect 165856 142656 165908 142708
rect 166592 142656 166644 142708
rect 182232 142656 182284 142708
rect 183244 142656 183296 142708
rect 189684 142656 189736 142708
rect 190788 142656 190840 142708
rect 191340 142656 191392 142708
rect 193088 142656 193140 142708
rect 194100 142656 194152 142708
rect 197136 142656 197188 142708
rect 201000 142656 201052 142708
rect 215904 142656 215956 142708
rect 81216 142588 81268 142640
rect 83516 142588 83568 142640
rect 86736 142588 86788 142640
rect 92808 142588 92860 142640
rect 118292 142588 118344 142640
rect 119948 142588 120000 142640
rect 125468 142588 125520 142640
rect 130436 142588 130488 142640
rect 165488 142588 165540 142640
rect 169352 142588 169404 142640
rect 189316 142588 189368 142640
rect 190236 142588 190288 142640
rect 196952 142588 197004 142640
rect 201092 142588 201144 142640
rect 71188 142520 71240 142572
rect 121052 142520 121104 142572
rect 124456 142520 124508 142572
rect 124640 142520 124692 142572
rect 129332 142520 129384 142572
rect 134484 142520 134536 142572
rect 143224 142520 143276 142572
rect 197320 142520 197372 142572
rect 201644 142520 201696 142572
rect 27580 142452 27632 142504
rect 37240 142384 37292 142436
rect 41012 142384 41064 142436
rect 39264 142316 39316 142368
rect 42208 142316 42260 142368
rect 48648 142452 48700 142504
rect 50212 142452 50264 142504
rect 50672 142452 50724 142504
rect 53616 142452 53668 142504
rect 87840 142452 87892 142504
rect 94740 142452 94792 142504
rect 102284 142452 102336 142504
rect 174320 142452 174372 142504
rect 190144 142452 190196 142504
rect 191432 142452 191484 142504
rect 194560 142452 194612 142504
rect 197688 142452 197740 142504
rect 51408 142384 51460 142436
rect 54996 142384 55048 142436
rect 69164 142384 69216 142436
rect 72292 142384 72344 142436
rect 101456 142384 101508 142436
rect 173216 142384 173268 142436
rect 192904 142384 192956 142436
rect 195388 142384 195440 142436
rect 195756 142384 195808 142436
rect 199068 142384 199120 142436
rect 54720 142316 54772 142368
rect 83424 142316 83476 142368
rect 87288 142316 87340 142368
rect 98972 142316 99024 142368
rect 102284 142316 102336 142368
rect 119488 142316 119540 142368
rect 121696 142316 121748 142368
rect 123904 142316 123956 142368
rect 128136 142316 128188 142368
rect 160980 142316 161032 142368
rect 168892 142316 168944 142368
rect 181680 142316 181732 142368
rect 182784 142316 182836 142368
rect 192444 142316 192496 142368
rect 194836 142316 194888 142368
rect 196124 142316 196176 142368
rect 199620 142316 199672 142368
rect 36596 142248 36648 142300
rect 40368 142248 40420 142300
rect 43404 142248 43456 142300
rect 44600 142248 44652 142300
rect 45428 142248 45480 142300
rect 45796 142248 45848 142300
rect 49752 142248 49804 142300
rect 51592 142248 51644 142300
rect 38620 142180 38672 142232
rect 41840 142180 41892 142232
rect 93452 142248 93504 142300
rect 98144 142248 98196 142300
rect 123720 142248 123772 142300
rect 127584 142248 127636 142300
rect 159876 142248 159928 142300
rect 167052 142248 167104 142300
rect 172112 142248 172164 142300
rect 174596 142248 174648 142300
rect 194652 142248 194704 142300
rect 198240 142248 198292 142300
rect 57480 142180 57532 142232
rect 92348 142180 92400 142232
rect 97224 142180 97276 142232
rect 121512 142180 121564 142232
rect 124640 142180 124692 142232
rect 168800 142180 168852 142232
rect 172756 142180 172808 142232
rect 195296 142180 195348 142232
rect 198792 142180 198844 142232
rect 37884 142112 37936 142164
rect 41472 142112 41524 142164
rect 49844 142112 49896 142164
rect 52236 142112 52288 142164
rect 52604 142112 52656 142164
rect 57020 142112 57072 142164
rect 62356 142112 62408 142164
rect 63460 142112 63512 142164
rect 117096 142112 117148 142164
rect 118200 142112 118252 142164
rect 123076 142112 123128 142164
rect 126940 142112 126992 142164
rect 158772 142112 158824 142164
rect 165120 142112 165172 142164
rect 190512 142112 190564 142164
rect 191984 142112 192036 142164
rect 193364 142112 193416 142164
rect 195940 142112 195992 142164
rect 196492 142112 196544 142164
rect 200540 142112 200592 142164
rect 51868 142044 51920 142096
rect 55364 142044 55416 142096
rect 182876 142044 182928 142096
rect 183612 142044 183664 142096
rect 222528 142044 222580 142096
rect 222804 142044 222856 142096
rect 53064 141976 53116 142028
rect 57664 141976 57716 142028
rect 63460 141976 63512 142028
rect 64564 141976 64616 142028
rect 88944 141976 88996 142028
rect 96856 141976 96908 142028
rect 110426 141976 110478 142028
rect 111484 141976 111536 142028
rect 113278 141976 113330 142028
rect 113508 141976 113560 142028
rect 116268 141976 116320 142028
rect 117418 141976 117470 142028
rect 117832 141976 117884 142028
rect 119718 141976 119770 142028
rect 120500 141976 120552 142028
rect 123214 141976 123266 142028
rect 124272 141976 124324 142028
rect 129010 141976 129062 142028
rect 164384 141976 164436 142028
rect 169260 141976 169312 142028
rect 193732 141976 193784 142028
rect 196492 141976 196544 142028
rect 207992 141976 208044 142028
rect 221240 141976 221292 142028
rect 109782 141908 109834 141960
rect 111116 141908 111168 141960
rect 116636 141908 116688 141960
rect 117970 141908 118022 141960
rect 119120 141908 119172 141960
rect 121466 141908 121518 141960
rect 121880 141908 121932 141960
rect 125514 141908 125566 141960
rect 153252 141908 153304 141960
rect 155828 141908 155880 141960
rect 207900 141908 207952 141960
rect 210568 141908 210620 141960
rect 222528 141908 222580 141960
rect 223540 141908 223592 141960
rect 71004 141840 71056 141892
rect 73396 141840 73448 141892
rect 84528 141840 84580 141892
rect 89128 141840 89180 141892
rect 132368 141883 132420 141892
rect 132368 141849 132377 141883
rect 132377 141849 132411 141883
rect 132411 141849 132420 141883
rect 132368 141840 132420 141849
rect 35584 141772 35636 141824
rect 39816 141772 39868 141824
rect 122892 141772 122944 141824
rect 126388 141772 126440 141824
rect 152148 141772 152200 141824
rect 153896 141772 153948 141824
rect 197412 141772 197464 141824
rect 201828 141772 201880 141824
rect 35952 141636 36004 141688
rect 40184 141636 40236 141688
rect 53432 141636 53484 141688
rect 53800 141636 53852 141688
rect 58676 141704 58728 141756
rect 122248 141704 122300 141756
rect 125836 141704 125888 141756
rect 58216 141636 58268 141688
rect 100076 141636 100128 141688
rect 103480 141636 103532 141688
rect 132092 141636 132144 141688
rect 132644 141636 132696 141688
rect 140832 141636 140884 141688
rect 144328 141636 144380 141688
rect 144512 141568 144564 141620
rect 146536 141568 146588 141620
rect 151044 141568 151096 141620
rect 152056 141568 152108 141620
rect 157944 141568 157996 141620
rect 163280 141568 163332 141620
rect 82320 141500 82372 141552
rect 85356 141500 85408 141552
rect 156564 141500 156616 141552
rect 161440 141500 161492 141552
rect 135128 141432 135180 141484
rect 137704 141432 137756 141484
rect 155460 141364 155512 141416
rect 159508 141364 159560 141416
rect 169904 141364 169956 141416
rect 97868 141296 97920 141348
rect 62816 141228 62868 141280
rect 69256 141228 69308 141280
rect 62724 141160 62776 141212
rect 68060 141160 68112 141212
rect 134576 141296 134628 141348
rect 136600 141296 136652 141348
rect 171008 141296 171060 141348
rect 102376 141160 102428 141212
rect 174228 141228 174280 141280
rect 174412 141160 174464 141212
rect 135312 141092 135364 141144
rect 141108 141092 141160 141144
rect 135312 140684 135364 140736
rect 141016 140684 141068 140736
rect 62816 139868 62868 139920
rect 66496 139868 66548 139920
rect 95476 139868 95528 139920
rect 102376 139868 102428 139920
rect 172756 139868 172808 139920
rect 174320 139868 174372 139920
rect 95568 139800 95620 139852
rect 102468 139800 102520 139852
rect 135312 139800 135364 139852
rect 139544 139800 139596 139852
rect 167236 139800 167288 139852
rect 174136 139800 174188 139852
rect 94096 139732 94148 139784
rect 102560 139732 102612 139784
rect 165856 139732 165908 139784
rect 174228 139732 174280 139784
rect 62356 139664 62408 139716
rect 66588 139664 66640 139716
rect 135312 139460 135364 139512
rect 138256 139460 138308 139512
rect 62816 139256 62868 139308
rect 65116 139256 65168 139308
rect 62908 138644 62960 138696
rect 66404 138644 66456 138696
rect 135404 138644 135456 138696
rect 136968 138644 137020 138696
rect 62816 138576 62868 138628
rect 66220 138576 66272 138628
rect 135312 138576 135364 138628
rect 136876 138576 136928 138628
rect 98144 138508 98196 138560
rect 102376 138508 102428 138560
rect 169260 138508 169312 138560
rect 174228 138508 174280 138560
rect 97224 138440 97276 138492
rect 102468 138440 102520 138492
rect 169352 138440 169404 138492
rect 174136 138440 174188 138492
rect 135220 137488 135272 137540
rect 136876 137488 136928 137540
rect 100076 137420 100128 137472
rect 102284 137420 102336 137472
rect 132644 137420 132696 137472
rect 62632 137216 62684 137268
rect 66404 137216 66456 137268
rect 99708 137216 99760 137268
rect 102192 137216 102244 137268
rect 135128 137216 135180 137268
rect 136876 137216 136928 137268
rect 172664 137216 172716 137268
rect 174044 137216 174096 137268
rect 62724 137148 62776 137200
rect 66312 137148 66364 137200
rect 101456 137148 101508 137200
rect 101916 137148 101968 137200
rect 132644 137148 132696 137200
rect 172572 137080 172624 137132
rect 174136 137080 174188 137132
rect 100628 137012 100680 137064
rect 102376 137012 102428 137064
rect 172204 137012 172256 137064
rect 174228 137012 174280 137064
rect 100536 136740 100588 136792
rect 102652 136740 102704 136792
rect 172664 135992 172716 136044
rect 173952 135992 174004 136044
rect 63000 135856 63052 135908
rect 65668 135856 65720 135908
rect 100904 135856 100956 135908
rect 102008 135856 102060 135908
rect 134300 135856 134352 135908
rect 136968 135856 137020 135908
rect 172664 135856 172716 135908
rect 173768 135856 173820 135908
rect 62908 135788 62960 135840
rect 66404 135788 66456 135840
rect 100628 135788 100680 135840
rect 135312 135788 135364 135840
rect 136876 135788 136928 135840
rect 172572 135788 172624 135840
rect 102376 135720 102428 135772
rect 174228 135720 174280 135772
rect 62816 135652 62868 135704
rect 65024 135652 65076 135704
rect 172756 135652 172808 135704
rect 174136 135652 174188 135704
rect 135220 135380 135272 135432
rect 136784 135380 136836 135432
rect 99892 134632 99944 134684
rect 102284 134632 102336 134684
rect 100904 134564 100956 134616
rect 102100 134564 102152 134616
rect 62724 134496 62776 134548
rect 66220 134496 66272 134548
rect 135128 134496 135180 134548
rect 136968 134496 137020 134548
rect 172664 134496 172716 134548
rect 174044 134496 174096 134548
rect 62816 134428 62868 134480
rect 65852 134428 65904 134480
rect 135404 134428 135456 134480
rect 136876 134428 136928 134480
rect 172572 134428 172624 134480
rect 173860 134428 173912 134480
rect 100996 134360 101048 134412
rect 102376 134360 102428 134412
rect 204772 134360 204824 134412
rect 204956 134360 205008 134412
rect 100904 133204 100956 133256
rect 102008 133204 102060 133256
rect 100260 133136 100312 133188
rect 102192 133136 102244 133188
rect 63460 133068 63512 133120
rect 65484 133068 65536 133120
rect 135220 133068 135272 133120
rect 136968 133068 137020 133120
rect 171652 133068 171704 133120
rect 173216 133068 173268 133120
rect 63552 133000 63604 133052
rect 66404 133000 66456 133052
rect 135312 133000 135364 133052
rect 136876 133000 136928 133052
rect 63092 131708 63144 131760
rect 65668 131708 65720 131760
rect 100904 131708 100956 131760
rect 102100 131708 102152 131760
rect 135036 131708 135088 131760
rect 136968 131708 137020 131760
rect 172020 131708 172072 131760
rect 172756 131708 172808 131760
rect 63644 131640 63696 131692
rect 66404 131640 66456 131692
rect 100260 131640 100312 131692
rect 102284 131640 102336 131692
rect 135404 131640 135456 131692
rect 136876 131640 136928 131692
rect 171652 131640 171704 131692
rect 173032 131640 173084 131692
rect 173124 131572 173176 131624
rect 174136 131572 174188 131624
rect 172940 131300 172992 131352
rect 175056 131300 175108 131352
rect 172756 131028 172808 131080
rect 174136 131028 174188 131080
rect 62816 130756 62868 130808
rect 65024 130756 65076 130808
rect 134300 130756 134352 130808
rect 136784 130756 136836 130808
rect 172388 130552 172440 130604
rect 174044 130552 174096 130604
rect 100260 130416 100312 130468
rect 102284 130416 102336 130468
rect 62908 130348 62960 130400
rect 66404 130348 66456 130400
rect 100904 130348 100956 130400
rect 102008 130348 102060 130400
rect 135128 130348 135180 130400
rect 136968 130348 137020 130400
rect 62724 130280 62776 130332
rect 66312 130280 66364 130332
rect 135312 130280 135364 130332
rect 136876 130280 136928 130332
rect 100996 130212 101048 130264
rect 102376 130212 102428 130264
rect 173032 130212 173084 130264
rect 174136 130212 174188 130264
rect 172848 130144 172900 130196
rect 174504 130144 174556 130196
rect 172664 129192 172716 129244
rect 173952 129192 174004 129244
rect 62632 128988 62684 129040
rect 66404 128988 66456 129040
rect 100260 128988 100312 129040
rect 102100 128988 102152 129040
rect 134300 128988 134352 129040
rect 136968 128988 137020 129040
rect 62816 128920 62868 128972
rect 65484 128920 65536 128972
rect 100904 128920 100956 128972
rect 102192 128920 102244 128972
rect 135220 128920 135272 128972
rect 136876 128920 136928 128972
rect 172664 128920 172716 128972
rect 173860 128920 173912 128972
rect 172756 128852 172808 128904
rect 174136 128852 174188 128904
rect 100076 127832 100128 127884
rect 102284 127832 102336 127884
rect 100812 127560 100864 127612
rect 102008 127560 102060 127612
rect 132644 127560 132696 127612
rect 135128 127560 135180 127612
rect 136876 127560 136928 127612
rect 62908 127492 62960 127544
rect 66404 127492 66456 127544
rect 171652 127492 171704 127544
rect 222804 127492 222856 127544
rect 174228 127424 174280 127476
rect 132644 127356 132696 127408
rect 132736 127399 132788 127408
rect 132736 127365 132745 127399
rect 132745 127365 132779 127399
rect 132779 127365 132788 127399
rect 132736 127356 132788 127365
rect 134668 127152 134720 127204
rect 136784 127152 136836 127204
rect 62816 126880 62868 126932
rect 65024 126880 65076 126932
rect 172388 126336 172440 126388
rect 174044 126336 174096 126388
rect 62724 126200 62776 126252
rect 66312 126200 66364 126252
rect 100628 126200 100680 126252
rect 102284 126200 102336 126252
rect 135404 126200 135456 126252
rect 136968 126200 137020 126252
rect 172664 126200 172716 126252
rect 173860 126200 173912 126252
rect 62632 126132 62684 126184
rect 66404 126132 66456 126184
rect 100536 126132 100588 126184
rect 135312 126132 135364 126184
rect 136876 126132 136928 126184
rect 172020 126132 172072 126184
rect 102376 126064 102428 126116
rect 134852 126064 134904 126116
rect 136784 126064 136836 126116
rect 174136 126064 174188 126116
rect 172756 125996 172808 126048
rect 174228 125996 174280 126048
rect 62816 125520 62868 125572
rect 65024 125520 65076 125572
rect 100628 125112 100680 125164
rect 102100 125112 102152 125164
rect 100628 124840 100680 124892
rect 102008 124840 102060 124892
rect 172664 124840 172716 124892
rect 173952 124840 174004 124892
rect 62908 124772 62960 124824
rect 65852 124772 65904 124824
rect 135128 124772 135180 124824
rect 136876 124772 136928 124824
rect 172020 124772 172072 124824
rect 222712 124815 222764 124824
rect 100996 124704 101048 124756
rect 102376 124704 102428 124756
rect 222712 124781 222721 124815
rect 222721 124781 222755 124815
rect 222755 124781 222764 124815
rect 222712 124772 222764 124781
rect 174228 124704 174280 124756
rect 135220 124364 135272 124416
rect 136784 124364 136836 124416
rect 62816 124092 62868 124144
rect 65024 124092 65076 124144
rect 100628 123616 100680 123668
rect 102284 123616 102336 123668
rect 63552 123344 63604 123396
rect 66404 123344 66456 123396
rect 99892 123344 99944 123396
rect 102192 123344 102244 123396
rect 135404 123344 135456 123396
rect 136876 123344 136928 123396
rect 172388 123344 172440 123396
rect 174044 123344 174096 123396
rect 135312 122868 135364 122920
rect 136784 122868 136836 122920
rect 62816 122596 62868 122648
rect 65024 122596 65076 122648
rect 100168 122188 100220 122240
rect 102284 122188 102336 122240
rect 135128 122120 135180 122172
rect 137060 122120 137112 122172
rect 63460 122052 63512 122104
rect 66312 122052 66364 122104
rect 100904 122052 100956 122104
rect 102100 122052 102152 122104
rect 135220 122052 135272 122104
rect 136968 122052 137020 122104
rect 63644 121984 63696 122036
rect 66404 121984 66456 122036
rect 135312 121916 135364 121968
rect 136876 121984 136928 122036
rect 171560 121984 171612 122036
rect 174136 121916 174188 121968
rect 172848 121780 172900 121832
rect 174320 121780 174372 121832
rect 62816 121440 62868 121492
rect 65024 121440 65076 121492
rect 100628 120896 100680 120948
rect 102284 120896 102336 120948
rect 171744 120896 171796 120948
rect 174044 120896 174096 120948
rect 100628 120624 100680 120676
rect 102192 120624 102244 120676
rect 172664 120624 172716 120676
rect 173952 120624 174004 120676
rect 100996 120556 101048 120608
rect 102376 120556 102428 120608
rect 172940 120556 172992 120608
rect 174136 120556 174188 120608
rect 172756 120488 172808 120540
rect 174320 120488 174372 120540
rect 134852 120216 134904 120268
rect 136784 120216 136836 120268
rect 62816 119944 62868 119996
rect 65024 119944 65076 119996
rect 172664 119536 172716 119588
rect 174044 119536 174096 119588
rect 100628 119400 100680 119452
rect 102284 119400 102336 119452
rect 62908 119264 62960 119316
rect 66404 119264 66456 119316
rect 135220 119264 135272 119316
rect 136968 119264 137020 119316
rect 62724 119128 62776 119180
rect 66220 119128 66272 119180
rect 135312 119060 135364 119112
rect 136876 119060 136928 119112
rect 62816 118720 62868 118772
rect 65024 118720 65076 118772
rect 135036 118652 135088 118704
rect 136784 118652 136836 118704
rect 100628 118312 100680 118364
rect 102192 118312 102244 118364
rect 132644 118244 132696 118296
rect 132736 118108 132788 118160
rect 172664 118040 172716 118092
rect 173952 118040 174004 118092
rect 100628 117904 100680 117956
rect 102284 117904 102336 117956
rect 132736 117947 132788 117956
rect 132736 117913 132745 117947
rect 132745 117913 132779 117947
rect 132779 117913 132788 117947
rect 132736 117904 132788 117913
rect 135312 117904 135364 117956
rect 136876 117904 136928 117956
rect 62724 117836 62776 117888
rect 66404 117836 66456 117888
rect 100996 117768 101048 117820
rect 102376 117768 102428 117820
rect 134116 117768 134168 117820
rect 136968 117836 137020 117888
rect 172020 117836 172072 117888
rect 174044 117836 174096 117888
rect 172756 117768 172808 117820
rect 174136 117768 174188 117820
rect 132644 117743 132696 117752
rect 132644 117709 132653 117743
rect 132653 117709 132687 117743
rect 132687 117709 132696 117743
rect 132644 117700 132696 117709
rect 62816 117292 62868 117344
rect 65024 117292 65076 117344
rect 62816 117156 62868 117208
rect 64932 117156 64984 117208
rect 134668 117156 134720 117208
rect 136784 117156 136836 117208
rect 100628 116612 100680 116664
rect 102192 116612 102244 116664
rect 172572 116544 172624 116596
rect 173860 116544 173912 116596
rect 100536 116476 100588 116528
rect 172664 116476 172716 116528
rect 102376 116408 102428 116460
rect 174228 116408 174280 116460
rect 100720 116340 100772 116392
rect 102468 116340 102520 116392
rect 172480 116340 172532 116392
rect 174136 116340 174188 116392
rect 62816 115728 62868 115780
rect 65024 115728 65076 115780
rect 134484 115728 134536 115780
rect 136784 115728 136836 115780
rect 172664 115592 172716 115644
rect 174044 115592 174096 115644
rect 100628 115184 100680 115236
rect 102284 115184 102336 115236
rect 144880 115116 144932 115168
rect 204772 115116 204824 115168
rect 132644 115048 132696 115100
rect 222620 115048 222672 115100
rect 222988 115048 223040 115100
rect 135312 114980 135364 115032
rect 136876 114980 136928 115032
rect 144880 114912 144932 114964
rect 62816 114844 62868 114896
rect 66404 114844 66456 114896
rect 62816 114572 62868 114624
rect 65024 114572 65076 114624
rect 134852 114436 134904 114488
rect 136784 114436 136836 114488
rect 30432 114300 30484 114352
rect 92716 114300 92768 114352
rect 132092 113756 132144 113808
rect 132460 113688 132512 113740
rect 73212 113620 73264 113672
rect 109460 113620 109512 113672
rect 113508 113620 113560 113672
rect 114382 113620 114434 113672
rect 114520 113620 114572 113672
rect 115486 113620 115538 113672
rect 116636 113620 116688 113672
rect 118798 113620 118850 113672
rect 120132 113620 120184 113672
rect 123122 113620 123174 113672
rect 126296 113620 126348 113672
rect 131954 113620 132006 113672
rect 154816 113620 154868 113672
rect 205048 113620 205100 113672
rect 122708 113552 122760 113604
rect 127032 113552 127084 113604
rect 123076 113416 123128 113468
rect 127492 113416 127544 113468
rect 123904 113348 123956 113400
rect 128596 113348 128648 113400
rect 124640 113280 124692 113332
rect 129700 113280 129752 113332
rect 122248 113212 122300 113264
rect 126388 113212 126440 113264
rect 81676 113144 81728 113196
rect 82504 113144 82556 113196
rect 116268 113144 116320 113196
rect 118200 113144 118252 113196
rect 125468 113144 125520 113196
rect 130804 113144 130856 113196
rect 188948 113144 189000 113196
rect 189684 113144 189736 113196
rect 113876 113076 113928 113128
rect 114888 113076 114940 113128
rect 115072 113076 115124 113128
rect 116544 113076 116596 113128
rect 121880 113076 121932 113128
rect 125836 113076 125888 113128
rect 183980 113076 184032 113128
rect 184440 113076 184492 113128
rect 188488 113076 188540 113128
rect 189132 113076 189184 113128
rect 195756 113076 195808 113128
rect 199344 113076 199396 113128
rect 115440 113008 115492 113060
rect 117096 113008 117148 113060
rect 125100 113008 125152 113060
rect 130252 113008 130304 113060
rect 193732 113008 193784 113060
rect 196492 113008 196544 113060
rect 125836 112940 125888 112992
rect 131356 112940 131408 112992
rect 196124 112940 196176 112992
rect 199988 112940 200040 112992
rect 114704 112872 114756 112924
rect 115992 112872 116044 112924
rect 124272 112872 124324 112924
rect 129148 112872 129200 112924
rect 191340 112872 191392 112924
rect 193088 112872 193140 112924
rect 123444 112804 123496 112856
rect 128044 112804 128096 112856
rect 117832 112736 117884 112788
rect 120224 112736 120276 112788
rect 126664 112736 126716 112788
rect 132552 112736 132604 112788
rect 188028 112736 188080 112788
rect 188580 112736 188632 112788
rect 192904 112736 192956 112788
rect 195388 112736 195440 112788
rect 196492 112736 196544 112788
rect 200540 112736 200592 112788
rect 197320 112668 197372 112720
rect 201644 112668 201696 112720
rect 189224 112600 189276 112652
rect 190236 112600 190288 112652
rect 192536 112600 192588 112652
rect 194744 112600 194796 112652
rect 196952 112600 197004 112652
rect 201092 112600 201144 112652
rect 121512 112532 121564 112584
rect 125284 112532 125336 112584
rect 197412 112532 197464 112584
rect 202196 112532 202248 112584
rect 121052 112464 121104 112516
rect 124732 112464 124784 112516
rect 189592 112464 189644 112516
rect 190788 112464 190840 112516
rect 198148 112464 198200 112516
rect 202840 112464 202892 112516
rect 120316 112396 120368 112448
rect 113048 112328 113100 112380
rect 113784 112328 113836 112380
rect 119120 112328 119172 112380
rect 81676 112260 81728 112312
rect 110472 112260 110524 112312
rect 121972 112260 122024 112312
rect 190512 112396 190564 112448
rect 191984 112396 192036 112448
rect 194560 112396 194612 112448
rect 197688 112396 197740 112448
rect 198884 112396 198936 112448
rect 190144 112328 190196 112380
rect 191432 112328 191484 112380
rect 191708 112328 191760 112380
rect 123628 112260 123680 112312
rect 193180 112328 193232 112380
rect 193640 112260 193692 112312
rect 194744 112328 194796 112380
rect 198240 112328 198292 112380
rect 198516 112328 198568 112380
rect 195940 112260 195992 112312
rect 203392 112260 203444 112312
rect 203944 112260 203996 112312
rect 109460 112192 109512 112244
rect 132460 112192 132512 112244
rect 34480 112124 34532 112176
rect 39448 112124 39500 112176
rect 52604 112124 52656 112176
rect 57020 112124 57072 112176
rect 110012 112124 110064 112176
rect 164476 112124 164528 112176
rect 51040 112056 51092 112108
rect 54260 112056 54312 112108
rect 116176 112056 116228 112108
rect 117648 112056 117700 112108
rect 120960 112056 121012 112108
rect 124180 112056 124232 112108
rect 190604 112056 190656 112108
rect 192444 112056 192496 112108
rect 53064 111988 53116 112040
rect 57664 111988 57716 112040
rect 51868 111920 51920 111972
rect 55640 111920 55692 111972
rect 35216 111852 35268 111904
rect 39816 111852 39868 111904
rect 52512 111852 52564 111904
rect 56376 111852 56428 111904
rect 53800 111784 53852 111836
rect 59044 111784 59096 111836
rect 54260 111716 54312 111768
rect 59780 111716 59832 111768
rect 35860 111648 35912 111700
rect 40276 111648 40328 111700
rect 53432 111648 53484 111700
rect 58400 111648 58452 111700
rect 33836 111580 33888 111632
rect 39080 111580 39132 111632
rect 54628 111580 54680 111632
rect 60424 111580 60476 111632
rect 37884 111512 37936 111564
rect 41472 111512 41524 111564
rect 39264 111444 39316 111496
rect 42208 111444 42260 111496
rect 118844 111444 118896 111496
rect 121420 111444 121472 111496
rect 40000 111376 40052 111428
rect 42300 111376 42352 111428
rect 48280 111376 48332 111428
rect 49476 111376 49528 111428
rect 50672 111376 50724 111428
rect 53616 111376 53668 111428
rect 117464 111376 117516 111428
rect 119764 111376 119816 111428
rect 182232 111376 182284 111428
rect 183244 111376 183296 111428
rect 194100 111376 194152 111428
rect 197136 111376 197188 111428
rect 40644 111308 40696 111360
rect 43036 111308 43088 111360
rect 43404 111308 43456 111360
rect 44600 111308 44652 111360
rect 47820 111308 47872 111360
rect 48832 111308 48884 111360
rect 49844 111308 49896 111360
rect 52236 111308 52288 111360
rect 117372 111308 117424 111360
rect 119212 111308 119264 111360
rect 182876 111308 182928 111360
rect 183796 111308 183848 111360
rect 191984 111308 192036 111360
rect 194284 111308 194336 111360
rect 195296 111308 195348 111360
rect 198792 111308 198844 111360
rect 37240 111240 37292 111292
rect 41012 111240 41064 111292
rect 48648 111240 48700 111292
rect 50212 111240 50264 111292
rect 51408 111240 51460 111292
rect 54996 111240 55048 111292
rect 118568 111240 118620 111292
rect 120868 111240 120920 111292
rect 36596 111172 36648 111224
rect 40644 111172 40696 111224
rect 41288 111172 41340 111224
rect 43404 111172 43456 111224
rect 44324 111172 44376 111224
rect 45060 111172 45112 111224
rect 49476 111172 49528 111224
rect 51592 111172 51644 111224
rect 105228 111172 105280 111224
rect 106608 111172 106660 111224
rect 119764 111172 119816 111224
rect 122524 111172 122576 111224
rect 177264 111172 177316 111224
rect 178276 111172 178328 111224
rect 42024 111104 42076 111156
rect 43864 111104 43916 111156
rect 50212 111104 50264 111156
rect 52972 111104 53024 111156
rect 105504 111104 105556 111156
rect 107160 111104 107212 111156
rect 177080 111104 177132 111156
rect 178828 111104 178880 111156
rect 38620 111036 38672 111088
rect 41840 111036 41892 111088
rect 49016 111036 49068 111088
rect 50856 111036 50908 111088
rect 105688 111036 105740 111088
rect 107712 111036 107764 111088
rect 176896 111036 176948 111088
rect 179380 111036 179432 111088
rect 42668 110968 42720 111020
rect 44232 110968 44284 111020
rect 105964 110900 106016 110952
rect 108816 110968 108868 111020
rect 176988 110968 177040 111020
rect 180024 110968 180076 111020
rect 181680 110968 181732 111020
rect 183106 110968 183158 111020
rect 183428 110968 183480 111020
rect 184302 110968 184354 111020
rect 177724 110900 177776 110952
rect 181128 110900 181180 110952
rect 132552 110220 132604 110272
rect 222712 110220 222764 110272
rect 105780 109472 105832 109524
rect 108264 109472 108316 109524
rect 177356 108996 177408 109048
rect 180576 108996 180628 109048
rect 222804 107951 222856 107960
rect 222804 107917 222813 107951
rect 222813 107917 222847 107951
rect 222847 107917 222856 107951
rect 222804 107908 222856 107917
rect 32640 104032 32692 104084
rect 37424 104032 37476 104084
rect 105688 104032 105740 104084
rect 107896 104032 107948 104084
rect 178184 104032 178236 104084
rect 179656 104032 179708 104084
rect 106332 101312 106384 101364
rect 107896 101312 107948 101364
rect 177632 101312 177684 101364
rect 179656 101312 179708 101364
rect 57572 100972 57624 101024
rect 60516 100972 60568 101024
rect 105964 100768 106016 100820
rect 108632 100768 108684 100820
rect 176988 100768 177040 100820
rect 180300 100768 180352 100820
rect 106424 99884 106476 99936
rect 107896 99884 107948 99936
rect 177724 99884 177776 99936
rect 179656 99884 179708 99936
rect 105596 99408 105648 99460
rect 108540 99408 108592 99460
rect 177356 99272 177408 99324
rect 180392 99272 180444 99324
rect 105780 97164 105832 97216
rect 107896 97164 107948 97216
rect 177540 97164 177592 97216
rect 179656 97164 179708 97216
rect 222988 97096 223040 97148
rect 223540 97096 223592 97148
rect 105780 94308 105832 94360
rect 107804 94308 107856 94360
rect 177356 93900 177408 93952
rect 179564 93900 179616 93952
rect 222804 92540 222856 92592
rect 223540 92540 223592 92592
rect 105228 92064 105280 92116
rect 107804 92064 107856 92116
rect 176988 91996 177040 92048
rect 179564 91996 179616 92048
rect 201092 91588 201144 91640
rect 204496 91588 204548 91640
rect 28868 90228 28920 90280
rect 36412 90228 36464 90280
rect 59596 90228 59648 90280
rect 105780 89208 105832 89260
rect 107804 89208 107856 89260
rect 132368 88868 132420 88920
rect 132552 88800 132604 88852
rect 105412 87848 105464 87900
rect 107896 87848 107948 87900
rect 177356 87508 177408 87560
rect 179656 87508 179708 87560
rect 106424 86352 106476 86404
rect 107988 86352 108040 86404
rect 54812 86123 54864 86132
rect 54812 86089 54821 86123
rect 54821 86089 54855 86123
rect 54855 86089 54864 86123
rect 54812 86080 54864 86089
rect 177540 86080 177592 86132
rect 179748 86080 179800 86132
rect 54812 85987 54864 85996
rect 54812 85953 54821 85987
rect 54821 85953 54855 85987
rect 54855 85953 54864 85987
rect 54812 85944 54864 85953
rect 105136 84788 105188 84840
rect 107804 84788 107856 84840
rect 176988 84788 177040 84840
rect 179564 84788 179616 84840
rect 222804 84788 222856 84840
rect 223540 84788 223592 84840
rect 105688 84720 105740 84772
rect 107620 84720 107672 84772
rect 178184 84720 178236 84772
rect 179656 84720 179708 84772
rect 178092 83428 178144 83480
rect 179472 83428 179524 83480
rect 105228 83360 105280 83412
rect 107712 83360 107764 83412
rect 177724 82272 177776 82324
rect 179748 82272 179800 82324
rect 106424 82136 106476 82188
rect 107896 82136 107948 82188
rect 105964 80776 106016 80828
rect 108540 80776 108592 80828
rect 178092 80572 178144 80624
rect 180300 80572 180352 80624
rect 132552 79280 132604 79332
rect 105412 79212 105464 79264
rect 108080 79212 108132 79264
rect 177632 79212 177684 79264
rect 180024 79212 180076 79264
rect 132552 79144 132604 79196
rect 105228 77852 105280 77904
rect 107528 77852 107580 77904
rect 176988 77852 177040 77904
rect 179380 77852 179432 77904
rect 30524 77784 30576 77836
rect 37424 77784 37476 77836
rect 57480 77580 57532 77632
rect 59596 77580 59648 77632
rect 54996 76424 55048 76476
rect 222988 75064 223040 75116
rect 223540 75064 223592 75116
rect 222804 73568 222856 73620
rect 223080 73568 223132 73620
rect 105872 72412 105924 72464
rect 109184 72412 109236 72464
rect 177632 72344 177684 72396
rect 180944 72344 180996 72396
rect 177356 70916 177408 70968
rect 180576 70848 180628 70900
rect 189822 70712 189874 70764
rect 191432 70712 191484 70764
rect 182876 70644 182928 70696
rect 183842 70644 183894 70696
rect 189454 70644 189506 70696
rect 190788 70644 190840 70696
rect 191846 70644 191898 70696
rect 194284 70644 194336 70696
rect 106516 70304 106568 70356
rect 108356 70304 108408 70356
rect 49476 69760 49528 69812
rect 51592 69760 51644 69812
rect 119856 69760 119908 69812
rect 122340 69760 122392 69812
rect 48648 69692 48700 69744
rect 50212 69692 50264 69744
rect 119488 69692 119540 69744
rect 121696 69692 121748 69744
rect 48280 69624 48332 69676
rect 49476 69624 49528 69676
rect 49844 69624 49896 69676
rect 52236 69624 52288 69676
rect 117096 69624 117148 69676
rect 118200 69624 118252 69676
rect 118660 69624 118712 69676
rect 120592 69624 120644 69676
rect 191708 69624 191760 69676
rect 193640 69624 193692 69676
rect 39264 69556 39316 69608
rect 22244 69488 22296 69540
rect 28684 69488 28736 69540
rect 16632 69420 16684 69472
rect 31904 69420 31956 69472
rect 36044 69488 36096 69540
rect 40276 69488 40328 69540
rect 47820 69556 47872 69608
rect 48832 69556 48884 69608
rect 49016 69556 49068 69608
rect 50856 69556 50908 69608
rect 42208 69488 42260 69540
rect 35584 69420 35636 69472
rect 39816 69420 39868 69472
rect 34664 69352 34716 69404
rect 39448 69352 39500 69404
rect 27580 69284 27632 69336
rect 54996 69556 55048 69608
rect 53800 69488 53852 69540
rect 59044 69556 59096 69608
rect 116636 69556 116688 69608
rect 117648 69556 117700 69608
rect 118292 69556 118344 69608
rect 120316 69556 120368 69608
rect 126296 69488 126348 69540
rect 131632 69556 131684 69608
rect 190420 69556 190472 69608
rect 191984 69556 192036 69608
rect 198884 69488 198936 69540
rect 203944 69556 203996 69608
rect 201000 69488 201052 69540
rect 215904 69488 215956 69540
rect 53432 69420 53484 69472
rect 58124 69420 58176 69472
rect 123444 69420 123496 69472
rect 127584 69420 127636 69472
rect 198516 69420 198568 69472
rect 203024 69420 203076 69472
rect 57480 69352 57532 69404
rect 124640 69352 124692 69404
rect 129332 69352 129384 69404
rect 196124 69352 196176 69404
rect 199988 69352 200040 69404
rect 51868 69284 51920 69336
rect 91244 69284 91296 69336
rect 132092 69284 132144 69336
rect 194560 69284 194612 69336
rect 197688 69284 197740 69336
rect 201092 69284 201144 69336
rect 210568 69284 210620 69336
rect 121880 69216 121932 69268
rect 125192 69216 125244 69268
rect 125468 69216 125520 69268
rect 130436 69216 130488 69268
rect 196492 69216 196544 69268
rect 200540 69216 200592 69268
rect 40184 69148 40236 69200
rect 42668 69148 42720 69200
rect 54628 69148 54680 69200
rect 60148 69148 60200 69200
rect 92348 69148 92400 69200
rect 97500 69148 97552 69200
rect 122248 69148 122300 69200
rect 34112 69080 34164 69132
rect 39080 69080 39132 69132
rect 40644 69080 40696 69132
rect 43036 69080 43088 69132
rect 52604 69080 52656 69132
rect 56744 69080 56796 69132
rect 110564 69080 110616 69132
rect 111484 69080 111536 69132
rect 121052 69080 121104 69132
rect 124456 69080 124508 69132
rect 125836 69148 125888 69200
rect 131264 69148 131316 69200
rect 125928 69080 125980 69132
rect 126664 69080 126716 69132
rect 132184 69080 132236 69132
rect 36596 69012 36648 69064
rect 40368 69012 40420 69064
rect 42024 69012 42076 69064
rect 43864 69012 43916 69064
rect 53064 69012 53116 69064
rect 57664 69012 57716 69064
rect 125100 69012 125152 69064
rect 129884 69012 129936 69064
rect 37240 68944 37292 68996
rect 41012 68944 41064 68996
rect 42668 68944 42720 68996
rect 44232 68944 44284 68996
rect 52512 68944 52564 68996
rect 41288 68876 41340 68928
rect 43404 68876 43456 68928
rect 50672 68876 50724 68928
rect 53616 68876 53668 68928
rect 54260 68944 54312 68996
rect 59504 68944 59556 68996
rect 62908 68944 62960 68996
rect 67876 68944 67928 68996
rect 88944 68944 88996 68996
rect 96856 68944 96908 68996
rect 122708 68944 122760 68996
rect 126388 68944 126440 68996
rect 160980 68944 161032 68996
rect 168892 69148 168944 69200
rect 192536 69148 192588 69200
rect 194836 69148 194888 69200
rect 196952 69148 197004 69200
rect 201092 69148 201144 69200
rect 192904 69080 192956 69132
rect 195388 69080 195440 69132
rect 197412 69080 197464 69132
rect 201828 69080 201880 69132
rect 167696 69012 167748 69064
rect 174136 69012 174188 69064
rect 194100 69012 194152 69064
rect 197136 69012 197188 69064
rect 197320 69012 197372 69064
rect 201644 69012 201696 69064
rect 166592 68944 166644 68996
rect 174228 68944 174280 68996
rect 181680 68944 181732 68996
rect 182784 68944 182836 68996
rect 193364 68944 193416 68996
rect 195940 68944 195992 68996
rect 198148 68944 198200 68996
rect 202840 68944 202892 68996
rect 38620 68808 38672 68860
rect 41840 68808 41892 68860
rect 51040 68808 51092 68860
rect 54260 68808 54312 68860
rect 37884 68740 37936 68792
rect 41472 68740 41524 68792
rect 51408 68740 51460 68792
rect 54996 68740 55048 68792
rect 83424 68876 83476 68928
rect 87196 68876 87248 68928
rect 87840 68876 87892 68928
rect 94740 68876 94792 68928
rect 120500 68876 120552 68928
rect 123076 68876 123128 68928
rect 124272 68876 124324 68928
rect 128688 68876 128740 68928
rect 151044 68876 151096 68928
rect 152056 68876 152108 68928
rect 159876 68876 159928 68928
rect 55640 68808 55692 68860
rect 62724 68808 62776 68860
rect 68980 68808 69032 68860
rect 82320 68808 82372 68860
rect 85356 68808 85408 68860
rect 93452 68808 93504 68860
rect 102560 68808 102612 68860
rect 110104 68808 110156 68860
rect 111116 68808 111168 68860
rect 116268 68808 116320 68860
rect 117096 68808 117148 68860
rect 117464 68808 117516 68860
rect 118936 68808 118988 68860
rect 123352 68808 123404 68860
rect 127308 68808 127360 68860
rect 140832 68808 140884 68860
rect 144328 68808 144380 68860
rect 158772 68808 158824 68860
rect 165120 68808 165172 68860
rect 168800 68876 168852 68928
rect 173860 68876 173912 68928
rect 193732 68876 193784 68928
rect 196492 68876 196544 68928
rect 167052 68808 167104 68860
rect 169904 68808 169956 68860
rect 173952 68808 174004 68860
rect 195756 68808 195808 68860
rect 199344 68808 199396 68860
rect 205140 68808 205192 68860
rect 221240 68808 221292 68860
rect 56376 68740 56428 68792
rect 120684 68740 120736 68792
rect 123444 68740 123496 68792
rect 132552 68740 132604 68792
rect 165488 68740 165540 68792
rect 174412 68740 174464 68792
rect 190604 68740 190656 68792
rect 192536 68740 192588 68792
rect 195296 68740 195348 68792
rect 198792 68740 198844 68792
rect 43404 68672 43456 68724
rect 44600 68672 44652 68724
rect 50488 68672 50540 68724
rect 52972 68672 53024 68724
rect 102284 68672 102336 68724
rect 174320 68672 174372 68724
rect 101180 68604 101232 68656
rect 173216 68604 173268 68656
rect 194652 68604 194704 68656
rect 198240 68604 198292 68656
rect 90140 68536 90192 68588
rect 123904 68536 123956 68588
rect 128136 68536 128188 68588
rect 182232 68536 182284 68588
rect 183244 68536 183296 68588
rect 97868 68468 97920 68520
rect 102376 68468 102428 68520
rect 121512 68468 121564 68520
rect 124640 68468 124692 68520
rect 74592 68400 74644 68452
rect 75604 68400 75656 68452
rect 94556 68400 94608 68452
rect 102652 68400 102704 68452
rect 86736 68332 86788 68384
rect 92808 68332 92860 68384
rect 95660 68332 95712 68384
rect 102744 68332 102796 68384
rect 155460 68332 155512 68384
rect 159508 68332 159560 68384
rect 63000 68264 63052 68316
rect 64564 68264 64616 68316
rect 71004 68264 71056 68316
rect 73396 68264 73448 68316
rect 81216 68264 81268 68316
rect 83516 68264 83568 68316
rect 85632 68264 85684 68316
rect 90968 68264 91020 68316
rect 96764 68264 96816 68316
rect 102468 68264 102520 68316
rect 144512 68264 144564 68316
rect 146536 68264 146588 68316
rect 153252 68264 153304 68316
rect 155828 68264 155880 68316
rect 156564 68264 156616 68316
rect 161440 68264 161492 68316
rect 62356 68196 62408 68248
rect 63460 68196 63512 68248
rect 69164 68196 69216 68248
rect 72292 68196 72344 68248
rect 72844 68196 72896 68248
rect 74500 68196 74552 68248
rect 80112 68196 80164 68248
rect 81676 68196 81728 68248
rect 84528 68196 84580 68248
rect 89128 68196 89180 68248
rect 98972 68196 99024 68248
rect 63368 68128 63420 68180
rect 71188 68128 71240 68180
rect 134484 68196 134536 68248
rect 136600 68196 136652 68248
rect 142672 68196 142724 68248
rect 145432 68196 145484 68248
rect 146444 68196 146496 68248
rect 147640 68196 147692 68248
rect 152148 68196 152200 68248
rect 153896 68196 153948 68248
rect 154356 68196 154408 68248
rect 157668 68196 157720 68248
rect 157944 68196 157996 68248
rect 163280 68264 163332 68316
rect 171008 68264 171060 68316
rect 174044 68264 174096 68316
rect 164384 68196 164436 68248
rect 169444 68196 169496 68248
rect 172112 68196 172164 68248
rect 102928 68128 102980 68180
rect 135312 68128 135364 68180
rect 143224 68128 143276 68180
rect 175056 68128 175108 68180
rect 135036 68060 135088 68112
rect 142120 68060 142172 68112
rect 100076 67652 100128 67704
rect 103480 67652 103532 67704
rect 62816 66700 62868 66752
rect 70084 66700 70136 66752
rect 134668 66700 134720 66752
rect 139912 66700 139964 66752
rect 135312 66428 135364 66480
rect 141016 66428 141068 66480
rect 63368 65544 63420 65596
rect 66404 65544 66456 65596
rect 172664 65544 172716 65596
rect 175332 65544 175384 65596
rect 100904 65408 100956 65460
rect 102376 65408 102428 65460
rect 134668 65408 134720 65460
rect 136876 65408 136928 65460
rect 62816 65340 62868 65392
rect 66312 65340 66364 65392
rect 134852 65340 134904 65392
rect 137704 65340 137756 65392
rect 62724 65272 62776 65324
rect 65668 65272 65720 65324
rect 135312 65204 135364 65256
rect 138164 65204 138216 65256
rect 100628 64456 100680 64508
rect 102744 64456 102796 64508
rect 63552 64320 63604 64372
rect 66404 64320 66456 64372
rect 172664 64320 172716 64372
rect 174228 64320 174280 64372
rect 63460 64184 63512 64236
rect 65668 64184 65720 64236
rect 135312 64116 135364 64168
rect 136968 64116 137020 64168
rect 100904 64048 100956 64100
rect 102468 64048 102520 64100
rect 134852 64048 134904 64100
rect 136876 64048 136928 64100
rect 171836 64048 171888 64100
rect 175240 64048 175292 64100
rect 169444 63980 169496 64032
rect 174136 63980 174188 64032
rect 97500 63776 97552 63828
rect 102560 63776 102612 63828
rect 172664 62960 172716 63012
rect 174136 62960 174188 63012
rect 100628 62824 100680 62876
rect 102376 62824 102428 62876
rect 62724 62688 62776 62740
rect 65668 62688 65720 62740
rect 100628 62688 100680 62740
rect 102560 62688 102612 62740
rect 134484 62688 134536 62740
rect 136968 62688 137020 62740
rect 172664 62688 172716 62740
rect 174320 62688 174372 62740
rect 13320 62620 13372 62672
rect 29236 62620 29288 62672
rect 62816 62620 62868 62672
rect 66404 62620 66456 62672
rect 135404 62620 135456 62672
rect 136876 62620 136928 62672
rect 62908 61464 62960 61516
rect 65668 61464 65720 61516
rect 172664 61464 172716 61516
rect 174228 61464 174280 61516
rect 100628 61328 100680 61380
rect 102468 61328 102520 61380
rect 63736 61260 63788 61312
rect 66404 61260 66456 61312
rect 100536 61260 100588 61312
rect 102744 61260 102796 61312
rect 135312 61260 135364 61312
rect 136876 61260 136928 61312
rect 171836 61260 171888 61312
rect 174412 61260 174464 61312
rect 135036 60920 135088 60972
rect 136784 60920 136836 60972
rect 63828 60580 63880 60632
rect 65484 60580 65536 60632
rect 100628 60376 100680 60428
rect 102652 60376 102704 60428
rect 100628 60240 100680 60292
rect 102376 60240 102428 60292
rect 172664 60240 172716 60292
rect 174320 60240 174372 60292
rect 62632 60104 62684 60156
rect 66404 60104 66456 60156
rect 172204 60104 172256 60156
rect 174136 60104 174188 60156
rect 134484 60036 134536 60088
rect 136968 60036 137020 60088
rect 100628 59968 100680 60020
rect 102560 59968 102612 60020
rect 172664 59968 172716 60020
rect 174504 59968 174556 60020
rect 62724 59900 62776 59952
rect 66312 59900 66364 59952
rect 135404 59900 135456 59952
rect 136876 59900 136928 59952
rect 135036 59832 135088 59884
rect 136784 59832 136836 59884
rect 172204 58880 172256 58932
rect 174596 58880 174648 58932
rect 100628 58744 100680 58796
rect 102468 58744 102520 58796
rect 171836 58744 171888 58796
rect 174228 58744 174280 58796
rect 62816 58608 62868 58660
rect 66312 58608 66364 58660
rect 100628 58608 100680 58660
rect 102652 58608 102704 58660
rect 62908 58540 62960 58592
rect 66404 58540 66456 58592
rect 135312 58540 135364 58592
rect 136876 58540 136928 58592
rect 135036 58404 135088 58456
rect 136784 58404 136836 58456
rect 62724 57384 62776 57436
rect 66404 57384 66456 57436
rect 100628 57384 100680 57436
rect 102376 57384 102428 57436
rect 172664 57384 172716 57436
rect 174320 57384 174372 57436
rect 172664 57248 172716 57300
rect 174412 57248 174464 57300
rect 100628 57180 100680 57232
rect 102468 57180 102520 57232
rect 135404 57180 135456 57232
rect 136968 57180 137020 57232
rect 62632 57112 62684 57164
rect 66404 57112 66456 57164
rect 100536 57112 100588 57164
rect 102560 57112 102612 57164
rect 134760 57112 134812 57164
rect 136876 57112 136928 57164
rect 172020 57112 172072 57164
rect 174136 57112 174188 57164
rect 135036 57044 135088 57096
rect 136784 57044 136836 57096
rect 62540 56976 62592 57028
rect 65024 56976 65076 57028
rect 63644 56296 63696 56348
rect 66404 56296 66456 56348
rect 172664 56024 172716 56076
rect 174228 56024 174280 56076
rect 63276 55888 63328 55940
rect 66404 55888 66456 55940
rect 100628 55888 100680 55940
rect 102376 55888 102428 55940
rect 100904 55752 100956 55804
rect 102652 55752 102704 55804
rect 134208 55752 134260 55804
rect 136876 55752 136928 55804
rect 172664 55752 172716 55804
rect 174964 55752 175016 55804
rect 135036 55412 135088 55464
rect 136784 55412 136836 55464
rect 100628 54800 100680 54852
rect 102468 54800 102520 54852
rect 63368 54664 63420 54716
rect 66404 54664 66456 54716
rect 100812 54528 100864 54580
rect 102560 54528 102612 54580
rect 134300 54528 134352 54580
rect 137152 54528 137204 54580
rect 172112 54528 172164 54580
rect 174780 54528 174832 54580
rect 172664 54460 172716 54512
rect 175332 54460 175384 54512
rect 63552 54392 63604 54444
rect 66312 54392 66364 54444
rect 135128 53916 135180 53968
rect 136784 53916 136836 53968
rect 62816 53304 62868 53356
rect 65300 53304 65352 53356
rect 100628 53236 100680 53288
rect 102744 53236 102796 53288
rect 171652 53168 171704 53220
rect 174136 53168 174188 53220
rect 100628 53032 100680 53084
rect 102376 53032 102428 53084
rect 172664 53032 172716 53084
rect 174504 53032 174556 53084
rect 63736 52964 63788 53016
rect 66404 52964 66456 53016
rect 135404 52964 135456 53016
rect 136876 52964 136928 53016
rect 135128 52556 135180 52608
rect 136784 52556 136836 52608
rect 100628 52216 100680 52268
rect 102652 52216 102704 52268
rect 63368 52080 63420 52132
rect 65300 52080 65352 52132
rect 172572 51944 172624 51996
rect 174320 51944 174372 51996
rect 172664 51808 172716 51860
rect 174412 51808 174464 51860
rect 62724 51672 62776 51724
rect 65668 51672 65720 51724
rect 100628 51672 100680 51724
rect 102468 51672 102520 51724
rect 63736 51604 63788 51656
rect 66312 51604 66364 51656
rect 100536 51604 100588 51656
rect 102560 51604 102612 51656
rect 135312 51604 135364 51656
rect 136876 51604 136928 51656
rect 172020 51604 172072 51656
rect 174228 51604 174280 51656
rect 135036 51332 135088 51384
rect 136784 51332 136836 51384
rect 135404 51060 135456 51112
rect 136692 51060 136744 51112
rect 63828 50584 63880 50636
rect 66404 50584 66456 50636
rect 62816 50448 62868 50500
rect 65668 50448 65720 50500
rect 100628 50448 100680 50500
rect 102652 50448 102704 50500
rect 100628 50312 100680 50364
rect 102376 50312 102428 50364
rect 172204 50312 172256 50364
rect 174136 50312 174188 50364
rect 135404 50244 135456 50296
rect 136876 50244 136928 50296
rect 172664 50244 172716 50296
rect 174320 50244 174372 50296
rect 134852 50176 134904 50228
rect 136784 50176 136836 50228
rect 100628 49224 100680 49276
rect 102468 49224 102520 49276
rect 172664 49224 172716 49276
rect 174228 49224 174280 49276
rect 171836 49088 171888 49140
rect 174412 49088 174464 49140
rect 63736 48952 63788 49004
rect 65484 48952 65536 49004
rect 100628 48952 100680 49004
rect 102560 48952 102612 49004
rect 63368 48884 63420 48936
rect 66404 48884 66456 48936
rect 135312 48816 135364 48868
rect 136876 48884 136928 48936
rect 134760 48408 134812 48460
rect 136784 48408 136836 48460
rect 100628 47864 100680 47916
rect 102652 47864 102704 47916
rect 172572 47864 172624 47916
rect 174228 47864 174280 47916
rect 172664 47728 172716 47780
rect 174136 47728 174188 47780
rect 100628 47592 100680 47644
rect 102376 47592 102428 47644
rect 172664 47592 172716 47644
rect 174320 47592 174372 47644
rect 62816 47456 62868 47508
rect 65668 47456 65720 47508
rect 100628 47456 100680 47508
rect 102468 47456 102520 47508
rect 135404 47456 135456 47508
rect 136876 47456 136928 47508
rect 62908 47388 62960 47440
rect 64932 47388 64984 47440
rect 134852 47320 134904 47372
rect 136784 47320 136836 47372
rect 135312 47116 135364 47168
rect 136692 47116 136744 47168
rect 62724 46912 62776 46964
rect 65024 46912 65076 46964
rect 172664 46504 172716 46556
rect 174228 46504 174280 46556
rect 63736 46368 63788 46420
rect 66404 46368 66456 46420
rect 100628 46232 100680 46284
rect 102560 46232 102612 46284
rect 100904 46096 100956 46148
rect 102376 46096 102428 46148
rect 172664 46096 172716 46148
rect 175332 46096 175384 46148
rect 134668 46028 134720 46080
rect 136784 46028 136836 46080
rect 100536 45212 100588 45264
rect 102468 45212 102520 45264
rect 99984 44940 100036 44992
rect 102560 44940 102612 44992
rect 171652 44940 171704 44992
rect 175424 44940 175476 44992
rect 63736 44804 63788 44856
rect 66312 44804 66364 44856
rect 63644 44736 63696 44788
rect 66404 44736 66456 44788
rect 171836 44736 171888 44788
rect 174780 44736 174832 44788
rect 62816 44668 62868 44720
rect 65208 44668 65260 44720
rect 135036 44668 135088 44720
rect 137520 44668 137572 44720
rect 135404 44396 135456 44448
rect 136692 44396 136744 44448
rect 135036 44260 135088 44312
rect 136784 44260 136836 44312
rect 99892 44056 99944 44108
rect 102284 44056 102336 44108
rect 172664 43580 172716 43632
rect 174044 43580 174096 43632
rect 63736 43512 63788 43564
rect 66220 43512 66272 43564
rect 63828 43308 63880 43360
rect 66404 43308 66456 43360
rect 100628 43308 100680 43360
rect 102376 43240 102428 43292
rect 134944 43240 134996 43292
rect 136876 43308 136928 43360
rect 172572 43308 172624 43360
rect 174136 43240 174188 43292
rect 135404 43036 135456 43088
rect 136784 43036 136836 43088
rect 100628 42628 100680 42680
rect 102560 42628 102612 42680
rect 63828 42288 63880 42340
rect 66404 42288 66456 42340
rect 172204 42288 172256 42340
rect 174228 42288 174280 42340
rect 100628 42152 100680 42204
rect 102468 42152 102520 42204
rect 172664 42152 172716 42204
rect 174320 42152 174372 42204
rect 100628 42016 100680 42068
rect 102376 42016 102428 42068
rect 172664 42016 172716 42068
rect 174136 42016 174188 42068
rect 63736 41948 63788 42000
rect 66312 41948 66364 42000
rect 135404 41880 135456 41932
rect 136876 41948 136928 42000
rect 135312 41812 135364 41864
rect 136692 41812 136744 41864
rect 134852 41472 134904 41524
rect 136784 41472 136836 41524
rect 63184 40520 63236 40572
rect 66404 40520 66456 40572
rect 71924 39908 71976 39960
rect 82504 39908 82556 39960
rect 143592 39908 143644 39960
rect 154816 39908 154868 39960
rect 66312 39840 66364 39892
rect 86276 39840 86328 39892
rect 138072 39840 138124 39892
rect 158588 39840 158640 39892
rect 62816 39160 62868 39212
rect 72568 39160 72620 39212
rect 93176 39160 93228 39212
rect 102376 39160 102428 39212
rect 134484 39160 134536 39212
rect 144880 39160 144932 39212
rect 164844 39160 164896 39212
rect 174136 39160 174188 39212
rect 79376 37732 79428 37784
rect 127768 37732 127820 37784
rect 151044 37732 151096 37784
rect 200080 37732 200132 37784
rect 222528 37775 222580 37784
rect 222528 37741 222537 37775
rect 222537 37741 222571 37775
rect 222571 37741 222580 37775
rect 222528 37732 222580 37741
rect 190788 37664 190840 37716
rect 205140 37664 205192 37716
rect 30524 33584 30576 33636
rect 66220 33584 66272 33636
rect 118844 33584 118896 33636
rect 136876 33584 136928 33636
rect 222712 28144 222764 28196
rect 77996 12572 78048 12624
rect 79054 12572 79106 12624
rect 86920 11688 86972 11740
rect 132552 11688 132604 11740
rect 166040 11688 166092 11740
rect 214248 11688 214300 11740
rect 94004 11620 94056 11672
rect 187016 11620 187068 11672
rect 23532 10940 23584 10992
rect 71280 10940 71332 10992
rect 105228 10940 105280 10992
rect 151044 10940 151096 10992
rect 50764 10872 50816 10924
rect 143592 10872 143644 10924
rect 158588 10396 158640 10448
rect 159784 10396 159836 10448
<< metal2 >>
rect 23530 246344 23586 246824
rect 50762 246344 50818 246824
rect 77994 246344 78050 246824
rect 105226 246344 105282 246824
rect 132550 246344 132606 246824
rect 159782 246344 159838 246824
rect 187014 246344 187070 246824
rect 214246 246344 214302 246824
rect 23544 244918 23572 246344
rect 23532 244912 23584 244918
rect 23532 244854 23584 244860
rect 50776 244850 50804 246344
rect 70544 244912 70596 244918
rect 70544 244854 70596 244860
rect 50764 244844 50816 244850
rect 50764 244786 50816 244792
rect 70556 242812 70584 244854
rect 78008 242812 78036 246344
rect 105240 244918 105268 246344
rect 105228 244912 105280 244918
rect 105228 244854 105280 244860
rect 85632 242464 85684 242470
rect 85566 242412 85632 242418
rect 85566 242406 85684 242412
rect 85566 242390 85672 242406
rect 93018 242390 93400 242418
rect 93372 242130 93400 242390
rect 132564 242198 132592 246344
rect 149664 244912 149716 244918
rect 149664 244854 149716 244860
rect 142396 244844 142448 244850
rect 142396 244786 142448 244792
rect 142408 242826 142436 244786
rect 149676 242826 149704 244854
rect 159796 244850 159824 246344
rect 157484 244844 157536 244850
rect 157484 244786 157536 244792
rect 159784 244844 159836 244850
rect 159784 244786 159836 244792
rect 157496 242826 157524 244786
rect 142408 242798 142560 242826
rect 149676 242798 150012 242826
rect 157496 242798 157556 242826
rect 165008 242390 165344 242418
rect 165316 242198 165344 242390
rect 132552 242192 132604 242198
rect 132552 242134 132604 242140
rect 165304 242192 165356 242198
rect 165304 242134 165356 242140
rect 187028 242130 187056 246344
rect 214260 242198 214288 246344
rect 214248 242192 214300 242198
rect 214248 242134 214300 242140
rect 93360 242124 93412 242130
rect 93360 242066 93412 242072
rect 187016 242124 187068 242130
rect 187016 242066 187068 242072
rect 98234 238760 98290 238769
rect 98234 238695 98290 238704
rect 169994 238760 170050 238769
rect 169994 238695 170050 238704
rect 12030 235904 12086 235913
rect 12030 235839 12086 235848
rect 11938 214280 11994 214289
rect 11938 214215 11994 214224
rect 11952 105761 11980 214215
rect 12044 179745 12072 235839
rect 71372 217984 71424 217990
rect 71372 217926 71424 217932
rect 46532 217916 46584 217922
rect 46532 217858 46584 217864
rect 37240 217236 37292 217242
rect 37240 217178 37292 217184
rect 37252 215748 37280 217178
rect 46544 215748 46572 217858
rect 55822 217272 55878 217281
rect 71384 217242 71412 217926
rect 55822 217207 55878 217216
rect 71372 217236 71424 217242
rect 55836 215748 55864 217207
rect 71372 217178 71424 217184
rect 62540 215808 62592 215814
rect 62540 215750 62592 215756
rect 62552 215377 62580 215750
rect 62538 215368 62594 215377
rect 62538 215303 62594 215312
rect 62630 214688 62686 214697
rect 62630 214623 62686 214632
rect 62644 214590 62672 214623
rect 62632 214584 62684 214590
rect 62632 214526 62684 214532
rect 65024 214584 65076 214590
rect 65024 214526 65076 214532
rect 63642 214008 63698 214017
rect 63698 213966 63776 213994
rect 63642 213943 63698 213952
rect 62538 213328 62594 213337
rect 62538 213263 62540 213272
rect 62592 213263 62594 213272
rect 62540 213234 62592 213240
rect 63748 213094 63776 213966
rect 65036 213473 65064 214526
rect 71384 213586 71412 217178
rect 71844 215814 71872 218876
rect 79376 217236 79428 217242
rect 79376 217178 79428 217184
rect 71832 215808 71884 215814
rect 71832 215750 71884 215756
rect 79388 213586 79416 217178
rect 81780 216630 81808 218876
rect 81768 216624 81820 216630
rect 81768 216566 81820 216572
rect 91808 216562 91836 218876
rect 98248 217922 98276 238695
rect 98326 230736 98382 230745
rect 98326 230671 98382 230680
rect 98236 217916 98288 217922
rect 98236 217858 98288 217864
rect 94004 216624 94056 216630
rect 94004 216566 94056 216572
rect 91796 216556 91848 216562
rect 91796 216498 91848 216504
rect 86920 216488 86972 216494
rect 86920 216430 86972 216436
rect 86932 213586 86960 216430
rect 71384 213558 71628 213586
rect 79080 213558 79416 213586
rect 86624 213558 86960 213586
rect 94016 213586 94044 216566
rect 98340 216494 98368 230671
rect 168522 230192 168578 230201
rect 168522 230127 168578 230136
rect 168536 229822 168564 230127
rect 167788 229816 167840 229822
rect 167708 229764 167788 229770
rect 167708 229758 167840 229764
rect 168524 229816 168576 229822
rect 168524 229758 168576 229764
rect 167708 229742 167828 229758
rect 98418 222848 98474 222857
rect 98418 222783 98474 222792
rect 98432 217922 98460 222783
rect 167708 218890 167736 229742
rect 143788 218862 143848 218890
rect 153784 218862 154120 218890
rect 163812 218862 164148 218890
rect 143684 217984 143736 217990
rect 143684 217926 143736 217932
rect 98420 217916 98472 217922
rect 98420 217858 98472 217864
rect 109276 217916 109328 217922
rect 109276 217858 109328 217864
rect 118844 217916 118896 217922
rect 118844 217858 118896 217864
rect 109288 217310 109316 217858
rect 109276 217304 109328 217310
rect 109276 217246 109328 217252
rect 102376 216556 102428 216562
rect 102376 216498 102428 216504
rect 98328 216488 98380 216494
rect 98328 216430 98380 216436
rect 102388 215377 102416 216498
rect 109288 215762 109316 217246
rect 118856 215762 118884 217858
rect 143696 217310 143724 217926
rect 143684 217304 143736 217310
rect 143684 217246 143736 217252
rect 127768 217236 127820 217242
rect 127768 217178 127820 217184
rect 109288 215734 109532 215762
rect 118824 215734 118884 215762
rect 127780 215762 127808 217178
rect 135404 215808 135456 215814
rect 127780 215734 128116 215762
rect 135404 215750 135456 215756
rect 135416 215649 135444 215750
rect 135402 215640 135458 215649
rect 135402 215575 135458 215584
rect 102374 215368 102430 215377
rect 102374 215303 102430 215312
rect 102558 214688 102614 214697
rect 100996 214652 101048 214658
rect 102558 214623 102560 214632
rect 100996 214594 101048 214600
rect 102612 214623 102614 214632
rect 135402 214688 135458 214697
rect 135402 214623 135404 214632
rect 102560 214594 102612 214600
rect 135456 214623 135458 214632
rect 136784 214652 136836 214658
rect 135404 214594 135456 214600
rect 136784 214594 136836 214600
rect 101008 213881 101036 214594
rect 103110 214008 103166 214017
rect 103110 213943 103166 213952
rect 135402 214008 135458 214017
rect 135402 213943 135458 213952
rect 100994 213872 101050 213881
rect 100994 213807 101050 213816
rect 94016 213558 94076 213586
rect 65022 213464 65078 213473
rect 65022 213399 65078 213408
rect 103124 213366 103152 213943
rect 135416 213706 135444 213943
rect 135404 213700 135456 213706
rect 135404 213642 135456 213648
rect 100996 213360 101048 213366
rect 103112 213360 103164 213366
rect 100996 213302 101048 213308
rect 102374 213328 102430 213337
rect 65024 213292 65076 213298
rect 65024 213234 65076 213240
rect 63736 213088 63788 213094
rect 63736 213030 63788 213036
rect 62354 212648 62410 212657
rect 62354 212583 62410 212592
rect 62368 211802 62396 212583
rect 62630 211968 62686 211977
rect 62630 211903 62686 211912
rect 62356 211796 62408 211802
rect 62356 211738 62408 211744
rect 62644 211734 62672 211903
rect 65036 211841 65064 213234
rect 66404 213088 66456 213094
rect 66404 213030 66456 213036
rect 100536 213088 100588 213094
rect 100536 213030 100588 213036
rect 66416 212793 66444 213030
rect 66402 212784 66458 212793
rect 66402 212719 66458 212728
rect 100548 212113 100576 213030
rect 101008 212793 101036 213302
rect 136796 213337 136824 214594
rect 136876 213700 136928 213706
rect 136876 213642 136928 213648
rect 103112 213302 103164 213308
rect 135034 213328 135090 213337
rect 102374 213263 102430 213272
rect 135034 213263 135036 213272
rect 102388 213162 102416 213263
rect 135088 213263 135090 213272
rect 136782 213328 136838 213337
rect 136782 213263 136838 213272
rect 135036 213234 135088 213240
rect 102376 213156 102428 213162
rect 102376 213098 102428 213104
rect 136888 212793 136916 213642
rect 143696 213586 143724 217246
rect 143788 215814 143816 218862
rect 154092 216494 154120 218862
rect 158588 216624 158640 216630
rect 158588 216566 158640 216572
rect 154080 216488 154132 216494
rect 154080 216430 154132 216436
rect 151042 215912 151098 215921
rect 151042 215847 151098 215856
rect 143776 215808 143828 215814
rect 143776 215750 143828 215756
rect 143618 213558 143724 213586
rect 151056 213572 151084 215847
rect 158600 213572 158628 216566
rect 164120 216562 164148 218862
rect 167432 218862 167736 218890
rect 167432 218618 167460 218862
rect 167248 218590 167460 218618
rect 167248 216630 167276 218590
rect 170008 217922 170036 238695
rect 223078 234952 223134 234961
rect 223078 234887 223134 234896
rect 223092 223430 223120 234887
rect 207256 223424 207308 223430
rect 207256 223366 207308 223372
rect 223080 223424 223132 223430
rect 223080 223366 223132 223372
rect 170086 222848 170142 222857
rect 207268 222818 207296 223366
rect 170086 222783 170088 222792
rect 170140 222783 170142 222792
rect 207256 222812 207308 222818
rect 170088 222754 170140 222760
rect 207256 222754 207308 222760
rect 170100 217990 170128 222754
rect 170088 217984 170140 217990
rect 170088 217926 170140 217932
rect 169996 217916 170048 217922
rect 169996 217858 170048 217864
rect 167236 216624 167288 216630
rect 167236 216566 167288 216572
rect 164108 216556 164160 216562
rect 164108 216498 164160 216504
rect 174228 216556 174280 216562
rect 174228 216498 174280 216504
rect 166040 216488 166092 216494
rect 166040 216430 166092 216436
rect 166052 213572 166080 216430
rect 174240 215785 174268 216498
rect 174226 215776 174282 215785
rect 174226 215711 174282 215720
rect 174042 214688 174098 214697
rect 174042 214623 174098 214632
rect 174056 214046 174084 214623
rect 172020 214040 172072 214046
rect 172020 213982 172072 213988
rect 174044 214040 174096 214046
rect 174044 213982 174096 213988
rect 174226 214008 174282 214017
rect 172032 213881 172060 213982
rect 174226 213943 174282 213952
rect 172018 213872 172074 213881
rect 172018 213807 172074 213816
rect 174042 213328 174098 213337
rect 137060 213292 137112 213298
rect 174042 213263 174098 213272
rect 137060 213234 137112 213240
rect 100994 212784 101050 212793
rect 100994 212719 101050 212728
rect 136874 212784 136930 212793
rect 136874 212719 136930 212728
rect 102466 212648 102522 212657
rect 102466 212583 102522 212592
rect 135402 212648 135458 212657
rect 135402 212583 135458 212592
rect 100534 212104 100590 212113
rect 100534 212039 100590 212048
rect 102374 211968 102430 211977
rect 100996 211932 101048 211938
rect 102374 211903 102376 211912
rect 100996 211874 101048 211880
rect 102428 211903 102430 211912
rect 102376 211874 102428 211880
rect 65022 211832 65078 211841
rect 64932 211796 64984 211802
rect 65022 211767 65078 211776
rect 64932 211738 64984 211744
rect 62632 211728 62684 211734
rect 62632 211670 62684 211676
rect 62538 211288 62594 211297
rect 62538 211223 62594 211232
rect 62552 210850 62580 211223
rect 62540 210844 62592 210850
rect 62540 210786 62592 210792
rect 62630 210608 62686 210617
rect 62630 210543 62686 210552
rect 62644 210442 62672 210543
rect 64944 210481 64972 211738
rect 65024 211728 65076 211734
rect 65024 211670 65076 211676
rect 65036 210617 65064 211670
rect 100812 211660 100864 211666
rect 100812 211602 100864 211608
rect 100824 211569 100852 211602
rect 65666 211560 65722 211569
rect 65666 211495 65722 211504
rect 100810 211560 100866 211569
rect 100810 211495 100866 211504
rect 65484 210844 65536 210850
rect 65484 210786 65536 210792
rect 65022 210608 65078 210617
rect 65022 210543 65078 210552
rect 64930 210472 64986 210481
rect 62632 210436 62684 210442
rect 64930 210407 64986 210416
rect 65024 210436 65076 210442
rect 62632 210378 62684 210384
rect 65024 210378 65076 210384
rect 62630 209928 62686 209937
rect 62630 209863 62632 209872
rect 62684 209863 62686 209872
rect 62632 209834 62684 209840
rect 65036 209393 65064 210378
rect 65496 210345 65524 210786
rect 65680 210481 65708 211495
rect 101008 211025 101036 211874
rect 102480 211734 102508 212583
rect 135416 212210 135444 212583
rect 135404 212204 135456 212210
rect 135404 212146 135456 212152
rect 136968 212204 137020 212210
rect 136968 212146 137020 212152
rect 135402 211968 135458 211977
rect 135402 211903 135404 211912
rect 135456 211903 135458 211912
rect 136876 211932 136928 211938
rect 135404 211874 135456 211880
rect 136876 211874 136928 211880
rect 102468 211728 102520 211734
rect 102468 211670 102520 211676
rect 136888 211025 136916 211874
rect 136980 211569 137008 212146
rect 137072 212113 137100 213234
rect 172664 213088 172716 213094
rect 172662 213056 172664 213065
rect 172716 213056 172718 213065
rect 172662 212991 172718 213000
rect 174056 212686 174084 213263
rect 174240 213162 174268 213943
rect 174228 213156 174280 213162
rect 174228 213098 174280 213104
rect 172664 212680 172716 212686
rect 172664 212622 172716 212628
rect 174044 212680 174096 212686
rect 174044 212622 174096 212628
rect 174226 212648 174282 212657
rect 172676 212521 172704 212622
rect 174226 212583 174282 212592
rect 172662 212512 172718 212521
rect 172662 212447 172718 212456
rect 137058 212104 137114 212113
rect 137058 212039 137114 212048
rect 174042 211968 174098 211977
rect 174042 211903 174098 211912
rect 172756 211728 172808 211734
rect 172662 211696 172718 211705
rect 172718 211676 172756 211682
rect 172718 211670 172808 211676
rect 172718 211654 172796 211670
rect 172662 211631 172718 211640
rect 136966 211560 137022 211569
rect 136966 211495 137022 211504
rect 174056 211326 174084 211903
rect 174240 211734 174268 212583
rect 174228 211728 174280 211734
rect 174228 211670 174280 211676
rect 172388 211320 172440 211326
rect 172386 211288 172388 211297
rect 174044 211320 174096 211326
rect 172440 211288 172442 211297
rect 174044 211262 174096 211268
rect 174226 211288 174282 211297
rect 172386 211223 172442 211232
rect 174226 211223 174282 211232
rect 100994 211016 101050 211025
rect 100994 210951 101050 210960
rect 136874 211016 136930 211025
rect 136874 210951 136930 210960
rect 103662 210880 103718 210889
rect 100904 210844 100956 210850
rect 103662 210815 103664 210824
rect 100904 210786 100956 210792
rect 103716 210815 103718 210824
rect 103664 210786 103716 210792
rect 65666 210472 65722 210481
rect 65666 210407 65722 210416
rect 100916 210345 100944 210786
rect 174240 210646 174268 211223
rect 172664 210640 172716 210646
rect 102374 210608 102430 210617
rect 100996 210572 101048 210578
rect 102374 210543 102376 210552
rect 100996 210514 101048 210520
rect 102428 210543 102430 210552
rect 134666 210608 134722 210617
rect 172662 210608 172664 210617
rect 174228 210640 174280 210646
rect 172716 210608 172718 210617
rect 134666 210543 134668 210552
rect 102376 210514 102428 210520
rect 134720 210543 134722 210552
rect 136876 210572 136928 210578
rect 134668 210514 134720 210520
rect 172662 210543 172718 210552
rect 174042 210608 174098 210617
rect 174228 210582 174280 210588
rect 174042 210543 174098 210552
rect 136876 210514 136928 210520
rect 65482 210336 65538 210345
rect 65482 210271 65538 210280
rect 100902 210336 100958 210345
rect 100902 210271 100958 210280
rect 66404 209892 66456 209898
rect 66404 209834 66456 209840
rect 65022 209384 65078 209393
rect 65022 209319 65078 209328
rect 62722 209248 62778 209257
rect 62722 209183 62778 209192
rect 62736 209082 62764 209183
rect 66416 209121 66444 209834
rect 101008 209801 101036 210514
rect 136888 209801 136916 210514
rect 174056 210102 174084 210543
rect 172664 210096 172716 210102
rect 172662 210064 172664 210073
rect 174044 210096 174096 210102
rect 172716 210064 172718 210073
rect 174044 210038 174096 210044
rect 172662 209999 172718 210008
rect 174134 209928 174190 209937
rect 174134 209863 174190 209872
rect 100994 209792 101050 209801
rect 100994 209727 101050 209736
rect 136874 209792 136930 209801
rect 136874 209727 136930 209736
rect 174148 209422 174176 209863
rect 171652 209416 171704 209422
rect 171650 209384 171652 209393
rect 174136 209416 174188 209422
rect 171704 209384 171706 209393
rect 174136 209358 174188 209364
rect 171650 209319 171706 209328
rect 135310 209248 135366 209257
rect 135310 209183 135366 209192
rect 174594 209248 174650 209257
rect 174594 209183 174650 209192
rect 66402 209112 66458 209121
rect 62724 209076 62776 209082
rect 62724 209018 62776 209024
rect 65024 209076 65076 209082
rect 135324 209082 135352 209183
rect 66402 209047 66458 209056
rect 135312 209076 135364 209082
rect 65024 209018 65076 209024
rect 135312 209018 135364 209024
rect 137704 209076 137756 209082
rect 137704 209018 137756 209024
rect 62630 208568 62686 208577
rect 62630 208503 62686 208512
rect 62644 208402 62672 208503
rect 62632 208396 62684 208402
rect 62632 208338 62684 208344
rect 63642 207888 63698 207897
rect 63698 207846 63776 207874
rect 63642 207823 63698 207832
rect 63748 207518 63776 207846
rect 65036 207625 65064 209018
rect 137716 208577 137744 209018
rect 174608 209014 174636 209183
rect 174596 209008 174648 209014
rect 174596 208950 174648 208956
rect 172112 208940 172164 208946
rect 172112 208882 172164 208888
rect 172124 208849 172152 208882
rect 172110 208840 172166 208849
rect 172110 208775 172166 208784
rect 65850 208568 65906 208577
rect 65850 208503 65906 208512
rect 137702 208568 137758 208577
rect 137702 208503 137758 208512
rect 65864 207625 65892 208503
rect 66404 208396 66456 208402
rect 66404 208338 66456 208344
rect 66416 208033 66444 208338
rect 66402 208024 66458 208033
rect 66402 207959 66458 207968
rect 135402 207888 135458 207897
rect 135402 207823 135404 207832
rect 135456 207823 135458 207832
rect 136876 207852 136928 207858
rect 135404 207794 135456 207800
rect 136876 207794 136928 207800
rect 65022 207616 65078 207625
rect 65022 207551 65078 207560
rect 65850 207616 65906 207625
rect 65850 207551 65906 207560
rect 63736 207512 63788 207518
rect 63736 207454 63788 207460
rect 65300 207512 65352 207518
rect 65300 207454 65352 207460
rect 65312 207353 65340 207454
rect 136888 207353 136916 207794
rect 65298 207344 65354 207353
rect 65298 207279 65354 207288
rect 136874 207344 136930 207353
rect 136874 207279 136930 207288
rect 62538 207208 62594 207217
rect 62538 207143 62594 207152
rect 174134 207208 174190 207217
rect 174134 207143 174190 207152
rect 62552 206770 62580 207143
rect 174148 206838 174176 207143
rect 171652 206832 171704 206838
rect 65666 206800 65722 206809
rect 62540 206764 62592 206770
rect 171652 206774 171704 206780
rect 174136 206832 174188 206838
rect 174136 206774 174188 206780
rect 65666 206735 65668 206744
rect 62540 206706 62592 206712
rect 65720 206735 65722 206744
rect 65668 206706 65720 206712
rect 171664 206673 171692 206774
rect 171650 206664 171706 206673
rect 171650 206599 171706 206608
rect 62630 206528 62686 206537
rect 62630 206463 62686 206472
rect 135402 206528 135458 206537
rect 135402 206463 135458 206472
rect 174042 206528 174098 206537
rect 174042 206463 174098 206472
rect 62644 206226 62672 206463
rect 135416 206362 135444 206463
rect 135404 206356 135456 206362
rect 135404 206298 135456 206304
rect 136876 206356 136928 206362
rect 136876 206298 136928 206304
rect 62632 206220 62684 206226
rect 62632 206162 62684 206168
rect 64932 206220 64984 206226
rect 64932 206162 64984 206168
rect 62630 205848 62686 205857
rect 62630 205783 62686 205792
rect 62644 205478 62672 205783
rect 62632 205472 62684 205478
rect 62632 205414 62684 205420
rect 64944 205313 64972 206162
rect 136888 206129 136916 206298
rect 136874 206120 136930 206129
rect 136874 206055 136930 206064
rect 174056 206022 174084 206463
rect 171836 206016 171888 206022
rect 171834 205984 171836 205993
rect 174044 206016 174096 206022
rect 171888 205984 171890 205993
rect 174044 205958 174096 205964
rect 171834 205919 171890 205928
rect 66402 205576 66458 205585
rect 66402 205511 66458 205520
rect 66416 205478 66444 205511
rect 66404 205472 66456 205478
rect 66404 205414 66456 205420
rect 64930 205304 64986 205313
rect 64930 205239 64986 205248
rect 62630 204488 62686 204497
rect 62630 204423 62686 204432
rect 62644 204390 62672 204423
rect 62632 204384 62684 204390
rect 65668 204384 65720 204390
rect 62632 204326 62684 204332
rect 65666 204352 65668 204361
rect 65720 204352 65722 204361
rect 65666 204287 65722 204296
rect 62540 204248 62592 204254
rect 62540 204190 62592 204196
rect 65484 204248 65536 204254
rect 65484 204190 65536 204196
rect 62552 203817 62580 204190
rect 65496 203817 65524 204190
rect 62538 203808 62594 203817
rect 62538 203743 62594 203752
rect 65482 203808 65538 203817
rect 65482 203743 65538 203752
rect 100904 200712 100956 200718
rect 100902 200680 100904 200689
rect 102376 200712 102428 200718
rect 100956 200680 100958 200689
rect 102376 200654 102428 200660
rect 136782 200680 136838 200689
rect 100902 200615 100958 200624
rect 102388 200417 102416 200654
rect 136782 200615 136838 200624
rect 136796 200514 136824 200615
rect 135404 200508 135456 200514
rect 135404 200450 135456 200456
rect 136784 200508 136836 200514
rect 136784 200450 136836 200456
rect 135416 200417 135444 200450
rect 65022 200408 65078 200417
rect 65022 200343 65078 200352
rect 66402 200408 66458 200417
rect 66402 200343 66458 200352
rect 102374 200408 102430 200417
rect 102374 200343 102430 200352
rect 135402 200408 135458 200417
rect 135402 200343 135458 200352
rect 65036 199154 65064 200343
rect 65114 200136 65170 200145
rect 65114 200071 65170 200080
rect 65128 199329 65156 200071
rect 66416 199601 66444 200343
rect 66402 199592 66458 199601
rect 66402 199527 66458 199536
rect 136782 199456 136838 199465
rect 136782 199391 136838 199400
rect 172202 199456 172258 199465
rect 172202 199391 172204 199400
rect 100904 199352 100956 199358
rect 65114 199320 65170 199329
rect 65114 199255 65170 199264
rect 100902 199320 100904 199329
rect 102376 199352 102428 199358
rect 100956 199320 100958 199329
rect 102376 199294 102428 199300
rect 100902 199255 100958 199264
rect 62356 199148 62408 199154
rect 62356 199090 62408 199096
rect 65024 199148 65076 199154
rect 65024 199090 65076 199096
rect 62368 199057 62396 199090
rect 102388 199057 102416 199294
rect 136796 199154 136824 199391
rect 172256 199391 172258 199400
rect 175240 199420 175292 199426
rect 172204 199362 172256 199368
rect 175240 199362 175292 199368
rect 134760 199148 134812 199154
rect 134760 199090 134812 199096
rect 136784 199148 136836 199154
rect 136784 199090 136836 199096
rect 134772 199057 134800 199090
rect 175252 199057 175280 199362
rect 62354 199048 62410 199057
rect 62354 198983 62410 198992
rect 102374 199048 102430 199057
rect 102374 198983 102430 198992
rect 134758 199048 134814 199057
rect 134758 198983 134814 198992
rect 175238 199048 175294 199057
rect 175238 198983 175294 198992
rect 172202 198096 172258 198105
rect 172202 198031 172204 198040
rect 172256 198031 172258 198040
rect 174228 198060 174280 198066
rect 172204 198002 172256 198008
rect 174228 198002 174280 198008
rect 65022 197960 65078 197969
rect 65022 197895 65078 197904
rect 100902 197960 100958 197969
rect 136782 197960 136838 197969
rect 100902 197895 100904 197904
rect 65036 197794 65064 197895
rect 100956 197895 100958 197904
rect 102376 197924 102428 197930
rect 100904 197866 100956 197872
rect 136782 197895 136838 197904
rect 102376 197866 102428 197872
rect 62632 197788 62684 197794
rect 62632 197730 62684 197736
rect 65024 197788 65076 197794
rect 65024 197730 65076 197736
rect 62644 197697 62672 197730
rect 102388 197697 102416 197866
rect 136796 197794 136824 197895
rect 135404 197788 135456 197794
rect 135404 197730 135456 197736
rect 136784 197788 136836 197794
rect 136784 197730 136836 197736
rect 135416 197697 135444 197730
rect 174240 197697 174268 198002
rect 62630 197688 62686 197697
rect 62630 197623 62686 197632
rect 102374 197688 102430 197697
rect 102374 197623 102430 197632
rect 135402 197688 135458 197697
rect 135402 197623 135458 197632
rect 174226 197688 174282 197697
rect 174226 197623 174282 197632
rect 65022 196872 65078 196881
rect 65022 196807 65078 196816
rect 172662 196872 172718 196881
rect 172662 196807 172664 196816
rect 63736 196564 63788 196570
rect 63736 196506 63788 196512
rect 62632 196496 62684 196502
rect 62632 196438 62684 196444
rect 62644 196337 62672 196438
rect 62630 196328 62686 196337
rect 62630 196263 62686 196272
rect 63642 195648 63698 195657
rect 63748 195634 63776 196506
rect 65036 196502 65064 196807
rect 172716 196807 172718 196816
rect 174136 196836 174188 196842
rect 172664 196778 172716 196784
rect 174136 196778 174188 196784
rect 100902 196736 100958 196745
rect 136782 196736 136838 196745
rect 100902 196671 100904 196680
rect 100956 196671 100958 196680
rect 102376 196700 102428 196706
rect 100904 196642 100956 196648
rect 136782 196671 136838 196680
rect 172202 196736 172258 196745
rect 172202 196671 172204 196680
rect 102376 196642 102428 196648
rect 66402 196600 66458 196609
rect 66402 196535 66404 196544
rect 66456 196535 66458 196544
rect 100902 196600 100958 196609
rect 100902 196535 100904 196544
rect 66404 196506 66456 196512
rect 100956 196535 100958 196544
rect 100904 196506 100956 196512
rect 65024 196496 65076 196502
rect 65024 196438 65076 196444
rect 102388 196337 102416 196642
rect 136690 196600 136746 196609
rect 102468 196564 102520 196570
rect 136690 196535 136746 196544
rect 102468 196506 102520 196512
rect 102374 196328 102430 196337
rect 102374 196263 102430 196272
rect 102480 195657 102508 196506
rect 135404 196428 135456 196434
rect 135404 196370 135456 196376
rect 135416 196337 135444 196370
rect 135402 196328 135458 196337
rect 135402 196263 135458 196272
rect 136704 196094 136732 196535
rect 136796 196434 136824 196671
rect 172256 196671 172258 196680
rect 172204 196642 172256 196648
rect 136784 196428 136836 196434
rect 136784 196370 136836 196376
rect 174148 196337 174176 196778
rect 174228 196700 174280 196706
rect 174228 196642 174280 196648
rect 174134 196328 174190 196337
rect 174134 196263 174190 196272
rect 174240 196201 174268 196642
rect 174226 196192 174282 196201
rect 174226 196127 174282 196136
rect 134300 196088 134352 196094
rect 134298 196056 134300 196065
rect 136692 196088 136744 196094
rect 134352 196056 134354 196065
rect 136692 196030 136744 196036
rect 134298 195991 134354 196000
rect 63698 195606 63776 195634
rect 65022 195648 65078 195657
rect 63642 195583 63698 195592
rect 65022 195583 65078 195592
rect 102466 195648 102522 195657
rect 102466 195583 102522 195592
rect 171466 195648 171522 195657
rect 171466 195583 171468 195592
rect 62540 195136 62592 195142
rect 62540 195078 62592 195084
rect 62552 194297 62580 195078
rect 65036 195006 65064 195583
rect 171520 195583 171522 195592
rect 174136 195612 174188 195618
rect 171468 195554 171520 195560
rect 174136 195554 174188 195560
rect 100718 195512 100774 195521
rect 100718 195447 100774 195456
rect 136874 195512 136930 195521
rect 136874 195447 136930 195456
rect 66402 195376 66458 195385
rect 100732 195346 100760 195447
rect 66402 195311 66458 195320
rect 100720 195340 100772 195346
rect 66416 195210 66444 195311
rect 100720 195282 100772 195288
rect 102468 195340 102520 195346
rect 102468 195282 102520 195288
rect 100902 195240 100958 195249
rect 66404 195204 66456 195210
rect 100902 195175 100904 195184
rect 66404 195146 66456 195152
rect 100956 195175 100958 195184
rect 102376 195204 102428 195210
rect 100904 195146 100956 195152
rect 102376 195146 102428 195152
rect 62632 195000 62684 195006
rect 62630 194968 62632 194977
rect 65024 195000 65076 195006
rect 62684 194968 62686 194977
rect 65024 194942 65076 194948
rect 62630 194903 62686 194912
rect 65114 194832 65170 194841
rect 65114 194767 65170 194776
rect 65022 194424 65078 194433
rect 65022 194359 65078 194368
rect 62538 194288 62594 194297
rect 62538 194223 62594 194232
rect 65036 193306 65064 194359
rect 65128 193889 65156 194767
rect 102388 194297 102416 195146
rect 102480 194977 102508 195282
rect 136782 195240 136838 195249
rect 136888 195210 136916 195447
rect 172662 195240 172718 195249
rect 136782 195175 136838 195184
rect 136876 195204 136928 195210
rect 135404 195136 135456 195142
rect 135404 195078 135456 195084
rect 135416 194977 135444 195078
rect 102466 194968 102522 194977
rect 102466 194903 102522 194912
rect 135402 194968 135458 194977
rect 135402 194903 135458 194912
rect 136796 194870 136824 195175
rect 172662 195175 172664 195184
rect 136876 195146 136928 195152
rect 172716 195175 172718 195184
rect 172664 195146 172716 195152
rect 174148 194977 174176 195554
rect 174228 195204 174280 195210
rect 174228 195146 174280 195152
rect 174134 194968 174190 194977
rect 174134 194903 174190 194912
rect 135404 194864 135456 194870
rect 135402 194832 135404 194841
rect 136784 194864 136836 194870
rect 135456 194832 135458 194841
rect 174240 194841 174268 195146
rect 136784 194806 136836 194812
rect 174226 194832 174282 194841
rect 135402 194767 135458 194776
rect 174226 194767 174282 194776
rect 100626 194288 100682 194297
rect 100626 194223 100628 194232
rect 100680 194223 100682 194232
rect 102374 194288 102430 194297
rect 136782 194288 136838 194297
rect 102374 194223 102430 194232
rect 102468 194252 102520 194258
rect 100628 194194 100680 194200
rect 136782 194223 136838 194232
rect 171558 194288 171614 194297
rect 171558 194223 171560 194232
rect 102468 194194 102520 194200
rect 65114 193880 65170 193889
rect 65114 193815 65170 193824
rect 100626 193880 100682 193889
rect 100626 193815 100628 193824
rect 100680 193815 100682 193824
rect 102376 193844 102428 193850
rect 100628 193786 100680 193792
rect 102376 193786 102428 193792
rect 66402 193608 66458 193617
rect 66402 193543 66458 193552
rect 62356 193300 62408 193306
rect 62356 193242 62408 193248
rect 65024 193300 65076 193306
rect 65024 193242 65076 193248
rect 62368 192937 62396 193242
rect 62354 192928 62410 192937
rect 62354 192863 62410 192872
rect 12214 192656 12270 192665
rect 12214 192591 12270 192600
rect 65022 192656 65078 192665
rect 65022 192591 65078 192600
rect 12030 179736 12086 179745
rect 12030 179671 12086 179680
rect 12122 171032 12178 171041
rect 12122 170967 12178 170976
rect 12030 149816 12086 149825
rect 12030 149751 12086 149760
rect 11938 105752 11994 105761
rect 11938 105687 11994 105696
rect 11938 75152 11994 75161
rect 11938 75087 11994 75096
rect 11952 41297 11980 75087
rect 12044 62921 12072 149751
rect 12136 95833 12164 170967
rect 12228 170089 12256 192591
rect 64930 192520 64986 192529
rect 64930 192455 64986 192464
rect 64944 192286 64972 192455
rect 62540 192280 62592 192286
rect 62538 192248 62540 192257
rect 64932 192280 64984 192286
rect 62592 192248 62594 192257
rect 64932 192222 64984 192228
rect 62538 192183 62594 192192
rect 65036 191606 65064 192591
rect 66416 192529 66444 193543
rect 99706 193200 99762 193209
rect 99706 193135 99762 193144
rect 99720 192898 99748 193135
rect 102388 192937 102416 193786
rect 102480 193617 102508 194194
rect 136690 193880 136746 193889
rect 136690 193815 136746 193824
rect 135404 193708 135456 193714
rect 135404 193650 135456 193656
rect 135416 193617 135444 193650
rect 102466 193608 102522 193617
rect 102466 193543 102522 193552
rect 135402 193608 135458 193617
rect 135402 193543 135458 193552
rect 136704 193510 136732 193815
rect 136796 193714 136824 194223
rect 171612 194223 171614 194232
rect 174136 194252 174188 194258
rect 171560 194194 171612 194200
rect 174136 194194 174188 194200
rect 172662 194016 172718 194025
rect 172662 193951 172718 193960
rect 172676 193850 172704 193951
rect 172664 193844 172716 193850
rect 172664 193786 172716 193792
rect 136784 193708 136836 193714
rect 136784 193650 136836 193656
rect 174148 193617 174176 194194
rect 174228 193844 174280 193850
rect 174228 193786 174280 193792
rect 174134 193608 174190 193617
rect 174134 193543 174190 193552
rect 135404 193504 135456 193510
rect 135402 193472 135404 193481
rect 136692 193504 136744 193510
rect 135456 193472 135458 193481
rect 174240 193481 174268 193786
rect 136692 193446 136744 193452
rect 174226 193472 174282 193481
rect 135402 193407 135458 193416
rect 174226 193407 174282 193416
rect 136782 193200 136838 193209
rect 136782 193135 136838 193144
rect 171650 193200 171706 193209
rect 171650 193135 171706 193144
rect 102374 192928 102430 192937
rect 99708 192892 99760 192898
rect 102374 192863 102430 192872
rect 102468 192892 102520 192898
rect 99708 192834 99760 192840
rect 102468 192834 102520 192840
rect 66402 192520 66458 192529
rect 66402 192455 66458 192464
rect 100626 192520 100682 192529
rect 100626 192455 100628 192464
rect 100680 192455 100682 192464
rect 102376 192484 102428 192490
rect 100628 192426 100680 192432
rect 102376 192426 102428 192432
rect 66402 192384 66458 192393
rect 66402 192319 66458 192328
rect 66310 191840 66366 191849
rect 66310 191775 66366 191784
rect 62356 191600 62408 191606
rect 62354 191568 62356 191577
rect 65024 191600 65076 191606
rect 62408 191568 62410 191577
rect 65024 191542 65076 191548
rect 62354 191503 62410 191512
rect 65022 191296 65078 191305
rect 65022 191231 65078 191240
rect 62448 190988 62500 190994
rect 62448 190930 62500 190936
rect 62460 190217 62488 190930
rect 65036 190926 65064 191231
rect 65206 191160 65262 191169
rect 65206 191095 65262 191104
rect 62632 190920 62684 190926
rect 62630 190888 62632 190897
rect 65024 190920 65076 190926
rect 62684 190888 62686 190897
rect 65024 190862 65076 190868
rect 62630 190823 62686 190832
rect 62446 190208 62502 190217
rect 62446 190143 62502 190152
rect 63644 189696 63696 189702
rect 63644 189638 63696 189644
rect 65022 189664 65078 189673
rect 62632 189560 62684 189566
rect 62630 189528 62632 189537
rect 62684 189528 62686 189537
rect 62630 189463 62686 189472
rect 62632 189084 62684 189090
rect 62632 189026 62684 189032
rect 62644 188857 62672 189026
rect 62630 188848 62686 188857
rect 62630 188783 62686 188792
rect 63656 188177 63684 189638
rect 65022 189599 65078 189608
rect 65036 189090 65064 189599
rect 65220 189566 65248 191095
rect 66324 191062 66352 191775
rect 66416 191305 66444 192319
rect 99890 191976 99946 191985
rect 99890 191911 99892 191920
rect 99944 191911 99946 191920
rect 102284 191940 102336 191946
rect 99892 191882 99944 191888
rect 102284 191882 102336 191888
rect 66402 191296 66458 191305
rect 66402 191231 66458 191240
rect 100626 191296 100682 191305
rect 100626 191231 100628 191240
rect 100680 191231 100682 191240
rect 102192 191260 102244 191266
rect 100628 191202 100680 191208
rect 102192 191202 102244 191208
rect 100902 191160 100958 191169
rect 100902 191095 100958 191104
rect 100916 191062 100944 191095
rect 66312 191056 66364 191062
rect 66312 190998 66364 191004
rect 100904 191056 100956 191062
rect 100904 190998 100956 191004
rect 66310 190616 66366 190625
rect 66310 190551 66366 190560
rect 66324 189673 66352 190551
rect 102204 190217 102232 191202
rect 102296 190897 102324 191882
rect 102388 191577 102416 192426
rect 102480 192257 102508 192834
rect 136690 192520 136746 192529
rect 136690 192455 136746 192464
rect 135404 192348 135456 192354
rect 135404 192290 135456 192296
rect 134300 192280 134352 192286
rect 102466 192248 102522 192257
rect 135416 192257 135444 192290
rect 136704 192286 136732 192455
rect 136796 192354 136824 193135
rect 171664 193034 171692 193135
rect 171652 193028 171704 193034
rect 171652 192970 171704 192976
rect 174228 193028 174280 193034
rect 174228 192970 174280 192976
rect 172202 192792 172258 192801
rect 172202 192727 172258 192736
rect 172216 192626 172244 192727
rect 172204 192620 172256 192626
rect 172204 192562 172256 192568
rect 174136 192620 174188 192626
rect 174136 192562 174188 192568
rect 136784 192348 136836 192354
rect 136784 192290 136836 192296
rect 136692 192280 136744 192286
rect 134300 192222 134352 192228
rect 135402 192248 135458 192257
rect 102466 192183 102522 192192
rect 134312 192121 134340 192222
rect 136692 192222 136744 192228
rect 135402 192183 135458 192192
rect 174148 192121 174176 192562
rect 174240 192257 174268 192970
rect 207268 192529 207296 222754
rect 223538 211152 223594 211161
rect 223538 211087 223594 211096
rect 223552 210374 223580 211087
rect 207900 210368 207952 210374
rect 207900 210310 207952 210316
rect 223540 210368 223592 210374
rect 223540 210310 223592 210316
rect 207912 201777 207940 210310
rect 207898 201768 207954 201777
rect 207898 201703 207954 201712
rect 207254 192520 207310 192529
rect 207254 192455 207310 192464
rect 207254 192384 207310 192393
rect 207254 192319 207310 192328
rect 174226 192248 174282 192257
rect 174226 192183 174282 192192
rect 134298 192112 134354 192121
rect 134298 192047 134354 192056
rect 174134 192112 174190 192121
rect 174134 192047 174190 192056
rect 136782 191976 136838 191985
rect 136782 191911 136838 191920
rect 172202 191976 172258 191985
rect 172202 191911 172258 191920
rect 102374 191568 102430 191577
rect 102374 191503 102430 191512
rect 136690 191296 136746 191305
rect 136690 191231 136746 191240
rect 102560 191056 102612 191062
rect 102560 190998 102612 191004
rect 134300 191056 134352 191062
rect 134300 190998 134352 191004
rect 102282 190888 102338 190897
rect 102282 190823 102338 190832
rect 100534 190208 100590 190217
rect 100534 190143 100590 190152
rect 102190 190208 102246 190217
rect 102190 190143 102246 190152
rect 100548 190110 100576 190143
rect 100536 190104 100588 190110
rect 66402 190072 66458 190081
rect 100536 190046 100588 190052
rect 102468 190104 102520 190110
rect 102468 190046 102520 190052
rect 66402 190007 66458 190016
rect 66416 189702 66444 190007
rect 99890 189936 99946 189945
rect 99890 189871 99946 189880
rect 99904 189838 99932 189871
rect 99892 189832 99944 189838
rect 99892 189774 99944 189780
rect 102376 189832 102428 189838
rect 102376 189774 102428 189780
rect 66404 189696 66456 189702
rect 66310 189664 66366 189673
rect 66404 189638 66456 189644
rect 66310 189599 66366 189608
rect 65208 189560 65260 189566
rect 65208 189502 65260 189508
rect 65024 189084 65076 189090
rect 65024 189026 65076 189032
rect 102388 188177 102416 189774
rect 102480 188857 102508 190046
rect 102572 189537 102600 190998
rect 134312 189537 134340 190998
rect 135404 190988 135456 190994
rect 135404 190930 135456 190936
rect 134760 190920 134812 190926
rect 135416 190897 135444 190930
rect 136704 190926 136732 191231
rect 136796 190994 136824 191911
rect 172216 191402 172244 191911
rect 172662 191432 172718 191441
rect 172204 191396 172256 191402
rect 172662 191367 172718 191376
rect 174044 191396 174096 191402
rect 172204 191338 172256 191344
rect 172676 191334 172704 191367
rect 174044 191338 174096 191344
rect 172664 191328 172716 191334
rect 172664 191270 172716 191276
rect 173952 191328 174004 191334
rect 173952 191270 174004 191276
rect 136966 191160 137022 191169
rect 136966 191095 137022 191104
rect 136980 191062 137008 191095
rect 136968 191056 137020 191062
rect 172664 191056 172716 191062
rect 136968 190998 137020 191004
rect 172662 191024 172664 191033
rect 172716 191024 172718 191033
rect 136784 190988 136836 190994
rect 172662 190959 172718 190968
rect 136784 190930 136836 190936
rect 136692 190920 136744 190926
rect 134760 190862 134812 190868
rect 135402 190888 135458 190897
rect 134772 190761 134800 190862
rect 136692 190862 136744 190868
rect 135402 190823 135458 190832
rect 173964 190761 173992 191270
rect 174056 190897 174084 191338
rect 174964 191056 175016 191062
rect 174964 190998 175016 191004
rect 174042 190888 174098 190897
rect 174042 190823 174098 190832
rect 134758 190752 134814 190761
rect 134758 190687 134814 190696
rect 173950 190752 174006 190761
rect 173950 190687 174006 190696
rect 136782 190208 136838 190217
rect 136782 190143 136838 190152
rect 172386 190208 172442 190217
rect 172386 190143 172388 190152
rect 102558 189528 102614 189537
rect 102558 189463 102614 189472
rect 134298 189528 134354 189537
rect 134298 189463 134354 189472
rect 136796 189294 136824 190143
rect 172440 190143 172442 190152
rect 174412 190172 174464 190178
rect 172388 190114 172440 190120
rect 174412 190114 174464 190120
rect 172018 189936 172074 189945
rect 172018 189871 172074 189880
rect 137426 189800 137482 189809
rect 172032 189770 172060 189871
rect 137426 189735 137482 189744
rect 172020 189764 172072 189770
rect 134760 189288 134812 189294
rect 134758 189256 134760 189265
rect 136784 189288 136836 189294
rect 134812 189256 134814 189265
rect 136784 189230 136836 189236
rect 134758 189191 134814 189200
rect 102466 188848 102522 188857
rect 102466 188783 102522 188792
rect 137440 188206 137468 189735
rect 172020 189706 172072 189712
rect 174424 189265 174452 190114
rect 174976 189537 175004 190998
rect 175424 189764 175476 189770
rect 175424 189706 175476 189712
rect 174962 189528 175018 189537
rect 174962 189463 175018 189472
rect 174410 189256 174466 189265
rect 174410 189191 174466 189200
rect 135036 188200 135088 188206
rect 63642 188168 63698 188177
rect 63642 188103 63698 188112
rect 102374 188168 102430 188177
rect 102374 188103 102430 188112
rect 135034 188168 135036 188177
rect 137428 188200 137480 188206
rect 135088 188168 135090 188177
rect 175436 188177 175464 189706
rect 137428 188142 137480 188148
rect 175422 188168 175478 188177
rect 135034 188103 135090 188112
rect 175422 188103 175478 188112
rect 177276 187990 177750 188018
rect 32008 187854 32942 187882
rect 32008 178249 32036 187854
rect 33572 184126 33600 187868
rect 34216 184262 34244 187868
rect 34952 184330 34980 187868
rect 35596 185486 35624 187868
rect 35584 185480 35636 185486
rect 35584 185422 35636 185428
rect 36332 185350 36360 187868
rect 36320 185344 36372 185350
rect 36320 185286 36372 185292
rect 36976 184942 37004 187868
rect 37620 185214 37648 187868
rect 37884 185480 37936 185486
rect 37884 185422 37936 185428
rect 37608 185208 37660 185214
rect 37608 185150 37660 185156
rect 37896 185049 37924 185422
rect 38356 185078 38384 187868
rect 39000 185146 39028 187868
rect 39736 185282 39764 187868
rect 40380 185418 40408 187868
rect 41024 185486 41052 187868
rect 41012 185480 41064 185486
rect 41012 185422 41064 185428
rect 40368 185412 40420 185418
rect 40368 185354 40420 185360
rect 41760 185350 41788 187868
rect 40644 185344 40696 185350
rect 40644 185286 40696 185292
rect 41748 185344 41800 185350
rect 41748 185286 41800 185292
rect 39724 185276 39776 185282
rect 39724 185218 39776 185224
rect 38988 185140 39040 185146
rect 38988 185082 39040 185088
rect 38344 185072 38396 185078
rect 37882 185040 37938 185049
rect 38344 185014 38396 185020
rect 40274 185040 40330 185049
rect 37882 184975 37938 184984
rect 40274 184975 40330 184984
rect 36964 184936 37016 184942
rect 36964 184878 37016 184884
rect 40288 184740 40316 184975
rect 40656 184740 40684 185286
rect 41472 185208 41524 185214
rect 41472 185150 41524 185156
rect 41012 184936 41064 184942
rect 41012 184878 41064 184884
rect 41024 184740 41052 184878
rect 41484 184740 41512 185150
rect 42404 185146 42432 187868
rect 43140 185418 43168 187868
rect 43784 185486 43812 187868
rect 44534 187854 45100 187882
rect 45178 187854 45652 187882
rect 45822 187854 46112 187882
rect 43404 185480 43456 185486
rect 43404 185422 43456 185428
rect 43772 185480 43824 185486
rect 43772 185422 43824 185428
rect 44692 185480 44744 185486
rect 44692 185422 44744 185428
rect 43036 185412 43088 185418
rect 43036 185354 43088 185360
rect 43128 185412 43180 185418
rect 43128 185354 43180 185360
rect 42668 185276 42720 185282
rect 42668 185218 42720 185224
rect 42208 185140 42260 185146
rect 42208 185082 42260 185088
rect 42392 185140 42444 185146
rect 42392 185082 42444 185088
rect 41840 185072 41892 185078
rect 41840 185014 41892 185020
rect 41852 184740 41880 185014
rect 42220 184740 42248 185082
rect 42680 184740 42708 185218
rect 43048 184740 43076 185354
rect 43416 184740 43444 185422
rect 44600 185412 44652 185418
rect 44600 185354 44652 185360
rect 43864 185344 43916 185350
rect 43864 185286 43916 185292
rect 43876 184740 43904 185286
rect 44232 185140 44284 185146
rect 44232 185082 44284 185088
rect 44244 184740 44272 185082
rect 44612 184740 44640 185354
rect 44704 184754 44732 185422
rect 45072 184890 45100 187854
rect 45072 184862 45192 184890
rect 45164 184754 45192 184862
rect 45624 184754 45652 187854
rect 46084 184754 46112 187854
rect 46544 184754 46572 187868
rect 47188 184754 47216 187868
rect 47648 187854 47938 187882
rect 48200 187854 48582 187882
rect 48660 187854 49226 187882
rect 47648 184754 47676 187854
rect 48200 184754 48228 187854
rect 48660 185162 48688 187854
rect 49016 185480 49068 185486
rect 49016 185422 49068 185428
rect 48568 185134 48688 185162
rect 48568 184754 48596 185134
rect 48648 185072 48700 185078
rect 48648 185014 48700 185020
rect 44704 184726 45086 184754
rect 45164 184726 45454 184754
rect 45624 184726 45822 184754
rect 46084 184726 46282 184754
rect 46544 184726 46650 184754
rect 47110 184726 47216 184754
rect 47478 184726 47676 184754
rect 47846 184726 48228 184754
rect 48306 184726 48596 184754
rect 48660 184740 48688 185014
rect 49028 184740 49056 185422
rect 49476 185276 49528 185282
rect 49476 185218 49528 185224
rect 49488 184740 49516 185218
rect 49844 185140 49896 185146
rect 49844 185082 49896 185088
rect 49856 184740 49884 185082
rect 49948 185078 49976 187868
rect 50592 185486 50620 187868
rect 50580 185480 50632 185486
rect 50580 185422 50632 185428
rect 50672 185480 50724 185486
rect 50672 185422 50724 185428
rect 50212 185412 50264 185418
rect 50212 185354 50264 185360
rect 49936 185072 49988 185078
rect 49936 185014 49988 185020
rect 50224 184740 50252 185354
rect 50684 184740 50712 185422
rect 51328 185282 51356 187868
rect 51316 185276 51368 185282
rect 51316 185218 51368 185224
rect 51040 185208 51092 185214
rect 51040 185150 51092 185156
rect 51052 184740 51080 185150
rect 51972 185146 52000 187868
rect 52708 185418 52736 187868
rect 53352 185486 53380 187868
rect 53340 185480 53392 185486
rect 53340 185422 53392 185428
rect 53432 185480 53484 185486
rect 53432 185422 53484 185428
rect 52696 185412 52748 185418
rect 52696 185354 52748 185360
rect 52236 185344 52288 185350
rect 52236 185286 52288 185292
rect 51960 185140 52012 185146
rect 51960 185082 52012 185088
rect 51408 185072 51460 185078
rect 51408 185014 51460 185020
rect 51420 184740 51448 185014
rect 51868 185004 51920 185010
rect 51868 184946 51920 184952
rect 51880 184740 51908 184946
rect 52248 184740 52276 185286
rect 53064 185276 53116 185282
rect 53064 185218 53116 185224
rect 52604 185140 52656 185146
rect 52604 185082 52656 185088
rect 52616 184740 52644 185082
rect 53076 184740 53104 185218
rect 53444 184740 53472 185422
rect 53996 185214 54024 187868
rect 53984 185208 54036 185214
rect 53984 185150 54036 185156
rect 54732 185078 54760 187868
rect 54720 185072 54772 185078
rect 54720 185014 54772 185020
rect 55376 185010 55404 187868
rect 56112 185350 56140 187868
rect 56100 185344 56152 185350
rect 56100 185286 56152 185292
rect 56756 185146 56784 187868
rect 57400 185282 57428 187868
rect 58136 185486 58164 187868
rect 58124 185480 58176 185486
rect 58124 185422 58176 185428
rect 57388 185276 57440 185282
rect 57388 185218 57440 185224
rect 56744 185140 56796 185146
rect 56744 185082 56796 185088
rect 55364 185004 55416 185010
rect 55364 184946 55416 184952
rect 53826 184602 54024 184618
rect 58780 184602 58808 187868
rect 53826 184596 54036 184602
rect 53826 184590 53984 184596
rect 53984 184538 54036 184544
rect 58768 184596 58820 184602
rect 58768 184538 58820 184544
rect 37974 184496 38030 184505
rect 39630 184496 39686 184505
rect 37974 184431 38030 184440
rect 38908 184454 39106 184482
rect 39276 184466 39474 184482
rect 39264 184460 39474 184466
rect 37988 184330 38016 184431
rect 34940 184324 34992 184330
rect 34940 184266 34992 184272
rect 37976 184324 38028 184330
rect 37976 184266 38028 184272
rect 34204 184256 34256 184262
rect 34204 184198 34256 184204
rect 38908 184126 38936 184454
rect 39316 184454 39474 184460
rect 39686 184454 39842 184482
rect 54286 184466 54576 184482
rect 54286 184460 54588 184466
rect 54286 184454 54536 184460
rect 39630 184431 39686 184440
rect 39264 184402 39316 184408
rect 54654 184454 54944 184482
rect 54536 184402 54588 184408
rect 54916 184233 54944 184454
rect 59516 184262 59544 187868
rect 59504 184256 59556 184262
rect 54902 184224 54958 184233
rect 60160 184233 60188 187868
rect 105194 187610 105222 187868
rect 105148 187582 105222 187610
rect 105332 187854 105760 187882
rect 105884 187854 106312 187882
rect 106620 187854 106956 187882
rect 107172 187854 107508 187882
rect 107908 187854 108060 187882
rect 108368 187854 108704 187882
rect 109256 187854 109316 187882
rect 109808 187854 110144 187882
rect 110452 187854 110788 187882
rect 111004 187854 111432 187882
rect 111556 187854 111984 187882
rect 112200 187854 112444 187882
rect 112752 187854 113088 187882
rect 113304 187854 113456 187882
rect 59504 184198 59556 184204
rect 60146 184224 60202 184233
rect 54902 184159 54958 184168
rect 60146 184159 60202 184168
rect 33560 184120 33612 184126
rect 33560 184062 33612 184068
rect 38896 184120 38948 184126
rect 38896 184062 38948 184068
rect 31994 178240 32050 178249
rect 31994 178175 32050 178184
rect 37422 178240 37478 178249
rect 37422 178175 37478 178184
rect 59594 178240 59650 178249
rect 59594 178175 59650 178184
rect 37436 177258 37464 178175
rect 59608 177258 59636 178175
rect 32640 177252 32692 177258
rect 32640 177194 32692 177200
rect 37424 177252 37476 177258
rect 37424 177194 37476 177200
rect 57572 177252 57624 177258
rect 57572 177194 57624 177200
rect 59596 177252 59648 177258
rect 59596 177194 59648 177200
rect 12214 170080 12270 170089
rect 12214 170015 12270 170024
rect 32652 164921 32680 177194
rect 57584 174849 57612 177194
rect 105148 175801 105176 187582
rect 105332 183938 105360 187854
rect 105596 185276 105648 185282
rect 105596 185218 105648 185224
rect 105608 184777 105636 185218
rect 105594 184768 105650 184777
rect 105594 184703 105650 184712
rect 105240 183910 105360 183938
rect 105240 177161 105268 183910
rect 105596 182420 105648 182426
rect 105596 182362 105648 182368
rect 105608 182329 105636 182362
rect 105594 182320 105650 182329
rect 105594 182255 105650 182264
rect 105884 181218 105912 187854
rect 106056 184256 106108 184262
rect 106056 184198 106108 184204
rect 105964 184120 106016 184126
rect 105964 184062 106016 184068
rect 105332 181190 105912 181218
rect 105332 178521 105360 181190
rect 105412 180380 105464 180386
rect 105412 180322 105464 180328
rect 105318 178512 105374 178521
rect 105318 178447 105374 178456
rect 105226 177152 105282 177161
rect 105226 177087 105282 177096
rect 105134 175792 105190 175801
rect 105134 175727 105190 175736
rect 57570 174840 57626 174849
rect 57570 174775 57626 174784
rect 105424 173761 105452 180322
rect 105976 179881 106004 184062
rect 106068 181105 106096 184198
rect 106620 184126 106648 187854
rect 107172 184262 107200 187854
rect 107160 184256 107212 184262
rect 107160 184198 107212 184204
rect 106608 184120 106660 184126
rect 106608 184062 106660 184068
rect 106148 184052 106200 184058
rect 106148 183994 106200 184000
rect 106160 183553 106188 183994
rect 106146 183544 106202 183553
rect 106146 183479 106202 183488
rect 107908 182426 107936 187854
rect 108368 184126 108396 187854
rect 109288 185282 109316 187854
rect 110116 185486 110144 187854
rect 110104 185480 110156 185486
rect 110104 185422 110156 185428
rect 110760 185418 110788 187854
rect 111404 185570 111432 187854
rect 111404 185542 111616 185570
rect 111116 185480 111168 185486
rect 111116 185422 111168 185428
rect 110748 185412 110800 185418
rect 110748 185354 110800 185360
rect 109276 185276 109328 185282
rect 109276 185218 109328 185224
rect 111128 184740 111156 185422
rect 111484 185412 111536 185418
rect 111484 185354 111536 185360
rect 111496 184740 111524 185354
rect 111588 184754 111616 185542
rect 111956 184754 111984 187854
rect 112416 184754 112444 187854
rect 111588 184726 111878 184754
rect 111956 184726 112338 184754
rect 112416 184726 112706 184754
rect 113060 184740 113088 187854
rect 113428 184754 113456 187854
rect 113934 187610 113962 187868
rect 113888 187582 113962 187610
rect 114256 187854 114500 187882
rect 114716 187854 115052 187882
rect 115360 187854 115696 187882
rect 115820 187854 116248 187882
rect 116372 187854 116800 187882
rect 113428 184726 113534 184754
rect 113888 184740 113916 187582
rect 114256 184740 114284 187854
rect 114716 184740 114744 187854
rect 115360 184754 115388 187854
rect 115820 184754 115848 187854
rect 116372 184890 116400 187854
rect 117430 187662 117458 187868
rect 117660 187854 117996 187882
rect 118212 187854 118548 187882
rect 118948 187854 119192 187882
rect 119592 187854 119744 187882
rect 120296 187854 120356 187882
rect 116452 187656 116504 187662
rect 116452 187598 116504 187604
rect 117418 187656 117470 187662
rect 117418 187598 117470 187604
rect 116188 184862 116400 184890
rect 116188 184754 116216 184862
rect 116464 184754 116492 187598
rect 117094 185448 117150 185457
rect 117094 185383 117150 185392
rect 116910 184768 116966 184777
rect 115098 184726 115388 184754
rect 115466 184726 115848 184754
rect 115926 184726 116216 184754
rect 116294 184726 116492 184754
rect 116662 184726 116910 184754
rect 117108 184740 117136 185383
rect 117462 185312 117518 185321
rect 117462 185247 117518 185256
rect 117476 184740 117504 185247
rect 117660 184777 117688 187854
rect 118212 185457 118240 187854
rect 118198 185448 118254 185457
rect 118198 185383 118254 185392
rect 118658 185448 118714 185457
rect 118658 185383 118714 185392
rect 118290 185176 118346 185185
rect 118290 185111 118346 185120
rect 117646 184768 117702 184777
rect 116910 184703 116966 184712
rect 118106 184768 118162 184777
rect 117858 184726 118106 184754
rect 117646 184703 117702 184712
rect 118304 184740 118332 185111
rect 118672 184740 118700 185383
rect 118948 185321 118976 187854
rect 118934 185312 118990 185321
rect 118934 185247 118990 185256
rect 119118 185040 119174 185049
rect 119118 184975 119174 184984
rect 119132 184740 119160 184975
rect 119592 184777 119620 187854
rect 120328 185185 120356 187854
rect 120604 187854 120940 187882
rect 121156 187854 121492 187882
rect 121708 187854 122044 187882
rect 122688 187854 122840 187882
rect 120604 185457 120632 187854
rect 120590 185448 120646 185457
rect 120590 185383 120646 185392
rect 120958 185448 121014 185457
rect 120958 185383 121014 185392
rect 120314 185176 120370 185185
rect 120314 185111 120370 185120
rect 120590 185176 120646 185185
rect 120590 185111 120646 185120
rect 119670 184904 119726 184913
rect 119670 184839 119726 184848
rect 119578 184768 119634 184777
rect 118106 184703 118162 184712
rect 119578 184703 119634 184712
rect 119684 184618 119712 184839
rect 120604 184754 120632 185111
rect 120972 184754 121000 185383
rect 121050 185312 121106 185321
rect 121050 185247 121106 185256
rect 120342 184726 120632 184754
rect 120710 184726 121000 184754
rect 121064 184740 121092 185247
rect 121156 185049 121184 187854
rect 121708 185049 121736 187854
rect 121880 186908 121932 186914
rect 121880 186850 121932 186856
rect 121142 185040 121198 185049
rect 121142 184975 121198 184984
rect 121694 185040 121750 185049
rect 121694 184975 121750 184984
rect 121602 184904 121658 184913
rect 121602 184839 121658 184848
rect 121616 184754 121644 184839
rect 121538 184726 121644 184754
rect 121892 184740 121920 186850
rect 122706 185040 122762 185049
rect 122706 184975 122762 184984
rect 122522 184768 122578 184777
rect 122274 184726 122522 184754
rect 122720 184740 122748 184975
rect 122522 184703 122578 184712
rect 122812 184641 122840 187854
rect 123088 187854 123240 187882
rect 123456 187854 123792 187882
rect 124436 187854 124496 187882
rect 123088 185185 123116 187854
rect 123456 185457 123484 187854
rect 123442 185448 123498 185457
rect 123442 185383 123498 185392
rect 123902 185448 123958 185457
rect 123902 185383 123958 185392
rect 123074 185176 123130 185185
rect 123074 185111 123130 185120
rect 123350 185176 123406 185185
rect 123350 185111 123406 185120
rect 123364 184754 123392 185111
rect 123102 184726 123392 184754
rect 123916 184740 123944 185383
rect 124362 185312 124418 185321
rect 124468 185298 124496 187854
rect 124418 185270 124496 185298
rect 124560 187854 124988 187882
rect 125204 187854 125540 187882
rect 125848 187854 126184 187882
rect 126400 187854 126736 187882
rect 127288 187854 127348 187882
rect 124362 185247 124418 185256
rect 124362 184904 124418 184913
rect 124560 184890 124588 187854
rect 125204 186914 125232 187854
rect 125192 186908 125244 186914
rect 125192 186850 125244 186856
rect 124824 185276 124876 185282
rect 124824 185218 124876 185224
rect 124836 185049 124864 185218
rect 125098 185176 125154 185185
rect 125098 185111 125154 185120
rect 124822 185040 124878 185049
rect 124822 184975 124878 184984
rect 124418 184862 124588 184890
rect 124914 184904 124970 184913
rect 124362 184839 124418 184848
rect 124914 184839 124970 184848
rect 124928 184754 124956 184839
rect 124666 184726 124956 184754
rect 125112 184740 125140 185111
rect 125466 185040 125522 185049
rect 125466 184975 125522 184984
rect 125480 184740 125508 184975
rect 125848 184890 125876 187854
rect 125928 185480 125980 185486
rect 125926 185448 125928 185457
rect 125980 185448 125982 185457
rect 125926 185383 125982 185392
rect 125928 185344 125980 185350
rect 125926 185312 125928 185321
rect 125980 185312 125982 185321
rect 125926 185247 125982 185256
rect 126110 185312 126166 185321
rect 126400 185282 126428 187854
rect 126662 185448 126718 185457
rect 126662 185383 126718 185392
rect 127216 185412 127268 185418
rect 126110 185247 126166 185256
rect 126388 185276 126440 185282
rect 125664 184862 125876 184890
rect 125664 184777 125692 184862
rect 125650 184768 125706 184777
rect 126124 184754 126152 185247
rect 126388 185218 126440 185224
rect 126478 184768 126534 184777
rect 125862 184726 126152 184754
rect 126322 184726 126478 184754
rect 125650 184703 125706 184712
rect 126676 184740 126704 185383
rect 127216 185354 127268 185360
rect 127228 185185 127256 185354
rect 127320 185350 127348 187854
rect 127596 187854 127932 187882
rect 128148 187854 128484 187882
rect 128700 187854 129036 187882
rect 129344 187854 129680 187882
rect 129988 187854 130232 187882
rect 130448 187854 130784 187882
rect 131428 187854 131488 187882
rect 127308 185344 127360 185350
rect 127308 185286 127360 185292
rect 127214 185176 127270 185185
rect 127214 185111 127270 185120
rect 127216 185072 127268 185078
rect 127214 185040 127216 185049
rect 127268 185040 127270 185049
rect 127214 184975 127270 184984
rect 127216 184936 127268 184942
rect 127214 184904 127216 184913
rect 127268 184904 127270 184913
rect 127214 184839 127270 184848
rect 126478 184703 126534 184712
rect 127032 184732 127084 184738
rect 127032 184674 127084 184680
rect 127044 184641 127072 184674
rect 120130 184632 120186 184641
rect 119514 184590 119712 184618
rect 119882 184590 120130 184618
rect 120130 184567 120186 184576
rect 122798 184632 122854 184641
rect 124362 184632 124418 184641
rect 124298 184590 124362 184618
rect 122798 184567 122854 184576
rect 124362 184567 124418 184576
rect 127030 184632 127086 184641
rect 127030 184567 127086 184576
rect 127596 184534 127624 187854
rect 128148 185486 128176 187854
rect 128136 185480 128188 185486
rect 128136 185422 128188 185428
rect 128700 184738 128728 187854
rect 129344 184942 129372 187854
rect 129988 185418 130016 187854
rect 129976 185412 130028 185418
rect 129976 185354 130028 185360
rect 130448 185078 130476 187854
rect 131460 185321 131488 187854
rect 131644 187854 131980 187882
rect 132196 187854 132532 187882
rect 176908 187854 177198 187882
rect 131446 185312 131502 185321
rect 131446 185247 131502 185256
rect 130436 185072 130488 185078
rect 130436 185014 130488 185020
rect 129332 184936 129384 184942
rect 129332 184878 129384 184884
rect 131644 184777 131672 187854
rect 132092 186908 132144 186914
rect 132092 186850 132144 186856
rect 131630 184768 131686 184777
rect 128688 184732 128740 184738
rect 131630 184703 131686 184712
rect 128688 184674 128740 184680
rect 127032 184528 127084 184534
rect 123718 184496 123774 184505
rect 123470 184454 123718 184482
rect 123718 184431 123774 184440
rect 127030 184496 127032 184505
rect 127584 184528 127636 184534
rect 127084 184496 127086 184505
rect 127584 184470 127636 184476
rect 127030 184431 127086 184440
rect 108356 184120 108408 184126
rect 108356 184062 108408 184068
rect 108538 183544 108594 183553
rect 108538 183479 108594 183488
rect 107896 182420 107948 182426
rect 107896 182362 107948 182368
rect 108078 181232 108134 181241
rect 108078 181167 108134 181176
rect 106054 181096 106110 181105
rect 106054 181031 106110 181040
rect 108092 180386 108120 181167
rect 108080 180380 108132 180386
rect 108080 180322 108132 180328
rect 105962 179872 106018 179881
rect 105962 179807 106018 179816
rect 107894 178920 107950 178929
rect 107894 178855 107950 178864
rect 107908 178618 107936 178855
rect 106332 178612 106384 178618
rect 106332 178554 106384 178560
rect 107896 178612 107948 178618
rect 107896 178554 107948 178560
rect 106146 174432 106202 174441
rect 106146 174367 106148 174376
rect 106200 174367 106202 174376
rect 106148 174338 106200 174344
rect 105410 173752 105466 173761
rect 105410 173687 105466 173696
rect 106056 173104 106108 173110
rect 106056 173046 106108 173052
rect 105228 171744 105280 171750
rect 105228 171686 105280 171692
rect 105240 168865 105268 171686
rect 106068 170225 106096 173046
rect 106344 172537 106372 178554
rect 107894 176472 107950 176481
rect 107894 176407 107950 176416
rect 107908 175898 107936 176407
rect 106424 175892 106476 175898
rect 106424 175834 106476 175840
rect 107896 175892 107948 175898
rect 107896 175834 107948 175840
rect 106330 172528 106386 172537
rect 106330 172463 106386 172472
rect 106436 171449 106464 175834
rect 108552 174402 108580 183479
rect 108540 174396 108592 174402
rect 108540 174338 108592 174344
rect 108170 174160 108226 174169
rect 108170 174095 108226 174104
rect 108184 173110 108212 174095
rect 108172 173104 108224 173110
rect 108172 173046 108224 173052
rect 107894 171848 107950 171857
rect 107894 171783 107950 171792
rect 107908 171750 107936 171783
rect 107896 171744 107948 171750
rect 107896 171686 107948 171692
rect 106422 171440 106478 171449
rect 106422 171375 106478 171384
rect 106054 170216 106110 170225
rect 106054 170151 106110 170160
rect 107894 169400 107950 169409
rect 107894 169335 107950 169344
rect 107908 168962 107936 169335
rect 105964 168956 106016 168962
rect 105964 168898 106016 168904
rect 107896 168956 107948 168962
rect 107896 168898 107948 168904
rect 105226 168856 105282 168865
rect 105226 168791 105282 168800
rect 105976 167505 106004 168898
rect 105962 167496 106018 167505
rect 105962 167431 106018 167440
rect 107802 167088 107858 167097
rect 107802 167023 107858 167032
rect 107816 166174 107844 167023
rect 106424 166168 106476 166174
rect 106422 166136 106424 166145
rect 107804 166168 107856 166174
rect 106476 166136 106478 166145
rect 107804 166110 107856 166116
rect 106422 166071 106478 166080
rect 32638 164912 32694 164921
rect 32638 164847 32694 164856
rect 37422 164912 37478 164921
rect 59594 164912 59650 164921
rect 37422 164847 37478 164856
rect 54732 164870 54944 164898
rect 37436 164814 37464 164847
rect 28868 164808 28920 164814
rect 28868 164750 28920 164756
rect 37424 164808 37476 164814
rect 37424 164750 37476 164756
rect 12214 159336 12270 159345
rect 12214 159271 12270 159280
rect 12228 106169 12256 159271
rect 28880 156466 28908 164750
rect 28788 156438 28908 156466
rect 12582 149408 12638 149417
rect 12582 149343 12638 149352
rect 12596 142617 12624 149343
rect 28788 146930 28816 156438
rect 31994 151584 32050 151593
rect 31994 151519 32050 151528
rect 28776 146924 28828 146930
rect 28776 146866 28828 146872
rect 22244 145224 22296 145230
rect 21948 145172 22244 145178
rect 21948 145166 22296 145172
rect 21948 145150 22284 145166
rect 16598 144634 16626 144892
rect 27284 144878 27620 144906
rect 16598 144606 16672 144634
rect 16644 142646 16672 144606
rect 16632 142640 16684 142646
rect 12582 142608 12638 142617
rect 16632 142582 16684 142588
rect 12582 142543 12638 142552
rect 27592 142510 27620 144878
rect 31812 142640 31864 142646
rect 31812 142582 31864 142588
rect 27580 142504 27632 142510
rect 27580 142446 27632 142452
rect 31824 141393 31852 142582
rect 32008 142322 32036 151519
rect 39092 142714 39120 144892
rect 34112 142708 34164 142714
rect 34112 142650 34164 142656
rect 39080 142708 39132 142714
rect 39080 142650 39132 142656
rect 32008 142294 32956 142322
rect 32928 141778 32956 142294
rect 34124 141778 34152 142650
rect 39460 142578 39488 144892
rect 34664 142572 34716 142578
rect 34664 142514 34716 142520
rect 39448 142572 39500 142578
rect 39448 142514 39500 142520
rect 34676 141778 34704 142514
rect 37240 142436 37292 142442
rect 37240 142378 37292 142384
rect 36596 142300 36648 142306
rect 36596 142242 36648 142248
rect 35584 141824 35636 141830
rect 32928 141750 33218 141778
rect 33862 141750 34152 141778
rect 34506 141750 34704 141778
rect 35242 141772 35584 141778
rect 35242 141766 35636 141772
rect 35242 141750 35624 141766
rect 36608 141764 36636 142242
rect 37252 141764 37280 142378
rect 39264 142368 39316 142374
rect 39264 142310 39316 142316
rect 38620 142232 38672 142238
rect 38620 142174 38672 142180
rect 37884 142164 37936 142170
rect 37884 142106 37936 142112
rect 37896 141764 37924 142106
rect 38632 141764 38660 142174
rect 39276 141764 39304 142310
rect 39828 141830 39856 144892
rect 40000 142708 40052 142714
rect 40000 142650 40052 142656
rect 39816 141824 39868 141830
rect 39816 141766 39868 141772
rect 40012 141764 40040 142650
rect 35952 141688 36004 141694
rect 35886 141636 35952 141642
rect 35886 141630 36004 141636
rect 40184 141688 40236 141694
rect 40288 141676 40316 144892
rect 40380 144878 40670 144906
rect 40380 142306 40408 144878
rect 40644 144204 40696 144210
rect 40644 144146 40696 144152
rect 40368 142300 40420 142306
rect 40368 142242 40420 142248
rect 40656 141764 40684 144146
rect 41024 142442 41052 144892
rect 41288 144136 41340 144142
rect 41288 144078 41340 144084
rect 41012 142436 41064 142442
rect 41012 142378 41064 142384
rect 41300 141764 41328 144078
rect 41484 142170 41512 144892
rect 41852 142238 41880 144892
rect 42024 142572 42076 142578
rect 42024 142514 42076 142520
rect 41840 142232 41892 142238
rect 41840 142174 41892 142180
rect 41472 142164 41524 142170
rect 41472 142106 41524 142112
rect 42036 141764 42064 142514
rect 42220 142374 42248 144892
rect 42312 144878 42694 144906
rect 42312 142714 42340 144878
rect 43048 144210 43076 144892
rect 43036 144204 43088 144210
rect 43036 144146 43088 144152
rect 43416 144142 43444 144892
rect 43404 144136 43456 144142
rect 43404 144078 43456 144084
rect 42300 142708 42352 142714
rect 42300 142650 42352 142656
rect 42668 142708 42720 142714
rect 42668 142650 42720 142656
rect 42208 142368 42260 142374
rect 42208 142310 42260 142316
rect 42680 141764 42708 142650
rect 43876 142578 43904 144892
rect 44244 142714 44272 144892
rect 44232 142708 44284 142714
rect 44232 142650 44284 142656
rect 43864 142572 43916 142578
rect 43864 142514 43916 142520
rect 44612 142306 44640 144892
rect 44704 144878 45086 144906
rect 45164 144878 45454 144906
rect 43404 142300 43456 142306
rect 43404 142242 43456 142248
rect 44600 142300 44652 142306
rect 44600 142242 44652 142248
rect 43416 141764 43444 142242
rect 44704 141914 44732 144878
rect 44520 141886 44732 141914
rect 44520 141778 44548 141886
rect 45164 141778 45192 144878
rect 45808 142306 45836 144892
rect 45428 142300 45480 142306
rect 45428 142242 45480 142248
rect 45796 142300 45848 142306
rect 45796 142242 45848 142248
rect 44074 141750 44548 141778
rect 44810 141750 45192 141778
rect 45440 141764 45468 142242
rect 46268 141778 46296 144892
rect 46098 141750 46296 141778
rect 46636 141778 46664 144892
rect 47096 141778 47124 144892
rect 47478 144878 47768 144906
rect 47740 141778 47768 144878
rect 47832 142714 47860 144892
rect 47820 142708 47872 142714
rect 47820 142650 47872 142656
rect 48292 142578 48320 144892
rect 48280 142572 48332 142578
rect 48280 142514 48332 142520
rect 48660 142510 48688 144892
rect 49028 142714 49056 144892
rect 49502 144878 49792 144906
rect 48832 142708 48884 142714
rect 48832 142650 48884 142656
rect 49016 142708 49068 142714
rect 49016 142650 49068 142656
rect 48648 142504 48700 142510
rect 48648 142446 48700 142452
rect 46636 141750 46834 141778
rect 47096 141750 47478 141778
rect 47740 141750 48214 141778
rect 48844 141764 48872 142650
rect 49476 142572 49528 142578
rect 49476 142514 49528 142520
rect 49488 141764 49516 142514
rect 49764 142306 49792 144878
rect 49752 142300 49804 142306
rect 49752 142242 49804 142248
rect 49856 142170 49884 144892
rect 50238 144878 50528 144906
rect 50500 142578 50528 144878
rect 50488 142572 50540 142578
rect 50488 142514 50540 142520
rect 50684 142510 50712 144892
rect 51052 142714 51080 144892
rect 50856 142708 50908 142714
rect 50856 142650 50908 142656
rect 51040 142708 51092 142714
rect 51040 142650 51092 142656
rect 50212 142504 50264 142510
rect 50212 142446 50264 142452
rect 50672 142504 50724 142510
rect 50672 142446 50724 142452
rect 49844 142164 49896 142170
rect 49844 142106 49896 142112
rect 50224 141764 50252 142446
rect 50868 141764 50896 142650
rect 51420 142442 51448 144892
rect 51408 142436 51460 142442
rect 51408 142378 51460 142384
rect 51592 142300 51644 142306
rect 51592 142242 51644 142248
rect 51604 141764 51632 142242
rect 51880 142102 51908 144892
rect 52262 144878 52552 144906
rect 52524 144550 52552 144878
rect 52512 144544 52564 144550
rect 52512 144486 52564 144492
rect 52616 142170 52644 144892
rect 52972 142572 53024 142578
rect 52972 142514 53024 142520
rect 52236 142164 52288 142170
rect 52236 142106 52288 142112
rect 52604 142164 52656 142170
rect 52604 142106 52656 142112
rect 51868 142096 51920 142102
rect 51868 142038 51920 142044
rect 52248 141764 52276 142106
rect 52984 141764 53012 142514
rect 53076 142034 53104 144892
rect 53064 142028 53116 142034
rect 53064 141970 53116 141976
rect 53444 141694 53472 144892
rect 53616 142504 53668 142510
rect 53616 142446 53668 142452
rect 53628 141764 53656 142446
rect 53812 141694 53840 144892
rect 54272 144210 54300 144892
rect 54640 144278 54668 144892
rect 54628 144272 54680 144278
rect 54628 144214 54680 144220
rect 54260 144204 54312 144210
rect 54260 144146 54312 144152
rect 54260 142708 54312 142714
rect 54260 142650 54312 142656
rect 54272 141764 54300 142650
rect 54732 142374 54760 164870
rect 54916 164814 54944 164870
rect 59594 164847 59650 164856
rect 59608 164814 59636 164847
rect 54904 164808 54956 164814
rect 54904 164750 54956 164756
rect 59596 164808 59648 164814
rect 59596 164750 59648 164756
rect 106422 163552 106478 163561
rect 106422 163487 106424 163496
rect 106476 163487 106478 163496
rect 107804 163516 107856 163522
rect 106424 163458 106476 163464
rect 107804 163458 107856 163464
rect 107816 162473 107844 163458
rect 107802 162464 107858 162473
rect 107802 162399 107858 162408
rect 106146 162192 106202 162201
rect 106146 162127 106148 162136
rect 106200 162127 106202 162136
rect 108540 162156 108592 162162
rect 106148 162098 106200 162104
rect 108540 162098 108592 162104
rect 105778 160696 105834 160705
rect 105778 160631 105780 160640
rect 105832 160631 105834 160640
rect 107804 160660 107856 160666
rect 105780 160602 105832 160608
rect 107804 160602 107856 160608
rect 106422 159336 106478 159345
rect 106422 159271 106424 159280
rect 106476 159271 106478 159280
rect 107712 159300 107764 159306
rect 106424 159242 106476 159248
rect 107712 159242 107764 159248
rect 105410 158384 105466 158393
rect 105410 158319 105466 158328
rect 105424 158218 105452 158319
rect 105412 158212 105464 158218
rect 105412 158154 105464 158160
rect 105410 157024 105466 157033
rect 105410 156959 105412 156968
rect 105464 156959 105466 156968
rect 107252 156988 107304 156994
rect 105412 156930 105464 156936
rect 107252 156930 107304 156936
rect 105226 155800 105282 155809
rect 105226 155735 105228 155744
rect 105280 155735 105282 155744
rect 107160 155764 107212 155770
rect 105228 155706 105280 155712
rect 107160 155706 107212 155712
rect 57478 154848 57534 154857
rect 57478 154783 57534 154792
rect 57492 151554 57520 154783
rect 105778 154576 105834 154585
rect 105778 154511 105834 154520
rect 105594 153896 105650 153905
rect 105594 153831 105596 153840
rect 105648 153831 105650 153840
rect 105596 153802 105648 153808
rect 105792 153798 105820 154511
rect 105780 153792 105832 153798
rect 105780 153734 105832 153740
rect 106422 152536 106478 152545
rect 106478 152494 106556 152522
rect 106422 152471 106478 152480
rect 59594 151584 59650 151593
rect 57480 151548 57532 151554
rect 59594 151519 59596 151528
rect 57480 151490 57532 151496
rect 59648 151519 59650 151528
rect 59596 151490 59648 151496
rect 55364 144544 55416 144550
rect 55364 144486 55416 144492
rect 55376 144142 55404 144486
rect 55364 144136 55416 144142
rect 55364 144078 55416 144084
rect 56376 144136 56428 144142
rect 56376 144078 56428 144084
rect 54996 142436 55048 142442
rect 54996 142378 55048 142384
rect 54720 142368 54772 142374
rect 54720 142310 54772 142316
rect 55008 141764 55036 142378
rect 55364 142096 55416 142102
rect 55364 142038 55416 142044
rect 55376 141778 55404 142038
rect 55376 141750 55666 141778
rect 56388 141764 56416 144078
rect 57492 142238 57520 151490
rect 105962 149680 106018 149689
rect 105962 149615 106018 149624
rect 105410 148456 105466 148465
rect 105410 148391 105466 148400
rect 105226 147232 105282 147241
rect 105226 147167 105282 147176
rect 60424 144272 60476 144278
rect 60424 144214 60476 144220
rect 59780 144204 59832 144210
rect 59780 144146 59832 144152
rect 57480 142232 57532 142238
rect 57480 142174 57532 142180
rect 57020 142164 57072 142170
rect 57020 142106 57072 142112
rect 57032 141764 57060 142106
rect 57664 142028 57716 142034
rect 57664 141970 57716 141976
rect 57676 141764 57704 141970
rect 58688 141762 59070 141778
rect 59792 141764 59820 144146
rect 60436 141764 60464 144214
rect 62816 142708 62868 142714
rect 62816 142650 62868 142656
rect 62356 142164 62408 142170
rect 62356 142106 62408 142112
rect 58676 141756 59070 141762
rect 58728 141750 59070 141756
rect 58676 141698 58728 141704
rect 40236 141648 40316 141676
rect 53432 141688 53484 141694
rect 40184 141630 40236 141636
rect 53432 141630 53484 141636
rect 53800 141688 53852 141694
rect 53800 141630 53852 141636
rect 58216 141688 58268 141694
rect 58268 141636 58426 141642
rect 58216 141630 58426 141636
rect 35886 141614 35992 141630
rect 58228 141614 58426 141630
rect 31810 141384 31866 141393
rect 31810 141319 31866 141328
rect 62368 139806 62396 142106
rect 62828 142073 62856 142650
rect 63472 142170 63500 144892
rect 63460 142164 63512 142170
rect 63460 142106 63512 142112
rect 62814 142064 62870 142073
rect 64576 142034 64604 144892
rect 65128 144878 65694 144906
rect 66600 144878 66798 144906
rect 62814 141999 62870 142008
rect 63460 142028 63512 142034
rect 63460 141970 63512 141976
rect 64564 142028 64616 142034
rect 64564 141970 64616 141976
rect 62816 141280 62868 141286
rect 62816 141222 62868 141228
rect 62724 141212 62776 141218
rect 62724 141154 62776 141160
rect 62736 140713 62764 141154
rect 62828 140985 62856 141222
rect 62814 140976 62870 140985
rect 62814 140911 62870 140920
rect 62722 140704 62778 140713
rect 62722 140639 62778 140648
rect 62816 139920 62868 139926
rect 62816 139862 62868 139868
rect 62368 139778 62580 139806
rect 62356 139716 62408 139722
rect 62356 139658 62408 139664
rect 62368 139489 62396 139658
rect 62354 139480 62410 139489
rect 62354 139415 62410 139424
rect 62552 137721 62580 139778
rect 62828 139761 62856 139862
rect 62814 139752 62870 139761
rect 62814 139687 62870 139696
rect 62816 139308 62868 139314
rect 62816 139250 62868 139256
rect 62828 138945 62856 139250
rect 62814 138936 62870 138945
rect 62814 138871 62870 138880
rect 62908 138696 62960 138702
rect 62908 138638 62960 138644
rect 62816 138628 62868 138634
rect 62816 138570 62868 138576
rect 62538 137712 62594 137721
rect 62538 137647 62594 137656
rect 62632 137268 62684 137274
rect 62632 137210 62684 137216
rect 30522 137168 30578 137177
rect 30522 137103 30578 137112
rect 30430 127784 30486 127793
rect 30430 127719 30486 127728
rect 30444 114358 30472 127719
rect 30432 114352 30484 114358
rect 30432 114294 30484 114300
rect 12214 106160 12270 106169
rect 12214 106095 12270 106104
rect 12122 95824 12178 95833
rect 12122 95759 12178 95768
rect 28512 90342 28908 90370
rect 28512 88874 28540 90342
rect 28880 90286 28908 90342
rect 28868 90280 28920 90286
rect 28868 90222 28920 90228
rect 28512 88846 28632 88874
rect 28604 79218 28632 88846
rect 28604 79190 28724 79218
rect 16598 70650 16626 70908
rect 21948 70894 22284 70922
rect 27284 70894 27620 70922
rect 16598 70622 16672 70650
rect 16644 69478 16672 70622
rect 22256 69546 22284 70894
rect 22244 69540 22296 69546
rect 22244 69482 22296 69488
rect 16632 69472 16684 69478
rect 16632 69414 16684 69420
rect 27592 69342 27620 70894
rect 28696 69546 28724 79190
rect 30536 77842 30564 137103
rect 62644 135409 62672 137210
rect 62724 137200 62776 137206
rect 62828 137177 62856 138570
rect 62724 137142 62776 137148
rect 62814 137168 62870 137177
rect 62736 135681 62764 137142
rect 62814 137103 62870 137112
rect 62920 136633 62948 138638
rect 63472 138401 63500 141970
rect 65128 139314 65156 144878
rect 66496 142708 66548 142714
rect 66496 142650 66548 142656
rect 66508 139926 66536 142650
rect 66496 139920 66548 139926
rect 66496 139862 66548 139868
rect 66600 139722 66628 144878
rect 67888 142714 67916 144892
rect 68072 144878 69006 144906
rect 69268 144878 70110 144906
rect 67876 142708 67928 142714
rect 67876 142650 67928 142656
rect 68072 141218 68100 144878
rect 69164 142436 69216 142442
rect 69164 142378 69216 142384
rect 68060 141212 68112 141218
rect 68060 141154 68112 141160
rect 69176 139738 69204 142378
rect 69268 141286 69296 144878
rect 71200 142578 71228 144892
rect 71188 142572 71240 142578
rect 71188 142514 71240 142520
rect 72304 142442 72332 144892
rect 72844 142708 72896 142714
rect 72844 142650 72896 142656
rect 72292 142436 72344 142442
rect 72292 142378 72344 142384
rect 71004 141892 71056 141898
rect 71004 141834 71056 141840
rect 69256 141280 69308 141286
rect 69256 141222 69308 141228
rect 71016 139738 71044 141834
rect 72856 139738 72884 142650
rect 73408 141898 73436 144892
rect 74512 142714 74540 144892
rect 75616 142714 75644 144892
rect 76260 144878 76826 144906
rect 77930 144878 78128 144906
rect 79034 144878 80060 144906
rect 74500 142708 74552 142714
rect 74500 142650 74552 142656
rect 74776 142708 74828 142714
rect 74776 142650 74828 142656
rect 75604 142708 75656 142714
rect 75604 142650 75656 142656
rect 73396 141892 73448 141898
rect 73396 141834 73448 141840
rect 74788 141370 74816 142650
rect 74696 141342 74816 141370
rect 74696 139738 74724 141342
rect 66588 139716 66640 139722
rect 68868 139710 69204 139738
rect 70708 139710 71044 139738
rect 72548 139710 72884 139738
rect 74480 139710 74724 139738
rect 76260 139738 76288 144878
rect 78100 139738 78128 144878
rect 80032 139738 80060 144878
rect 80124 142714 80152 144892
rect 80112 142708 80164 142714
rect 80112 142650 80164 142656
rect 81228 142646 81256 144892
rect 81676 142708 81728 142714
rect 81676 142650 81728 142656
rect 81216 142640 81268 142646
rect 81216 142582 81268 142588
rect 81688 139738 81716 142650
rect 82332 141558 82360 144892
rect 83436 142374 83464 144892
rect 83516 142640 83568 142646
rect 83516 142582 83568 142588
rect 83424 142368 83476 142374
rect 83424 142310 83476 142316
rect 82320 141552 82372 141558
rect 82320 141494 82372 141500
rect 83528 139738 83556 142582
rect 84540 141898 84568 144892
rect 85644 142714 85672 144892
rect 85632 142708 85684 142714
rect 85632 142650 85684 142656
rect 86748 142646 86776 144892
rect 86736 142640 86788 142646
rect 86736 142582 86788 142588
rect 87852 142510 87880 144892
rect 87840 142504 87892 142510
rect 87840 142446 87892 142452
rect 87288 142368 87340 142374
rect 87288 142310 87340 142316
rect 84528 141892 84580 141898
rect 84528 141834 84580 141840
rect 85356 141552 85408 141558
rect 85356 141494 85408 141500
rect 85368 139738 85396 141494
rect 87300 139738 87328 142310
rect 88956 142034 88984 144892
rect 88944 142028 88996 142034
rect 88944 141970 88996 141976
rect 90152 141937 90180 144892
rect 90968 142708 91020 142714
rect 90968 142650 91020 142656
rect 90138 141928 90194 141937
rect 89128 141892 89180 141898
rect 90138 141863 90194 141872
rect 89128 141834 89180 141840
rect 89140 139738 89168 141834
rect 90980 139738 91008 142650
rect 91256 141393 91284 144892
rect 92360 142238 92388 144892
rect 92808 142640 92860 142646
rect 92808 142582 92860 142588
rect 92348 142232 92400 142238
rect 92348 142174 92400 142180
rect 91242 141384 91298 141393
rect 91242 141319 91298 141328
rect 92820 139738 92848 142582
rect 93464 142306 93492 144892
rect 94108 144878 94582 144906
rect 95580 144878 95686 144906
rect 93452 142300 93504 142306
rect 93452 142242 93504 142248
rect 94108 139790 94136 144878
rect 95476 142708 95528 142714
rect 95476 142650 95528 142656
rect 94740 142504 94792 142510
rect 94740 142446 94792 142452
rect 94096 139784 94148 139790
rect 76260 139710 76320 139738
rect 78100 139710 78160 139738
rect 80032 139710 80092 139738
rect 81688 139710 81932 139738
rect 83528 139710 83864 139738
rect 85368 139710 85704 139738
rect 87300 139710 87544 139738
rect 89140 139710 89476 139738
rect 90980 139710 91316 139738
rect 92820 139710 93156 139738
rect 94096 139726 94148 139732
rect 94752 139738 94780 142446
rect 95488 139926 95516 142650
rect 95476 139920 95528 139926
rect 95476 139862 95528 139868
rect 95580 139858 95608 144878
rect 96776 142714 96804 144892
rect 96764 142708 96816 142714
rect 96764 142650 96816 142656
rect 97224 142232 97276 142238
rect 97224 142174 97276 142180
rect 96856 142028 96908 142034
rect 96856 141970 96908 141976
rect 95568 139852 95620 139858
rect 95568 139794 95620 139800
rect 96868 139738 96896 141970
rect 94752 139710 95088 139738
rect 96868 139710 96928 139738
rect 66588 139658 66640 139664
rect 66218 139480 66274 139489
rect 66218 139415 66274 139424
rect 65116 139308 65168 139314
rect 65116 139250 65168 139256
rect 66232 138634 66260 139415
rect 66402 138936 66458 138945
rect 66402 138871 66458 138880
rect 66416 138702 66444 138871
rect 66404 138696 66456 138702
rect 66404 138638 66456 138644
rect 66220 138628 66272 138634
rect 66220 138570 66272 138576
rect 97236 138498 97264 142174
rect 97880 141354 97908 144892
rect 98984 142374 99012 144892
rect 98972 142368 99024 142374
rect 98972 142310 99024 142316
rect 98144 142300 98196 142306
rect 98144 142242 98196 142248
rect 97868 141348 97920 141354
rect 97868 141290 97920 141296
rect 98156 138566 98184 142242
rect 100088 141694 100116 144892
rect 101206 144878 101496 144906
rect 101468 142442 101496 144878
rect 102296 142617 102324 144892
rect 102282 142608 102338 142617
rect 102282 142543 102338 142552
rect 102296 142510 102324 142543
rect 102284 142504 102336 142510
rect 102284 142446 102336 142452
rect 101456 142436 101508 142442
rect 101456 142378 101508 142384
rect 100076 141688 100128 141694
rect 100076 141630 100128 141636
rect 100626 139072 100682 139081
rect 100626 139007 100682 139016
rect 100534 138664 100590 138673
rect 100534 138599 100590 138608
rect 98144 138560 98196 138566
rect 98144 138502 98196 138508
rect 97224 138492 97276 138498
rect 97224 138434 97276 138440
rect 63458 138392 63514 138401
rect 63458 138327 63514 138336
rect 66310 138256 66366 138265
rect 66310 138191 66366 138200
rect 66324 137206 66352 138191
rect 100074 137848 100130 137857
rect 100074 137783 100130 137792
rect 66402 137712 66458 137721
rect 66402 137647 66458 137656
rect 66416 137274 66444 137647
rect 100088 137478 100116 137783
rect 100076 137472 100128 137478
rect 100076 137414 100128 137420
rect 99706 137304 99762 137313
rect 66404 137268 66456 137274
rect 99706 137239 99708 137248
rect 66404 137210 66456 137216
rect 99760 137239 99762 137248
rect 99708 137210 99760 137216
rect 66312 137200 66364 137206
rect 66312 137142 66364 137148
rect 100548 136798 100576 138599
rect 100640 137070 100668 139007
rect 101468 137206 101496 142378
rect 102284 142368 102336 142374
rect 102284 142310 102336 142316
rect 102296 140985 102324 142310
rect 105240 141778 105268 147167
rect 105208 141750 105268 141778
rect 105424 141778 105452 148391
rect 105870 146008 105926 146017
rect 105870 145943 105926 145952
rect 105884 145502 105912 145943
rect 105872 145496 105924 145502
rect 105872 145438 105924 145444
rect 105976 141778 106004 149615
rect 106422 144920 106478 144929
rect 106422 144855 106478 144864
rect 106436 144210 106464 144855
rect 106424 144204 106476 144210
rect 106424 144146 106476 144152
rect 106528 144142 106556 152494
rect 106606 151040 106662 151049
rect 106606 150975 106662 150984
rect 106516 144136 106568 144142
rect 106516 144078 106568 144084
rect 106620 141778 106648 150975
rect 107172 148329 107200 155706
rect 107264 150641 107292 156930
rect 107724 155401 107752 159242
rect 107816 157713 107844 160602
rect 108552 160025 108580 162098
rect 108538 160016 108594 160025
rect 108538 159951 108594 159960
rect 107896 158212 107948 158218
rect 107896 158154 107948 158160
rect 107802 157704 107858 157713
rect 107802 157639 107858 157648
rect 107710 155392 107766 155401
rect 107710 155327 107766 155336
rect 107908 152953 107936 158154
rect 107988 153860 108040 153866
rect 107988 153802 108040 153808
rect 107894 152944 107950 152953
rect 107894 152879 107950 152888
rect 107250 150632 107306 150641
rect 107250 150567 107306 150576
rect 107158 148320 107214 148329
rect 107158 148255 107214 148264
rect 107160 144136 107212 144142
rect 107160 144078 107212 144084
rect 107172 141778 107200 144078
rect 108000 142050 108028 153802
rect 108540 153792 108592 153798
rect 108540 153734 108592 153740
rect 108552 146017 108580 153734
rect 108538 146008 108594 146017
rect 108538 145943 108594 145952
rect 109276 145428 109328 145434
rect 109276 145370 109328 145376
rect 108356 144204 108408 144210
rect 108356 144146 108408 144152
rect 108000 142022 108074 142050
rect 105424 141750 105760 141778
rect 105976 141750 106312 141778
rect 106620 141750 106956 141778
rect 107172 141750 107508 141778
rect 108046 141764 108074 142022
rect 108368 141778 108396 144146
rect 109288 141778 109316 145370
rect 110426 142028 110478 142034
rect 110426 141970 110478 141976
rect 109782 141960 109834 141966
rect 109782 141902 109834 141908
rect 108368 141750 108704 141778
rect 109256 141750 109316 141778
rect 109794 141764 109822 141902
rect 110438 141764 110466 141970
rect 111128 141966 111156 144892
rect 111496 142034 111524 144892
rect 111588 144878 111878 144906
rect 111956 144878 112338 144906
rect 112416 144878 112706 144906
rect 111484 142028 111536 142034
rect 111484 141970 111536 141976
rect 111116 141960 111168 141966
rect 111588 141914 111616 144878
rect 111116 141902 111168 141908
rect 111404 141886 111616 141914
rect 111404 141778 111432 141886
rect 111956 141778 111984 144878
rect 112416 141778 112444 144878
rect 113060 141778 113088 144892
rect 113520 142034 113548 144892
rect 113902 144878 114008 144906
rect 113278 142028 113330 142034
rect 113278 141970 113330 141976
rect 113508 142028 113560 142034
rect 113508 141970 113560 141976
rect 111004 141750 111432 141778
rect 111556 141750 111984 141778
rect 112200 141750 112444 141778
rect 112752 141750 113088 141778
rect 113290 141764 113318 141970
rect 103480 141688 103532 141694
rect 113980 141642 114008 144878
rect 114256 141778 114284 144892
rect 114716 141778 114744 144892
rect 115098 144878 115388 144906
rect 115466 144878 115848 144906
rect 115926 144878 116216 144906
rect 115360 141778 115388 144878
rect 115820 141778 115848 144878
rect 116188 141914 116216 144878
rect 116280 142034 116308 144892
rect 116268 142028 116320 142034
rect 116268 141970 116320 141976
rect 116648 141966 116676 144892
rect 117108 142170 117136 144892
rect 117476 142714 117504 144892
rect 117464 142708 117516 142714
rect 117464 142650 117516 142656
rect 117096 142164 117148 142170
rect 117096 142106 117148 142112
rect 117844 142034 117872 144892
rect 118304 142646 118332 144892
rect 118686 144878 118976 144906
rect 118948 144142 118976 144878
rect 118936 144136 118988 144142
rect 118936 144078 118988 144084
rect 118844 142708 118896 142714
rect 118844 142650 118896 142656
rect 118292 142640 118344 142646
rect 118292 142582 118344 142588
rect 118200 142164 118252 142170
rect 118200 142106 118252 142112
rect 117418 142028 117470 142034
rect 117418 141970 117470 141976
rect 117832 142028 117884 142034
rect 117832 141970 117884 141976
rect 116636 141960 116688 141966
rect 116188 141886 116400 141914
rect 116636 141902 116688 141908
rect 116372 141778 116400 141886
rect 114256 141750 114500 141778
rect 114716 141750 115052 141778
rect 115360 141750 115696 141778
rect 115820 141750 116248 141778
rect 116372 141750 116800 141778
rect 117430 141764 117458 141970
rect 117970 141960 118022 141966
rect 117970 141902 118022 141908
rect 117982 141764 118010 141902
rect 118212 141778 118240 142106
rect 118856 141778 118884 142650
rect 119132 141966 119160 144892
rect 119500 142374 119528 144892
rect 119882 144878 120264 144906
rect 120342 144878 120540 144906
rect 120236 144226 120264 144878
rect 120236 144210 120356 144226
rect 120236 144204 120368 144210
rect 120236 144198 120316 144204
rect 120316 144146 120368 144152
rect 119948 142640 120000 142646
rect 119948 142582 120000 142588
rect 119488 142368 119540 142374
rect 119488 142310 119540 142316
rect 119718 142028 119770 142034
rect 119718 141970 119770 141976
rect 119120 141960 119172 141966
rect 119120 141902 119172 141908
rect 118212 141750 118548 141778
rect 118856 141750 119192 141778
rect 119730 141764 119758 141970
rect 119960 141778 119988 142582
rect 120512 142034 120540 144878
rect 120592 144136 120644 144142
rect 120592 144078 120644 144084
rect 120500 142028 120552 142034
rect 120500 141970 120552 141976
rect 120604 141778 120632 144078
rect 120696 142714 120724 144892
rect 120684 142708 120736 142714
rect 120684 142650 120736 142656
rect 121064 142578 121092 144892
rect 121052 142572 121104 142578
rect 121052 142514 121104 142520
rect 121524 142238 121552 144892
rect 121696 142368 121748 142374
rect 121696 142310 121748 142316
rect 121512 142232 121564 142238
rect 121512 142174 121564 142180
rect 121466 141960 121518 141966
rect 121466 141902 121518 141908
rect 119960 141750 120296 141778
rect 120604 141750 120940 141778
rect 121478 141764 121506 141902
rect 121708 141778 121736 142310
rect 121892 141966 121920 144892
rect 121880 141960 121932 141966
rect 121880 141902 121932 141908
rect 121708 141750 122044 141778
rect 122260 141762 122288 144892
rect 122734 144878 122932 144906
rect 122340 144204 122392 144210
rect 122340 144146 122392 144152
rect 122352 141778 122380 144146
rect 122904 141830 122932 144878
rect 123088 142170 123116 144892
rect 123470 144878 123760 144906
rect 123444 142708 123496 142714
rect 123444 142650 123496 142656
rect 123076 142164 123128 142170
rect 123076 142106 123128 142112
rect 123214 142028 123266 142034
rect 123214 141970 123266 141976
rect 122892 141824 122944 141830
rect 122248 141756 122300 141762
rect 122352 141750 122688 141778
rect 122892 141766 122944 141772
rect 123226 141764 123254 141970
rect 123456 141778 123484 142650
rect 123732 142306 123760 144878
rect 123916 142374 123944 144892
rect 123904 142368 123956 142374
rect 123904 142310 123956 142316
rect 123720 142300 123772 142306
rect 123720 142242 123772 142248
rect 124284 142034 124312 144892
rect 124652 142578 124680 144892
rect 125112 142714 125140 144892
rect 125100 142708 125152 142714
rect 125100 142650 125152 142656
rect 125480 142646 125508 144892
rect 125848 144278 125876 144892
rect 125836 144272 125888 144278
rect 125836 144214 125888 144220
rect 126308 144142 126336 144892
rect 126676 144210 126704 144892
rect 131448 144272 131500 144278
rect 131448 144214 131500 144220
rect 126664 144204 126716 144210
rect 126664 144146 126716 144152
rect 126296 144136 126348 144142
rect 126296 144078 126348 144084
rect 129884 142708 129936 142714
rect 129884 142650 129936 142656
rect 125468 142640 125520 142646
rect 125468 142582 125520 142588
rect 124456 142572 124508 142578
rect 124456 142514 124508 142520
rect 124640 142572 124692 142578
rect 124640 142514 124692 142520
rect 129332 142572 129384 142578
rect 129332 142514 129384 142520
rect 124272 142028 124324 142034
rect 124272 141970 124324 141976
rect 124468 141778 124496 142514
rect 128136 142368 128188 142374
rect 128136 142310 128188 142316
rect 127584 142300 127636 142306
rect 127584 142242 127636 142248
rect 124640 142232 124692 142238
rect 124640 142174 124692 142180
rect 123456 141750 123792 141778
rect 124436 141750 124496 141778
rect 124652 141778 124680 142174
rect 126940 142164 126992 142170
rect 126940 142106 126992 142112
rect 125514 141960 125566 141966
rect 125514 141902 125566 141908
rect 124652 141750 124988 141778
rect 125526 141764 125554 141902
rect 126388 141824 126440 141830
rect 125848 141762 126184 141778
rect 126952 141778 126980 142106
rect 127596 141778 127624 142242
rect 128148 141778 128176 142310
rect 129010 142028 129062 142034
rect 129010 141970 129062 141976
rect 126440 141772 126736 141778
rect 126388 141766 126736 141772
rect 125836 141756 126184 141762
rect 122248 141698 122300 141704
rect 125888 141750 126184 141756
rect 126400 141750 126736 141766
rect 126952 141750 127288 141778
rect 127596 141750 127932 141778
rect 128148 141750 128484 141778
rect 129022 141764 129050 141970
rect 129344 141778 129372 142514
rect 129896 141778 129924 142650
rect 130436 142640 130488 142646
rect 130436 142582 130488 142588
rect 130448 141778 130476 142582
rect 131460 141778 131488 144214
rect 131632 144136 131684 144142
rect 131632 144078 131684 144084
rect 129344 141750 129680 141778
rect 129896 141750 130232 141778
rect 130448 141750 130784 141778
rect 131428 141750 131488 141778
rect 131644 141778 131672 144078
rect 131644 141750 131980 141778
rect 125836 141698 125888 141704
rect 132104 141694 132132 186850
rect 132196 185457 132224 187854
rect 132644 186976 132696 186982
rect 132644 186918 132696 186924
rect 144880 186976 144932 186982
rect 144880 186918 144932 186924
rect 132182 185448 132238 185457
rect 132182 185383 132238 185392
rect 132366 151584 132422 151593
rect 132366 151519 132422 151528
rect 132184 144204 132236 144210
rect 132184 144146 132236 144152
rect 132196 141778 132224 144146
rect 132380 141898 132408 151519
rect 132368 141892 132420 141898
rect 132368 141834 132420 141840
rect 132656 141778 132684 186918
rect 144892 184740 144920 186918
rect 164844 186908 164896 186914
rect 164844 186850 164896 186856
rect 164856 184740 164884 186850
rect 176908 175665 176936 187854
rect 177080 184256 177132 184262
rect 177080 184198 177132 184204
rect 176988 182488 177040 182494
rect 176988 182430 177040 182436
rect 177000 181785 177028 182430
rect 176986 181776 177042 181785
rect 176986 181711 177042 181720
rect 177092 180561 177120 184198
rect 177078 180552 177134 180561
rect 177078 180487 177134 180496
rect 177276 180402 177304 187990
rect 177724 185004 177776 185010
rect 177724 184946 177776 184952
rect 177736 184233 177764 184946
rect 177722 184224 177778 184233
rect 177632 184188 177684 184194
rect 177722 184159 177778 184168
rect 177632 184130 177684 184136
rect 177540 184120 177592 184126
rect 177540 184062 177592 184068
rect 177448 184052 177500 184058
rect 177448 183994 177500 184000
rect 177460 183009 177488 183994
rect 177446 183000 177502 183009
rect 177446 182935 177502 182944
rect 177000 180374 177304 180402
rect 177000 176889 177028 180374
rect 177552 178113 177580 184062
rect 177644 179337 177672 184130
rect 178288 184126 178316 187868
rect 178840 184194 178868 187868
rect 179392 184262 179420 187868
rect 179380 184256 179432 184262
rect 179380 184198 179432 184204
rect 178828 184188 178880 184194
rect 178828 184130 178880 184136
rect 178276 184120 178328 184126
rect 178276 184062 178328 184068
rect 180036 182494 180064 187868
rect 180588 184126 180616 187868
rect 181140 185010 181168 187868
rect 181692 185010 181720 187868
rect 181128 185004 181180 185010
rect 181128 184946 181180 184952
rect 181680 185004 181732 185010
rect 181680 184946 181732 184952
rect 182244 184942 182272 187868
rect 182888 185486 182916 187868
rect 183454 187854 183744 187882
rect 184006 187854 184480 187882
rect 184558 187854 184848 187882
rect 185110 187854 185308 187882
rect 182876 185480 182928 185486
rect 182876 185422 182928 185428
rect 183612 185480 183664 185486
rect 183612 185422 183664 185428
rect 183106 185004 183158 185010
rect 183106 184946 183158 184952
rect 182232 184936 182284 184942
rect 182232 184878 182284 184884
rect 183118 184740 183146 184946
rect 183474 184936 183526 184942
rect 183474 184878 183526 184884
rect 183486 184740 183514 184878
rect 183624 184754 183652 185422
rect 183716 184890 183744 187854
rect 183716 184862 184020 184890
rect 183992 184754 184020 184862
rect 184452 184754 184480 187854
rect 184820 184754 184848 187854
rect 185280 184754 185308 187854
rect 185740 184754 185768 187868
rect 186200 187854 186306 187882
rect 183624 184726 183868 184754
rect 183992 184726 184328 184754
rect 184452 184726 184696 184754
rect 184820 184726 185064 184754
rect 185280 184726 185524 184754
rect 185740 184726 185892 184754
rect 186200 184618 186228 187854
rect 186844 184754 186872 187868
rect 187212 187854 187410 187882
rect 187672 187854 187962 187882
rect 188132 187854 188606 187882
rect 188684 187854 189158 187882
rect 189236 187854 189710 187882
rect 187212 184754 187240 187854
rect 187672 184754 187700 187854
rect 188132 184754 188160 187854
rect 188684 184890 188712 187854
rect 189236 185298 189264 187854
rect 190144 185480 190196 185486
rect 190144 185422 190196 185428
rect 188500 184862 188712 184890
rect 188960 185270 189264 185298
rect 188500 184754 188528 184862
rect 188960 184754 188988 185270
rect 189086 185004 189138 185010
rect 189086 184946 189138 184952
rect 186720 184726 186872 184754
rect 187088 184726 187240 184754
rect 187456 184726 187700 184754
rect 187916 184726 188160 184754
rect 188284 184726 188528 184754
rect 188652 184726 188988 184754
rect 189098 184740 189126 184946
rect 189454 184936 189506 184942
rect 189454 184878 189506 184884
rect 189466 184740 189494 184878
rect 190156 184754 190184 185422
rect 190248 185010 190276 187868
rect 190604 185412 190656 185418
rect 190604 185354 190656 185360
rect 190420 185140 190472 185146
rect 190420 185082 190472 185088
rect 190236 185004 190288 185010
rect 190236 184946 190288 184952
rect 190432 184754 190460 185082
rect 189848 184726 190184 184754
rect 190308 184726 190460 184754
rect 190616 184754 190644 185354
rect 190800 184942 190828 187868
rect 191444 185486 191472 187868
rect 191432 185480 191484 185486
rect 191432 185422 191484 185428
rect 191996 185146 192024 187868
rect 192548 185418 192576 187868
rect 192536 185412 192588 185418
rect 192536 185354 192588 185360
rect 192904 185412 192956 185418
rect 192904 185354 192956 185360
rect 192536 185276 192588 185282
rect 192536 185218 192588 185224
rect 191984 185140 192036 185146
rect 191984 185082 192036 185088
rect 191110 185004 191162 185010
rect 191110 184946 191162 184952
rect 190788 184936 190840 184942
rect 190788 184878 190840 184884
rect 190616 184726 190676 184754
rect 191122 184740 191150 184946
rect 191478 184936 191530 184942
rect 191478 184878 191530 184884
rect 191490 184740 191518 184878
rect 191984 184868 192036 184874
rect 191984 184810 192036 184816
rect 191996 184618 192024 184810
rect 192548 184754 192576 185218
rect 192916 184754 192944 185354
rect 193100 185010 193128 187868
rect 193364 185344 193416 185350
rect 193364 185286 193416 185292
rect 193088 185004 193140 185010
rect 193088 184946 193140 184952
rect 193376 184754 193404 185286
rect 193502 185004 193554 185010
rect 193502 184946 193554 184952
rect 192332 184726 192576 184754
rect 192700 184726 192944 184754
rect 193068 184726 193404 184754
rect 193514 184740 193542 184946
rect 193652 184942 193680 187868
rect 194020 187854 194310 187882
rect 193640 184936 193692 184942
rect 193640 184878 193692 184884
rect 194020 184874 194048 187854
rect 194848 185282 194876 187868
rect 195400 185418 195428 187868
rect 195388 185412 195440 185418
rect 195388 185354 195440 185360
rect 195756 185412 195808 185418
rect 195756 185354 195808 185360
rect 194836 185276 194888 185282
rect 194836 185218 194888 185224
rect 195296 185276 195348 185282
rect 195296 185218 195348 185224
rect 194100 185208 194152 185214
rect 194100 185150 194152 185156
rect 194008 184868 194060 184874
rect 194008 184810 194060 184816
rect 194112 184754 194140 185150
rect 194560 185140 194612 185146
rect 194560 185082 194612 185088
rect 194572 184754 194600 185082
rect 194652 185072 194704 185078
rect 194652 185014 194704 185020
rect 193896 184726 194140 184754
rect 194264 184726 194600 184754
rect 186200 184590 186260 184618
rect 191872 184590 192024 184618
rect 194664 184618 194692 185014
rect 195308 184754 195336 185218
rect 195768 184754 195796 185354
rect 195952 185350 195980 187868
rect 195940 185344 195992 185350
rect 195940 185286 195992 185292
rect 196124 185344 196176 185350
rect 196124 185286 196176 185292
rect 196136 184754 196164 185286
rect 196504 185010 196532 187868
rect 197148 185214 197176 187868
rect 197320 185480 197372 185486
rect 197320 185422 197372 185428
rect 197136 185208 197188 185214
rect 197136 185150 197188 185156
rect 196492 185004 196544 185010
rect 196492 184946 196544 184952
rect 196630 184936 196682 184942
rect 196630 184878 196682 184884
rect 196492 184868 196544 184874
rect 196492 184810 196544 184816
rect 196504 184754 196532 184810
rect 195092 184726 195336 184754
rect 195460 184726 195796 184754
rect 195920 184726 196164 184754
rect 196288 184726 196532 184754
rect 196642 184740 196670 184878
rect 197332 184754 197360 185422
rect 197700 185146 197728 187868
rect 197688 185140 197740 185146
rect 197688 185082 197740 185088
rect 198252 185078 198280 187868
rect 198804 185282 198832 187868
rect 199356 185418 199384 187868
rect 199344 185412 199396 185418
rect 199344 185354 199396 185360
rect 200000 185350 200028 187868
rect 199988 185344 200040 185350
rect 199988 185286 200040 185292
rect 198792 185276 198844 185282
rect 198792 185218 198844 185224
rect 198240 185072 198292 185078
rect 197456 185040 197512 185049
rect 198240 185014 198292 185020
rect 197456 184975 197512 184984
rect 197826 185004 197878 185010
rect 197116 184726 197360 184754
rect 197470 184740 197498 184975
rect 197826 184946 197878 184952
rect 197838 184740 197866 184946
rect 200552 184874 200580 187868
rect 201104 184942 201132 187868
rect 201656 185486 201684 187868
rect 201644 185480 201696 185486
rect 201644 185422 201696 185428
rect 202208 185049 202236 187868
rect 202194 185040 202250 185049
rect 202852 185010 202880 187868
rect 202194 184975 202250 184984
rect 202840 185004 202892 185010
rect 202840 184946 202892 184952
rect 201092 184936 201144 184942
rect 201092 184878 201144 184884
rect 200540 184868 200592 184874
rect 200540 184810 200592 184816
rect 194664 184590 194724 184618
rect 198514 184496 198570 184505
rect 198312 184454 198514 184482
rect 198882 184496 198938 184505
rect 198680 184454 198882 184482
rect 198514 184431 198570 184440
rect 198882 184431 198938 184440
rect 203404 184369 203432 187868
rect 203956 184505 203984 187868
rect 203942 184496 203998 184505
rect 203942 184431 203998 184440
rect 203390 184360 203446 184369
rect 203390 184295 203446 184304
rect 180576 184120 180628 184126
rect 180576 184062 180628 184068
rect 180298 183544 180354 183553
rect 180298 183479 180354 183488
rect 180024 182488 180076 182494
rect 180024 182430 180076 182436
rect 179746 181232 179802 181241
rect 179746 181167 179802 181176
rect 177630 179328 177686 179337
rect 177630 179263 177686 179272
rect 179760 179042 179788 181167
rect 179760 179014 179972 179042
rect 179746 178920 179802 178929
rect 179746 178855 179802 178864
rect 177538 178104 177594 178113
rect 177538 178039 177594 178048
rect 176986 176880 177042 176889
rect 176986 176815 177042 176824
rect 179654 176472 179710 176481
rect 179654 176407 179710 176416
rect 179668 175898 179696 176407
rect 177724 175892 177776 175898
rect 177724 175834 177776 175840
rect 179656 175892 179708 175898
rect 179656 175834 179708 175840
rect 176894 175656 176950 175665
rect 176894 175591 176950 175600
rect 177354 174432 177410 174441
rect 177354 174367 177356 174376
rect 177408 174367 177410 174376
rect 177356 174338 177408 174344
rect 176988 174328 177040 174334
rect 176988 174270 177040 174276
rect 177000 173217 177028 174270
rect 176986 173208 177042 173217
rect 176986 173143 177042 173152
rect 177632 173104 177684 173110
rect 177632 173046 177684 173052
rect 177540 172968 177592 172974
rect 177540 172910 177592 172916
rect 177552 172129 177580 172910
rect 177538 172120 177594 172129
rect 177538 172055 177594 172064
rect 177644 169681 177672 173046
rect 177736 170905 177764 175834
rect 179654 174160 179710 174169
rect 179654 174095 179710 174104
rect 179668 173110 179696 174095
rect 179656 173104 179708 173110
rect 179656 173046 179708 173052
rect 179760 172974 179788 178855
rect 179944 174334 179972 179014
rect 180312 174402 180340 183479
rect 204508 178249 204536 187868
rect 207268 183009 207296 192319
rect 225194 187352 225250 187361
rect 225194 187287 225250 187296
rect 207254 183000 207310 183009
rect 207254 182935 207310 182944
rect 225208 179745 225236 187287
rect 225194 179736 225250 179745
rect 225194 179671 225250 179680
rect 201090 178240 201146 178249
rect 201090 178175 201146 178184
rect 204494 178240 204550 178249
rect 204494 178175 204550 178184
rect 180300 174396 180352 174402
rect 180300 174338 180352 174344
rect 179932 174328 179984 174334
rect 179932 174270 179984 174276
rect 179748 172968 179800 172974
rect 179748 172910 179800 172916
rect 179654 171848 179710 171857
rect 179654 171783 179710 171792
rect 179668 171750 179696 171783
rect 178092 171744 178144 171750
rect 178092 171686 178144 171692
rect 179656 171744 179708 171750
rect 179656 171686 179708 171692
rect 177722 170896 177778 170905
rect 177722 170831 177778 170840
rect 177630 169672 177686 169681
rect 177630 169607 177686 169616
rect 177540 168956 177592 168962
rect 177540 168898 177592 168904
rect 177552 167233 177580 168898
rect 178104 168457 178132 171686
rect 179654 169400 179710 169409
rect 179654 169335 179710 169344
rect 179668 168962 179696 169335
rect 179656 168956 179708 168962
rect 179656 168898 179708 168904
rect 178090 168448 178146 168457
rect 178090 168383 178146 168392
rect 177538 167224 177594 167233
rect 177538 167159 177594 167168
rect 179562 167088 179618 167097
rect 179562 167023 179618 167032
rect 179576 166174 179604 167023
rect 201104 166174 201132 178175
rect 223538 169264 223594 169273
rect 223538 169199 223594 169208
rect 223552 169166 223580 169199
rect 222804 169160 222856 169166
rect 222724 169120 222804 169148
rect 177540 166168 177592 166174
rect 177540 166110 177592 166116
rect 179564 166168 179616 166174
rect 179564 166110 179616 166116
rect 201092 166168 201144 166174
rect 201092 166110 201144 166116
rect 204496 166168 204548 166174
rect 222724 166122 222752 169120
rect 222804 169102 222856 169108
rect 223540 169160 223592 169166
rect 223540 169102 223592 169108
rect 204496 166110 204548 166116
rect 177552 166009 177580 166110
rect 177538 166000 177594 166009
rect 177538 165935 177594 165944
rect 204508 164921 204536 166110
rect 222632 166094 222752 166122
rect 200998 164912 201054 164921
rect 200998 164847 201054 164856
rect 204494 164912 204550 164921
rect 204494 164847 204550 164856
rect 177722 163552 177778 163561
rect 177722 163487 177724 163496
rect 177776 163487 177778 163496
rect 179564 163516 179616 163522
rect 177724 163458 177776 163464
rect 179564 163458 179616 163464
rect 179576 162473 179604 163458
rect 179562 162464 179618 162473
rect 179562 162399 179618 162408
rect 176986 162328 177042 162337
rect 176986 162263 177042 162272
rect 177000 162094 177028 162263
rect 176988 162088 177040 162094
rect 176988 162030 177040 162036
rect 179656 162088 179708 162094
rect 179656 162030 179708 162036
rect 176986 161104 177042 161113
rect 176986 161039 177042 161048
rect 177000 160870 177028 161039
rect 176988 160864 177040 160870
rect 176988 160806 177040 160812
rect 179564 160864 179616 160870
rect 179564 160806 179616 160812
rect 177538 159880 177594 159889
rect 177538 159815 177594 159824
rect 177552 159306 177580 159815
rect 177540 159300 177592 159306
rect 177540 159242 177592 159248
rect 179472 159300 179524 159306
rect 179472 159242 179524 159248
rect 177354 158792 177410 158801
rect 177354 158727 177410 158736
rect 177368 157946 177396 158727
rect 177356 157940 177408 157946
rect 177356 157882 177408 157888
rect 177538 157568 177594 157577
rect 177538 157503 177594 157512
rect 177552 156518 177580 157503
rect 177540 156512 177592 156518
rect 177540 156454 177592 156460
rect 177538 156344 177594 156353
rect 177538 156279 177594 156288
rect 177552 155158 177580 156279
rect 179484 155401 179512 159242
rect 179576 157713 179604 160806
rect 179668 160025 179696 162030
rect 179654 160016 179710 160025
rect 179654 159951 179710 159960
rect 179656 157940 179708 157946
rect 179656 157882 179708 157888
rect 179562 157704 179618 157713
rect 179562 157639 179618 157648
rect 179470 155392 179526 155401
rect 179470 155327 179526 155336
rect 177540 155152 177592 155158
rect 177354 155120 177410 155129
rect 177540 155094 177592 155100
rect 177354 155055 177410 155064
rect 177368 153866 177396 155055
rect 178182 153896 178238 153905
rect 177356 153860 177408 153866
rect 178182 153831 178238 153840
rect 177356 153802 177408 153808
rect 178196 153798 178224 153831
rect 178184 153792 178236 153798
rect 178184 153734 178236 153740
rect 179668 152953 179696 157882
rect 180484 156512 180536 156518
rect 180484 156454 180536 156460
rect 180392 155152 180444 155158
rect 180392 155094 180444 155100
rect 180300 153860 180352 153866
rect 180300 153802 180352 153808
rect 179748 153792 179800 153798
rect 179748 153734 179800 153740
rect 179654 152944 179710 152953
rect 179654 152879 179710 152888
rect 178274 152672 178330 152681
rect 178274 152607 178330 152616
rect 177722 149000 177778 149009
rect 177722 148935 177778 148944
rect 177170 147776 177226 147785
rect 177170 147711 177226 147720
rect 134484 142572 134536 142578
rect 134484 142514 134536 142520
rect 134496 142073 134524 142514
rect 134482 142064 134538 142073
rect 134482 141999 134538 142008
rect 132196 141750 132532 141778
rect 132656 141750 132776 141778
rect 103480 141630 103532 141636
rect 103492 141529 103520 141630
rect 113948 141614 114008 141642
rect 132092 141688 132144 141694
rect 132092 141630 132144 141636
rect 132644 141688 132696 141694
rect 132644 141630 132696 141636
rect 103478 141520 103534 141529
rect 103478 141455 103534 141464
rect 102376 141212 102428 141218
rect 102376 141154 102428 141160
rect 102282 140976 102338 140985
rect 102282 140911 102338 140920
rect 102388 140441 102416 141154
rect 102374 140432 102430 140441
rect 102374 140367 102430 140376
rect 102376 139920 102428 139926
rect 102376 139862 102428 139868
rect 102388 139761 102416 139862
rect 102468 139852 102520 139858
rect 102468 139794 102520 139800
rect 102374 139752 102430 139761
rect 102374 139687 102430 139696
rect 102480 139217 102508 139794
rect 102560 139784 102612 139790
rect 102560 139726 102612 139732
rect 102466 139208 102522 139217
rect 102466 139143 102522 139152
rect 102572 138673 102600 139726
rect 102558 138664 102614 138673
rect 102558 138599 102614 138608
rect 102376 138560 102428 138566
rect 102376 138502 102428 138508
rect 102388 137993 102416 138502
rect 102468 138492 102520 138498
rect 102468 138434 102520 138440
rect 102374 137984 102430 137993
rect 102374 137919 102430 137928
rect 102284 137472 102336 137478
rect 102480 137449 102508 138434
rect 132656 137478 132684 141630
rect 132644 137472 132696 137478
rect 102284 137414 102336 137420
rect 102466 137440 102522 137449
rect 102192 137268 102244 137274
rect 102192 137210 102244 137216
rect 101456 137200 101508 137206
rect 101456 137142 101508 137148
rect 101916 137200 101968 137206
rect 101916 137142 101968 137148
rect 100628 137064 100680 137070
rect 100628 137006 100680 137012
rect 100536 136792 100588 136798
rect 65022 136760 65078 136769
rect 100536 136734 100588 136740
rect 65022 136695 65078 136704
rect 62906 136624 62962 136633
rect 62906 136559 62962 136568
rect 63000 135908 63052 135914
rect 63000 135850 63052 135856
rect 62908 135840 62960 135846
rect 62908 135782 62960 135788
rect 62816 135704 62868 135710
rect 62722 135672 62778 135681
rect 62816 135646 62868 135652
rect 62722 135607 62778 135616
rect 62630 135400 62686 135409
rect 62630 135335 62686 135344
rect 62828 134865 62856 135646
rect 62814 134856 62870 134865
rect 62814 134791 62870 134800
rect 62724 134548 62776 134554
rect 62724 134490 62776 134496
rect 62736 132553 62764 134490
rect 62816 134480 62868 134486
rect 62816 134422 62868 134428
rect 62828 132825 62856 134422
rect 62920 134321 62948 135782
rect 62906 134312 62962 134321
rect 62906 134247 62962 134256
rect 63012 133641 63040 135850
rect 65036 135710 65064 136695
rect 100626 136624 100682 136633
rect 100626 136559 100682 136568
rect 66402 136488 66458 136497
rect 66402 136423 66458 136432
rect 65666 135944 65722 135953
rect 65666 135879 65668 135888
rect 65720 135879 65722 135888
rect 65668 135850 65720 135856
rect 66416 135846 66444 136423
rect 100640 135846 100668 136559
rect 100902 136080 100958 136089
rect 100958 136038 101036 136066
rect 100902 136015 100958 136024
rect 100902 135944 100958 135953
rect 100902 135879 100904 135888
rect 100956 135879 100958 135888
rect 100904 135850 100956 135856
rect 66404 135840 66456 135846
rect 66404 135782 66456 135788
rect 100628 135840 100680 135846
rect 100628 135782 100680 135788
rect 65024 135704 65076 135710
rect 65024 135646 65076 135652
rect 65850 135264 65906 135273
rect 65850 135199 65906 135208
rect 65864 134486 65892 135199
rect 99890 134856 99946 134865
rect 99890 134791 99946 134800
rect 66218 134720 66274 134729
rect 99904 134690 99932 134791
rect 100902 134720 100958 134729
rect 66218 134655 66274 134664
rect 99892 134684 99944 134690
rect 66232 134554 66260 134655
rect 100902 134655 100958 134664
rect 99892 134626 99944 134632
rect 100916 134622 100944 134655
rect 100904 134616 100956 134622
rect 100904 134558 100956 134564
rect 66220 134548 66272 134554
rect 66220 134490 66272 134496
rect 65852 134480 65904 134486
rect 65852 134422 65904 134428
rect 101008 134418 101036 136038
rect 100996 134412 101048 134418
rect 100996 134354 101048 134360
rect 65482 134176 65538 134185
rect 65482 134111 65538 134120
rect 62998 133632 63054 133641
rect 62998 133567 63054 133576
rect 65496 133126 65524 134111
rect 100902 133632 100958 133641
rect 100902 133567 100958 133576
rect 66402 133496 66458 133505
rect 66402 133431 66458 133440
rect 63460 133120 63512 133126
rect 63460 133062 63512 133068
rect 65484 133120 65536 133126
rect 65484 133062 65536 133068
rect 62814 132816 62870 132825
rect 62814 132751 62870 132760
rect 62722 132544 62778 132553
rect 62722 132479 62778 132488
rect 63092 131760 63144 131766
rect 63092 131702 63144 131708
rect 62816 130808 62868 130814
rect 62814 130776 62816 130785
rect 62868 130776 62870 130785
rect 62814 130711 62870 130720
rect 62908 130400 62960 130406
rect 62908 130342 62960 130348
rect 62724 130332 62776 130338
rect 62724 130274 62776 130280
rect 62632 129040 62684 129046
rect 62632 128982 62684 128988
rect 62644 127249 62672 128982
rect 62736 128745 62764 130274
rect 62816 128972 62868 128978
rect 62816 128914 62868 128920
rect 62722 128736 62778 128745
rect 62722 128671 62778 128680
rect 62828 127521 62856 128914
rect 62920 128473 62948 130342
rect 63104 129561 63132 131702
rect 63472 131601 63500 133062
rect 66416 133058 66444 133431
rect 100916 133262 100944 133567
rect 100904 133256 100956 133262
rect 100258 133224 100314 133233
rect 100904 133198 100956 133204
rect 100258 133159 100260 133168
rect 100312 133159 100314 133168
rect 100260 133130 100312 133136
rect 63552 133052 63604 133058
rect 63552 132994 63604 133000
rect 66404 133052 66456 133058
rect 66404 132994 66456 133000
rect 63458 131592 63514 131601
rect 63458 131527 63514 131536
rect 63564 131329 63592 132994
rect 65022 132544 65078 132553
rect 65022 132479 65078 132488
rect 63644 131692 63696 131698
rect 63644 131634 63696 131640
rect 63550 131320 63606 131329
rect 63550 131255 63606 131264
rect 63656 130241 63684 131634
rect 65036 130814 65064 132479
rect 100258 132408 100314 132417
rect 100258 132343 100314 132352
rect 66402 132272 66458 132281
rect 66402 132207 66458 132216
rect 65668 131760 65720 131766
rect 65666 131728 65668 131737
rect 65720 131728 65722 131737
rect 66416 131698 66444 132207
rect 100272 131698 100300 132343
rect 100902 132000 100958 132009
rect 100958 131958 101036 131986
rect 100902 131935 100958 131944
rect 100904 131760 100956 131766
rect 100902 131728 100904 131737
rect 100956 131728 100958 131737
rect 65666 131663 65722 131672
rect 66404 131692 66456 131698
rect 66404 131634 66456 131640
rect 100260 131692 100312 131698
rect 100902 131663 100958 131672
rect 100260 131634 100312 131640
rect 66310 131184 66366 131193
rect 66310 131119 66366 131128
rect 65024 130808 65076 130814
rect 65024 130750 65076 130756
rect 66324 130338 66352 131119
rect 100258 130640 100314 130649
rect 100258 130575 100314 130584
rect 66402 130504 66458 130513
rect 100272 130474 100300 130575
rect 100902 130504 100958 130513
rect 66402 130439 66458 130448
rect 100260 130468 100312 130474
rect 66416 130406 66444 130439
rect 100902 130439 100958 130448
rect 100260 130410 100312 130416
rect 100916 130406 100944 130439
rect 66404 130400 66456 130406
rect 66404 130342 66456 130348
rect 100904 130400 100956 130406
rect 100904 130342 100956 130348
rect 66312 130332 66364 130338
rect 66312 130274 66364 130280
rect 101008 130270 101036 131958
rect 101928 131465 101956 137142
rect 102008 135908 102060 135914
rect 102008 135850 102060 135856
rect 102020 133369 102048 135850
rect 102204 135137 102232 137210
rect 102296 135681 102324 137414
rect 132644 137414 132696 137420
rect 102466 137375 102522 137384
rect 132644 137200 132696 137206
rect 132644 137142 132696 137148
rect 102376 137064 102428 137070
rect 102376 137006 102428 137012
rect 102388 136905 102416 137006
rect 102374 136896 102430 136905
rect 102374 136831 102430 136840
rect 102652 136792 102704 136798
rect 102652 136734 102704 136740
rect 102664 136361 102692 136734
rect 102650 136352 102706 136361
rect 102650 136287 102706 136296
rect 102376 135772 102428 135778
rect 102376 135714 102428 135720
rect 102282 135672 102338 135681
rect 102282 135607 102338 135616
rect 102190 135128 102246 135137
rect 102190 135063 102246 135072
rect 102284 134684 102336 134690
rect 102284 134626 102336 134632
rect 102100 134616 102152 134622
rect 102100 134558 102152 134564
rect 102006 133360 102062 133369
rect 102006 133295 102062 133304
rect 102008 133256 102060 133262
rect 102008 133198 102060 133204
rect 102020 131601 102048 133198
rect 102112 132281 102140 134558
rect 102192 133188 102244 133194
rect 102192 133130 102244 133136
rect 102098 132272 102154 132281
rect 102098 132207 102154 132216
rect 102100 131760 102152 131766
rect 102100 131702 102152 131708
rect 102006 131592 102062 131601
rect 102006 131527 102062 131536
rect 101914 131456 101970 131465
rect 101914 131391 101970 131400
rect 102008 130400 102060 130406
rect 102008 130342 102060 130348
rect 100996 130264 101048 130270
rect 63642 130232 63698 130241
rect 100996 130206 101048 130212
rect 63642 130167 63698 130176
rect 65482 129960 65538 129969
rect 65482 129895 65538 129904
rect 63090 129552 63146 129561
rect 63090 129487 63146 129496
rect 65496 128978 65524 129895
rect 100258 129416 100314 129425
rect 100258 129351 100314 129360
rect 66402 129280 66458 129289
rect 66402 129215 66458 129224
rect 66416 129046 66444 129215
rect 100272 129046 100300 129351
rect 66404 129040 66456 129046
rect 66404 128982 66456 128988
rect 100260 129040 100312 129046
rect 100260 128982 100312 128988
rect 100902 129008 100958 129017
rect 65484 128972 65536 128978
rect 100902 128943 100904 128952
rect 65484 128914 65536 128920
rect 100956 128943 100958 128952
rect 100904 128914 100956 128920
rect 62906 128464 62962 128473
rect 62906 128399 62962 128408
rect 100074 128328 100130 128337
rect 100074 128263 100130 128272
rect 66402 128192 66458 128201
rect 66402 128127 66458 128136
rect 65022 127920 65078 127929
rect 65022 127855 65078 127864
rect 62908 127544 62960 127550
rect 62814 127512 62870 127521
rect 62908 127486 62960 127492
rect 62814 127447 62870 127456
rect 62630 127240 62686 127249
rect 62630 127175 62686 127184
rect 62816 126932 62868 126938
rect 62816 126874 62868 126880
rect 62828 126705 62856 126874
rect 62814 126696 62870 126705
rect 62814 126631 62870 126640
rect 62724 126252 62776 126258
rect 62724 126194 62776 126200
rect 62632 126184 62684 126190
rect 62632 126126 62684 126132
rect 62644 124393 62672 126126
rect 62736 124665 62764 126194
rect 62920 126025 62948 127486
rect 65036 126938 65064 127855
rect 66416 127550 66444 128127
rect 100088 127890 100116 128263
rect 102020 128201 102048 130342
rect 102112 129289 102140 131702
rect 102204 131057 102232 133130
rect 102296 132825 102324 134626
rect 102388 134593 102416 135714
rect 102374 134584 102430 134593
rect 102374 134519 102430 134528
rect 102376 134412 102428 134418
rect 102376 134354 102428 134360
rect 102388 133913 102416 134354
rect 102374 133904 102430 133913
rect 102374 133839 102430 133848
rect 102282 132816 102338 132825
rect 102282 132751 102338 132760
rect 102284 131692 102336 131698
rect 102284 131634 102336 131640
rect 102190 131048 102246 131057
rect 102190 130983 102246 130992
rect 102296 130785 102324 131634
rect 102282 130776 102338 130785
rect 102282 130711 102338 130720
rect 102284 130468 102336 130474
rect 102284 130410 102336 130416
rect 102098 129280 102154 129289
rect 102098 129215 102154 129224
rect 102100 129040 102152 129046
rect 102100 128982 102152 128988
rect 102006 128192 102062 128201
rect 102006 128127 102062 128136
rect 100076 127884 100128 127890
rect 100076 127826 100128 127832
rect 100810 127648 100866 127657
rect 100810 127583 100812 127592
rect 100864 127583 100866 127592
rect 102008 127612 102060 127618
rect 100812 127554 100864 127560
rect 102008 127554 102060 127560
rect 66404 127544 66456 127550
rect 66404 127486 66456 127492
rect 100534 127104 100590 127113
rect 100534 127039 100590 127048
rect 66310 126968 66366 126977
rect 65024 126932 65076 126938
rect 66310 126903 66366 126912
rect 65024 126874 65076 126880
rect 65022 126560 65078 126569
rect 65022 126495 65078 126504
rect 62906 126016 62962 126025
rect 62906 125951 62962 125960
rect 65036 125578 65064 126495
rect 66324 126258 66352 126903
rect 66402 126288 66458 126297
rect 66312 126252 66364 126258
rect 66402 126223 66458 126232
rect 66312 126194 66364 126200
rect 66416 126190 66444 126223
rect 100548 126190 100576 127039
rect 100626 126424 100682 126433
rect 100626 126359 100682 126368
rect 100640 126258 100668 126359
rect 100902 126288 100958 126297
rect 100628 126252 100680 126258
rect 100958 126246 101036 126274
rect 100902 126223 100958 126232
rect 100628 126194 100680 126200
rect 66404 126184 66456 126190
rect 66404 126126 66456 126132
rect 100536 126184 100588 126190
rect 100536 126126 100588 126132
rect 66402 125744 66458 125753
rect 66402 125679 66458 125688
rect 62816 125572 62868 125578
rect 62816 125514 62868 125520
rect 65024 125572 65076 125578
rect 65024 125514 65076 125520
rect 62828 125481 62856 125514
rect 62814 125472 62870 125481
rect 62814 125407 62870 125416
rect 65850 125200 65906 125209
rect 65850 125135 65906 125144
rect 65022 124928 65078 124937
rect 65022 124863 65078 124872
rect 62908 124824 62960 124830
rect 62908 124766 62960 124772
rect 62722 124656 62778 124665
rect 62722 124591 62778 124600
rect 62630 124384 62686 124393
rect 62630 124319 62686 124328
rect 62816 124144 62868 124150
rect 62816 124086 62868 124092
rect 62828 123713 62856 124086
rect 62814 123704 62870 123713
rect 62814 123639 62870 123648
rect 62920 123169 62948 124766
rect 65036 124150 65064 124863
rect 65864 124830 65892 125135
rect 66416 124937 66444 125679
rect 100626 125336 100682 125345
rect 100626 125271 100682 125280
rect 100640 125170 100668 125271
rect 100628 125164 100680 125170
rect 100628 125106 100680 125112
rect 66402 124928 66458 124937
rect 66402 124863 66458 124872
rect 100626 124928 100682 124937
rect 100626 124863 100628 124872
rect 100680 124863 100682 124872
rect 100628 124834 100680 124840
rect 65852 124824 65904 124830
rect 65852 124766 65904 124772
rect 101008 124762 101036 126246
rect 102020 125753 102048 127554
rect 102112 127521 102140 128982
rect 102192 128972 102244 128978
rect 102192 128914 102244 128920
rect 102098 127512 102154 127521
rect 102098 127447 102154 127456
rect 102204 126977 102232 128914
rect 102296 128745 102324 130410
rect 102376 130264 102428 130270
rect 102376 130206 102428 130212
rect 102388 129833 102416 130206
rect 102374 129824 102430 129833
rect 102374 129759 102430 129768
rect 102282 128736 102338 128745
rect 102282 128671 102338 128680
rect 102284 127884 102336 127890
rect 102284 127826 102336 127832
rect 102190 126968 102246 126977
rect 102190 126903 102246 126912
rect 102296 126433 102324 127826
rect 132656 127618 132684 137142
rect 132644 127612 132696 127618
rect 132644 127554 132696 127560
rect 132748 127414 132776 141750
rect 135128 141484 135180 141490
rect 135128 141426 135180 141432
rect 134576 141348 134628 141354
rect 134576 141290 134628 141296
rect 134588 138401 134616 141290
rect 135140 138945 135168 141426
rect 135508 141370 135536 144892
rect 135232 141342 135536 141370
rect 136612 141354 136640 144892
rect 137716 141490 137744 144892
rect 138268 144878 138834 144906
rect 139648 144878 139938 144906
rect 137704 141484 137756 141490
rect 137704 141426 137756 141432
rect 136600 141348 136652 141354
rect 135126 138936 135182 138945
rect 135126 138871 135182 138880
rect 134574 138392 134630 138401
rect 134574 138327 134630 138336
rect 135232 137721 135260 141342
rect 136600 141290 136652 141296
rect 135312 141144 135364 141150
rect 135312 141086 135364 141092
rect 135324 140985 135352 141086
rect 135310 140976 135366 140985
rect 135310 140911 135366 140920
rect 135312 140736 135364 140742
rect 135312 140678 135364 140684
rect 135324 140441 135352 140678
rect 135310 140432 135366 140441
rect 135310 140367 135366 140376
rect 135312 139852 135364 139858
rect 135312 139794 135364 139800
rect 135324 139761 135352 139794
rect 135310 139752 135366 139761
rect 135310 139687 135366 139696
rect 138268 139518 138296 144878
rect 139648 142696 139676 144878
rect 139556 142668 139676 142696
rect 139556 139858 139584 142668
rect 140832 141688 140884 141694
rect 140832 141630 140884 141636
rect 139544 139852 139596 139858
rect 139544 139794 139596 139800
rect 140844 139724 140872 141630
rect 141028 140742 141056 144892
rect 141120 144878 142146 144906
rect 141120 141150 141148 144878
rect 142672 142708 142724 142714
rect 142672 142650 142724 142656
rect 141108 141144 141160 141150
rect 141108 141086 141160 141092
rect 141016 140736 141068 140742
rect 141016 140678 141068 140684
rect 142684 139724 142712 142650
rect 143236 142578 143264 144892
rect 143224 142572 143276 142578
rect 143224 142514 143276 142520
rect 144340 141694 144368 144892
rect 145444 142714 145472 144892
rect 145432 142708 145484 142714
rect 145432 142650 145484 142656
rect 146444 142708 146496 142714
rect 146444 142650 146496 142656
rect 144328 141688 144380 141694
rect 144328 141630 144380 141636
rect 144512 141620 144564 141626
rect 144512 141562 144564 141568
rect 144524 139724 144552 141562
rect 146456 139724 146484 142650
rect 146548 141626 146576 144892
rect 147652 142714 147680 144892
rect 148296 144878 148862 144906
rect 149966 144878 150164 144906
rect 147640 142708 147692 142714
rect 147640 142650 147692 142656
rect 146536 141620 146588 141626
rect 146536 141562 146588 141568
rect 148296 139724 148324 144878
rect 150136 139724 150164 144878
rect 151056 141626 151084 144892
rect 152160 141830 152188 144892
rect 153264 141966 153292 144892
rect 154368 142714 154396 144892
rect 154356 142708 154408 142714
rect 154356 142650 154408 142656
rect 153252 141960 153304 141966
rect 153252 141902 153304 141908
rect 152148 141824 152200 141830
rect 152148 141766 152200 141772
rect 153896 141824 153948 141830
rect 153896 141766 153948 141772
rect 151044 141620 151096 141626
rect 151044 141562 151096 141568
rect 152056 141620 152108 141626
rect 152056 141562 152108 141568
rect 152068 139724 152096 141562
rect 153908 139724 153936 141766
rect 155472 141422 155500 144892
rect 155828 141960 155880 141966
rect 155828 141902 155880 141908
rect 155460 141416 155512 141422
rect 155460 141358 155512 141364
rect 155840 139724 155868 141902
rect 156576 141558 156604 144892
rect 157694 144878 157984 144906
rect 157668 142708 157720 142714
rect 157668 142650 157720 142656
rect 156564 141552 156616 141558
rect 156564 141494 156616 141500
rect 157680 139724 157708 142650
rect 157956 141626 157984 144878
rect 158784 142170 158812 144892
rect 159888 142306 159916 144892
rect 160992 142374 161020 144892
rect 160980 142368 161032 142374
rect 160980 142310 161032 142316
rect 159876 142300 159928 142306
rect 159876 142242 159928 142248
rect 158772 142164 158824 142170
rect 158772 142106 158824 142112
rect 162188 141937 162216 144892
rect 163292 142617 163320 144892
rect 163278 142608 163334 142617
rect 163278 142543 163334 142552
rect 164396 142034 164424 144892
rect 165500 142646 165528 144892
rect 166604 142714 166632 144892
rect 167248 144878 167722 144906
rect 165856 142708 165908 142714
rect 165856 142650 165908 142656
rect 166592 142708 166644 142714
rect 166592 142650 166644 142656
rect 165488 142640 165540 142646
rect 165488 142582 165540 142588
rect 165120 142164 165172 142170
rect 165120 142106 165172 142112
rect 164384 142028 164436 142034
rect 164384 141970 164436 141976
rect 162174 141928 162230 141937
rect 162174 141863 162230 141872
rect 157944 141620 157996 141626
rect 157944 141562 157996 141568
rect 163280 141620 163332 141626
rect 163280 141562 163332 141568
rect 161440 141552 161492 141558
rect 161440 141494 161492 141500
rect 159508 141416 159560 141422
rect 159508 141358 159560 141364
rect 159520 139724 159548 141358
rect 161452 139724 161480 141494
rect 163292 139724 163320 141562
rect 165132 139724 165160 142106
rect 165868 139790 165896 142650
rect 167052 142300 167104 142306
rect 167052 142242 167104 142248
rect 165856 139784 165908 139790
rect 165856 139726 165908 139732
rect 167064 139724 167092 142242
rect 167248 139858 167276 144878
rect 168812 142238 168840 144892
rect 169352 142640 169404 142646
rect 169352 142582 169404 142588
rect 168892 142368 168944 142374
rect 168892 142310 168944 142316
rect 168800 142232 168852 142238
rect 168800 142174 168852 142180
rect 167236 139852 167288 139858
rect 167236 139794 167288 139800
rect 168904 139724 168932 142310
rect 169260 142028 169312 142034
rect 169260 141970 169312 141976
rect 135312 139512 135364 139518
rect 135312 139454 135364 139460
rect 138256 139512 138308 139518
rect 138256 139454 138308 139460
rect 135324 139217 135352 139454
rect 135310 139208 135366 139217
rect 135310 139143 135366 139152
rect 136966 139072 137022 139081
rect 136966 139007 137022 139016
rect 136874 138936 136930 138945
rect 136874 138871 136930 138880
rect 135404 138696 135456 138702
rect 135404 138638 135456 138644
rect 135312 138628 135364 138634
rect 135312 138570 135364 138576
rect 135218 137712 135274 137721
rect 135218 137647 135274 137656
rect 135220 137540 135272 137546
rect 135220 137482 135272 137488
rect 135128 137268 135180 137274
rect 135128 137210 135180 137216
rect 134300 135908 134352 135914
rect 134300 135850 134352 135856
rect 134312 133641 134340 135850
rect 135140 135409 135168 137210
rect 135232 135681 135260 137482
rect 135324 136633 135352 138570
rect 135416 136905 135444 138638
rect 136888 138634 136916 138871
rect 136980 138702 137008 139007
rect 136968 138696 137020 138702
rect 136968 138638 137020 138644
rect 136876 138628 136928 138634
rect 136876 138570 136928 138576
rect 169272 138566 169300 141970
rect 169260 138560 169312 138566
rect 169260 138502 169312 138508
rect 169364 138498 169392 142582
rect 169916 141422 169944 144892
rect 169904 141416 169956 141422
rect 169904 141358 169956 141364
rect 171020 141354 171048 144892
rect 172124 142306 172152 144892
rect 173228 142442 173256 144892
rect 174332 142510 174360 144892
rect 174320 142504 174372 142510
rect 174320 142446 174372 142452
rect 173216 142436 173268 142442
rect 173216 142378 173268 142384
rect 172112 142300 172164 142306
rect 172112 142242 172164 142248
rect 174596 142300 174648 142306
rect 174596 142242 174648 142248
rect 172756 142232 172808 142238
rect 174608 142209 174636 142242
rect 172756 142174 172808 142180
rect 174594 142200 174650 142209
rect 171008 141348 171060 141354
rect 171008 141290 171060 141296
rect 172768 139926 172796 142174
rect 174594 142135 174650 142144
rect 177184 141764 177212 147711
rect 177446 145464 177502 145473
rect 177446 145399 177502 145408
rect 177460 145094 177488 145399
rect 177448 145088 177500 145094
rect 177448 145030 177500 145036
rect 177736 141764 177764 148935
rect 178288 146658 178316 152607
rect 178366 151448 178422 151457
rect 178366 151383 178422 151392
rect 178380 150346 178408 151383
rect 178380 150318 178776 150346
rect 178458 150224 178514 150233
rect 178458 150159 178514 150168
rect 178276 146652 178328 146658
rect 178276 146594 178328 146600
rect 178182 146552 178238 146561
rect 178238 146510 178316 146538
rect 178182 146487 178238 146496
rect 178288 145298 178316 146510
rect 178276 145292 178328 145298
rect 178276 145234 178328 145240
rect 178472 145178 178500 150159
rect 178288 145150 178500 145178
rect 178288 141764 178316 145150
rect 178748 141778 178776 150318
rect 179012 146652 179064 146658
rect 179012 146594 179064 146600
rect 179024 141778 179052 146594
rect 179760 141778 179788 153734
rect 180312 146017 180340 153802
rect 180404 148329 180432 155094
rect 180496 150641 180524 156454
rect 200538 151584 200594 151593
rect 200538 151519 200540 151528
rect 200592 151519 200594 151528
rect 200540 151490 200592 151496
rect 180482 150632 180538 150641
rect 180482 150567 180538 150576
rect 180390 148320 180446 148329
rect 180390 148255 180446 148264
rect 180298 146008 180354 146017
rect 180298 145943 180354 145952
rect 181128 145292 181180 145298
rect 181128 145234 181180 145240
rect 180576 145088 180628 145094
rect 180576 145030 180628 145036
rect 178748 141750 178854 141778
rect 179024 141750 179406 141778
rect 179760 141750 180050 141778
rect 180588 141764 180616 145030
rect 181140 141764 181168 145234
rect 182796 144878 183132 144906
rect 183256 144878 183500 144906
rect 183624 144878 183868 144906
rect 183992 144878 184328 144906
rect 184452 144878 184696 144906
rect 184820 144878 185064 144906
rect 185280 144878 185524 144906
rect 185740 144878 185892 144906
rect 182232 142708 182284 142714
rect 182232 142650 182284 142656
rect 181680 142368 181732 142374
rect 181680 142310 181732 142316
rect 181692 141764 181720 142310
rect 182244 141764 182272 142650
rect 182796 142374 182824 144878
rect 183256 142714 183284 144878
rect 183244 142708 183296 142714
rect 183244 142650 183296 142656
rect 182784 142368 182836 142374
rect 182784 142310 182836 142316
rect 183624 142102 183652 144878
rect 183992 142186 184020 144878
rect 183808 142158 184020 142186
rect 182876 142096 182928 142102
rect 182876 142038 182928 142044
rect 183612 142096 183664 142102
rect 183612 142038 183664 142044
rect 182888 141764 182916 142038
rect 183808 141778 183836 142158
rect 184452 141778 184480 144878
rect 184820 141778 184848 144878
rect 185280 141778 185308 144878
rect 183454 141750 183836 141778
rect 184006 141750 184480 141778
rect 184558 141750 184848 141778
rect 185110 141750 185308 141778
rect 185740 141764 185768 144878
rect 186246 144634 186274 144892
rect 186720 144878 186872 144906
rect 187088 144878 187240 144906
rect 187456 144878 187700 144906
rect 187916 144878 188160 144906
rect 188284 144878 188528 144906
rect 188652 144878 188988 144906
rect 189112 144878 189356 144906
rect 189480 144878 189724 144906
rect 189848 144878 190184 144906
rect 190308 144878 190552 144906
rect 186246 144606 186320 144634
rect 186292 141764 186320 144606
rect 186844 141764 186872 144878
rect 187212 141778 187240 144878
rect 187672 141778 187700 144878
rect 188132 141778 188160 144878
rect 188500 141914 188528 144878
rect 188960 141914 188988 144878
rect 189328 142646 189356 144878
rect 189696 142714 189724 144878
rect 189684 142708 189736 142714
rect 189684 142650 189736 142656
rect 189316 142640 189368 142646
rect 189316 142582 189368 142588
rect 190156 142510 190184 144878
rect 190236 142640 190288 142646
rect 190236 142582 190288 142588
rect 190144 142504 190196 142510
rect 190144 142446 190196 142452
rect 188500 141886 188804 141914
rect 188960 141886 189264 141914
rect 188776 141778 188804 141886
rect 189236 141778 189264 141886
rect 187212 141750 187410 141778
rect 187672 141750 187962 141778
rect 188132 141750 188606 141778
rect 188776 141750 189158 141778
rect 189236 141750 189710 141778
rect 190248 141764 190276 142582
rect 190524 142170 190552 144878
rect 190616 144878 190676 144906
rect 191136 144878 191380 144906
rect 190616 144278 190644 144878
rect 190604 144272 190656 144278
rect 190604 144214 190656 144220
rect 191352 142714 191380 144878
rect 191490 144686 191518 144892
rect 191858 144754 191886 144892
rect 192332 144878 192484 144906
rect 192700 144878 192944 144906
rect 193068 144878 193404 144906
rect 193528 144878 193772 144906
rect 193896 144878 194140 144906
rect 194264 144878 194600 144906
rect 191846 144748 191898 144754
rect 191846 144690 191898 144696
rect 191478 144680 191530 144686
rect 191478 144622 191530 144628
rect 190788 142708 190840 142714
rect 190788 142650 190840 142656
rect 191340 142708 191392 142714
rect 191340 142650 191392 142656
rect 190512 142164 190564 142170
rect 190512 142106 190564 142112
rect 190800 141764 190828 142650
rect 191432 142504 191484 142510
rect 191432 142446 191484 142452
rect 191444 141764 191472 142446
rect 192456 142374 192484 144878
rect 192536 144272 192588 144278
rect 192536 144214 192588 144220
rect 192444 142368 192496 142374
rect 192444 142310 192496 142316
rect 191984 142164 192036 142170
rect 191984 142106 192036 142112
rect 191996 141764 192024 142106
rect 192548 141764 192576 144214
rect 192916 142442 192944 144878
rect 193088 142708 193140 142714
rect 193088 142650 193140 142656
rect 192904 142436 192956 142442
rect 192904 142378 192956 142384
rect 193100 141764 193128 142650
rect 193376 142170 193404 144878
rect 193640 144680 193692 144686
rect 193640 144622 193692 144628
rect 193364 142164 193416 142170
rect 193364 142106 193416 142112
rect 193652 141764 193680 144622
rect 193744 142034 193772 144878
rect 194112 142714 194140 144878
rect 194284 144748 194336 144754
rect 194284 144690 194336 144696
rect 194100 142708 194152 142714
rect 194100 142650 194152 142656
rect 193732 142028 193784 142034
rect 193732 141970 193784 141976
rect 194296 141764 194324 144690
rect 194572 142510 194600 144878
rect 194664 144878 194724 144906
rect 195092 144878 195336 144906
rect 195460 144878 195796 144906
rect 195920 144878 196164 144906
rect 196288 144878 196532 144906
rect 196656 144878 196992 144906
rect 197116 144878 197360 144906
rect 194560 142504 194612 142510
rect 194560 142446 194612 142452
rect 194664 142306 194692 144878
rect 194836 142368 194888 142374
rect 194836 142310 194888 142316
rect 194652 142300 194704 142306
rect 194652 142242 194704 142248
rect 194848 141764 194876 142310
rect 195308 142238 195336 144878
rect 195768 142442 195796 144878
rect 195388 142436 195440 142442
rect 195388 142378 195440 142384
rect 195756 142436 195808 142442
rect 195756 142378 195808 142384
rect 195296 142232 195348 142238
rect 195296 142174 195348 142180
rect 195400 141764 195428 142378
rect 196136 142374 196164 144878
rect 196124 142368 196176 142374
rect 196124 142310 196176 142316
rect 196504 142170 196532 144878
rect 196964 142646 196992 144878
rect 197136 142708 197188 142714
rect 197136 142650 197188 142656
rect 196952 142640 197004 142646
rect 196952 142582 197004 142588
rect 195940 142164 195992 142170
rect 195940 142106 195992 142112
rect 196492 142164 196544 142170
rect 196492 142106 196544 142112
rect 195952 141764 195980 142106
rect 196492 142028 196544 142034
rect 196492 141970 196544 141976
rect 196504 141764 196532 141970
rect 197148 141764 197176 142650
rect 197332 142578 197360 144878
rect 197424 144878 197484 144906
rect 197320 142572 197372 142578
rect 197320 142514 197372 142520
rect 197424 141830 197452 144878
rect 197838 144686 197866 144892
rect 198312 144878 198556 144906
rect 198680 144878 198924 144906
rect 197826 144680 197878 144686
rect 197826 144622 197878 144628
rect 198528 144278 198556 144878
rect 198516 144272 198568 144278
rect 198516 144214 198568 144220
rect 198896 144210 198924 144878
rect 198884 144204 198936 144210
rect 198884 144146 198936 144152
rect 201012 142714 201040 164847
rect 222632 163402 222660 166094
rect 224458 163552 224514 163561
rect 224458 163487 224514 163496
rect 222632 163374 222752 163402
rect 207438 163280 207494 163289
rect 207438 163215 207494 163224
rect 207452 153769 207480 163215
rect 222724 159594 222752 163374
rect 222632 159566 222752 159594
rect 222632 158098 222660 159566
rect 223538 159200 223594 159209
rect 223538 159135 223594 159144
rect 222632 158070 222936 158098
rect 222804 156920 222856 156926
rect 222540 156868 222804 156874
rect 222540 156862 222856 156868
rect 222540 156846 222844 156862
rect 207438 153760 207494 153769
rect 207438 153695 207494 153704
rect 207438 152264 207494 152273
rect 207438 152199 207494 152208
rect 204494 151584 204550 151593
rect 207452 151554 207480 152199
rect 204494 151519 204550 151528
rect 207440 151548 207492 151554
rect 202840 144680 202892 144686
rect 202840 144622 202892 144628
rect 201000 142708 201052 142714
rect 201000 142650 201052 142656
rect 201092 142640 201144 142646
rect 201092 142582 201144 142588
rect 197688 142504 197740 142510
rect 197688 142446 197740 142452
rect 197412 141824 197464 141830
rect 197412 141766 197464 141772
rect 197700 141764 197728 142446
rect 199068 142436 199120 142442
rect 199068 142378 199120 142384
rect 198240 142300 198292 142306
rect 198240 142242 198292 142248
rect 198252 141764 198280 142242
rect 198792 142232 198844 142238
rect 198792 142174 198844 142180
rect 198804 141764 198832 142174
rect 199080 141778 199108 142378
rect 199620 142368 199672 142374
rect 199620 142310 199672 142316
rect 199632 141778 199660 142310
rect 200540 142164 200592 142170
rect 200540 142106 200592 142112
rect 199080 141750 199370 141778
rect 199632 141750 200014 141778
rect 200552 141764 200580 142106
rect 201104 141764 201132 142582
rect 201644 142572 201696 142578
rect 201644 142514 201696 142520
rect 201656 141764 201684 142514
rect 201828 141824 201880 141830
rect 201880 141772 202222 141778
rect 201828 141766 202222 141772
rect 201840 141750 202222 141766
rect 202852 141764 202880 144622
rect 203392 144272 203444 144278
rect 203392 144214 203444 144220
rect 203404 141764 203432 144214
rect 203944 144204 203996 144210
rect 203944 144146 203996 144152
rect 203956 141764 203984 144146
rect 204508 141764 204536 151519
rect 207440 151490 207492 151496
rect 207452 142753 207480 151490
rect 207438 142744 207494 142753
rect 207438 142679 207494 142688
rect 207898 142608 207954 142617
rect 207898 142543 207954 142552
rect 207912 141966 207940 142543
rect 207992 142028 208044 142034
rect 207992 141970 208044 141976
rect 207900 141960 207952 141966
rect 207900 141902 207952 141908
rect 174228 141280 174280 141286
rect 174228 141222 174280 141228
rect 174240 140441 174268 141222
rect 174412 141212 174464 141218
rect 174412 141154 174464 141160
rect 174424 140985 174452 141154
rect 174410 140976 174466 140985
rect 174410 140911 174466 140920
rect 174226 140432 174282 140441
rect 174226 140367 174282 140376
rect 172756 139920 172808 139926
rect 172756 139862 172808 139868
rect 174320 139920 174372 139926
rect 174320 139862 174372 139868
rect 174136 139852 174188 139858
rect 174136 139794 174188 139800
rect 174148 139217 174176 139794
rect 174228 139784 174280 139790
rect 174332 139761 174360 139862
rect 174228 139726 174280 139732
rect 174318 139752 174374 139761
rect 174134 139208 174190 139217
rect 174134 139143 174190 139152
rect 172570 139072 172626 139081
rect 172570 139007 172626 139016
rect 172202 138664 172258 138673
rect 172202 138599 172258 138608
rect 169352 138492 169404 138498
rect 169352 138434 169404 138440
rect 136874 137848 136930 137857
rect 136874 137783 136930 137792
rect 136888 137546 136916 137783
rect 136876 137540 136928 137546
rect 136876 137482 136928 137488
rect 136874 137304 136930 137313
rect 136874 137239 136876 137248
rect 136928 137239 136930 137248
rect 136876 137210 136928 137216
rect 172216 137070 172244 138599
rect 172584 137138 172612 139007
rect 174240 138673 174268 139726
rect 174318 139687 174374 139696
rect 174226 138664 174282 138673
rect 174226 138599 174282 138608
rect 174228 138560 174280 138566
rect 174228 138502 174280 138508
rect 174136 138492 174188 138498
rect 174136 138434 174188 138440
rect 174148 137993 174176 138434
rect 174134 137984 174190 137993
rect 174134 137919 174190 137928
rect 172662 137848 172718 137857
rect 172718 137806 172796 137834
rect 172662 137783 172718 137792
rect 172662 137304 172718 137313
rect 172662 137239 172664 137248
rect 172716 137239 172718 137248
rect 172664 137210 172716 137216
rect 172572 137132 172624 137138
rect 172572 137074 172624 137080
rect 172204 137064 172256 137070
rect 172204 137006 172256 137012
rect 135402 136896 135458 136905
rect 135402 136831 135458 136840
rect 135310 136624 135366 136633
rect 135310 136559 135366 136568
rect 136782 136624 136838 136633
rect 136782 136559 136838 136568
rect 172570 136624 172626 136633
rect 172570 136559 172626 136568
rect 135312 135840 135364 135846
rect 135312 135782 135364 135788
rect 135218 135672 135274 135681
rect 135218 135607 135274 135616
rect 135220 135432 135272 135438
rect 135126 135400 135182 135409
rect 135220 135374 135272 135380
rect 135126 135335 135182 135344
rect 135232 134865 135260 135374
rect 135218 134856 135274 134865
rect 135218 134791 135274 134800
rect 135128 134548 135180 134554
rect 135128 134490 135180 134496
rect 134298 133632 134354 133641
rect 134298 133567 134354 133576
rect 135140 132553 135168 134490
rect 135324 134321 135352 135782
rect 136796 135438 136824 136559
rect 136874 136080 136930 136089
rect 136874 136015 136930 136024
rect 136888 135846 136916 136015
rect 136966 135944 137022 135953
rect 136966 135879 136968 135888
rect 137020 135879 137022 135888
rect 136968 135850 137020 135856
rect 172584 135846 172612 136559
rect 172662 136080 172718 136089
rect 172662 136015 172664 136024
rect 172716 136015 172718 136024
rect 172664 135986 172716 135992
rect 172662 135944 172718 135953
rect 172662 135879 172664 135888
rect 172716 135879 172718 135888
rect 172664 135850 172716 135856
rect 136876 135840 136928 135846
rect 136876 135782 136928 135788
rect 172572 135840 172624 135846
rect 172572 135782 172624 135788
rect 172768 135710 172796 137806
rect 174240 137449 174268 138502
rect 174226 137440 174282 137449
rect 174226 137375 174282 137384
rect 174044 137268 174096 137274
rect 174044 137210 174096 137216
rect 173952 136044 174004 136050
rect 173952 135986 174004 135992
rect 173768 135908 173820 135914
rect 173768 135850 173820 135856
rect 172756 135704 172808 135710
rect 172756 135646 172808 135652
rect 136784 135432 136836 135438
rect 136784 135374 136836 135380
rect 136874 134856 136930 134865
rect 136874 134791 136930 134800
rect 172662 134856 172718 134865
rect 172662 134791 172718 134800
rect 136888 134486 136916 134791
rect 136966 134720 137022 134729
rect 136966 134655 137022 134664
rect 136980 134554 137008 134655
rect 172570 134584 172626 134593
rect 136968 134548 137020 134554
rect 172676 134554 172704 134791
rect 172570 134519 172626 134528
rect 172664 134548 172716 134554
rect 136968 134490 137020 134496
rect 172584 134486 172612 134519
rect 172664 134490 172716 134496
rect 135404 134480 135456 134486
rect 135404 134422 135456 134428
rect 136876 134480 136928 134486
rect 136876 134422 136928 134428
rect 172572 134480 172624 134486
rect 172572 134422 172624 134428
rect 135310 134312 135366 134321
rect 135310 134247 135366 134256
rect 135220 133120 135272 133126
rect 135220 133062 135272 133068
rect 135126 132544 135182 132553
rect 135126 132479 135182 132488
rect 135036 131760 135088 131766
rect 135036 131702 135088 131708
rect 134300 130808 134352 130814
rect 134298 130776 134300 130785
rect 134352 130776 134354 130785
rect 134298 130711 134354 130720
rect 135048 129561 135076 131702
rect 135232 131601 135260 133062
rect 135312 133052 135364 133058
rect 135312 132994 135364 133000
rect 135218 131592 135274 131601
rect 135218 131527 135274 131536
rect 135324 131329 135352 132994
rect 135416 132825 135444 134422
rect 136966 133632 137022 133641
rect 136966 133567 137022 133576
rect 171650 133632 171706 133641
rect 171650 133567 171706 133576
rect 136980 133126 137008 133567
rect 171664 133126 171692 133567
rect 173780 133369 173808 135850
rect 173860 134480 173912 134486
rect 173860 134422 173912 134428
rect 173766 133360 173822 133369
rect 173766 133295 173822 133304
rect 136968 133120 137020 133126
rect 136874 133088 136930 133097
rect 136968 133062 137020 133068
rect 171652 133120 171704 133126
rect 173216 133120 173268 133126
rect 171652 133062 171704 133068
rect 172662 133088 172718 133097
rect 136874 133023 136876 133032
rect 136928 133023 136930 133032
rect 172718 133046 172796 133074
rect 173216 133062 173268 133068
rect 172662 133023 172718 133032
rect 136876 132994 136928 133000
rect 135402 132816 135458 132825
rect 172768 132802 172796 133046
rect 172768 132774 172980 132802
rect 135402 132751 135458 132760
rect 136782 132408 136838 132417
rect 136782 132343 136838 132352
rect 172018 132408 172074 132417
rect 172018 132343 172074 132352
rect 135404 131692 135456 131698
rect 135404 131634 135456 131640
rect 135310 131320 135366 131329
rect 135310 131255 135366 131264
rect 135128 130400 135180 130406
rect 135128 130342 135180 130348
rect 135034 129552 135090 129561
rect 135034 129487 135090 129496
rect 134300 129040 134352 129046
rect 134300 128982 134352 128988
rect 132644 127408 132696 127414
rect 132644 127350 132696 127356
rect 132736 127408 132788 127414
rect 132736 127350 132788 127356
rect 102282 126424 102338 126433
rect 102282 126359 102338 126368
rect 102284 126252 102336 126258
rect 102284 126194 102336 126200
rect 102006 125744 102062 125753
rect 102006 125679 102062 125688
rect 102100 125164 102152 125170
rect 102100 125106 102152 125112
rect 102008 124892 102060 124898
rect 102008 124834 102060 124840
rect 100996 124756 101048 124762
rect 100996 124698 101048 124704
rect 65024 124144 65076 124150
rect 65024 124086 65076 124092
rect 100626 124112 100682 124121
rect 100626 124047 100682 124056
rect 66402 123976 66458 123985
rect 66402 123911 66458 123920
rect 65022 123568 65078 123577
rect 65022 123503 65078 123512
rect 63552 123396 63604 123402
rect 63552 123338 63604 123344
rect 62906 123160 62962 123169
rect 62906 123095 62962 123104
rect 62816 122648 62868 122654
rect 62814 122616 62816 122625
rect 62868 122616 62870 122625
rect 62814 122551 62870 122560
rect 63460 122104 63512 122110
rect 63460 122046 63512 122052
rect 62816 121492 62868 121498
rect 62816 121434 62868 121440
rect 62828 121401 62856 121434
rect 62814 121392 62870 121401
rect 62814 121327 62870 121336
rect 63472 120585 63500 122046
rect 63564 121673 63592 123338
rect 65036 122654 65064 123503
rect 66416 123402 66444 123911
rect 100640 123674 100668 124047
rect 100628 123668 100680 123674
rect 100628 123610 100680 123616
rect 99890 123432 99946 123441
rect 66404 123396 66456 123402
rect 99890 123367 99892 123376
rect 66404 123338 66456 123344
rect 99944 123367 99946 123376
rect 99892 123338 99944 123344
rect 102020 122897 102048 124834
rect 102112 123441 102140 125106
rect 102296 124665 102324 126194
rect 102376 126116 102428 126122
rect 102376 126058 102428 126064
rect 102388 125209 102416 126058
rect 102374 125200 102430 125209
rect 102374 125135 102430 125144
rect 102376 124756 102428 124762
rect 102376 124698 102428 124704
rect 102282 124656 102338 124665
rect 102282 124591 102338 124600
rect 102388 123985 102416 124698
rect 102374 123976 102430 123985
rect 102374 123911 102430 123920
rect 102284 123668 102336 123674
rect 102284 123610 102336 123616
rect 102098 123432 102154 123441
rect 102098 123367 102154 123376
rect 102192 123396 102244 123402
rect 102192 123338 102244 123344
rect 100166 122888 100222 122897
rect 100166 122823 100222 122832
rect 102006 122888 102062 122897
rect 102006 122823 102062 122832
rect 66310 122752 66366 122761
rect 66310 122687 66366 122696
rect 65024 122648 65076 122654
rect 65024 122590 65076 122596
rect 65022 122480 65078 122489
rect 65022 122415 65078 122424
rect 63644 122036 63696 122042
rect 63644 121978 63696 121984
rect 63550 121664 63606 121673
rect 63550 121599 63606 121608
rect 63458 120576 63514 120585
rect 63458 120511 63514 120520
rect 63656 120313 63684 121978
rect 65036 121498 65064 122415
rect 66324 122110 66352 122687
rect 100180 122246 100208 122823
rect 100994 122344 101050 122353
rect 100994 122279 101050 122288
rect 100168 122240 100220 122246
rect 66402 122208 66458 122217
rect 100168 122182 100220 122188
rect 100902 122208 100958 122217
rect 66402 122143 66458 122152
rect 100902 122143 100958 122152
rect 66312 122104 66364 122110
rect 66312 122046 66364 122052
rect 66416 122042 66444 122143
rect 100916 122110 100944 122143
rect 100904 122104 100956 122110
rect 100904 122046 100956 122052
rect 66404 122036 66456 122042
rect 66404 121978 66456 121984
rect 65024 121492 65076 121498
rect 65024 121434 65076 121440
rect 100626 121120 100682 121129
rect 100626 121055 100682 121064
rect 66218 120984 66274 120993
rect 100640 120954 100668 121055
rect 66218 120919 66274 120928
rect 100628 120948 100680 120954
rect 65022 120712 65078 120721
rect 65022 120647 65078 120656
rect 63642 120304 63698 120313
rect 63642 120239 63698 120248
rect 65036 120002 65064 120647
rect 62816 119996 62868 120002
rect 62816 119938 62868 119944
rect 65024 119996 65076 120002
rect 65024 119938 65076 119944
rect 62828 119633 62856 119938
rect 62814 119624 62870 119633
rect 62814 119559 62870 119568
rect 65022 119488 65078 119497
rect 65022 119423 65078 119432
rect 62908 119316 62960 119322
rect 62908 119258 62960 119264
rect 62724 119180 62776 119186
rect 62724 119122 62776 119128
rect 62736 118817 62764 119122
rect 62722 118808 62778 118817
rect 62722 118743 62778 118752
rect 62816 118772 62868 118778
rect 62816 118714 62868 118720
rect 62828 118545 62856 118714
rect 62814 118536 62870 118545
rect 62814 118471 62870 118480
rect 62724 117888 62776 117894
rect 62920 117865 62948 119258
rect 65036 118778 65064 119423
rect 66232 119186 66260 120919
rect 100628 120890 100680 120896
rect 100626 120712 100682 120721
rect 100626 120647 100628 120656
rect 100680 120647 100682 120656
rect 100628 120618 100680 120624
rect 101008 120614 101036 122279
rect 102100 122104 102152 122110
rect 102100 122046 102152 122052
rect 100996 120608 101048 120614
rect 100996 120550 101048 120556
rect 102112 119905 102140 122046
rect 102204 121673 102232 123338
rect 102296 122353 102324 123610
rect 102282 122344 102338 122353
rect 102282 122279 102338 122288
rect 102284 122240 102336 122246
rect 102284 122182 102336 122188
rect 102190 121664 102246 121673
rect 102190 121599 102246 121608
rect 102296 121129 102324 122182
rect 102282 121120 102338 121129
rect 102282 121055 102338 121064
rect 102284 120948 102336 120954
rect 102284 120890 102336 120896
rect 102192 120676 102244 120682
rect 102192 120618 102244 120624
rect 100626 119896 100682 119905
rect 100626 119831 100682 119840
rect 102098 119896 102154 119905
rect 102098 119831 102154 119840
rect 66402 119760 66458 119769
rect 66402 119695 66458 119704
rect 66416 119322 66444 119695
rect 100640 119458 100668 119831
rect 100628 119452 100680 119458
rect 100628 119394 100680 119400
rect 100902 119352 100958 119361
rect 66404 119316 66456 119322
rect 100958 119310 101036 119338
rect 100902 119287 100958 119296
rect 66404 119258 66456 119264
rect 66402 119216 66458 119225
rect 66220 119180 66272 119186
rect 66402 119151 66458 119160
rect 66220 119122 66272 119128
rect 65024 118772 65076 118778
rect 65024 118714 65076 118720
rect 64930 118536 64986 118545
rect 64930 118471 64986 118480
rect 62724 117830 62776 117836
rect 62906 117856 62962 117865
rect 62736 116233 62764 117830
rect 62906 117791 62962 117800
rect 62816 117344 62868 117350
rect 62814 117312 62816 117321
rect 62868 117312 62870 117321
rect 62814 117247 62870 117256
rect 64944 117214 64972 118471
rect 66416 118273 66444 119151
rect 100626 118672 100682 118681
rect 100626 118607 100682 118616
rect 100640 118370 100668 118607
rect 100628 118364 100680 118370
rect 100628 118306 100680 118312
rect 65022 118264 65078 118273
rect 65022 118199 65078 118208
rect 66402 118264 66458 118273
rect 66402 118199 66458 118208
rect 65036 117350 65064 118199
rect 100626 118128 100682 118137
rect 100626 118063 100682 118072
rect 66402 117992 66458 118001
rect 100640 117962 100668 118063
rect 100718 117992 100774 118001
rect 66402 117927 66458 117936
rect 100628 117956 100680 117962
rect 66416 117894 66444 117927
rect 100718 117927 100774 117936
rect 100628 117898 100680 117904
rect 66404 117888 66456 117894
rect 66404 117830 66456 117836
rect 65024 117344 65076 117350
rect 65024 117286 65076 117292
rect 62816 117208 62868 117214
rect 62816 117150 62868 117156
rect 64932 117208 64984 117214
rect 64932 117150 64984 117156
rect 62828 116777 62856 117150
rect 100534 116904 100590 116913
rect 100534 116839 100590 116848
rect 62814 116768 62870 116777
rect 62814 116703 62870 116712
rect 66402 116768 66458 116777
rect 66402 116703 66458 116712
rect 65022 116496 65078 116505
rect 65022 116431 65078 116440
rect 62722 116224 62778 116233
rect 62722 116159 62778 116168
rect 65036 115786 65064 116431
rect 62816 115780 62868 115786
rect 62816 115722 62868 115728
rect 65024 115780 65076 115786
rect 65024 115722 65076 115728
rect 62828 115553 62856 115722
rect 62814 115544 62870 115553
rect 62814 115479 62870 115488
rect 65022 115136 65078 115145
rect 65022 115071 65078 115080
rect 62816 114896 62868 114902
rect 62816 114838 62868 114844
rect 62828 114737 62856 114838
rect 62814 114728 62870 114737
rect 62814 114663 62870 114672
rect 65036 114630 65064 115071
rect 66416 114902 66444 116703
rect 100548 116534 100576 116839
rect 100626 116768 100682 116777
rect 100626 116703 100682 116712
rect 100640 116670 100668 116703
rect 100628 116664 100680 116670
rect 100628 116606 100680 116612
rect 100536 116528 100588 116534
rect 100536 116470 100588 116476
rect 100732 116398 100760 117927
rect 101008 117826 101036 119310
rect 102204 118817 102232 120618
rect 102296 119633 102324 120890
rect 102376 120608 102428 120614
rect 102374 120576 102376 120585
rect 102428 120576 102430 120585
rect 102374 120511 102430 120520
rect 102282 119624 102338 119633
rect 102282 119559 102338 119568
rect 102284 119452 102336 119458
rect 102284 119394 102336 119400
rect 102190 118808 102246 118817
rect 102190 118743 102246 118752
rect 102192 118364 102244 118370
rect 102192 118306 102244 118312
rect 100996 117820 101048 117826
rect 100996 117762 101048 117768
rect 102204 117049 102232 118306
rect 102296 118273 102324 119394
rect 132656 118302 132684 127350
rect 134312 127249 134340 128982
rect 135140 128473 135168 130342
rect 135312 130332 135364 130338
rect 135312 130274 135364 130280
rect 135220 128972 135272 128978
rect 135220 128914 135272 128920
rect 135126 128464 135182 128473
rect 135126 128399 135182 128408
rect 135128 127612 135180 127618
rect 135128 127554 135180 127560
rect 134298 127240 134354 127249
rect 134298 127175 134354 127184
rect 134668 127204 134720 127210
rect 134668 127146 134720 127152
rect 134680 126705 134708 127146
rect 134666 126696 134722 126705
rect 134666 126631 134722 126640
rect 134852 126116 134904 126122
rect 134852 126058 134904 126064
rect 134864 125481 134892 126058
rect 135140 126025 135168 127554
rect 135232 127521 135260 128914
rect 135324 128745 135352 130274
rect 135416 130241 135444 131634
rect 136796 130814 136824 132343
rect 136874 132000 136930 132009
rect 136874 131935 136930 131944
rect 171650 132000 171706 132009
rect 171650 131935 171706 131944
rect 136888 131698 136916 131935
rect 136968 131760 137020 131766
rect 136966 131728 136968 131737
rect 137020 131728 137022 131737
rect 136876 131692 136928 131698
rect 171664 131698 171692 131935
rect 172032 131766 172060 132343
rect 172662 131864 172718 131873
rect 172718 131822 172888 131850
rect 172662 131799 172718 131808
rect 172020 131760 172072 131766
rect 172020 131702 172072 131708
rect 172756 131760 172808 131766
rect 172756 131702 172808 131708
rect 136966 131663 137022 131672
rect 171652 131692 171704 131698
rect 136876 131634 136928 131640
rect 171652 131634 171704 131640
rect 172768 131086 172796 131702
rect 172756 131080 172808 131086
rect 172756 131022 172808 131028
rect 136784 130808 136836 130814
rect 136784 130750 136836 130756
rect 136874 130640 136930 130649
rect 136874 130575 136930 130584
rect 172386 130640 172442 130649
rect 172386 130575 172388 130584
rect 136888 130338 136916 130575
rect 172440 130575 172442 130584
rect 172388 130546 172440 130552
rect 136966 130504 137022 130513
rect 136966 130439 137022 130448
rect 136980 130406 137008 130439
rect 136968 130400 137020 130406
rect 136968 130342 137020 130348
rect 172662 130368 172718 130377
rect 136876 130332 136928 130338
rect 172718 130326 172796 130354
rect 172662 130303 172718 130312
rect 136876 130274 136928 130280
rect 135402 130232 135458 130241
rect 135402 130167 135458 130176
rect 136874 129416 136930 129425
rect 136874 129351 136930 129360
rect 172662 129416 172718 129425
rect 172662 129351 172718 129360
rect 136888 128978 136916 129351
rect 172676 129250 172704 129351
rect 172664 129244 172716 129250
rect 172664 129186 172716 129192
rect 136968 129040 137020 129046
rect 136966 129008 136968 129017
rect 137020 129008 137022 129017
rect 136876 128972 136928 128978
rect 136966 128943 137022 128952
rect 172662 129008 172718 129017
rect 172662 128943 172664 128952
rect 136876 128914 136928 128920
rect 172716 128943 172718 128952
rect 172664 128914 172716 128920
rect 172768 128910 172796 130326
rect 172860 130202 172888 131822
rect 172952 131358 172980 132774
rect 173228 131714 173256 133062
rect 173872 132281 173900 134422
rect 173964 133913 173992 135986
rect 174056 135137 174084 137210
rect 174136 137132 174188 137138
rect 174136 137074 174188 137080
rect 174148 136905 174176 137074
rect 174228 137064 174280 137070
rect 174228 137006 174280 137012
rect 174134 136896 174190 136905
rect 174134 136831 174190 136840
rect 174240 136361 174268 137006
rect 204770 136624 204826 136633
rect 204770 136559 204826 136568
rect 174226 136352 174282 136361
rect 174226 136287 174282 136296
rect 174228 135772 174280 135778
rect 174228 135714 174280 135720
rect 174136 135704 174188 135710
rect 174134 135672 174136 135681
rect 174188 135672 174190 135681
rect 174134 135607 174190 135616
rect 174042 135128 174098 135137
rect 174042 135063 174098 135072
rect 174240 134593 174268 135714
rect 174226 134584 174282 134593
rect 174044 134548 174096 134554
rect 174226 134519 174282 134528
rect 174044 134490 174096 134496
rect 173950 133904 174006 133913
rect 173950 133839 174006 133848
rect 174056 132825 174084 134490
rect 204784 134418 204812 136559
rect 204772 134412 204824 134418
rect 204772 134354 204824 134360
rect 204956 134412 205008 134418
rect 204956 134354 205008 134360
rect 174042 132816 174098 132825
rect 174042 132751 174098 132760
rect 173858 132272 173914 132281
rect 173858 132207 173914 132216
rect 173032 131692 173084 131698
rect 173032 131634 173084 131640
rect 173136 131686 173256 131714
rect 172940 131352 172992 131358
rect 172940 131294 172992 131300
rect 173044 130270 173072 131634
rect 173136 131630 173164 131686
rect 173124 131624 173176 131630
rect 174136 131624 174188 131630
rect 173124 131566 173176 131572
rect 174134 131592 174136 131601
rect 174188 131592 174190 131601
rect 174134 131527 174190 131536
rect 175056 131352 175108 131358
rect 175056 131294 175108 131300
rect 174136 131080 174188 131086
rect 175068 131057 175096 131294
rect 174136 131022 174188 131028
rect 175054 131048 175110 131057
rect 174044 130604 174096 130610
rect 174044 130546 174096 130552
rect 173032 130264 173084 130270
rect 173032 130206 173084 130212
rect 172848 130196 172900 130202
rect 172848 130138 172900 130144
rect 173952 129244 174004 129250
rect 173952 129186 174004 129192
rect 173860 128972 173912 128978
rect 173860 128914 173912 128920
rect 172756 128904 172808 128910
rect 172756 128846 172808 128852
rect 135310 128736 135366 128745
rect 135310 128671 135366 128680
rect 136782 128328 136838 128337
rect 136782 128263 136838 128272
rect 171650 128328 171706 128337
rect 171650 128263 171706 128272
rect 135218 127512 135274 127521
rect 135218 127447 135274 127456
rect 136796 127210 136824 128263
rect 136874 127648 136930 127657
rect 136874 127583 136876 127592
rect 136928 127583 136930 127592
rect 136876 127554 136928 127560
rect 171664 127550 171692 128263
rect 172662 127648 172718 127657
rect 172718 127606 172796 127634
rect 172662 127583 172718 127592
rect 171652 127544 171704 127550
rect 171652 127486 171704 127492
rect 136784 127204 136836 127210
rect 136784 127146 136836 127152
rect 136782 127104 136838 127113
rect 136782 127039 136838 127048
rect 172018 127104 172074 127113
rect 172018 127039 172074 127048
rect 135404 126252 135456 126258
rect 135404 126194 135456 126200
rect 135312 126184 135364 126190
rect 135312 126126 135364 126132
rect 135126 126016 135182 126025
rect 135126 125951 135182 125960
rect 134850 125472 134906 125481
rect 134850 125407 134906 125416
rect 135128 124824 135180 124830
rect 135128 124766 135180 124772
rect 135140 123169 135168 124766
rect 135324 124665 135352 126126
rect 135310 124656 135366 124665
rect 135310 124591 135366 124600
rect 135220 124416 135272 124422
rect 135416 124393 135444 126194
rect 136796 126122 136824 127039
rect 136874 126424 136930 126433
rect 136874 126359 136930 126368
rect 136888 126190 136916 126359
rect 136966 126288 137022 126297
rect 136966 126223 136968 126232
rect 137020 126223 137022 126232
rect 136968 126194 137020 126200
rect 172032 126190 172060 127039
rect 172386 126424 172442 126433
rect 172386 126359 172388 126368
rect 172440 126359 172442 126368
rect 172388 126330 172440 126336
rect 172664 126252 172716 126258
rect 172664 126194 172716 126200
rect 136876 126184 136928 126190
rect 136876 126126 136928 126132
rect 172020 126184 172072 126190
rect 172676 126161 172704 126194
rect 172020 126126 172072 126132
rect 172662 126152 172718 126161
rect 136784 126116 136836 126122
rect 172662 126087 172718 126096
rect 136784 126058 136836 126064
rect 172768 126054 172796 127606
rect 173872 126977 173900 128914
rect 173964 127521 173992 129186
rect 174056 128745 174084 130546
rect 174148 130513 174176 131022
rect 175054 130983 175110 130992
rect 174134 130504 174190 130513
rect 174134 130439 174190 130448
rect 174136 130264 174188 130270
rect 174136 130206 174188 130212
rect 174148 129833 174176 130206
rect 174504 130196 174556 130202
rect 174504 130138 174556 130144
rect 174134 129824 174190 129833
rect 174134 129759 174190 129768
rect 174516 129289 174544 130138
rect 174502 129280 174558 129289
rect 174502 129215 174558 129224
rect 174136 128904 174188 128910
rect 174136 128846 174188 128852
rect 174042 128736 174098 128745
rect 174042 128671 174098 128680
rect 174148 128201 174176 128846
rect 174134 128192 174190 128201
rect 174134 128127 174190 128136
rect 173950 127512 174006 127521
rect 173950 127447 174006 127456
rect 174228 127476 174280 127482
rect 174228 127418 174280 127424
rect 173858 126968 173914 126977
rect 173858 126903 173914 126912
rect 174240 126433 174268 127418
rect 174226 126424 174282 126433
rect 174044 126388 174096 126394
rect 174226 126359 174282 126368
rect 174044 126330 174096 126336
rect 173860 126252 173912 126258
rect 173860 126194 173912 126200
rect 172756 126048 172808 126054
rect 172756 125990 172808 125996
rect 136782 125336 136838 125345
rect 136782 125271 136838 125280
rect 172018 125336 172074 125345
rect 172018 125271 172074 125280
rect 136796 124422 136824 125271
rect 136874 124928 136930 124937
rect 136874 124863 136930 124872
rect 136888 124830 136916 124863
rect 172032 124830 172060 125271
rect 172662 124928 172718 124937
rect 172662 124863 172664 124872
rect 172716 124863 172718 124872
rect 172664 124834 172716 124840
rect 136876 124824 136928 124830
rect 136876 124766 136928 124772
rect 172020 124824 172072 124830
rect 172020 124766 172072 124772
rect 136784 124416 136836 124422
rect 135220 124358 135272 124364
rect 135402 124384 135458 124393
rect 135232 123713 135260 124358
rect 136784 124358 136836 124364
rect 135402 124319 135458 124328
rect 136782 124112 136838 124121
rect 136782 124047 136838 124056
rect 172386 124112 172442 124121
rect 172386 124047 172442 124056
rect 135218 123704 135274 123713
rect 135218 123639 135274 123648
rect 135404 123396 135456 123402
rect 135404 123338 135456 123344
rect 135126 123160 135182 123169
rect 135126 123095 135182 123104
rect 135312 122920 135364 122926
rect 135312 122862 135364 122868
rect 135324 122625 135352 122862
rect 135310 122616 135366 122625
rect 135310 122551 135366 122560
rect 135128 122172 135180 122178
rect 135128 122114 135180 122120
rect 135140 120313 135168 122114
rect 135220 122104 135272 122110
rect 135220 122046 135272 122052
rect 135232 120585 135260 122046
rect 135312 121968 135364 121974
rect 135416 121945 135444 123338
rect 136796 122926 136824 124047
rect 136874 123432 136930 123441
rect 172400 123402 172428 124047
rect 173872 123985 173900 126194
rect 173952 124892 174004 124898
rect 173952 124834 174004 124840
rect 173858 123976 173914 123985
rect 173858 123911 173914 123920
rect 172662 123432 172718 123441
rect 136874 123367 136876 123376
rect 136928 123367 136930 123376
rect 172388 123396 172440 123402
rect 136876 123338 136928 123344
rect 172718 123390 172888 123418
rect 172662 123367 172718 123376
rect 172388 123338 172440 123344
rect 136784 122920 136836 122926
rect 136784 122862 136836 122868
rect 136874 122888 136930 122897
rect 136874 122823 136930 122832
rect 171558 122888 171614 122897
rect 171558 122823 171614 122832
rect 136888 122042 136916 122823
rect 136966 122480 137022 122489
rect 136966 122415 137022 122424
rect 136980 122110 137008 122415
rect 137058 122208 137114 122217
rect 137058 122143 137060 122152
rect 137112 122143 137114 122152
rect 137060 122114 137112 122120
rect 136968 122104 137020 122110
rect 136968 122046 137020 122052
rect 171572 122042 171600 122823
rect 172662 122072 172718 122081
rect 136876 122036 136928 122042
rect 136876 121978 136928 121984
rect 171560 122036 171612 122042
rect 172718 122030 172796 122058
rect 172662 122007 172718 122016
rect 171560 121978 171612 121984
rect 135312 121910 135364 121916
rect 135402 121936 135458 121945
rect 135324 121401 135352 121910
rect 135402 121871 135458 121880
rect 135310 121392 135366 121401
rect 135310 121327 135366 121336
rect 136782 121120 136838 121129
rect 136782 121055 136838 121064
rect 171742 121120 171798 121129
rect 171742 121055 171798 121064
rect 135218 120576 135274 120585
rect 135218 120511 135274 120520
rect 135126 120304 135182 120313
rect 134852 120268 134904 120274
rect 136796 120274 136824 121055
rect 171756 120954 171784 121055
rect 171744 120948 171796 120954
rect 171744 120890 171796 120896
rect 136874 120712 136930 120721
rect 136874 120647 136930 120656
rect 172662 120712 172718 120721
rect 172662 120647 172664 120656
rect 135126 120239 135182 120248
rect 136784 120268 136836 120274
rect 134852 120210 134904 120216
rect 136784 120210 136836 120216
rect 134864 119633 134892 120210
rect 136782 119896 136838 119905
rect 136782 119831 136838 119840
rect 134850 119624 134906 119633
rect 134850 119559 134906 119568
rect 135220 119316 135272 119322
rect 135220 119258 135272 119264
rect 135036 118704 135088 118710
rect 135036 118646 135088 118652
rect 135048 118545 135076 118646
rect 135034 118536 135090 118545
rect 135034 118471 135090 118480
rect 132644 118296 132696 118302
rect 102282 118264 102338 118273
rect 132644 118238 132696 118244
rect 102282 118199 102338 118208
rect 132736 118160 132788 118166
rect 132656 118108 132736 118114
rect 132656 118102 132788 118108
rect 132656 118086 132776 118102
rect 102284 117956 102336 117962
rect 102284 117898 102336 117904
rect 102190 117040 102246 117049
rect 102190 116975 102246 116984
rect 102192 116664 102244 116670
rect 102192 116606 102244 116612
rect 100720 116392 100772 116398
rect 100720 116334 100772 116340
rect 72916 115910 73252 115938
rect 66404 114896 66456 114902
rect 66404 114838 66456 114844
rect 62816 114624 62868 114630
rect 62816 114566 62868 114572
rect 65024 114624 65076 114630
rect 65024 114566 65076 114572
rect 62828 114465 62856 114566
rect 62814 114456 62870 114465
rect 62814 114391 62870 114400
rect 32008 113870 33218 113898
rect 32008 104265 32036 113870
rect 33848 111638 33876 113884
rect 34492 112182 34520 113884
rect 34480 112176 34532 112182
rect 34480 112118 34532 112124
rect 35228 111910 35256 113884
rect 35216 111904 35268 111910
rect 35216 111846 35268 111852
rect 35872 111706 35900 113884
rect 35860 111700 35912 111706
rect 35860 111642 35912 111648
rect 33836 111632 33888 111638
rect 33836 111574 33888 111580
rect 36608 111230 36636 113884
rect 37252 111298 37280 113884
rect 37896 111570 37924 113884
rect 37884 111564 37936 111570
rect 37884 111506 37936 111512
rect 37240 111292 37292 111298
rect 37240 111234 37292 111240
rect 36596 111224 36648 111230
rect 36596 111166 36648 111172
rect 38632 111094 38660 113884
rect 39080 111632 39132 111638
rect 39080 111574 39132 111580
rect 38620 111088 38672 111094
rect 38620 111030 38672 111036
rect 39092 110756 39120 111574
rect 39276 111502 39304 113884
rect 39448 112176 39500 112182
rect 39448 112118 39500 112124
rect 39264 111496 39316 111502
rect 39264 111438 39316 111444
rect 39460 110756 39488 112118
rect 39816 111904 39868 111910
rect 39816 111846 39868 111852
rect 39828 110756 39856 111846
rect 40012 111434 40040 113884
rect 40276 111700 40328 111706
rect 40276 111642 40328 111648
rect 40000 111428 40052 111434
rect 40000 111370 40052 111376
rect 40288 110756 40316 111642
rect 40656 111366 40684 113884
rect 40644 111360 40696 111366
rect 40644 111302 40696 111308
rect 41012 111292 41064 111298
rect 41012 111234 41064 111240
rect 40644 111224 40696 111230
rect 40644 111166 40696 111172
rect 40656 110756 40684 111166
rect 41024 110756 41052 111234
rect 41300 111230 41328 113884
rect 41472 111564 41524 111570
rect 41472 111506 41524 111512
rect 41288 111224 41340 111230
rect 41288 111166 41340 111172
rect 41484 110756 41512 111506
rect 42036 111162 42064 113884
rect 42208 111496 42260 111502
rect 42208 111438 42260 111444
rect 42024 111156 42076 111162
rect 42024 111098 42076 111104
rect 41840 111088 41892 111094
rect 41840 111030 41892 111036
rect 41852 110756 41880 111030
rect 42220 110756 42248 111438
rect 42300 111428 42352 111434
rect 42300 111370 42352 111376
rect 42312 110770 42340 111370
rect 42680 111026 42708 113884
rect 43416 111366 43444 113884
rect 44074 113870 44364 113898
rect 44810 113870 45192 113898
rect 45454 113870 45744 113898
rect 43036 111360 43088 111366
rect 43036 111302 43088 111308
rect 43404 111360 43456 111366
rect 43404 111302 43456 111308
rect 42668 111020 42720 111026
rect 42668 110962 42720 110968
rect 42312 110742 42694 110770
rect 43048 110756 43076 111302
rect 44336 111230 44364 113870
rect 44600 111360 44652 111366
rect 44600 111302 44652 111308
rect 43404 111224 43456 111230
rect 43404 111166 43456 111172
rect 44324 111224 44376 111230
rect 44324 111166 44376 111172
rect 43416 110756 43444 111166
rect 43864 111156 43916 111162
rect 43864 111098 43916 111104
rect 43876 110756 43904 111098
rect 44232 111020 44284 111026
rect 44232 110962 44284 110968
rect 44244 110756 44272 110962
rect 44612 110756 44640 111302
rect 45060 111224 45112 111230
rect 45060 111166 45112 111172
rect 45072 110756 45100 111166
rect 45164 110770 45192 113870
rect 45716 112130 45744 113870
rect 45716 112102 45836 112130
rect 45164 110742 45454 110770
rect 45808 110756 45836 112102
rect 46084 110770 46112 113884
rect 46820 110770 46848 113884
rect 46084 110742 46282 110770
rect 46650 110742 46848 110770
rect 47188 113870 47478 113898
rect 47740 113870 48214 113898
rect 47188 110634 47216 113870
rect 47740 110770 47768 113870
rect 48280 111428 48332 111434
rect 48280 111370 48332 111376
rect 47820 111360 47872 111366
rect 47820 111302 47872 111308
rect 47478 110742 47768 110770
rect 47832 110756 47860 111302
rect 48292 110756 48320 111370
rect 48844 111366 48872 113884
rect 49488 111434 49516 113884
rect 49476 111428 49528 111434
rect 49476 111370 49528 111376
rect 48832 111360 48884 111366
rect 48832 111302 48884 111308
rect 49844 111360 49896 111366
rect 49844 111302 49896 111308
rect 48648 111292 48700 111298
rect 48648 111234 48700 111240
rect 48660 110756 48688 111234
rect 49476 111224 49528 111230
rect 49476 111166 49528 111172
rect 49016 111088 49068 111094
rect 49016 111030 49068 111036
rect 49028 110756 49056 111030
rect 49488 110756 49516 111166
rect 49856 110756 49884 111302
rect 50224 111298 50252 113884
rect 50672 111428 50724 111434
rect 50672 111370 50724 111376
rect 50212 111292 50264 111298
rect 50212 111234 50264 111240
rect 50212 111156 50264 111162
rect 50212 111098 50264 111104
rect 50224 110756 50252 111098
rect 50684 110756 50712 111370
rect 50868 111094 50896 113884
rect 51040 112108 51092 112114
rect 51040 112050 51092 112056
rect 50856 111088 50908 111094
rect 50856 111030 50908 111036
rect 51052 110756 51080 112050
rect 51408 111292 51460 111298
rect 51408 111234 51460 111240
rect 51420 110756 51448 111234
rect 51604 111230 51632 113884
rect 51868 111972 51920 111978
rect 51868 111914 51920 111920
rect 51592 111224 51644 111230
rect 51592 111166 51644 111172
rect 51880 110756 51908 111914
rect 52248 111366 52276 113884
rect 52604 112176 52656 112182
rect 52604 112118 52656 112124
rect 52512 111904 52564 111910
rect 52512 111846 52564 111852
rect 52236 111360 52288 111366
rect 52236 111302 52288 111308
rect 52524 110770 52552 111846
rect 52262 110742 52552 110770
rect 52616 110756 52644 112118
rect 52984 111162 53012 113884
rect 53064 112040 53116 112046
rect 53064 111982 53116 111988
rect 52972 111156 53024 111162
rect 52972 111098 53024 111104
rect 53076 110756 53104 111982
rect 53432 111700 53484 111706
rect 53432 111642 53484 111648
rect 53444 110756 53472 111642
rect 53628 111434 53656 113884
rect 54272 112114 54300 113884
rect 54260 112108 54312 112114
rect 54260 112050 54312 112056
rect 53800 111836 53852 111842
rect 53800 111778 53852 111784
rect 53616 111428 53668 111434
rect 53616 111370 53668 111376
rect 53812 110756 53840 111778
rect 54260 111768 54312 111774
rect 54260 111710 54312 111716
rect 54272 110756 54300 111710
rect 54628 111632 54680 111638
rect 54628 111574 54680 111580
rect 54640 110756 54668 111574
rect 55008 111298 55036 113884
rect 55652 111978 55680 113884
rect 55640 111972 55692 111978
rect 55640 111914 55692 111920
rect 56388 111910 56416 113884
rect 56926 113232 56982 113241
rect 56926 113167 56982 113176
rect 56376 111904 56428 111910
rect 56376 111846 56428 111852
rect 54996 111292 55048 111298
rect 54996 111234 55048 111240
rect 47110 110606 47216 110634
rect 31994 104256 32050 104265
rect 31994 104191 32050 104200
rect 37422 104256 37478 104265
rect 37422 104191 37478 104200
rect 37436 104090 37464 104191
rect 32640 104084 32692 104090
rect 32640 104026 32692 104032
rect 37424 104084 37476 104090
rect 37424 104026 37476 104032
rect 32652 90937 32680 104026
rect 32638 90928 32694 90937
rect 32638 90863 32694 90872
rect 36410 90928 36466 90937
rect 36410 90863 36466 90872
rect 36424 90286 36452 90863
rect 36412 90280 36464 90286
rect 36412 90222 36464 90228
rect 54812 86132 54864 86138
rect 54812 86074 54864 86080
rect 54824 86002 54852 86074
rect 54812 85996 54864 86002
rect 54812 85938 54864 85944
rect 56940 81961 56968 113167
rect 57032 112182 57060 113884
rect 57020 112176 57072 112182
rect 57020 112118 57072 112124
rect 57676 112046 57704 113884
rect 57664 112040 57716 112046
rect 57664 111982 57716 111988
rect 58412 111706 58440 113884
rect 59056 111842 59084 113884
rect 59044 111836 59096 111842
rect 59044 111778 59096 111784
rect 59792 111774 59820 113884
rect 59780 111768 59832 111774
rect 59780 111710 59832 111716
rect 58400 111700 58452 111706
rect 58400 111642 58452 111648
rect 60436 111638 60464 113884
rect 73224 113678 73252 115910
rect 82516 115910 82852 115938
rect 92728 115910 92880 115938
rect 73212 113672 73264 113678
rect 72842 113640 72898 113649
rect 73212 113614 73264 113620
rect 72842 113575 72898 113584
rect 60424 111632 60476 111638
rect 60424 111574 60476 111580
rect 72856 110756 72884 113575
rect 73224 113241 73252 113614
rect 73210 113232 73266 113241
rect 82516 113202 82544 115910
rect 92728 114358 92756 115910
rect 100626 115544 100682 115553
rect 100626 115479 100682 115488
rect 100640 115242 100668 115479
rect 100628 115236 100680 115242
rect 100628 115178 100680 115184
rect 102204 114737 102232 116606
rect 102296 116505 102324 117898
rect 102376 117820 102428 117826
rect 102376 117762 102428 117768
rect 102388 117593 102416 117762
rect 132656 117758 132684 118086
rect 132736 117956 132788 117962
rect 132736 117898 132788 117904
rect 132644 117752 132696 117758
rect 132644 117694 132696 117700
rect 132748 117638 132776 117898
rect 134116 117820 134168 117826
rect 134116 117762 134168 117768
rect 132656 117610 132776 117638
rect 102374 117584 102430 117593
rect 102374 117519 102430 117528
rect 102282 116496 102338 116505
rect 102282 116431 102338 116440
rect 102376 116460 102428 116466
rect 102376 116402 102428 116408
rect 102388 115281 102416 116402
rect 102468 116392 102520 116398
rect 102468 116334 102520 116340
rect 102480 115825 102508 116334
rect 102466 115816 102522 115825
rect 102466 115751 102522 115760
rect 102374 115272 102430 115281
rect 102284 115236 102336 115242
rect 102374 115207 102430 115216
rect 102284 115178 102336 115184
rect 102190 114728 102246 114737
rect 102190 114663 102246 114672
rect 92716 114352 92768 114358
rect 92716 114294 92768 114300
rect 102296 114193 102324 115178
rect 132656 115106 132684 117610
rect 134128 117321 134156 117762
rect 135232 117593 135260 119258
rect 135312 119112 135364 119118
rect 135310 119080 135312 119089
rect 135364 119080 135366 119089
rect 135310 119015 135366 119024
rect 136796 118710 136824 119831
rect 136888 119118 136916 120647
rect 172716 120647 172718 120656
rect 172664 120618 172716 120624
rect 172768 120546 172796 122030
rect 172860 121838 172888 123390
rect 173964 122897 173992 124834
rect 174056 124665 174084 126330
rect 174136 126116 174188 126122
rect 174136 126058 174188 126064
rect 174148 125209 174176 126058
rect 174228 126048 174280 126054
rect 174228 125990 174280 125996
rect 174240 125753 174268 125990
rect 174226 125744 174282 125753
rect 174226 125679 174282 125688
rect 174134 125200 174190 125209
rect 174134 125135 174190 125144
rect 204968 124778 204996 134354
rect 174228 124756 174280 124762
rect 204968 124750 205088 124778
rect 174228 124698 174280 124704
rect 174042 124656 174098 124665
rect 174042 124591 174098 124600
rect 174240 123441 174268 124698
rect 174226 123432 174282 123441
rect 174044 123396 174096 123402
rect 174226 123367 174282 123376
rect 174044 123338 174096 123344
rect 173950 122888 174006 122897
rect 173950 122823 174006 122832
rect 174056 122353 174084 123338
rect 172938 122344 172994 122353
rect 172938 122279 172994 122288
rect 174042 122344 174098 122353
rect 174042 122279 174098 122288
rect 172848 121832 172900 121838
rect 172848 121774 172900 121780
rect 172952 120614 172980 122279
rect 174136 121968 174188 121974
rect 174136 121910 174188 121916
rect 174148 121129 174176 121910
rect 174320 121832 174372 121838
rect 174320 121774 174372 121780
rect 174332 121673 174360 121774
rect 174318 121664 174374 121673
rect 174318 121599 174374 121608
rect 174134 121120 174190 121129
rect 174134 121055 174190 121064
rect 174044 120948 174096 120954
rect 174044 120890 174096 120896
rect 173952 120676 174004 120682
rect 173952 120618 174004 120624
rect 172940 120608 172992 120614
rect 172940 120550 172992 120556
rect 172756 120540 172808 120546
rect 172756 120482 172808 120488
rect 172662 119896 172718 119905
rect 172662 119831 172718 119840
rect 172676 119594 172704 119831
rect 172664 119588 172716 119594
rect 172664 119530 172716 119536
rect 136966 119352 137022 119361
rect 136966 119287 136968 119296
rect 137020 119287 137022 119296
rect 172662 119352 172718 119361
rect 172718 119310 172796 119338
rect 172662 119287 172718 119296
rect 136968 119258 137020 119264
rect 136876 119112 136928 119118
rect 136876 119054 136928 119060
rect 136784 118704 136836 118710
rect 136784 118646 136836 118652
rect 136966 118672 137022 118681
rect 136966 118607 137022 118616
rect 172018 118672 172074 118681
rect 172018 118607 172074 118616
rect 136782 118128 136838 118137
rect 136782 118063 136838 118072
rect 135312 117956 135364 117962
rect 135312 117898 135364 117904
rect 135218 117584 135274 117593
rect 135218 117519 135274 117528
rect 134114 117312 134170 117321
rect 134114 117247 134170 117256
rect 134668 117208 134720 117214
rect 134668 117150 134720 117156
rect 134680 116777 134708 117150
rect 134666 116768 134722 116777
rect 134666 116703 134722 116712
rect 135324 116233 135352 117898
rect 136796 117214 136824 118063
rect 136874 117992 136930 118001
rect 136874 117927 136876 117936
rect 136928 117927 136930 117936
rect 136876 117898 136928 117904
rect 136980 117894 137008 118607
rect 172032 117894 172060 118607
rect 172662 118128 172718 118137
rect 172662 118063 172664 118072
rect 172716 118063 172718 118072
rect 172664 118034 172716 118040
rect 172478 117992 172534 118001
rect 172478 117927 172534 117936
rect 136968 117888 137020 117894
rect 136968 117830 137020 117836
rect 172020 117888 172072 117894
rect 172020 117830 172072 117836
rect 136784 117208 136836 117214
rect 136784 117150 136836 117156
rect 136782 116904 136838 116913
rect 136782 116839 136838 116848
rect 135310 116224 135366 116233
rect 135310 116159 135366 116168
rect 136796 115786 136824 116839
rect 136874 116496 136930 116505
rect 136874 116431 136930 116440
rect 134484 115780 134536 115786
rect 134484 115722 134536 115728
rect 136784 115780 136836 115786
rect 136784 115722 136836 115728
rect 134496 115553 134524 115722
rect 134482 115544 134538 115553
rect 134482 115479 134538 115488
rect 136782 115544 136838 115553
rect 136782 115479 136838 115488
rect 132644 115100 132696 115106
rect 132644 115042 132696 115048
rect 135312 115032 135364 115038
rect 135310 115000 135312 115009
rect 135364 115000 135366 115009
rect 135310 114935 135366 114944
rect 136796 114494 136824 115479
rect 136888 115038 136916 116431
rect 172492 116398 172520 117927
rect 172768 117826 172796 119310
rect 173964 118817 173992 120618
rect 174056 120426 174084 120890
rect 174136 120608 174188 120614
rect 174134 120576 174136 120585
rect 174188 120576 174190 120585
rect 174134 120511 174190 120520
rect 174320 120540 174372 120546
rect 174320 120482 174372 120488
rect 174056 120398 174176 120426
rect 174044 119588 174096 119594
rect 174044 119530 174096 119536
rect 173950 118808 174006 118817
rect 173950 118743 174006 118752
rect 174056 118273 174084 119530
rect 174148 119361 174176 120398
rect 174332 119905 174360 120482
rect 174318 119896 174374 119905
rect 174318 119831 174374 119840
rect 174134 119352 174190 119361
rect 174134 119287 174190 119296
rect 174042 118264 174098 118273
rect 174042 118199 174098 118208
rect 173952 118092 174004 118098
rect 173952 118034 174004 118040
rect 172756 117820 172808 117826
rect 172756 117762 172808 117768
rect 172662 116904 172718 116913
rect 172662 116839 172718 116848
rect 172572 116596 172624 116602
rect 172572 116538 172624 116544
rect 172584 116505 172612 116538
rect 172676 116534 172704 116839
rect 173860 116596 173912 116602
rect 173860 116538 173912 116544
rect 172664 116528 172716 116534
rect 172570 116496 172626 116505
rect 172664 116470 172716 116476
rect 172570 116431 172626 116440
rect 172480 116392 172532 116398
rect 172480 116334 172532 116340
rect 144892 115174 144920 115924
rect 144880 115168 144932 115174
rect 144880 115110 144932 115116
rect 136876 115032 136928 115038
rect 136876 114974 136928 114980
rect 144892 114970 144920 115110
rect 144880 114964 144932 114970
rect 144880 114906 144932 114912
rect 134852 114488 134904 114494
rect 134850 114456 134852 114465
rect 136784 114488 136836 114494
rect 134904 114456 134906 114465
rect 136784 114430 136836 114436
rect 134850 114391 134906 114400
rect 102282 114184 102338 114193
rect 102282 114119 102338 114128
rect 105102 113626 105130 113884
rect 105562 113626 105590 113884
rect 106114 113626 106142 113884
rect 106666 113626 106694 113884
rect 107218 113626 107246 113884
rect 107770 113626 107798 113884
rect 108322 113626 108350 113884
rect 108874 113626 108902 113884
rect 109426 113762 109454 113884
rect 109426 113734 109500 113762
rect 109472 113678 109500 113734
rect 105102 113598 105176 113626
rect 105562 113598 105636 113626
rect 106114 113598 106188 113626
rect 73210 113167 73266 113176
rect 81676 113196 81728 113202
rect 81676 113138 81728 113144
rect 82504 113196 82556 113202
rect 82504 113138 82556 113144
rect 81688 112318 81716 113138
rect 92806 112688 92862 112697
rect 92806 112623 92862 112632
rect 81676 112312 81728 112318
rect 81676 112254 81728 112260
rect 92820 110756 92848 112623
rect 60514 104256 60570 104265
rect 60514 104191 60570 104200
rect 60528 101030 60556 104191
rect 105148 101681 105176 113598
rect 105228 111224 105280 111230
rect 105228 111166 105280 111172
rect 105240 105353 105268 111166
rect 105504 111156 105556 111162
rect 105504 111098 105556 111104
rect 105516 106577 105544 111098
rect 105502 106568 105558 106577
rect 105502 106503 105558 106512
rect 105226 105344 105282 105353
rect 105226 105279 105282 105288
rect 105608 102905 105636 113598
rect 105688 111088 105740 111094
rect 105688 111030 105740 111036
rect 105700 107801 105728 111030
rect 105964 110952 106016 110958
rect 105964 110894 106016 110900
rect 105976 110249 106004 110894
rect 105962 110240 106018 110249
rect 105962 110175 106018 110184
rect 105780 109524 105832 109530
rect 105780 109466 105832 109472
rect 105792 109025 105820 109466
rect 105778 109016 105834 109025
rect 105778 108951 105834 108960
rect 105686 107792 105742 107801
rect 105686 107727 105742 107736
rect 106160 104129 106188 113598
rect 106620 113598 106694 113626
rect 107172 113598 107246 113626
rect 107724 113598 107798 113626
rect 108276 113598 108350 113626
rect 108828 113598 108902 113626
rect 109460 113672 109512 113678
rect 109460 113614 109512 113620
rect 109978 113626 110006 113884
rect 110530 113626 110558 113884
rect 106620 111230 106648 113598
rect 106608 111224 106660 111230
rect 106608 111166 106660 111172
rect 107172 111162 107200 113598
rect 107160 111156 107212 111162
rect 107160 111098 107212 111104
rect 107724 111094 107752 113598
rect 107712 111088 107764 111094
rect 107712 111030 107764 111036
rect 108276 109530 108304 113598
rect 108828 111026 108856 113598
rect 109472 112250 109500 113614
rect 109978 113598 110052 113626
rect 109460 112244 109512 112250
rect 109460 112186 109512 112192
rect 110024 112182 110052 113598
rect 110484 113598 110558 113626
rect 111082 113626 111110 113884
rect 111634 113626 111662 113884
rect 112186 113626 112214 113884
rect 112738 113626 112766 113884
rect 113290 113626 113318 113884
rect 111082 113598 111156 113626
rect 110484 112318 110512 113598
rect 110472 112312 110524 112318
rect 110472 112254 110524 112260
rect 110012 112176 110064 112182
rect 110012 112118 110064 112124
rect 108816 111020 108868 111026
rect 108816 110962 108868 110968
rect 111128 110756 111156 113598
rect 111588 113598 111662 113626
rect 112140 113598 112214 113626
rect 112600 113598 112766 113626
rect 112968 113598 113318 113626
rect 113508 113672 113560 113678
rect 113842 113626 113870 113884
rect 114394 113678 114422 113884
rect 113508 113614 113560 113620
rect 111588 110770 111616 113598
rect 112140 110770 112168 113598
rect 112600 110770 112628 113598
rect 112968 110770 112996 113598
rect 113048 112380 113100 112386
rect 113048 112322 113100 112328
rect 111510 110742 111616 110770
rect 111878 110742 112168 110770
rect 112338 110742 112628 110770
rect 112706 110742 112996 110770
rect 113060 110756 113088 112322
rect 113520 110756 113548 113614
rect 113796 113598 113870 113626
rect 114382 113672 114434 113678
rect 114382 113614 114434 113620
rect 114520 113672 114572 113678
rect 114946 113626 114974 113884
rect 115498 113678 115526 113884
rect 114520 113614 114572 113620
rect 113796 112386 113824 113598
rect 113876 113128 113928 113134
rect 113876 113070 113928 113076
rect 113784 112380 113836 112386
rect 113784 112322 113836 112328
rect 113888 110756 113916 113070
rect 114532 110770 114560 113614
rect 114900 113598 114974 113626
rect 115486 113672 115538 113678
rect 116050 113626 116078 113884
rect 116602 113762 116630 113884
rect 115486 113614 115538 113620
rect 116004 113598 116078 113626
rect 116556 113734 116630 113762
rect 114900 113134 114928 113598
rect 114888 113128 114940 113134
rect 114888 113070 114940 113076
rect 115072 113128 115124 113134
rect 115072 113070 115124 113076
rect 114704 112924 114756 112930
rect 114704 112866 114756 112872
rect 114270 110742 114560 110770
rect 114716 110756 114744 112866
rect 115084 110756 115112 113070
rect 115440 113060 115492 113066
rect 115440 113002 115492 113008
rect 115452 110756 115480 113002
rect 116004 112930 116032 113598
rect 116268 113196 116320 113202
rect 116268 113138 116320 113144
rect 115992 112924 116044 112930
rect 115992 112866 116044 112872
rect 115912 112340 116216 112368
rect 115912 110756 115940 112340
rect 116188 112114 116216 112340
rect 116176 112108 116228 112114
rect 116176 112050 116228 112056
rect 116280 110756 116308 113138
rect 116556 113134 116584 113734
rect 116636 113672 116688 113678
rect 117154 113626 117182 113884
rect 117706 113626 117734 113884
rect 118258 113626 118286 113884
rect 118810 113678 118838 113884
rect 116636 113614 116688 113620
rect 116544 113128 116596 113134
rect 116544 113070 116596 113076
rect 116648 110756 116676 113614
rect 117108 113598 117182 113626
rect 117660 113598 117734 113626
rect 118212 113598 118286 113626
rect 118798 113672 118850 113678
rect 119270 113626 119298 113884
rect 119822 113626 119850 113884
rect 118798 113614 118850 113620
rect 119224 113598 119298 113626
rect 119776 113598 119850 113626
rect 120132 113672 120184 113678
rect 120374 113626 120402 113884
rect 120926 113626 120954 113884
rect 121478 113626 121506 113884
rect 122030 113626 122058 113884
rect 122582 113626 122610 113884
rect 123134 113678 123162 113884
rect 120132 113614 120184 113620
rect 117108 113066 117136 113598
rect 117096 113060 117148 113066
rect 117096 113002 117148 113008
rect 117660 112114 117688 113598
rect 118212 113202 118240 113598
rect 118200 113196 118252 113202
rect 118200 113138 118252 113144
rect 117832 112788 117884 112794
rect 117832 112730 117884 112736
rect 117648 112108 117700 112114
rect 117648 112050 117700 112056
rect 117464 111428 117516 111434
rect 117464 111370 117516 111376
rect 117372 111360 117424 111366
rect 117372 111302 117424 111308
rect 117384 110770 117412 111302
rect 117122 110742 117412 110770
rect 117476 110756 117504 111370
rect 117844 110756 117872 112730
rect 119120 112380 119172 112386
rect 119120 112322 119172 112328
rect 118844 111496 118896 111502
rect 118844 111438 118896 111444
rect 118568 111292 118620 111298
rect 118568 111234 118620 111240
rect 118580 110770 118608 111234
rect 118856 110770 118884 111438
rect 118318 110742 118608 110770
rect 118686 110742 118884 110770
rect 119132 110756 119160 112322
rect 119224 111366 119252 113598
rect 119776 111434 119804 113598
rect 119764 111428 119816 111434
rect 119764 111370 119816 111376
rect 119212 111360 119264 111366
rect 119212 111302 119264 111308
rect 119764 111224 119816 111230
rect 119764 111166 119816 111172
rect 119776 110770 119804 111166
rect 120144 110770 120172 113614
rect 120236 113598 120402 113626
rect 120880 113598 120954 113626
rect 121432 113598 121506 113626
rect 121984 113598 122058 113626
rect 122536 113598 122610 113626
rect 123122 113672 123174 113678
rect 123122 113614 123174 113620
rect 122708 113604 122760 113610
rect 120236 112794 120264 113598
rect 120224 112788 120276 112794
rect 120224 112730 120276 112736
rect 120316 112448 120368 112454
rect 120316 112390 120368 112396
rect 119514 110742 119804 110770
rect 119882 110742 120172 110770
rect 120328 110756 120356 112390
rect 120880 111298 120908 113598
rect 121052 112516 121104 112522
rect 121052 112458 121104 112464
rect 120960 112108 121012 112114
rect 120960 112050 121012 112056
rect 120868 111292 120920 111298
rect 120868 111234 120920 111240
rect 120972 110770 121000 112050
rect 120710 110742 121000 110770
rect 121064 110756 121092 112458
rect 121432 111502 121460 113598
rect 121880 113128 121932 113134
rect 121880 113070 121932 113076
rect 121512 112584 121564 112590
rect 121512 112526 121564 112532
rect 121420 111496 121472 111502
rect 121420 111438 121472 111444
rect 121524 110756 121552 112526
rect 121892 110756 121920 113070
rect 121984 112318 122012 113598
rect 122248 113264 122300 113270
rect 122248 113206 122300 113212
rect 121972 112312 122024 112318
rect 121972 112254 122024 112260
rect 122260 110756 122288 113206
rect 122536 111230 122564 113598
rect 123686 113592 123714 113884
rect 124238 113592 124266 113884
rect 124790 113592 124818 113884
rect 125342 113592 125370 113884
rect 125894 113592 125922 113884
rect 126296 113672 126348 113678
rect 126296 113614 126348 113620
rect 122708 113546 122760 113552
rect 123640 113564 123714 113592
rect 124192 113564 124266 113592
rect 124744 113564 124818 113592
rect 125296 113564 125370 113592
rect 125848 113564 125922 113592
rect 122524 111224 122576 111230
rect 122524 111166 122576 111172
rect 122720 110756 122748 113546
rect 123076 113468 123128 113474
rect 123076 113410 123128 113416
rect 123088 110756 123116 113410
rect 123444 112856 123496 112862
rect 123444 112798 123496 112804
rect 123456 110756 123484 112798
rect 123640 112318 123668 113564
rect 123904 113400 123956 113406
rect 123904 113342 123956 113348
rect 123628 112312 123680 112318
rect 123628 112254 123680 112260
rect 123916 110756 123944 113342
rect 124192 112114 124220 113564
rect 124640 113332 124692 113338
rect 124640 113274 124692 113280
rect 124272 112924 124324 112930
rect 124272 112866 124324 112872
rect 124180 112108 124232 112114
rect 124180 112050 124232 112056
rect 124284 110756 124312 112866
rect 124652 110756 124680 113274
rect 124744 112522 124772 113564
rect 125100 113060 125152 113066
rect 125100 113002 125152 113008
rect 124732 112516 124784 112522
rect 124732 112458 124784 112464
rect 125112 110756 125140 113002
rect 125296 112590 125324 113564
rect 125468 113196 125520 113202
rect 125468 113138 125520 113144
rect 125284 112584 125336 112590
rect 125284 112526 125336 112532
rect 125480 110756 125508 113138
rect 125848 113134 125876 113564
rect 125836 113128 125888 113134
rect 125836 113070 125888 113076
rect 125836 112992 125888 112998
rect 125836 112934 125888 112940
rect 125848 110756 125876 112934
rect 126308 110756 126336 113614
rect 126446 113592 126474 113884
rect 126998 113762 127026 113884
rect 126998 113734 127072 113762
rect 127044 113610 127072 113734
rect 126400 113564 126474 113592
rect 127032 113604 127084 113610
rect 126400 113270 126428 113564
rect 127550 113592 127578 113884
rect 128102 113592 128130 113884
rect 128654 113626 128682 113884
rect 129206 113626 129234 113884
rect 129758 113626 129786 113884
rect 130310 113626 130338 113884
rect 130862 113626 130890 113884
rect 131414 113626 131442 113884
rect 131966 113678 131994 113884
rect 132532 113870 132592 113898
rect 132092 113808 132144 113814
rect 132092 113750 132144 113756
rect 127032 113546 127084 113552
rect 127504 113564 127578 113592
rect 128056 113564 128130 113592
rect 128608 113598 128682 113626
rect 129160 113598 129234 113626
rect 129712 113598 129786 113626
rect 130264 113598 130338 113626
rect 130816 113598 130890 113626
rect 131368 113598 131442 113626
rect 131954 113672 132006 113678
rect 131954 113614 132006 113620
rect 127504 113474 127532 113564
rect 127492 113468 127544 113474
rect 127492 113410 127544 113416
rect 126388 113264 126440 113270
rect 126388 113206 126440 113212
rect 128056 112862 128084 113564
rect 128608 113406 128636 113598
rect 128596 113400 128648 113406
rect 128596 113342 128648 113348
rect 129160 112930 129188 113598
rect 129712 113338 129740 113598
rect 129700 113332 129752 113338
rect 129700 113274 129752 113280
rect 130264 113066 130292 113598
rect 130816 113202 130844 113598
rect 130804 113196 130856 113202
rect 130804 113138 130856 113144
rect 130252 113060 130304 113066
rect 130252 113002 130304 113008
rect 131368 112998 131396 113598
rect 131356 112992 131408 112998
rect 131356 112934 131408 112940
rect 129148 112924 129200 112930
rect 129148 112866 129200 112872
rect 128044 112856 128096 112862
rect 128044 112798 128096 112804
rect 126664 112788 126716 112794
rect 126664 112730 126716 112736
rect 126676 110756 126704 112730
rect 108630 109560 108686 109569
rect 108264 109524 108316 109530
rect 108630 109495 108686 109504
rect 108264 109466 108316 109472
rect 108538 107248 108594 107257
rect 108538 107183 108594 107192
rect 107894 104936 107950 104945
rect 107894 104871 107950 104880
rect 106146 104120 106202 104129
rect 105688 104084 105740 104090
rect 107908 104090 107936 104871
rect 106146 104055 106202 104064
rect 107896 104084 107948 104090
rect 105688 104026 105740 104032
rect 107896 104026 107948 104032
rect 105594 102896 105650 102905
rect 105594 102831 105650 102840
rect 105134 101672 105190 101681
rect 105134 101607 105190 101616
rect 57572 101024 57624 101030
rect 57572 100966 57624 100972
rect 60516 101024 60568 101030
rect 60516 100966 60568 100972
rect 57584 100865 57612 100966
rect 57570 100856 57626 100865
rect 57570 100791 57626 100800
rect 105596 99460 105648 99466
rect 105596 99402 105648 99408
rect 105608 99233 105636 99402
rect 105594 99224 105650 99233
rect 105594 99159 105650 99168
rect 105700 98145 105728 104026
rect 107894 102488 107950 102497
rect 107894 102423 107950 102432
rect 107908 101370 107936 102423
rect 106332 101364 106384 101370
rect 106332 101306 106384 101312
rect 107896 101364 107948 101370
rect 107896 101306 107948 101312
rect 105964 100820 106016 100826
rect 105964 100762 106016 100768
rect 105976 100457 106004 100762
rect 105962 100448 106018 100457
rect 105962 100383 106018 100392
rect 105686 98136 105742 98145
rect 105686 98071 105742 98080
rect 105780 97216 105832 97222
rect 105780 97158 105832 97164
rect 105792 94473 105820 97158
rect 106344 96921 106372 101306
rect 107894 100176 107950 100185
rect 107894 100111 107950 100120
rect 107908 99942 107936 100111
rect 106424 99936 106476 99942
rect 106424 99878 106476 99884
rect 107896 99936 107948 99942
rect 107896 99878 107948 99884
rect 106330 96912 106386 96921
rect 106330 96847 106386 96856
rect 106436 95697 106464 99878
rect 108552 99466 108580 107183
rect 108644 100826 108672 109495
rect 108632 100820 108684 100826
rect 108632 100762 108684 100768
rect 108540 99460 108592 99466
rect 108540 99402 108592 99408
rect 107894 97864 107950 97873
rect 107894 97799 107950 97808
rect 107908 97222 107936 97799
rect 107896 97216 107948 97222
rect 107896 97158 107948 97164
rect 106422 95688 106478 95697
rect 106422 95623 106478 95632
rect 107802 95416 107858 95425
rect 107802 95351 107858 95360
rect 105778 94464 105834 94473
rect 105778 94399 105834 94408
rect 107816 94366 107844 95351
rect 105780 94360 105832 94366
rect 105780 94302 105832 94308
rect 107804 94360 107856 94366
rect 107804 94302 107856 94308
rect 105792 93249 105820 94302
rect 105778 93240 105834 93249
rect 105778 93175 105834 93184
rect 107802 93104 107858 93113
rect 107802 93039 107858 93048
rect 107816 92122 107844 93039
rect 105228 92116 105280 92122
rect 105228 92058 105280 92064
rect 107804 92116 107856 92122
rect 107804 92058 107856 92064
rect 105240 92025 105268 92058
rect 105226 92016 105282 92025
rect 105226 91951 105282 91960
rect 59594 90928 59650 90937
rect 59594 90863 59650 90872
rect 59608 90286 59636 90863
rect 59596 90280 59648 90286
rect 59596 90222 59648 90228
rect 105778 89296 105834 89305
rect 105778 89231 105780 89240
rect 105832 89231 105834 89240
rect 107804 89260 107856 89266
rect 105780 89202 105832 89208
rect 107804 89202 107856 89208
rect 107816 88489 107844 89202
rect 107802 88480 107858 88489
rect 107802 88415 107858 88424
rect 105410 87936 105466 87945
rect 105410 87871 105412 87880
rect 105464 87871 105466 87880
rect 107896 87900 107948 87906
rect 105412 87842 105464 87848
rect 107896 87842 107948 87848
rect 106422 86576 106478 86585
rect 106422 86511 106478 86520
rect 106436 86410 106464 86511
rect 106424 86404 106476 86410
rect 106424 86346 106476 86352
rect 107908 86041 107936 87842
rect 107988 86404 108040 86410
rect 107988 86346 108040 86352
rect 107894 86032 107950 86041
rect 107894 85967 107950 85976
rect 105134 85352 105190 85361
rect 105134 85287 105190 85296
rect 105148 84846 105176 85287
rect 105136 84840 105188 84846
rect 107804 84840 107856 84846
rect 105136 84782 105188 84788
rect 105686 84808 105742 84817
rect 107804 84782 107856 84788
rect 105686 84743 105688 84752
rect 105740 84743 105742 84752
rect 107620 84772 107672 84778
rect 105688 84714 105740 84720
rect 107620 84714 107672 84720
rect 105226 83448 105282 83457
rect 105226 83383 105228 83392
rect 105280 83383 105282 83392
rect 105228 83354 105280 83360
rect 106422 82224 106478 82233
rect 106422 82159 106424 82168
rect 106476 82159 106478 82168
rect 106424 82130 106476 82136
rect 56926 81952 56982 81961
rect 56926 81887 56982 81896
rect 57478 81952 57534 81961
rect 57478 81887 57534 81896
rect 57492 80873 57520 81887
rect 57478 80864 57534 80873
rect 57478 80799 57534 80808
rect 105962 80864 106018 80873
rect 105962 80799 105964 80808
rect 30524 77836 30576 77842
rect 30524 77778 30576 77784
rect 37424 77836 37476 77842
rect 37424 77778 37476 77784
rect 37436 77609 37464 77778
rect 57492 77638 57520 80799
rect 106016 80799 106018 80808
rect 105964 80770 106016 80776
rect 105410 79640 105466 79649
rect 105410 79575 105466 79584
rect 105424 79270 105452 79575
rect 105412 79264 105464 79270
rect 105412 79206 105464 79212
rect 107632 78969 107660 84714
rect 107712 83412 107764 83418
rect 107712 83354 107764 83360
rect 107618 78960 107674 78969
rect 107618 78895 107674 78904
rect 105226 78008 105282 78017
rect 105226 77943 105282 77952
rect 105240 77910 105268 77943
rect 105228 77904 105280 77910
rect 105228 77846 105280 77852
rect 107528 77904 107580 77910
rect 107528 77846 107580 77852
rect 57480 77632 57532 77638
rect 31994 77600 32050 77609
rect 31994 77535 32050 77544
rect 37422 77600 37478 77609
rect 59596 77632 59648 77638
rect 57480 77574 57532 77580
rect 59594 77600 59596 77609
rect 59648 77600 59650 77609
rect 37422 77535 37478 77544
rect 28684 69540 28736 69546
rect 28684 69482 28736 69488
rect 31904 69472 31956 69478
rect 31902 69440 31904 69449
rect 31956 69440 31958 69449
rect 31902 69375 31958 69384
rect 27580 69336 27632 69342
rect 27580 69278 27632 69284
rect 32008 67658 32036 77535
rect 54996 76476 55048 76482
rect 54996 76418 55048 76424
rect 36044 69540 36096 69546
rect 36044 69482 36096 69488
rect 35584 69472 35636 69478
rect 35584 69414 35636 69420
rect 34664 69404 34716 69410
rect 34664 69346 34716 69352
rect 34112 69132 34164 69138
rect 34112 69074 34164 69080
rect 32008 67630 32956 67658
rect 32928 67522 32956 67630
rect 34124 67522 34152 69074
rect 34676 67522 34704 69346
rect 35596 67522 35624 69414
rect 36056 67522 36084 69482
rect 39092 69138 39120 70908
rect 39264 69608 39316 69614
rect 39264 69550 39316 69556
rect 39080 69132 39132 69138
rect 39080 69074 39132 69080
rect 36596 69064 36648 69070
rect 36596 69006 36648 69012
rect 32928 67494 33218 67522
rect 33862 67494 34152 67522
rect 34506 67494 34704 67522
rect 35242 67494 35624 67522
rect 35886 67494 36084 67522
rect 36608 67508 36636 69006
rect 37240 68996 37292 69002
rect 37240 68938 37292 68944
rect 37252 67508 37280 68938
rect 38620 68860 38672 68866
rect 38620 68802 38672 68808
rect 37884 68792 37936 68798
rect 37884 68734 37936 68740
rect 37896 67508 37924 68734
rect 38632 67508 38660 68802
rect 39276 67508 39304 69550
rect 39460 69410 39488 70908
rect 39828 69478 39856 70908
rect 40288 69546 40316 70908
rect 40380 70894 40670 70922
rect 40276 69540 40328 69546
rect 40276 69482 40328 69488
rect 39816 69472 39868 69478
rect 39816 69414 39868 69420
rect 39448 69404 39500 69410
rect 39448 69346 39500 69352
rect 40184 69200 40236 69206
rect 40184 69142 40236 69148
rect 40196 67522 40224 69142
rect 40380 69070 40408 70894
rect 40644 69132 40696 69138
rect 40644 69074 40696 69080
rect 40368 69064 40420 69070
rect 40368 69006 40420 69012
rect 40026 67494 40224 67522
rect 40656 67508 40684 69074
rect 41024 69002 41052 70908
rect 41012 68996 41064 69002
rect 41012 68938 41064 68944
rect 41288 68928 41340 68934
rect 41288 68870 41340 68876
rect 41300 67508 41328 68870
rect 41484 68798 41512 70908
rect 41852 68866 41880 70908
rect 42220 69546 42248 70908
rect 42208 69540 42260 69546
rect 42208 69482 42260 69488
rect 42680 69206 42708 70908
rect 42668 69200 42720 69206
rect 42668 69142 42720 69148
rect 43048 69138 43076 70908
rect 43036 69132 43088 69138
rect 43036 69074 43088 69080
rect 42024 69064 42076 69070
rect 42024 69006 42076 69012
rect 41840 68860 41892 68866
rect 41840 68802 41892 68808
rect 41472 68792 41524 68798
rect 41472 68734 41524 68740
rect 42036 67508 42064 69006
rect 42668 68996 42720 69002
rect 42668 68938 42720 68944
rect 42680 67508 42708 68938
rect 43416 68934 43444 70908
rect 43876 69070 43904 70908
rect 43864 69064 43916 69070
rect 43864 69006 43916 69012
rect 44244 69002 44272 70908
rect 44232 68996 44284 69002
rect 44232 68938 44284 68944
rect 43404 68928 43456 68934
rect 43404 68870 43456 68876
rect 44612 68730 44640 70908
rect 44704 70894 45086 70922
rect 45164 70894 45454 70922
rect 45716 70894 45822 70922
rect 43404 68724 43456 68730
rect 43404 68666 43456 68672
rect 44600 68724 44652 68730
rect 44600 68666 44652 68672
rect 43416 67508 43444 68666
rect 44704 68338 44732 70894
rect 44336 68310 44732 68338
rect 44336 67522 44364 68310
rect 45164 67522 45192 70894
rect 45716 67522 45744 70894
rect 46268 67522 46296 70908
rect 44074 67494 44364 67522
rect 44810 67494 45192 67522
rect 45454 67494 45744 67522
rect 46098 67494 46296 67522
rect 46636 67522 46664 70908
rect 47110 70894 47308 70922
rect 47478 70894 47768 70922
rect 47280 67522 47308 70894
rect 47740 67522 47768 70894
rect 47832 69614 47860 70908
rect 48292 69682 48320 70908
rect 48660 69750 48688 70908
rect 48648 69744 48700 69750
rect 48648 69686 48700 69692
rect 48280 69676 48332 69682
rect 48280 69618 48332 69624
rect 49028 69614 49056 70908
rect 49488 69818 49516 70908
rect 49476 69812 49528 69818
rect 49476 69754 49528 69760
rect 49856 69682 49884 70908
rect 50238 70894 50528 70922
rect 50212 69744 50264 69750
rect 50212 69686 50264 69692
rect 49476 69676 49528 69682
rect 49476 69618 49528 69624
rect 49844 69676 49896 69682
rect 49844 69618 49896 69624
rect 47820 69608 47872 69614
rect 47820 69550 47872 69556
rect 48832 69608 48884 69614
rect 48832 69550 48884 69556
rect 49016 69608 49068 69614
rect 49016 69550 49068 69556
rect 46636 67494 46834 67522
rect 47280 67494 47478 67522
rect 47740 67494 48214 67522
rect 48844 67508 48872 69550
rect 49488 67508 49516 69618
rect 50224 67508 50252 69686
rect 50500 68730 50528 70894
rect 50684 68934 50712 70908
rect 50856 69608 50908 69614
rect 50856 69550 50908 69556
rect 50672 68928 50724 68934
rect 50672 68870 50724 68876
rect 50488 68724 50540 68730
rect 50488 68666 50540 68672
rect 50868 67508 50896 69550
rect 51052 68866 51080 70908
rect 51040 68860 51092 68866
rect 51040 68802 51092 68808
rect 51420 68798 51448 70908
rect 51592 69812 51644 69818
rect 51592 69754 51644 69760
rect 51408 68792 51460 68798
rect 51408 68734 51460 68740
rect 51604 67508 51632 69754
rect 51880 69342 51908 70908
rect 52262 70894 52552 70922
rect 52236 69676 52288 69682
rect 52236 69618 52288 69624
rect 51868 69336 51920 69342
rect 51868 69278 51920 69284
rect 52248 67508 52276 69618
rect 52524 69002 52552 70894
rect 52616 69138 52644 70908
rect 52604 69132 52656 69138
rect 52604 69074 52656 69080
rect 53076 69070 53104 70908
rect 53444 69478 53472 70908
rect 53812 69546 53840 70908
rect 53800 69540 53852 69546
rect 53800 69482 53852 69488
rect 53432 69472 53484 69478
rect 53432 69414 53484 69420
rect 53064 69064 53116 69070
rect 53064 69006 53116 69012
rect 54272 69002 54300 70908
rect 54640 69206 54668 70908
rect 55008 69614 55036 76418
rect 54996 69608 55048 69614
rect 54996 69550 55048 69556
rect 57492 69410 57520 77574
rect 59594 77535 59650 77544
rect 106974 76784 107030 76793
rect 106974 76719 107030 76728
rect 105962 75560 106018 75569
rect 105962 75495 106018 75504
rect 105410 74336 105466 74345
rect 105410 74271 105466 74280
rect 105226 73792 105282 73801
rect 105226 73727 105282 73736
rect 101362 71208 101418 71217
rect 101206 71180 101362 71194
rect 101192 71166 101362 71180
rect 59044 69608 59096 69614
rect 59044 69550 59096 69556
rect 58124 69472 58176 69478
rect 58176 69420 58256 69426
rect 58124 69414 58256 69420
rect 57480 69404 57532 69410
rect 58136 69398 58256 69414
rect 57480 69346 57532 69352
rect 54628 69200 54680 69206
rect 54628 69142 54680 69148
rect 56744 69132 56796 69138
rect 56744 69074 56796 69080
rect 56756 69018 56784 69074
rect 57664 69064 57716 69070
rect 52512 68996 52564 69002
rect 52512 68938 52564 68944
rect 54260 68996 54312 69002
rect 56756 68990 56876 69018
rect 57664 69006 57716 69012
rect 54260 68938 54312 68944
rect 53616 68928 53668 68934
rect 53616 68870 53668 68876
rect 52972 68724 53024 68730
rect 52972 68666 53024 68672
rect 52984 67508 53012 68666
rect 53628 67508 53656 68870
rect 54260 68860 54312 68866
rect 54260 68802 54312 68808
rect 55640 68860 55692 68866
rect 55640 68802 55692 68808
rect 54272 67508 54300 68802
rect 54996 68792 55048 68798
rect 54996 68734 55048 68740
rect 55008 67508 55036 68734
rect 55652 67508 55680 68802
rect 56376 68792 56428 68798
rect 56376 68734 56428 68740
rect 56388 67508 56416 68734
rect 56848 67522 56876 68990
rect 56848 67494 57046 67522
rect 57676 67508 57704 69006
rect 58228 67522 58256 69398
rect 58228 67494 58426 67522
rect 59056 67508 59084 69550
rect 60148 69200 60200 69206
rect 60148 69142 60200 69148
rect 59504 68996 59556 69002
rect 59504 68938 59556 68944
rect 59516 68882 59544 68938
rect 59516 68854 59636 68882
rect 59608 67522 59636 68854
rect 60160 67522 60188 69142
rect 62908 68996 62960 69002
rect 62908 68938 62960 68944
rect 62724 68860 62776 68866
rect 62724 68802 62776 68808
rect 62356 68248 62408 68254
rect 62356 68190 62408 68196
rect 59608 67494 59806 67522
rect 60160 67494 60450 67522
rect 62368 63329 62396 68190
rect 62736 66185 62764 68802
rect 62816 66752 62868 66758
rect 62814 66720 62816 66729
rect 62868 66720 62870 66729
rect 62814 66655 62870 66664
rect 62722 66176 62778 66185
rect 62722 66111 62778 66120
rect 62920 65641 62948 68938
rect 63000 68316 63052 68322
rect 63000 68258 63052 68264
rect 62906 65632 62962 65641
rect 62906 65567 62962 65576
rect 62816 65392 62868 65398
rect 62816 65334 62868 65340
rect 62724 65324 62776 65330
rect 62724 65266 62776 65272
rect 62736 64417 62764 65266
rect 62828 64961 62856 65334
rect 62814 64952 62870 64961
rect 62814 64887 62870 64896
rect 62722 64408 62778 64417
rect 62722 64343 62778 64352
rect 63012 63873 63040 68258
rect 63472 68254 63500 70908
rect 64576 68322 64604 70908
rect 64564 68316 64616 68322
rect 64564 68258 64616 68264
rect 63460 68248 63512 68254
rect 63460 68190 63512 68196
rect 63368 68180 63420 68186
rect 63368 68122 63420 68128
rect 63380 67273 63408 68122
rect 63366 67264 63422 67273
rect 63366 67199 63422 67208
rect 63368 65596 63420 65602
rect 63368 65538 63420 65544
rect 62998 63864 63054 63873
rect 62998 63799 63054 63808
rect 62354 63320 62410 63329
rect 62354 63255 62410 63264
rect 12030 62912 12086 62921
rect 12030 62847 12086 62856
rect 29234 62912 29290 62921
rect 29234 62847 29290 62856
rect 29248 62678 29276 62847
rect 63380 62785 63408 65538
rect 65680 65330 65708 70908
rect 66508 70894 66798 70922
rect 66508 68202 66536 70894
rect 67888 69002 67916 70908
rect 67876 68996 67928 69002
rect 67876 68938 67928 68944
rect 68992 68866 69020 70908
rect 68980 68860 69032 68866
rect 68980 68802 69032 68808
rect 66324 68174 66536 68202
rect 69164 68248 69216 68254
rect 69164 68190 69216 68196
rect 66324 65398 66352 68174
rect 69176 65754 69204 68190
rect 70096 66758 70124 70908
rect 71004 68316 71056 68322
rect 71004 68258 71056 68264
rect 70084 66752 70136 66758
rect 70084 66694 70136 66700
rect 71016 65754 71044 68258
rect 71200 68186 71228 70908
rect 72304 68254 72332 70908
rect 73408 68322 73436 70908
rect 73396 68316 73448 68322
rect 73396 68258 73448 68264
rect 74512 68254 74540 70908
rect 75616 68458 75644 70908
rect 76536 70894 76826 70922
rect 74592 68452 74644 68458
rect 74592 68394 74644 68400
rect 75604 68452 75656 68458
rect 75604 68394 75656 68400
rect 72292 68248 72344 68254
rect 72292 68190 72344 68196
rect 72844 68248 72896 68254
rect 72844 68190 72896 68196
rect 74500 68248 74552 68254
rect 74500 68190 74552 68196
rect 71188 68180 71240 68186
rect 71188 68122 71240 68128
rect 72856 65754 72884 68190
rect 74604 65754 74632 68394
rect 76536 65754 76564 70894
rect 68868 65726 69204 65754
rect 70708 65726 71044 65754
rect 72548 65726 72884 65754
rect 74480 65726 74632 65754
rect 76320 65726 76564 65754
rect 77916 65754 77944 70908
rect 79034 70894 79692 70922
rect 79664 65754 79692 70894
rect 80124 68254 80152 70908
rect 81228 68322 81256 70908
rect 82332 68866 82360 70908
rect 83436 68934 83464 70908
rect 83424 68928 83476 68934
rect 83424 68870 83476 68876
rect 82320 68860 82372 68866
rect 82320 68802 82372 68808
rect 81216 68316 81268 68322
rect 81216 68258 81268 68264
rect 83516 68316 83568 68322
rect 83516 68258 83568 68264
rect 80112 68248 80164 68254
rect 80112 68190 80164 68196
rect 81676 68248 81728 68254
rect 81676 68190 81728 68196
rect 81688 65754 81716 68190
rect 83528 65754 83556 68258
rect 84540 68254 84568 70908
rect 85356 68860 85408 68866
rect 85356 68802 85408 68808
rect 84528 68248 84580 68254
rect 84528 68190 84580 68196
rect 85368 65754 85396 68802
rect 85644 68322 85672 70908
rect 86748 68390 86776 70908
rect 87852 68934 87880 70908
rect 88956 69002 88984 70908
rect 88944 68996 88996 69002
rect 88944 68938 88996 68944
rect 87196 68928 87248 68934
rect 87196 68870 87248 68876
rect 87840 68928 87892 68934
rect 87840 68870 87892 68876
rect 86736 68384 86788 68390
rect 86736 68326 86788 68332
rect 85632 68316 85684 68322
rect 85632 68258 85684 68264
rect 87208 65754 87236 68870
rect 90152 68594 90180 70908
rect 91256 69342 91284 70908
rect 91244 69336 91296 69342
rect 91244 69278 91296 69284
rect 92360 69206 92388 70908
rect 92348 69200 92400 69206
rect 92348 69142 92400 69148
rect 93464 68866 93492 70908
rect 93452 68860 93504 68866
rect 93452 68802 93504 68808
rect 90140 68588 90192 68594
rect 90140 68530 90192 68536
rect 94568 68458 94596 70908
rect 94740 68928 94792 68934
rect 94740 68870 94792 68876
rect 94556 68452 94608 68458
rect 94556 68394 94608 68400
rect 92808 68384 92860 68390
rect 92808 68326 92860 68332
rect 90968 68316 91020 68322
rect 90968 68258 91020 68264
rect 89128 68248 89180 68254
rect 89128 68190 89180 68196
rect 89140 65754 89168 68190
rect 90980 65754 91008 68258
rect 92820 65754 92848 68326
rect 94752 65754 94780 68870
rect 95672 68390 95700 70908
rect 95660 68384 95712 68390
rect 95660 68326 95712 68332
rect 96776 68322 96804 70908
rect 97500 69200 97552 69206
rect 97500 69142 97552 69148
rect 96856 68996 96908 69002
rect 96856 68938 96908 68944
rect 96764 68316 96816 68322
rect 96764 68258 96816 68264
rect 96868 65754 96896 68938
rect 77916 65726 78160 65754
rect 79664 65726 80092 65754
rect 81688 65726 81932 65754
rect 83528 65726 83864 65754
rect 85368 65726 85704 65754
rect 87208 65726 87544 65754
rect 89140 65726 89476 65754
rect 90980 65726 91316 65754
rect 92820 65726 93156 65754
rect 94752 65726 95088 65754
rect 96868 65726 96928 65754
rect 66404 65596 66456 65602
rect 66404 65538 66456 65544
rect 66416 65505 66444 65538
rect 66402 65496 66458 65505
rect 66402 65431 66458 65440
rect 66312 65392 66364 65398
rect 66312 65334 66364 65340
rect 65668 65324 65720 65330
rect 65668 65266 65720 65272
rect 66402 64952 66458 64961
rect 66402 64887 66458 64896
rect 66416 64378 66444 64887
rect 63552 64372 63604 64378
rect 63552 64314 63604 64320
rect 66404 64372 66456 64378
rect 66404 64314 66456 64320
rect 63460 64236 63512 64242
rect 63460 64178 63512 64184
rect 63366 62776 63422 62785
rect 62724 62740 62776 62746
rect 63366 62711 63422 62720
rect 62724 62682 62776 62688
rect 13320 62672 13372 62678
rect 13320 62614 13372 62620
rect 29236 62672 29288 62678
rect 29236 62614 29288 62620
rect 11938 41288 11994 41297
rect 11938 41223 11994 41232
rect 13332 19673 13360 62614
rect 62736 60473 62764 62682
rect 62816 62672 62868 62678
rect 62816 62614 62868 62620
rect 62828 61017 62856 62614
rect 63472 61561 63500 64178
rect 63564 62105 63592 64314
rect 65666 64272 65722 64281
rect 65666 64207 65668 64216
rect 65720 64207 65722 64216
rect 65668 64178 65720 64184
rect 97512 63834 97540 69142
rect 97880 68526 97908 70908
rect 97868 68520 97920 68526
rect 97868 68462 97920 68468
rect 98984 68254 99012 70908
rect 98972 68248 99024 68254
rect 98972 68190 99024 68196
rect 100088 67710 100116 70908
rect 101192 68662 101220 71166
rect 101362 71143 101418 71152
rect 101914 71072 101970 71081
rect 101970 71044 102310 71058
rect 101970 71030 102324 71044
rect 101914 71007 101970 71016
rect 102296 68730 102324 71030
rect 102560 68860 102612 68866
rect 102560 68802 102612 68808
rect 102284 68724 102336 68730
rect 102284 68666 102336 68672
rect 101180 68656 101232 68662
rect 101180 68598 101232 68604
rect 102376 68520 102428 68526
rect 102376 68462 102428 68468
rect 100076 67704 100128 67710
rect 100076 67646 100128 67652
rect 102388 66457 102416 68462
rect 102468 68316 102520 68322
rect 102468 68258 102520 68264
rect 102374 66448 102430 66457
rect 102374 66383 102430 66392
rect 102480 65913 102508 68258
rect 102466 65904 102522 65913
rect 102466 65839 102522 65848
rect 100902 65496 100958 65505
rect 100902 65431 100904 65440
rect 100956 65431 100958 65440
rect 102376 65460 102428 65466
rect 100904 65402 100956 65408
rect 102376 65402 102428 65408
rect 100626 64544 100682 64553
rect 100626 64479 100628 64488
rect 100680 64479 100682 64488
rect 100628 64450 100680 64456
rect 100902 64136 100958 64145
rect 100902 64071 100904 64080
rect 100956 64071 100958 64080
rect 100904 64042 100956 64048
rect 97500 63828 97552 63834
rect 97500 63770 97552 63776
rect 66402 63728 66458 63737
rect 66402 63663 66458 63672
rect 65666 63184 65722 63193
rect 65666 63119 65722 63128
rect 65680 62746 65708 63119
rect 65668 62740 65720 62746
rect 65668 62682 65720 62688
rect 66416 62678 66444 63663
rect 100626 63320 100682 63329
rect 100626 63255 100682 63264
rect 100640 62882 100668 63255
rect 102388 63057 102416 65402
rect 102572 64145 102600 68802
rect 102652 68452 102704 68458
rect 102652 68394 102704 68400
rect 102664 64689 102692 68394
rect 102744 68384 102796 68390
rect 102744 68326 102796 68332
rect 102756 65233 102784 68326
rect 102928 68180 102980 68186
rect 102928 68122 102980 68128
rect 102940 67001 102968 68122
rect 105240 67794 105268 73727
rect 105208 67766 105268 67794
rect 105424 67794 105452 74271
rect 105870 72568 105926 72577
rect 105870 72503 105926 72512
rect 105884 72470 105912 72503
rect 105872 72464 105924 72470
rect 105872 72406 105924 72412
rect 105976 67794 106004 75495
rect 106514 71072 106570 71081
rect 106514 71007 106570 71016
rect 106528 70362 106556 71007
rect 106516 70356 106568 70362
rect 106516 70298 106568 70304
rect 106988 67794 107016 76719
rect 107540 67794 107568 77846
rect 107724 76657 107752 83354
rect 107816 81417 107844 84782
rect 108000 83729 108028 86346
rect 107986 83720 108042 83729
rect 107986 83655 108042 83664
rect 107896 82188 107948 82194
rect 107896 82130 107948 82136
rect 107802 81408 107858 81417
rect 107802 81343 107858 81352
rect 107710 76648 107766 76657
rect 107710 76583 107766 76592
rect 107908 74345 107936 82130
rect 108540 80828 108592 80834
rect 108540 80770 108592 80776
rect 108080 79264 108132 79270
rect 108080 79206 108132 79212
rect 107894 74336 107950 74345
rect 107894 74271 107950 74280
rect 108092 67794 108120 79206
rect 108552 72033 108580 80770
rect 109184 72464 109236 72470
rect 109184 72406 109236 72412
rect 108538 72024 108594 72033
rect 108538 71959 108594 71968
rect 109196 70922 109224 72406
rect 109196 70894 109316 70922
rect 108356 70356 108408 70362
rect 108356 70298 108408 70304
rect 105424 67766 105760 67794
rect 105976 67766 106312 67794
rect 106956 67766 107016 67794
rect 107508 67766 107568 67794
rect 108060 67766 108120 67794
rect 108368 67794 108396 70298
rect 109288 67794 109316 70894
rect 110564 69132 110616 69138
rect 110564 69074 110616 69080
rect 110104 68860 110156 68866
rect 110104 68802 110156 68808
rect 110116 67794 110144 68802
rect 110576 67794 110604 69074
rect 111128 68866 111156 70908
rect 111496 69138 111524 70908
rect 111588 70894 111878 70922
rect 111956 70894 112338 70922
rect 112416 70894 112706 70922
rect 111484 69132 111536 69138
rect 111484 69074 111536 69080
rect 111116 68860 111168 68866
rect 111116 68802 111168 68808
rect 111588 67930 111616 70894
rect 111404 67902 111616 67930
rect 111404 67794 111432 67902
rect 111956 67794 111984 70894
rect 112416 67794 112444 70894
rect 113060 67794 113088 70908
rect 113336 70894 113534 70922
rect 113902 70894 114008 70922
rect 113336 67794 113364 70894
rect 108368 67766 108704 67794
rect 109256 67766 109316 67794
rect 109808 67766 110144 67794
rect 110452 67766 110604 67794
rect 111004 67766 111432 67794
rect 111556 67766 111984 67794
rect 112200 67766 112444 67794
rect 112752 67766 113088 67794
rect 113304 67766 113364 67794
rect 103480 67704 103532 67710
rect 113980 67658 114008 70894
rect 114256 67794 114284 70908
rect 114730 70894 114928 70922
rect 115098 70894 115388 70922
rect 115466 70894 115848 70922
rect 115926 70894 116216 70922
rect 114900 67794 114928 70894
rect 115360 67794 115388 70894
rect 115820 68202 115848 70894
rect 116188 68474 116216 70894
rect 116280 68866 116308 70908
rect 116648 69614 116676 70908
rect 117108 69682 117136 70908
rect 117096 69676 117148 69682
rect 117096 69618 117148 69624
rect 116636 69608 116688 69614
rect 116636 69550 116688 69556
rect 117476 68866 117504 70908
rect 117648 69608 117700 69614
rect 117648 69550 117700 69556
rect 116268 68860 116320 68866
rect 116268 68802 116320 68808
rect 117096 68860 117148 68866
rect 117096 68802 117148 68808
rect 117464 68860 117516 68866
rect 117464 68802 117516 68808
rect 116188 68446 116400 68474
rect 115820 68174 115940 68202
rect 114256 67766 114500 67794
rect 114900 67766 115052 67794
rect 115360 67766 115696 67794
rect 103480 67646 103532 67652
rect 103492 67545 103520 67646
rect 113948 67630 114008 67658
rect 115912 67658 115940 68174
rect 116372 67794 116400 68446
rect 117108 67794 117136 68802
rect 117660 67794 117688 69550
rect 117844 69177 117872 70908
rect 118200 69676 118252 69682
rect 118200 69618 118252 69624
rect 117830 69168 117886 69177
rect 117830 69103 117886 69112
rect 118212 67794 118240 69618
rect 118304 69614 118332 70908
rect 118672 69682 118700 70908
rect 118660 69676 118712 69682
rect 118660 69618 118712 69624
rect 118292 69608 118344 69614
rect 118292 69550 118344 69556
rect 119132 69041 119160 70908
rect 119500 69750 119528 70908
rect 119868 69818 119896 70908
rect 120342 70894 120540 70922
rect 119856 69812 119908 69818
rect 119856 69754 119908 69760
rect 119488 69744 119540 69750
rect 119488 69686 119540 69692
rect 120316 69608 120368 69614
rect 120316 69550 120368 69556
rect 119394 69168 119450 69177
rect 119394 69103 119450 69112
rect 119118 69032 119174 69041
rect 119118 68967 119174 68976
rect 118936 68860 118988 68866
rect 118936 68802 118988 68808
rect 118948 67794 118976 68802
rect 119408 67794 119436 69103
rect 120328 67794 120356 69550
rect 120512 68934 120540 70894
rect 120592 69676 120644 69682
rect 120592 69618 120644 69624
rect 120500 68928 120552 68934
rect 120500 68870 120552 68876
rect 116372 67766 116800 67794
rect 117108 67766 117444 67794
rect 117660 67766 117996 67794
rect 118212 67766 118548 67794
rect 118948 67766 119192 67794
rect 119408 67766 119744 67794
rect 120296 67766 120356 67794
rect 120604 67794 120632 69618
rect 120696 68798 120724 70908
rect 121064 69138 121092 70908
rect 121052 69132 121104 69138
rect 121052 69074 121104 69080
rect 121142 69032 121198 69041
rect 121142 68967 121198 68976
rect 120684 68792 120736 68798
rect 120684 68734 120736 68740
rect 121156 67794 121184 68967
rect 121524 68526 121552 70908
rect 121696 69744 121748 69750
rect 121696 69686 121748 69692
rect 121512 68520 121564 68526
rect 121512 68462 121564 68468
rect 121708 67794 121736 69686
rect 121892 69274 121920 70908
rect 121880 69268 121932 69274
rect 121880 69210 121932 69216
rect 122260 69206 122288 70908
rect 122340 69812 122392 69818
rect 122340 69754 122392 69760
rect 122248 69200 122300 69206
rect 122248 69142 122300 69148
rect 122352 67794 122380 69754
rect 122720 69002 122748 70908
rect 123102 70894 123392 70922
rect 122708 68996 122760 69002
rect 122708 68938 122760 68944
rect 123076 68928 123128 68934
rect 123076 68870 123128 68876
rect 123088 67794 123116 68870
rect 123364 68866 123392 70894
rect 123456 69478 123484 70908
rect 123444 69472 123496 69478
rect 123444 69414 123496 69420
rect 123352 68860 123404 68866
rect 123352 68802 123404 68808
rect 123444 68792 123496 68798
rect 123444 68734 123496 68740
rect 123456 67794 123484 68734
rect 123916 68594 123944 70908
rect 124284 68934 124312 70908
rect 124652 69410 124680 70908
rect 124640 69404 124692 69410
rect 124640 69346 124692 69352
rect 124456 69132 124508 69138
rect 124456 69074 124508 69080
rect 124272 68928 124324 68934
rect 124272 68870 124324 68876
rect 123904 68588 123956 68594
rect 123904 68530 123956 68536
rect 124468 67794 124496 69074
rect 125112 69070 125140 70908
rect 125480 69274 125508 70908
rect 125192 69268 125244 69274
rect 125192 69210 125244 69216
rect 125468 69268 125520 69274
rect 125468 69210 125520 69216
rect 125100 69064 125152 69070
rect 125100 69006 125152 69012
rect 124640 68520 124692 68526
rect 124640 68462 124692 68468
rect 120604 67766 120940 67794
rect 121156 67766 121492 67794
rect 121708 67766 122044 67794
rect 122352 67766 122688 67794
rect 123088 67766 123240 67794
rect 123456 67766 123792 67794
rect 124436 67766 124496 67794
rect 124652 67794 124680 68462
rect 125204 67794 125232 69210
rect 125848 69206 125876 70908
rect 126308 69546 126336 70908
rect 126296 69540 126348 69546
rect 126296 69482 126348 69488
rect 125836 69200 125888 69206
rect 125836 69142 125888 69148
rect 126676 69138 126704 70908
rect 131632 69608 131684 69614
rect 131632 69550 131684 69556
rect 127584 69472 127636 69478
rect 127584 69414 127636 69420
rect 125928 69132 125980 69138
rect 125928 69074 125980 69080
rect 126664 69132 126716 69138
rect 126664 69074 126716 69080
rect 125940 67794 125968 69074
rect 126388 68996 126440 69002
rect 126388 68938 126440 68944
rect 126400 67794 126428 68938
rect 127308 68860 127360 68866
rect 127308 68802 127360 68808
rect 124652 67766 124988 67794
rect 125204 67766 125540 67794
rect 125940 67766 126184 67794
rect 126400 67766 126736 67794
rect 127320 67658 127348 68802
rect 127596 67794 127624 69414
rect 129332 69404 129384 69410
rect 129332 69346 129384 69352
rect 128688 68928 128740 68934
rect 128688 68870 128740 68876
rect 128136 68588 128188 68594
rect 128136 68530 128188 68536
rect 128148 67794 128176 68530
rect 128700 67794 128728 68870
rect 129344 67794 129372 69346
rect 130436 69268 130488 69274
rect 130436 69210 130488 69216
rect 129884 69064 129936 69070
rect 129936 69012 130016 69018
rect 129884 69006 130016 69012
rect 129896 68990 130016 69006
rect 129988 67794 130016 68990
rect 130448 67794 130476 69210
rect 131264 69200 131316 69206
rect 131316 69148 131396 69154
rect 131264 69142 131396 69148
rect 131276 69126 131396 69142
rect 131368 68066 131396 69126
rect 131368 68038 131442 68066
rect 127596 67766 127932 67794
rect 128148 67766 128484 67794
rect 128700 67766 129036 67794
rect 129344 67766 129680 67794
rect 129988 67766 130232 67794
rect 130448 67766 130784 67794
rect 131414 67780 131442 68038
rect 115912 67630 116248 67658
rect 127288 67630 127348 67658
rect 131644 67658 131672 69550
rect 132104 69342 132132 113750
rect 132460 113740 132512 113746
rect 132460 113682 132512 113688
rect 132472 112250 132500 113682
rect 132564 112794 132592 113870
rect 154828 113678 154856 115924
rect 164488 115910 164870 115938
rect 154816 113672 154868 113678
rect 144878 113640 144934 113649
rect 154816 113614 154868 113620
rect 144878 113575 144934 113584
rect 132552 112788 132604 112794
rect 132552 112730 132604 112736
rect 132460 112244 132512 112250
rect 132460 112186 132512 112192
rect 144892 110756 144920 113575
rect 164488 112182 164516 115910
rect 172662 115680 172718 115689
rect 172662 115615 172664 115624
rect 172716 115615 172718 115624
rect 172664 115586 172716 115592
rect 173872 114737 173900 116538
rect 173964 116505 173992 118034
rect 204770 117992 204826 118001
rect 204770 117927 204826 117936
rect 174044 117888 174096 117894
rect 174044 117830 174096 117836
rect 174056 117049 174084 117830
rect 174136 117820 174188 117826
rect 174136 117762 174188 117768
rect 174148 117593 174176 117762
rect 174134 117584 174190 117593
rect 174134 117519 174190 117528
rect 174042 117040 174098 117049
rect 174042 116975 174098 116984
rect 173950 116496 174006 116505
rect 173950 116431 174006 116440
rect 174228 116460 174280 116466
rect 174228 116402 174280 116408
rect 174136 116392 174188 116398
rect 174136 116334 174188 116340
rect 174148 115825 174176 116334
rect 174134 115816 174190 115825
rect 174134 115751 174190 115760
rect 174044 115644 174096 115650
rect 174044 115586 174096 115592
rect 173858 114728 173914 114737
rect 173858 114663 173914 114672
rect 174056 114193 174084 115586
rect 174240 115281 174268 116402
rect 174226 115272 174282 115281
rect 174226 115207 174282 115216
rect 204784 115174 204812 117927
rect 204772 115168 204824 115174
rect 204772 115110 204824 115116
rect 174042 114184 174098 114193
rect 174042 114119 174098 114128
rect 164842 113640 164898 113649
rect 164842 113575 164898 113584
rect 164476 112176 164528 112182
rect 164476 112118 164528 112124
rect 164856 110756 164884 113575
rect 177080 111156 177132 111162
rect 177080 111098 177132 111104
rect 176896 111088 176948 111094
rect 176896 111030 176948 111036
rect 132552 110272 132604 110278
rect 132552 110214 132604 110220
rect 132564 95833 132592 110214
rect 176908 106577 176936 111030
rect 176988 111020 177040 111026
rect 176988 110962 177040 110968
rect 177000 107801 177028 110962
rect 176986 107792 177042 107801
rect 176986 107727 177042 107736
rect 176894 106568 176950 106577
rect 176894 106503 176950 106512
rect 177092 105353 177120 111098
rect 177078 105344 177134 105353
rect 177078 105279 177134 105288
rect 177184 105194 177212 113884
rect 177736 113762 177764 113884
rect 177552 113734 177764 113762
rect 177264 111224 177316 111230
rect 177264 111166 177316 111172
rect 176908 105166 177212 105194
rect 176908 101681 176936 105166
rect 177276 104129 177304 111166
rect 177356 109048 177408 109054
rect 177354 109016 177356 109025
rect 177408 109016 177410 109025
rect 177354 108951 177410 108960
rect 177262 104120 177318 104129
rect 177262 104055 177318 104064
rect 177552 102905 177580 113734
rect 178288 111230 178316 113884
rect 178276 111224 178328 111230
rect 178276 111166 178328 111172
rect 178840 111162 178868 113884
rect 178828 111156 178880 111162
rect 178828 111098 178880 111104
rect 179392 111094 179420 113884
rect 179380 111088 179432 111094
rect 179380 111030 179432 111036
rect 180036 111026 180064 113884
rect 180024 111020 180076 111026
rect 180024 110962 180076 110968
rect 177724 110952 177776 110958
rect 177724 110894 177776 110900
rect 177736 110249 177764 110894
rect 177722 110240 177778 110249
rect 177722 110175 177778 110184
rect 180298 109560 180354 109569
rect 180298 109495 180354 109504
rect 179654 104936 179710 104945
rect 179654 104871 179710 104880
rect 179668 104090 179696 104871
rect 178184 104084 178236 104090
rect 178184 104026 178236 104032
rect 179656 104084 179708 104090
rect 179656 104026 179708 104032
rect 177538 102896 177594 102905
rect 177538 102831 177594 102840
rect 176894 101672 176950 101681
rect 176894 101607 176950 101616
rect 177632 101364 177684 101370
rect 177632 101306 177684 101312
rect 176988 100820 177040 100826
rect 176988 100762 177040 100768
rect 177000 100457 177028 100762
rect 176986 100448 177042 100457
rect 176986 100383 177042 100392
rect 177356 99324 177408 99330
rect 177356 99266 177408 99272
rect 177368 99233 177396 99266
rect 177354 99224 177410 99233
rect 177354 99159 177410 99168
rect 177540 97216 177592 97222
rect 177540 97158 177592 97164
rect 132366 95824 132422 95833
rect 132366 95759 132422 95768
rect 132550 95824 132606 95833
rect 132550 95759 132606 95768
rect 132380 88926 132408 95759
rect 177552 94473 177580 97158
rect 177644 96921 177672 101306
rect 177724 99936 177776 99942
rect 177724 99878 177776 99884
rect 177630 96912 177686 96921
rect 177630 96847 177686 96856
rect 177736 95697 177764 99878
rect 178196 98145 178224 104026
rect 179654 102488 179710 102497
rect 179654 102423 179710 102432
rect 179668 101370 179696 102423
rect 179656 101364 179708 101370
rect 179656 101306 179708 101312
rect 180312 100826 180340 109495
rect 180588 109054 180616 113884
rect 181140 110958 181168 113884
rect 181692 111026 181720 113884
rect 182244 111434 182272 113884
rect 182232 111428 182284 111434
rect 182232 111370 182284 111376
rect 182888 111366 182916 113884
rect 183244 111428 183296 111434
rect 183244 111370 183296 111376
rect 182876 111360 182928 111366
rect 182876 111302 182928 111308
rect 181680 111020 181732 111026
rect 181680 110962 181732 110968
rect 183106 111020 183158 111026
rect 183106 110962 183158 110968
rect 181128 110952 181180 110958
rect 181128 110894 181180 110900
rect 183118 110756 183146 110962
rect 183256 110770 183284 111370
rect 183440 111026 183468 113884
rect 183992 113134 184020 113884
rect 183980 113128 184032 113134
rect 183980 113070 184032 113076
rect 184440 113128 184492 113134
rect 184440 113070 184492 113076
rect 183796 111360 183848 111366
rect 183796 111302 183848 111308
rect 183428 111020 183480 111026
rect 183428 110962 183480 110968
rect 183808 110770 183836 111302
rect 184302 111020 184354 111026
rect 184302 110962 184354 110968
rect 183256 110742 183500 110770
rect 183808 110742 183868 110770
rect 184314 110756 184342 110962
rect 184452 110770 184480 113070
rect 184544 110906 184572 113884
rect 185096 111042 185124 113884
rect 185096 111014 185216 111042
rect 184544 110878 184848 110906
rect 184820 110770 184848 110878
rect 185188 110770 185216 111014
rect 185740 110770 185768 113884
rect 186292 111042 186320 113884
rect 186246 111014 186320 111042
rect 184452 110742 184696 110770
rect 184820 110742 185064 110770
rect 185188 110742 185524 110770
rect 185740 110742 185892 110770
rect 186246 110756 186274 111014
rect 186844 110770 186872 113884
rect 187396 110906 187424 113884
rect 187948 111042 187976 113884
rect 188488 113128 188540 113134
rect 188488 113070 188540 113076
rect 188028 112788 188080 112794
rect 188028 112730 188080 112736
rect 187304 110878 187424 110906
rect 187764 111014 187976 111042
rect 187304 110770 187332 110878
rect 187764 110770 187792 111014
rect 188040 110770 188068 112730
rect 188500 110770 188528 113070
rect 188592 112794 188620 113884
rect 188948 113196 189000 113202
rect 188948 113138 189000 113144
rect 188580 112788 188632 112794
rect 188580 112730 188632 112736
rect 188960 110770 188988 113138
rect 189144 113134 189172 113884
rect 189696 113202 189724 113884
rect 189684 113196 189736 113202
rect 189684 113138 189736 113144
rect 189132 113128 189184 113134
rect 189132 113070 189184 113076
rect 190248 112658 190276 113884
rect 189224 112652 189276 112658
rect 189224 112594 189276 112600
rect 190236 112652 190288 112658
rect 190236 112594 190288 112600
rect 189236 110770 189264 112594
rect 190800 112522 190828 113884
rect 191340 112924 191392 112930
rect 191340 112866 191392 112872
rect 189592 112516 189644 112522
rect 189592 112458 189644 112464
rect 190788 112516 190840 112522
rect 190788 112458 190840 112464
rect 189604 110770 189632 112458
rect 190512 112448 190564 112454
rect 190512 112390 190564 112396
rect 190144 112380 190196 112386
rect 190144 112322 190196 112328
rect 190156 110770 190184 112322
rect 190524 110770 190552 112390
rect 190604 112108 190656 112114
rect 190604 112050 190656 112056
rect 186720 110742 186872 110770
rect 187088 110742 187332 110770
rect 187456 110742 187792 110770
rect 187916 110742 188068 110770
rect 188284 110742 188528 110770
rect 188652 110742 188988 110770
rect 189112 110742 189264 110770
rect 189480 110742 189632 110770
rect 189848 110742 190184 110770
rect 190308 110742 190552 110770
rect 190616 110770 190644 112050
rect 191352 110770 191380 112866
rect 191444 112386 191472 113884
rect 191996 112454 192024 113884
rect 192548 113082 192576 113884
rect 192456 113054 192576 113082
rect 191984 112448 192036 112454
rect 191984 112390 192036 112396
rect 191432 112380 191484 112386
rect 191432 112322 191484 112328
rect 191708 112380 191760 112386
rect 191708 112322 191760 112328
rect 191720 110770 191748 112322
rect 192456 112114 192484 113054
rect 193100 112930 193128 113884
rect 193088 112924 193140 112930
rect 193088 112866 193140 112872
rect 192904 112788 192956 112794
rect 192904 112730 192956 112736
rect 192536 112652 192588 112658
rect 192536 112594 192588 112600
rect 192444 112108 192496 112114
rect 192444 112050 192496 112056
rect 191984 111360 192036 111366
rect 191984 111302 192036 111308
rect 191996 110770 192024 111302
rect 192548 110770 192576 112594
rect 192916 110770 192944 112730
rect 193180 112380 193232 112386
rect 193180 112322 193232 112328
rect 193192 110770 193220 112322
rect 193652 112318 193680 113884
rect 193732 113060 193784 113066
rect 193732 113002 193784 113008
rect 193640 112312 193692 112318
rect 193640 112254 193692 112260
rect 193744 110770 193772 113002
rect 194100 111428 194152 111434
rect 194100 111370 194152 111376
rect 194112 110770 194140 111370
rect 194296 111366 194324 113884
rect 194744 112652 194796 112658
rect 194848 112640 194876 113884
rect 195400 112794 195428 113884
rect 195756 113128 195808 113134
rect 195756 113070 195808 113076
rect 195388 112788 195440 112794
rect 195388 112730 195440 112736
rect 194796 112612 194876 112640
rect 194744 112594 194796 112600
rect 194560 112448 194612 112454
rect 194560 112390 194612 112396
rect 194284 111360 194336 111366
rect 194284 111302 194336 111308
rect 194572 110770 194600 112390
rect 194744 112380 194796 112386
rect 194744 112322 194796 112328
rect 194756 111042 194784 112322
rect 195296 111360 195348 111366
rect 195296 111302 195348 111308
rect 190616 110742 190676 110770
rect 191136 110742 191380 110770
rect 191504 110742 191748 110770
rect 191872 110742 192024 110770
rect 192332 110742 192576 110770
rect 192700 110742 192944 110770
rect 193068 110742 193220 110770
rect 193528 110742 193772 110770
rect 193896 110742 194140 110770
rect 194264 110742 194600 110770
rect 194710 111014 194784 111042
rect 194710 110756 194738 111014
rect 195308 110770 195336 111302
rect 195768 110770 195796 113070
rect 195952 112318 195980 113884
rect 196504 113066 196532 113884
rect 196492 113060 196544 113066
rect 196492 113002 196544 113008
rect 196124 112992 196176 112998
rect 196124 112934 196176 112940
rect 195940 112312 195992 112318
rect 195940 112254 195992 112260
rect 196136 110770 196164 112934
rect 196492 112788 196544 112794
rect 196492 112730 196544 112736
rect 196504 110770 196532 112730
rect 196952 112652 197004 112658
rect 196952 112594 197004 112600
rect 196964 110770 196992 112594
rect 197148 111434 197176 113884
rect 197320 112720 197372 112726
rect 197320 112662 197372 112668
rect 197136 111428 197188 111434
rect 197136 111370 197188 111376
rect 197332 110770 197360 112662
rect 197412 112584 197464 112590
rect 197412 112526 197464 112532
rect 195092 110742 195336 110770
rect 195460 110742 195796 110770
rect 195920 110742 196164 110770
rect 196288 110742 196532 110770
rect 196656 110742 196992 110770
rect 197116 110742 197360 110770
rect 197424 110634 197452 112526
rect 197700 112454 197728 113884
rect 198148 112516 198200 112522
rect 198148 112458 198200 112464
rect 197688 112448 197740 112454
rect 197688 112390 197740 112396
rect 198160 110770 198188 112458
rect 198252 112386 198280 113884
rect 198240 112380 198292 112386
rect 198240 112322 198292 112328
rect 198516 112380 198568 112386
rect 198516 112322 198568 112328
rect 198528 110770 198556 112322
rect 198804 111366 198832 113884
rect 199356 113134 199384 113884
rect 199344 113128 199396 113134
rect 199344 113070 199396 113076
rect 200000 112998 200028 113884
rect 199988 112992 200040 112998
rect 199988 112934 200040 112940
rect 200552 112794 200580 113884
rect 200540 112788 200592 112794
rect 200540 112730 200592 112736
rect 201104 112658 201132 113884
rect 201656 112726 201684 113884
rect 201644 112720 201696 112726
rect 201644 112662 201696 112668
rect 201092 112652 201144 112658
rect 201092 112594 201144 112600
rect 202208 112590 202236 113884
rect 202196 112584 202248 112590
rect 202196 112526 202248 112532
rect 202852 112522 202880 113884
rect 202840 112516 202892 112522
rect 202840 112458 202892 112464
rect 198884 112448 198936 112454
rect 198884 112390 198936 112396
rect 198792 111360 198844 111366
rect 198792 111302 198844 111308
rect 198896 110770 198924 112390
rect 203404 112318 203432 113884
rect 203956 112318 203984 113884
rect 204522 113870 204720 113898
rect 203392 112312 203444 112318
rect 203392 112254 203444 112260
rect 203944 112312 203996 112318
rect 203944 112254 203996 112260
rect 197852 110742 198188 110770
rect 198312 110742 198556 110770
rect 198680 110742 198924 110770
rect 197424 110606 197484 110634
rect 180576 109048 180628 109054
rect 180576 108990 180628 108996
rect 180390 107248 180446 107257
rect 180390 107183 180446 107192
rect 180300 100820 180352 100826
rect 180300 100762 180352 100768
rect 179654 100176 179710 100185
rect 179654 100111 179710 100120
rect 179668 99942 179696 100111
rect 179656 99936 179708 99942
rect 179656 99878 179708 99884
rect 180404 99330 180432 107183
rect 204692 104265 204720 113870
rect 205060 113678 205088 124750
rect 207912 118545 207940 141902
rect 208004 127793 208032 141970
rect 210580 141966 210608 144892
rect 215916 142714 215944 144892
rect 215904 142708 215956 142714
rect 215904 142650 215956 142656
rect 221252 142034 221280 144892
rect 222540 142102 222568 156846
rect 222908 156602 222936 158070
rect 223552 156926 223580 159135
rect 223540 156920 223592 156926
rect 223540 156862 223592 156868
rect 222724 156574 222936 156602
rect 222724 146946 222752 156574
rect 223538 149544 223594 149553
rect 223538 149479 223594 149488
rect 222632 146918 222752 146946
rect 222632 146810 222660 146918
rect 222632 146782 222936 146810
rect 222528 142096 222580 142102
rect 222528 142038 222580 142044
rect 222804 142096 222856 142102
rect 222804 142038 222856 142044
rect 221240 142028 221292 142034
rect 221240 141970 221292 141976
rect 210568 141960 210620 141966
rect 210568 141902 210620 141908
rect 222528 141960 222580 141966
rect 222528 141902 222580 141908
rect 207990 127784 208046 127793
rect 207990 127719 208046 127728
rect 207898 118536 207954 118545
rect 207898 118471 207954 118480
rect 205048 113672 205100 113678
rect 205048 113614 205100 113620
rect 201090 104256 201146 104265
rect 201090 104191 201146 104200
rect 204678 104256 204734 104265
rect 204678 104191 204734 104200
rect 180392 99324 180444 99330
rect 180392 99266 180444 99272
rect 178182 98136 178238 98145
rect 178182 98071 178238 98080
rect 179654 97864 179710 97873
rect 179654 97799 179710 97808
rect 179668 97222 179696 97799
rect 179656 97216 179708 97222
rect 179656 97158 179708 97164
rect 177722 95688 177778 95697
rect 177722 95623 177778 95632
rect 179562 95416 179618 95425
rect 179562 95351 179618 95360
rect 177538 94464 177594 94473
rect 177538 94399 177594 94408
rect 179576 93958 179604 95351
rect 177356 93952 177408 93958
rect 177356 93894 177408 93900
rect 179564 93952 179616 93958
rect 179564 93894 179616 93900
rect 177368 93249 177396 93894
rect 177354 93240 177410 93249
rect 177354 93175 177410 93184
rect 179562 93104 179618 93113
rect 179562 93039 179618 93048
rect 179576 92054 179604 93039
rect 176988 92048 177040 92054
rect 176986 92016 176988 92025
rect 179564 92048 179616 92054
rect 177040 92016 177042 92025
rect 179564 91990 179616 91996
rect 176986 91951 177042 91960
rect 201104 91646 201132 104191
rect 201092 91640 201144 91646
rect 201092 91582 201144 91588
rect 204496 91640 204548 91646
rect 204496 91582 204548 91588
rect 204508 90937 204536 91582
rect 200998 90928 201054 90937
rect 200998 90863 201054 90872
rect 204494 90928 204550 90937
rect 204494 90863 204550 90872
rect 132368 88920 132420 88926
rect 132368 88862 132420 88868
rect 132552 88852 132604 88858
rect 132552 88794 132604 88800
rect 132564 79338 132592 88794
rect 177354 88344 177410 88353
rect 177354 88279 177410 88288
rect 177368 87566 177396 88279
rect 177356 87560 177408 87566
rect 177356 87502 177408 87508
rect 179656 87560 179708 87566
rect 179656 87502 179708 87508
rect 177538 87120 177594 87129
rect 177538 87055 177594 87064
rect 177552 86138 177580 87055
rect 177540 86132 177592 86138
rect 177540 86074 177592 86080
rect 179668 86041 179696 87502
rect 179748 86132 179800 86138
rect 179748 86074 179800 86080
rect 179654 86032 179710 86041
rect 179654 85967 179710 85976
rect 176986 85896 177042 85905
rect 176986 85831 177042 85840
rect 177000 84846 177028 85831
rect 176988 84840 177040 84846
rect 179564 84840 179616 84846
rect 176988 84782 177040 84788
rect 178182 84808 178238 84817
rect 179564 84782 179616 84788
rect 178182 84743 178184 84752
rect 178236 84743 178238 84752
rect 178184 84714 178236 84720
rect 178090 83584 178146 83593
rect 178090 83519 178146 83528
rect 178104 83486 178132 83519
rect 178092 83480 178144 83486
rect 178092 83422 178144 83428
rect 179472 83480 179524 83486
rect 179472 83422 179524 83428
rect 177722 82360 177778 82369
rect 177722 82295 177724 82304
rect 177776 82295 177778 82304
rect 177724 82266 177776 82272
rect 178090 81136 178146 81145
rect 178090 81071 178146 81080
rect 178104 80630 178132 81071
rect 178092 80624 178144 80630
rect 178092 80566 178144 80572
rect 177630 79912 177686 79921
rect 177630 79847 177686 79856
rect 132552 79332 132604 79338
rect 132552 79274 132604 79280
rect 177644 79270 177672 79847
rect 177632 79264 177684 79270
rect 177632 79206 177684 79212
rect 132552 79196 132604 79202
rect 132552 79138 132604 79144
rect 132092 69336 132144 69342
rect 132092 69278 132144 69284
rect 132184 69132 132236 69138
rect 132184 69074 132236 69080
rect 132196 67794 132224 69074
rect 132564 68798 132592 79138
rect 176986 78688 177042 78697
rect 176986 78623 177042 78632
rect 177000 77910 177028 78623
rect 176988 77904 177040 77910
rect 176988 77846 177040 77852
rect 179380 77904 179432 77910
rect 179380 77846 179432 77852
rect 178826 77464 178882 77473
rect 178826 77399 178882 77408
rect 178274 76240 178330 76249
rect 178274 76175 178330 76184
rect 177722 75016 177778 75025
rect 177722 74951 177778 74960
rect 177170 73792 177226 73801
rect 177170 73727 177226 73736
rect 135522 70894 135628 70922
rect 132552 68792 132604 68798
rect 132552 68734 132604 68740
rect 134484 68248 134536 68254
rect 134484 68190 134536 68196
rect 132196 67766 132532 67794
rect 131644 67630 131980 67658
rect 103478 67536 103534 67545
rect 103478 67471 103534 67480
rect 102926 66992 102982 67001
rect 102926 66927 102982 66936
rect 102742 65224 102798 65233
rect 102742 65159 102798 65168
rect 102650 64680 102706 64689
rect 102650 64615 102706 64624
rect 102744 64508 102796 64514
rect 102744 64450 102796 64456
rect 102558 64136 102614 64145
rect 102468 64100 102520 64106
rect 102558 64071 102614 64080
rect 102468 64042 102520 64048
rect 102374 63048 102430 63057
rect 102374 62983 102430 62992
rect 100628 62876 100680 62882
rect 100628 62818 100680 62824
rect 102376 62876 102428 62882
rect 102376 62818 102428 62824
rect 100626 62776 100682 62785
rect 100626 62711 100628 62720
rect 100680 62711 100682 62720
rect 100628 62682 100680 62688
rect 66404 62672 66456 62678
rect 66404 62614 66456 62620
rect 66402 62504 66458 62513
rect 66402 62439 66458 62448
rect 63550 62096 63606 62105
rect 63550 62031 63606 62040
rect 65666 61960 65722 61969
rect 65666 61895 65722 61904
rect 63458 61552 63514 61561
rect 62908 61516 62960 61522
rect 65680 61522 65708 61895
rect 63458 61487 63514 61496
rect 65668 61516 65720 61522
rect 62908 61458 62960 61464
rect 65668 61458 65720 61464
rect 62814 61008 62870 61017
rect 62814 60943 62870 60952
rect 62722 60464 62778 60473
rect 62722 60399 62778 60408
rect 62632 60156 62684 60162
rect 62632 60098 62684 60104
rect 62644 57617 62672 60098
rect 62724 59952 62776 59958
rect 62724 59894 62776 59900
rect 62736 58161 62764 59894
rect 62920 59249 62948 61458
rect 66416 61318 66444 62439
rect 100626 62096 100682 62105
rect 100626 62031 100682 62040
rect 100534 61416 100590 61425
rect 100640 61386 100668 62031
rect 100534 61351 100590 61360
rect 100628 61380 100680 61386
rect 100548 61318 100576 61351
rect 100628 61322 100680 61328
rect 63736 61312 63788 61318
rect 66404 61312 66456 61318
rect 63736 61254 63788 61260
rect 65482 61280 65538 61289
rect 63748 59929 63776 61254
rect 66404 61254 66456 61260
rect 100536 61312 100588 61318
rect 102388 61289 102416 62818
rect 102480 61833 102508 64042
rect 102560 63828 102612 63834
rect 102560 63770 102612 63776
rect 102572 63601 102600 63770
rect 102558 63592 102614 63601
rect 102558 63527 102614 63536
rect 102560 62740 102612 62746
rect 102560 62682 102612 62688
rect 102466 61824 102522 61833
rect 102466 61759 102522 61768
rect 102468 61380 102520 61386
rect 102468 61322 102520 61328
rect 100536 61254 100588 61260
rect 102374 61280 102430 61289
rect 65482 61215 65538 61224
rect 102374 61215 102430 61224
rect 65496 60638 65524 61215
rect 100626 60872 100682 60881
rect 100626 60807 100682 60816
rect 66310 60736 66366 60745
rect 66310 60671 66366 60680
rect 63828 60632 63880 60638
rect 63828 60574 63880 60580
rect 65484 60632 65536 60638
rect 65484 60574 65536 60580
rect 63734 59920 63790 59929
rect 63734 59855 63790 59864
rect 62906 59240 62962 59249
rect 62906 59175 62962 59184
rect 63840 58705 63868 60574
rect 66324 59958 66352 60671
rect 100640 60434 100668 60807
rect 100628 60428 100680 60434
rect 100628 60370 100680 60376
rect 100626 60328 100682 60337
rect 100626 60263 100628 60272
rect 100680 60263 100682 60272
rect 102376 60292 102428 60298
rect 100628 60234 100680 60240
rect 102376 60234 102428 60240
rect 66402 60192 66458 60201
rect 66402 60127 66404 60136
rect 66456 60127 66458 60136
rect 66404 60098 66456 60104
rect 100626 60056 100682 60065
rect 100626 59991 100628 60000
rect 100680 59991 100682 60000
rect 100628 59962 100680 59968
rect 66312 59952 66364 59958
rect 66312 59894 66364 59900
rect 66310 59512 66366 59521
rect 66310 59447 66366 59456
rect 63826 58696 63882 58705
rect 62816 58660 62868 58666
rect 66324 58666 66352 59447
rect 100626 59104 100682 59113
rect 100626 59039 100682 59048
rect 66402 58968 66458 58977
rect 66402 58903 66458 58912
rect 63826 58631 63882 58640
rect 66312 58660 66364 58666
rect 62816 58602 62868 58608
rect 66312 58602 66364 58608
rect 62722 58152 62778 58161
rect 62722 58087 62778 58096
rect 62630 57608 62686 57617
rect 62630 57543 62686 57552
rect 62724 57436 62776 57442
rect 62724 57378 62776 57384
rect 62632 57164 62684 57170
rect 62632 57106 62684 57112
rect 62540 57028 62592 57034
rect 62540 56970 62592 56976
rect 62552 55849 62580 56970
rect 62538 55840 62594 55849
rect 62538 55775 62594 55784
rect 62644 54761 62672 57106
rect 62736 55305 62764 57378
rect 62828 57073 62856 58602
rect 66416 58598 66444 58903
rect 100640 58802 100668 59039
rect 100628 58796 100680 58802
rect 100628 58738 100680 58744
rect 100626 58696 100682 58705
rect 100626 58631 100628 58640
rect 100680 58631 100682 58640
rect 100628 58602 100680 58608
rect 62908 58592 62960 58598
rect 62908 58534 62960 58540
rect 66404 58592 66456 58598
rect 66404 58534 66456 58540
rect 62814 57064 62870 57073
rect 62814 56999 62870 57008
rect 62920 56393 62948 58534
rect 102388 58433 102416 60234
rect 102480 60201 102508 61322
rect 102572 60745 102600 62682
rect 102756 62377 102784 64450
rect 134496 64145 134524 68190
rect 135312 68180 135364 68186
rect 135312 68122 135364 68128
rect 135036 68112 135088 68118
rect 135036 68054 135088 68060
rect 135048 67001 135076 68054
rect 135324 67545 135352 68122
rect 135310 67536 135366 67545
rect 135310 67471 135366 67480
rect 135034 66992 135090 67001
rect 135034 66927 135090 66936
rect 134668 66752 134720 66758
rect 134668 66694 134720 66700
rect 134680 65913 134708 66694
rect 135312 66480 135364 66486
rect 135310 66448 135312 66457
rect 135364 66448 135366 66457
rect 135310 66383 135366 66392
rect 134666 65904 134722 65913
rect 134666 65839 134722 65848
rect 134668 65460 134720 65466
rect 134668 65402 134720 65408
rect 134482 64136 134538 64145
rect 134482 64071 134538 64080
rect 134680 63057 134708 65402
rect 134852 65392 134904 65398
rect 134852 65334 134904 65340
rect 134864 64689 134892 65334
rect 135312 65256 135364 65262
rect 135310 65224 135312 65233
rect 135364 65224 135366 65233
rect 135310 65159 135366 65168
rect 134850 64680 134906 64689
rect 134850 64615 134906 64624
rect 135312 64168 135364 64174
rect 135312 64110 135364 64116
rect 134852 64100 134904 64106
rect 134852 64042 134904 64048
rect 134666 63048 134722 63057
rect 134666 62983 134722 62992
rect 134484 62740 134536 62746
rect 134484 62682 134536 62688
rect 102742 62368 102798 62377
rect 102742 62303 102798 62312
rect 102744 61312 102796 61318
rect 102744 61254 102796 61260
rect 102558 60736 102614 60745
rect 102558 60671 102614 60680
rect 102652 60428 102704 60434
rect 102652 60370 102704 60376
rect 102466 60192 102522 60201
rect 102466 60127 102522 60136
rect 102560 60020 102612 60026
rect 102560 59962 102612 59968
rect 102468 58796 102520 58802
rect 102468 58738 102520 58744
rect 102374 58424 102430 58433
rect 102374 58359 102430 58368
rect 65022 58288 65078 58297
rect 65022 58223 65078 58232
rect 65036 57034 65064 58223
rect 100626 57880 100682 57889
rect 100626 57815 100682 57824
rect 66402 57744 66458 57753
rect 66402 57679 66458 57688
rect 66416 57442 66444 57679
rect 100640 57442 100668 57815
rect 66404 57436 66456 57442
rect 66404 57378 66456 57384
rect 100628 57436 100680 57442
rect 100628 57378 100680 57384
rect 102376 57436 102428 57442
rect 102376 57378 102428 57384
rect 100626 57336 100682 57345
rect 100626 57271 100682 57280
rect 100640 57238 100668 57271
rect 100628 57232 100680 57238
rect 66402 57200 66458 57209
rect 66402 57135 66404 57144
rect 66456 57135 66458 57144
rect 100534 57200 100590 57209
rect 100628 57174 100680 57180
rect 100534 57135 100536 57144
rect 66404 57106 66456 57112
rect 100588 57135 100590 57144
rect 100536 57106 100588 57112
rect 65024 57028 65076 57034
rect 65024 56970 65076 56976
rect 66402 56520 66458 56529
rect 66402 56455 66458 56464
rect 62906 56384 62962 56393
rect 66416 56354 66444 56455
rect 62906 56319 62962 56328
rect 63644 56348 63696 56354
rect 63644 56290 63696 56296
rect 66404 56348 66456 56354
rect 66404 56290 66456 56296
rect 63276 55940 63328 55946
rect 63276 55882 63328 55888
rect 62722 55296 62778 55305
rect 62722 55231 62778 55240
rect 62630 54752 62686 54761
rect 62630 54687 62686 54696
rect 63288 53537 63316 55882
rect 63368 54716 63420 54722
rect 63368 54658 63420 54664
rect 30522 53528 30578 53537
rect 30522 53463 30578 53472
rect 63274 53528 63330 53537
rect 63274 53463 63330 53472
rect 30536 33642 30564 53463
rect 62816 53356 62868 53362
rect 62816 53298 62868 53304
rect 62724 51724 62776 51730
rect 62724 51666 62776 51672
rect 62736 49593 62764 51666
rect 62828 51361 62856 53298
rect 63380 52449 63408 54658
rect 63552 54444 63604 54450
rect 63552 54386 63604 54392
rect 63564 52993 63592 54386
rect 63656 54217 63684 56290
rect 102388 56121 102416 57378
rect 102480 57345 102508 58738
rect 102572 57889 102600 59962
rect 102664 58977 102692 60370
rect 102756 59521 102784 61254
rect 134496 60745 134524 62682
rect 134864 62377 134892 64042
rect 134850 62368 134906 62377
rect 134850 62303 134906 62312
rect 135324 61833 135352 64110
rect 135402 63592 135458 63601
rect 135600 63578 135628 70894
rect 136612 68254 136640 70908
rect 136600 68248 136652 68254
rect 136600 68190 136652 68196
rect 136874 65496 136930 65505
rect 136874 65431 136876 65440
rect 136928 65431 136930 65440
rect 136876 65402 136928 65408
rect 137716 65398 137744 70908
rect 138268 70894 138834 70922
rect 138268 68202 138296 70894
rect 138176 68174 138296 68202
rect 137704 65392 137756 65398
rect 137704 65334 137756 65340
rect 138176 65262 138204 68174
rect 139924 66758 139952 70908
rect 140832 68860 140884 68866
rect 140832 68802 140884 68808
rect 139912 66752 139964 66758
rect 139912 66694 139964 66700
rect 140844 65740 140872 68802
rect 141028 66486 141056 70908
rect 142132 68118 142160 70908
rect 142672 68248 142724 68254
rect 142672 68190 142724 68196
rect 142120 68112 142172 68118
rect 142120 68054 142172 68060
rect 141016 66480 141068 66486
rect 141016 66422 141068 66428
rect 142684 65740 142712 68190
rect 143236 68186 143264 70908
rect 144340 68866 144368 70908
rect 144328 68860 144380 68866
rect 144328 68802 144380 68808
rect 144512 68316 144564 68322
rect 144512 68258 144564 68264
rect 143224 68180 143276 68186
rect 143224 68122 143276 68128
rect 144524 65740 144552 68258
rect 145444 68254 145472 70908
rect 146548 68322 146576 70908
rect 146536 68316 146588 68322
rect 146536 68258 146588 68264
rect 147652 68254 147680 70908
rect 148572 70894 148862 70922
rect 145432 68248 145484 68254
rect 145432 68190 145484 68196
rect 146444 68248 146496 68254
rect 146444 68190 146496 68196
rect 147640 68248 147692 68254
rect 147640 68190 147692 68196
rect 146456 65740 146484 68190
rect 148572 65754 148600 70894
rect 148310 65726 148600 65754
rect 149952 65754 149980 70908
rect 151056 68934 151084 70908
rect 151044 68928 151096 68934
rect 151044 68870 151096 68876
rect 152056 68928 152108 68934
rect 152056 68870 152108 68876
rect 149952 65726 150150 65754
rect 152068 65740 152096 68870
rect 152160 68254 152188 70908
rect 153264 68322 153292 70908
rect 153252 68316 153304 68322
rect 153252 68258 153304 68264
rect 154368 68254 154396 70908
rect 155472 68390 155500 70908
rect 155460 68384 155512 68390
rect 155460 68326 155512 68332
rect 156576 68322 156604 70908
rect 157694 70894 157984 70922
rect 155828 68316 155880 68322
rect 155828 68258 155880 68264
rect 156564 68316 156616 68322
rect 156564 68258 156616 68264
rect 152148 68248 152200 68254
rect 152148 68190 152200 68196
rect 153896 68248 153948 68254
rect 153896 68190 153948 68196
rect 154356 68248 154408 68254
rect 154356 68190 154408 68196
rect 153908 65740 153936 68190
rect 155840 65740 155868 68258
rect 157956 68254 157984 70894
rect 158784 68866 158812 70908
rect 159888 68934 159916 70908
rect 160992 69002 161020 70908
rect 160980 68996 161032 69002
rect 160980 68938 161032 68944
rect 159876 68928 159928 68934
rect 159876 68870 159928 68876
rect 158772 68860 158824 68866
rect 158772 68802 158824 68808
rect 159508 68384 159560 68390
rect 159508 68326 159560 68332
rect 157668 68248 157720 68254
rect 157668 68190 157720 68196
rect 157944 68248 157996 68254
rect 157944 68190 157996 68196
rect 157680 65740 157708 68190
rect 159520 65740 159548 68326
rect 161440 68316 161492 68322
rect 161440 68258 161492 68264
rect 163280 68316 163332 68322
rect 163280 68258 163332 68264
rect 161452 65740 161480 68258
rect 163292 65740 163320 68258
rect 164396 68254 164424 70908
rect 165120 68860 165172 68866
rect 165120 68802 165172 68808
rect 164384 68248 164436 68254
rect 164384 68190 164436 68196
rect 165132 65740 165160 68802
rect 165500 68798 165528 70908
rect 166604 69002 166632 70908
rect 167708 69070 167736 70908
rect 167696 69064 167748 69070
rect 167696 69006 167748 69012
rect 166592 68996 166644 69002
rect 166592 68938 166644 68944
rect 168812 68934 168840 70908
rect 168892 69200 168944 69206
rect 168892 69142 168944 69148
rect 168800 68928 168852 68934
rect 168800 68870 168852 68876
rect 167052 68860 167104 68866
rect 167052 68802 167104 68808
rect 165488 68792 165540 68798
rect 165488 68734 165540 68740
rect 167064 65740 167092 68802
rect 168904 65740 168932 69142
rect 169916 68866 169944 70908
rect 169904 68860 169956 68866
rect 169904 68802 169956 68808
rect 171020 68322 171048 70908
rect 171008 68316 171060 68322
rect 171008 68258 171060 68264
rect 172124 68254 172152 70908
rect 173228 68662 173256 70908
rect 174136 69064 174188 69070
rect 174136 69006 174188 69012
rect 173860 68928 173912 68934
rect 173860 68870 173912 68876
rect 173216 68656 173268 68662
rect 173216 68598 173268 68604
rect 169444 68248 169496 68254
rect 169444 68190 169496 68196
rect 172112 68248 172164 68254
rect 172112 68190 172164 68196
rect 138164 65256 138216 65262
rect 138164 65198 138216 65204
rect 136874 64544 136930 64553
rect 136874 64479 136930 64488
rect 136888 64106 136916 64479
rect 136968 64168 137020 64174
rect 136966 64136 136968 64145
rect 137020 64136 137022 64145
rect 136876 64100 136928 64106
rect 136966 64071 137022 64080
rect 136876 64042 136928 64048
rect 169456 64038 169484 68190
rect 173872 65913 173900 68870
rect 173952 68860 174004 68866
rect 173952 68802 174004 68808
rect 173964 66457 173992 68802
rect 174044 68316 174096 68322
rect 174044 68258 174096 68264
rect 174056 67001 174084 68258
rect 174042 66992 174098 67001
rect 174042 66927 174098 66936
rect 173950 66448 174006 66457
rect 173950 66383 174006 66392
rect 173858 65904 173914 65913
rect 173858 65839 173914 65848
rect 172662 65632 172718 65641
rect 172662 65567 172664 65576
rect 172716 65567 172718 65576
rect 172664 65538 172716 65544
rect 174148 65233 174176 69006
rect 174228 68996 174280 69002
rect 174228 68938 174280 68944
rect 174134 65224 174190 65233
rect 174134 65159 174190 65168
rect 174240 64689 174268 68938
rect 174332 68730 174360 70908
rect 174412 68792 174464 68798
rect 174412 68734 174464 68740
rect 174320 68724 174372 68730
rect 174320 68666 174372 68672
rect 174226 64680 174282 64689
rect 174226 64615 174282 64624
rect 172662 64544 172718 64553
rect 172662 64479 172718 64488
rect 172676 64378 172704 64479
rect 172664 64372 172716 64378
rect 172664 64314 172716 64320
rect 174228 64372 174280 64378
rect 174228 64314 174280 64320
rect 171834 64136 171890 64145
rect 171834 64071 171836 64080
rect 171888 64071 171890 64080
rect 171836 64042 171888 64048
rect 169444 64032 169496 64038
rect 169444 63974 169496 63980
rect 174136 64032 174188 64038
rect 174136 63974 174188 63980
rect 174148 63601 174176 63974
rect 135458 63550 135628 63578
rect 174134 63592 174190 63601
rect 135402 63527 135458 63536
rect 174134 63527 174190 63536
rect 136874 63320 136930 63329
rect 136874 63255 136930 63264
rect 172662 63320 172718 63329
rect 172662 63255 172718 63264
rect 136888 62678 136916 63255
rect 172676 63018 172704 63255
rect 172664 63012 172716 63018
rect 172664 62954 172716 62960
rect 174136 63012 174188 63018
rect 174136 62954 174188 62960
rect 172662 62912 172718 62921
rect 172662 62847 172718 62856
rect 136966 62776 137022 62785
rect 172676 62746 172704 62847
rect 136966 62711 136968 62720
rect 137020 62711 137022 62720
rect 172664 62740 172716 62746
rect 136968 62682 137020 62688
rect 172664 62682 172716 62688
rect 135404 62672 135456 62678
rect 135404 62614 135456 62620
rect 136876 62672 136928 62678
rect 136876 62614 136928 62620
rect 135310 61824 135366 61833
rect 135310 61759 135366 61768
rect 135312 61312 135364 61318
rect 135416 61289 135444 62614
rect 136782 62096 136838 62105
rect 136782 62031 136838 62040
rect 172662 62096 172718 62105
rect 172662 62031 172718 62040
rect 135312 61254 135364 61260
rect 135402 61280 135458 61289
rect 135036 60972 135088 60978
rect 135036 60914 135088 60920
rect 134482 60736 134538 60745
rect 134482 60671 134538 60680
rect 135048 60201 135076 60914
rect 135034 60192 135090 60201
rect 135034 60127 135090 60136
rect 134484 60088 134536 60094
rect 134484 60030 134536 60036
rect 102742 59512 102798 59521
rect 102742 59447 102798 59456
rect 102650 58968 102706 58977
rect 102650 58903 102706 58912
rect 102652 58660 102704 58666
rect 102652 58602 102704 58608
rect 102558 57880 102614 57889
rect 102558 57815 102614 57824
rect 102466 57336 102522 57345
rect 102466 57271 102522 57280
rect 102468 57232 102520 57238
rect 102468 57174 102520 57180
rect 100626 56112 100682 56121
rect 100626 56047 100682 56056
rect 102374 56112 102430 56121
rect 102374 56047 102430 56056
rect 66402 55976 66458 55985
rect 100640 55946 100668 56047
rect 66402 55911 66404 55920
rect 66456 55911 66458 55920
rect 100628 55940 100680 55946
rect 66404 55882 66456 55888
rect 100628 55882 100680 55888
rect 102376 55940 102428 55946
rect 102376 55882 102428 55888
rect 100902 55840 100958 55849
rect 100902 55775 100904 55784
rect 100956 55775 100958 55784
rect 100904 55746 100956 55752
rect 66310 55296 66366 55305
rect 66310 55231 66366 55240
rect 66324 54450 66352 55231
rect 100626 54888 100682 54897
rect 100626 54823 100628 54832
rect 100680 54823 100682 54832
rect 100628 54794 100680 54800
rect 66402 54752 66458 54761
rect 66402 54687 66404 54696
rect 66456 54687 66458 54696
rect 66404 54658 66456 54664
rect 100810 54616 100866 54625
rect 100810 54551 100812 54560
rect 100864 54551 100866 54560
rect 100812 54522 100864 54528
rect 102388 54489 102416 55882
rect 102480 55577 102508 57174
rect 102560 57164 102612 57170
rect 102560 57106 102612 57112
rect 102466 55568 102522 55577
rect 102466 55503 102522 55512
rect 102572 55033 102600 57106
rect 102664 56665 102692 58602
rect 134496 58433 134524 60030
rect 135036 59884 135088 59890
rect 135036 59826 135088 59832
rect 135048 58977 135076 59826
rect 135324 59521 135352 61254
rect 135402 61215 135458 61224
rect 136796 60978 136824 62031
rect 171834 61688 171890 61697
rect 171834 61623 171890 61632
rect 136874 61416 136930 61425
rect 136874 61351 136930 61360
rect 136888 61318 136916 61351
rect 171848 61318 171876 61623
rect 172676 61522 172704 62031
rect 172664 61516 172716 61522
rect 172664 61458 172716 61464
rect 136876 61312 136928 61318
rect 136876 61254 136928 61260
rect 171836 61312 171888 61318
rect 174148 61289 174176 62954
rect 174240 62377 174268 64314
rect 174424 64145 174452 68734
rect 175056 68180 175108 68186
rect 175056 68122 175108 68128
rect 175068 67545 175096 68122
rect 177184 67780 177212 73727
rect 177630 72568 177686 72577
rect 177630 72503 177686 72512
rect 177644 72402 177672 72503
rect 177632 72396 177684 72402
rect 177632 72338 177684 72344
rect 177354 71480 177410 71489
rect 177354 71415 177410 71424
rect 177368 70974 177396 71415
rect 177356 70968 177408 70974
rect 177356 70910 177408 70916
rect 177736 67780 177764 74951
rect 178288 67780 178316 76175
rect 178840 67780 178868 77399
rect 179392 67780 179420 77846
rect 179484 76657 179512 83422
rect 179576 81417 179604 84782
rect 179656 84772 179708 84778
rect 179656 84714 179708 84720
rect 179562 81408 179618 81417
rect 179562 81343 179618 81352
rect 179668 78969 179696 84714
rect 179760 83729 179788 86074
rect 179746 83720 179802 83729
rect 179746 83655 179802 83664
rect 179748 82324 179800 82330
rect 179748 82266 179800 82272
rect 179654 78960 179710 78969
rect 179654 78895 179710 78904
rect 179470 76648 179526 76657
rect 179470 76583 179526 76592
rect 179760 74345 179788 82266
rect 180300 80624 180352 80630
rect 180300 80566 180352 80572
rect 180024 79264 180076 79270
rect 180024 79206 180076 79212
rect 179746 74336 179802 74345
rect 179746 74271 179802 74280
rect 180036 67780 180064 79206
rect 180312 72033 180340 80566
rect 180944 72396 180996 72402
rect 180944 72338 180996 72344
rect 180298 72024 180354 72033
rect 180298 71959 180354 71968
rect 180956 70922 180984 72338
rect 180576 70900 180628 70906
rect 180956 70894 181076 70922
rect 180576 70842 180628 70848
rect 180588 67780 180616 70842
rect 181048 67794 181076 70894
rect 182796 70894 183132 70922
rect 183256 70894 183500 70922
rect 182796 69002 182824 70894
rect 182876 70696 182928 70702
rect 182876 70638 182928 70644
rect 181680 68996 181732 69002
rect 181680 68938 181732 68944
rect 182784 68996 182836 69002
rect 182784 68938 182836 68944
rect 181048 67766 181154 67794
rect 181692 67780 181720 68938
rect 182232 68588 182284 68594
rect 182232 68530 182284 68536
rect 182244 67780 182272 68530
rect 182888 67780 182916 70638
rect 183256 68594 183284 70894
rect 183854 70702 183882 70908
rect 183992 70894 184328 70922
rect 184452 70894 184696 70922
rect 184820 70894 185064 70922
rect 185188 70894 185524 70922
rect 185740 70894 185892 70922
rect 183842 70696 183894 70702
rect 183842 70638 183894 70644
rect 183244 68588 183296 68594
rect 183244 68530 183296 68536
rect 183992 68338 184020 70894
rect 183716 68310 184020 68338
rect 183716 67794 183744 68310
rect 184452 67794 184480 70894
rect 184820 67794 184848 70894
rect 185188 69154 185216 70894
rect 183454 67766 183744 67794
rect 184006 67766 184480 67794
rect 184558 67766 184848 67794
rect 185096 69126 185216 69154
rect 185096 67780 185124 69126
rect 185740 67780 185768 70894
rect 186246 70650 186274 70908
rect 186720 70894 186872 70922
rect 187088 70894 187240 70922
rect 187456 70894 187792 70922
rect 187916 70894 188160 70922
rect 188284 70894 188528 70922
rect 188652 70894 188988 70922
rect 189112 70894 189356 70922
rect 186246 70622 186320 70650
rect 186292 67780 186320 70622
rect 186844 67780 186872 70894
rect 187212 67794 187240 70894
rect 187764 69154 187792 70894
rect 187764 69126 187976 69154
rect 187212 67766 187410 67794
rect 187948 67780 187976 69126
rect 188132 67794 188160 70894
rect 188500 67930 188528 70894
rect 188960 68338 188988 70894
rect 189328 69177 189356 70894
rect 189466 70702 189494 70908
rect 189834 70770 189862 70908
rect 190308 70894 190460 70922
rect 189822 70764 189874 70770
rect 189822 70706 189874 70712
rect 189454 70696 189506 70702
rect 189454 70638 189506 70644
rect 190432 69614 190460 70894
rect 190616 70894 190676 70922
rect 191136 70894 191380 70922
rect 191504 70894 191748 70922
rect 190420 69608 190472 69614
rect 190420 69550 190472 69556
rect 189314 69168 189370 69177
rect 189314 69103 189370 69112
rect 190234 69168 190290 69177
rect 190234 69103 190290 69112
rect 188960 68310 189356 68338
rect 188500 67902 188804 67930
rect 188776 67794 188804 67902
rect 189328 67794 189356 68310
rect 188132 67766 188606 67794
rect 188776 67766 189158 67794
rect 189328 67766 189710 67794
rect 190248 67780 190276 69103
rect 190616 68798 190644 70894
rect 190788 70696 190840 70702
rect 190788 70638 190840 70644
rect 190604 68792 190656 68798
rect 190604 68734 190656 68740
rect 190800 67780 190828 70638
rect 191352 69177 191380 70894
rect 191432 70764 191484 70770
rect 191432 70706 191484 70712
rect 191338 69168 191394 69177
rect 191338 69103 191394 69112
rect 191444 67780 191472 70706
rect 191720 69682 191748 70894
rect 191858 70702 191886 70908
rect 192332 70894 192576 70922
rect 192700 70894 192944 70922
rect 193068 70894 193404 70922
rect 193528 70894 193772 70922
rect 193896 70894 194140 70922
rect 194264 70894 194600 70922
rect 191846 70696 191898 70702
rect 191846 70638 191898 70644
rect 191708 69676 191760 69682
rect 191708 69618 191760 69624
rect 191984 69608 192036 69614
rect 191984 69550 192036 69556
rect 191996 67780 192024 69550
rect 192548 69206 192576 70894
rect 192536 69200 192588 69206
rect 192536 69142 192588 69148
rect 192916 69138 192944 70894
rect 193086 69168 193142 69177
rect 192904 69132 192956 69138
rect 193086 69103 193142 69112
rect 192904 69074 192956 69080
rect 192536 68792 192588 68798
rect 192536 68734 192588 68740
rect 192548 67780 192576 68734
rect 193100 67780 193128 69103
rect 193376 69002 193404 70894
rect 193640 69676 193692 69682
rect 193640 69618 193692 69624
rect 193364 68996 193416 69002
rect 193364 68938 193416 68944
rect 193652 67780 193680 69618
rect 193744 68934 193772 70894
rect 194112 69070 194140 70894
rect 194284 70696 194336 70702
rect 194284 70638 194336 70644
rect 194100 69064 194152 69070
rect 194100 69006 194152 69012
rect 193732 68928 193784 68934
rect 193732 68870 193784 68876
rect 194296 67780 194324 70638
rect 194572 69342 194600 70894
rect 194664 70894 194724 70922
rect 195092 70894 195336 70922
rect 195460 70894 195796 70922
rect 195920 70894 196164 70922
rect 196288 70894 196532 70922
rect 196656 70894 196992 70922
rect 197116 70894 197360 70922
rect 194560 69336 194612 69342
rect 194560 69278 194612 69284
rect 194664 68662 194692 70894
rect 194836 69200 194888 69206
rect 194836 69142 194888 69148
rect 194652 68656 194704 68662
rect 194652 68598 194704 68604
rect 194848 67780 194876 69142
rect 195308 68798 195336 70894
rect 195388 69132 195440 69138
rect 195388 69074 195440 69080
rect 195296 68792 195348 68798
rect 195296 68734 195348 68740
rect 195400 67780 195428 69074
rect 195768 68866 195796 70894
rect 196136 69410 196164 70894
rect 196124 69404 196176 69410
rect 196124 69346 196176 69352
rect 196504 69274 196532 70894
rect 196492 69268 196544 69274
rect 196492 69210 196544 69216
rect 196964 69206 196992 70894
rect 196952 69200 197004 69206
rect 196952 69142 197004 69148
rect 197332 69070 197360 70894
rect 197424 70894 197484 70922
rect 197852 70894 198188 70922
rect 198312 70894 198556 70922
rect 198680 70894 198924 70922
rect 197424 69138 197452 70894
rect 197688 69336 197740 69342
rect 197688 69278 197740 69284
rect 197412 69132 197464 69138
rect 197412 69074 197464 69080
rect 197136 69064 197188 69070
rect 197136 69006 197188 69012
rect 197320 69064 197372 69070
rect 197320 69006 197372 69012
rect 195940 68996 195992 69002
rect 195940 68938 195992 68944
rect 195756 68860 195808 68866
rect 195756 68802 195808 68808
rect 195952 67780 195980 68938
rect 196492 68928 196544 68934
rect 196492 68870 196544 68876
rect 196504 67780 196532 68870
rect 197148 67780 197176 69006
rect 197700 67780 197728 69278
rect 198160 69002 198188 70894
rect 198528 69478 198556 70894
rect 198896 69546 198924 70894
rect 201012 69546 201040 90863
rect 201090 77600 201146 77609
rect 201090 77535 201146 77544
rect 204494 77600 204550 77609
rect 204494 77535 204550 77544
rect 198884 69540 198936 69546
rect 198884 69482 198936 69488
rect 201000 69540 201052 69546
rect 201000 69482 201052 69488
rect 198516 69472 198568 69478
rect 198516 69414 198568 69420
rect 199988 69404 200040 69410
rect 199988 69346 200040 69352
rect 198148 68996 198200 69002
rect 198148 68938 198200 68944
rect 199344 68860 199396 68866
rect 199344 68802 199396 68808
rect 198792 68792 198844 68798
rect 198792 68734 198844 68740
rect 198240 68656 198292 68662
rect 198240 68598 198292 68604
rect 198252 67780 198280 68598
rect 198804 67780 198832 68734
rect 199356 67780 199384 68802
rect 200000 67780 200028 69346
rect 201104 69342 201132 77535
rect 203944 69608 203996 69614
rect 203944 69550 203996 69556
rect 203024 69472 203076 69478
rect 203076 69420 203156 69426
rect 203024 69414 203156 69420
rect 203036 69398 203156 69414
rect 201092 69336 201144 69342
rect 201090 69304 201092 69313
rect 201144 69304 201146 69313
rect 200540 69268 200592 69274
rect 201090 69239 201146 69248
rect 200540 69210 200592 69216
rect 200552 67780 200580 69210
rect 201092 69200 201144 69206
rect 201092 69142 201144 69148
rect 201104 67780 201132 69142
rect 201828 69132 201880 69138
rect 201828 69074 201880 69080
rect 201644 69064 201696 69070
rect 201644 69006 201696 69012
rect 201656 67780 201684 69006
rect 201840 67794 201868 69074
rect 202840 68996 202892 69002
rect 202840 68938 202892 68944
rect 201840 67766 202222 67794
rect 202852 67780 202880 68938
rect 203128 67794 203156 69398
rect 203128 67766 203418 67794
rect 203956 67780 203984 69550
rect 204508 67780 204536 77535
rect 210580 69342 210608 70908
rect 215916 69546 215944 70908
rect 215904 69540 215956 69546
rect 215904 69482 215956 69488
rect 210568 69336 210620 69342
rect 210568 69278 210620 69284
rect 221252 68866 221280 70908
rect 205140 68860 205192 68866
rect 205140 68802 205192 68808
rect 221240 68860 221292 68866
rect 221240 68802 221292 68808
rect 175054 67536 175110 67545
rect 175054 67471 175110 67480
rect 175332 65596 175384 65602
rect 175332 65538 175384 65544
rect 174410 64136 174466 64145
rect 174410 64071 174466 64080
rect 175240 64100 175292 64106
rect 175240 64042 175292 64048
rect 174320 62740 174372 62746
rect 174320 62682 174372 62688
rect 174226 62368 174282 62377
rect 174226 62303 174282 62312
rect 174228 61516 174280 61522
rect 174228 61458 174280 61464
rect 171836 61254 171888 61260
rect 174134 61280 174190 61289
rect 174134 61215 174190 61224
rect 136784 60972 136836 60978
rect 136784 60914 136836 60920
rect 136782 60872 136838 60881
rect 136782 60807 136838 60816
rect 172202 60872 172258 60881
rect 172202 60807 172258 60816
rect 135404 59952 135456 59958
rect 135404 59894 135456 59900
rect 135310 59512 135366 59521
rect 135310 59447 135366 59456
rect 135034 58968 135090 58977
rect 135034 58903 135090 58912
rect 135312 58592 135364 58598
rect 135312 58534 135364 58540
rect 135036 58456 135088 58462
rect 134482 58424 134538 58433
rect 135036 58398 135088 58404
rect 134482 58359 134538 58368
rect 135048 57345 135076 58398
rect 135034 57336 135090 57345
rect 135034 57271 135090 57280
rect 134760 57164 134812 57170
rect 134760 57106 134812 57112
rect 102650 56656 102706 56665
rect 102650 56591 102706 56600
rect 102652 55804 102704 55810
rect 102652 55746 102704 55752
rect 134208 55804 134260 55810
rect 134208 55746 134260 55752
rect 102558 55024 102614 55033
rect 102558 54959 102614 54968
rect 102468 54852 102520 54858
rect 102468 54794 102520 54800
rect 102374 54480 102430 54489
rect 66312 54444 66364 54450
rect 102374 54415 102430 54424
rect 66312 54386 66364 54392
rect 63642 54208 63698 54217
rect 63642 54143 63698 54152
rect 66402 54208 66458 54217
rect 66402 54143 66458 54152
rect 65298 53528 65354 53537
rect 65298 53463 65354 53472
rect 65312 53362 65340 53463
rect 65300 53356 65352 53362
rect 65300 53298 65352 53304
rect 66416 53022 66444 54143
rect 100626 53664 100682 53673
rect 100626 53599 100682 53608
rect 100640 53294 100668 53599
rect 100628 53288 100680 53294
rect 102480 53265 102508 54794
rect 102560 54580 102612 54586
rect 102560 54522 102612 54528
rect 100628 53230 100680 53236
rect 102466 53256 102522 53265
rect 102466 53191 102522 53200
rect 100626 53120 100682 53129
rect 100626 53055 100628 53064
rect 100680 53055 100682 53064
rect 102376 53084 102428 53090
rect 100628 53026 100680 53032
rect 102376 53026 102428 53032
rect 63736 53016 63788 53022
rect 63550 52984 63606 52993
rect 66404 53016 66456 53022
rect 63736 52958 63788 52964
rect 66310 52984 66366 52993
rect 63550 52919 63606 52928
rect 63366 52440 63422 52449
rect 63366 52375 63422 52384
rect 63368 52132 63420 52138
rect 63368 52074 63420 52080
rect 62814 51352 62870 51361
rect 62814 51287 62870 51296
rect 62816 50500 62868 50506
rect 62816 50442 62868 50448
rect 62722 49584 62778 49593
rect 62722 49519 62778 49528
rect 62828 48505 62856 50442
rect 63380 50137 63408 52074
rect 63748 51905 63776 52958
rect 66404 52958 66456 52964
rect 66310 52919 66366 52928
rect 65298 52304 65354 52313
rect 65298 52239 65354 52248
rect 65312 52138 65340 52239
rect 65300 52132 65352 52138
rect 65300 52074 65352 52080
rect 63734 51896 63790 51905
rect 63734 51831 63790 51840
rect 65666 51760 65722 51769
rect 65666 51695 65668 51704
rect 65720 51695 65722 51704
rect 65668 51666 65720 51672
rect 66324 51662 66352 52919
rect 100626 52440 100682 52449
rect 100626 52375 100682 52384
rect 100640 52274 100668 52375
rect 100628 52268 100680 52274
rect 100628 52210 100680 52216
rect 100626 51896 100682 51905
rect 100626 51831 100682 51840
rect 100534 51760 100590 51769
rect 100640 51730 100668 51831
rect 100534 51695 100590 51704
rect 100628 51724 100680 51730
rect 100548 51662 100576 51695
rect 100628 51666 100680 51672
rect 63736 51656 63788 51662
rect 63736 51598 63788 51604
rect 66312 51656 66364 51662
rect 66312 51598 66364 51604
rect 100536 51656 100588 51662
rect 102388 51633 102416 53026
rect 102572 52721 102600 54522
rect 102664 53809 102692 55746
rect 134220 53809 134248 55746
rect 134772 55577 134800 57106
rect 135036 57096 135088 57102
rect 135036 57038 135088 57044
rect 135048 56121 135076 57038
rect 135324 56665 135352 58534
rect 135416 57889 135444 59894
rect 136796 59890 136824 60807
rect 136966 60328 137022 60337
rect 136966 60263 137022 60272
rect 136980 60094 137008 60263
rect 172216 60162 172244 60807
rect 172662 60328 172718 60337
rect 172662 60263 172664 60272
rect 172716 60263 172718 60272
rect 172664 60234 172716 60240
rect 174240 60201 174268 61458
rect 174332 60745 174360 62682
rect 175252 61833 175280 64042
rect 175344 63057 175372 65538
rect 175330 63048 175386 63057
rect 175330 62983 175386 62992
rect 175238 61824 175294 61833
rect 175238 61759 175294 61768
rect 174412 61312 174464 61318
rect 174412 61254 174464 61260
rect 174318 60736 174374 60745
rect 174318 60671 174374 60680
rect 174320 60292 174372 60298
rect 174320 60234 174372 60240
rect 174226 60192 174282 60201
rect 172204 60156 172256 60162
rect 172204 60098 172256 60104
rect 174136 60156 174188 60162
rect 174226 60127 174282 60136
rect 174136 60098 174188 60104
rect 136968 60088 137020 60094
rect 136874 60056 136930 60065
rect 136968 60030 137020 60036
rect 172662 60056 172718 60065
rect 136874 59991 136930 60000
rect 172662 59991 172664 60000
rect 136888 59958 136916 59991
rect 172716 59991 172718 60000
rect 172664 59962 172716 59968
rect 136876 59952 136928 59958
rect 136876 59894 136928 59900
rect 136784 59884 136836 59890
rect 136784 59826 136836 59832
rect 136782 59104 136838 59113
rect 136782 59039 136838 59048
rect 172202 59104 172258 59113
rect 172202 59039 172258 59048
rect 136796 58462 136824 59039
rect 172216 58938 172244 59039
rect 174148 58977 174176 60098
rect 174134 58968 174190 58977
rect 172204 58932 172256 58938
rect 174134 58903 174190 58912
rect 172204 58874 172256 58880
rect 171834 58832 171890 58841
rect 171834 58767 171836 58776
rect 171888 58767 171890 58776
rect 174228 58796 174280 58802
rect 171836 58738 171888 58744
rect 174228 58738 174280 58744
rect 136874 58696 136930 58705
rect 136874 58631 136930 58640
rect 136888 58598 136916 58631
rect 136876 58592 136928 58598
rect 136876 58534 136928 58540
rect 136784 58456 136836 58462
rect 136784 58398 136836 58404
rect 135402 57880 135458 57889
rect 135402 57815 135458 57824
rect 136782 57880 136838 57889
rect 136782 57815 136838 57824
rect 172018 57880 172074 57889
rect 172018 57815 172074 57824
rect 135404 57232 135456 57238
rect 135404 57174 135456 57180
rect 135310 56656 135366 56665
rect 135310 56591 135366 56600
rect 135034 56112 135090 56121
rect 135034 56047 135090 56056
rect 134758 55568 134814 55577
rect 134758 55503 134814 55512
rect 135036 55464 135088 55470
rect 135036 55406 135088 55412
rect 134300 54580 134352 54586
rect 134300 54522 134352 54528
rect 102650 53800 102706 53809
rect 102650 53735 102706 53744
rect 134206 53800 134262 53809
rect 134206 53735 134262 53744
rect 102744 53288 102796 53294
rect 102744 53230 102796 53236
rect 102558 52712 102614 52721
rect 102558 52647 102614 52656
rect 102652 52268 102704 52274
rect 102652 52210 102704 52216
rect 102468 51724 102520 51730
rect 102468 51666 102520 51672
rect 100536 51598 100588 51604
rect 102374 51624 102430 51633
rect 63748 50681 63776 51598
rect 102374 51559 102430 51568
rect 66402 51216 66458 51225
rect 66402 51151 66458 51160
rect 63734 50672 63790 50681
rect 66416 50642 66444 51151
rect 100626 50672 100682 50681
rect 63734 50607 63790 50616
rect 63828 50636 63880 50642
rect 63828 50578 63880 50584
rect 66404 50636 66456 50642
rect 100626 50607 100682 50616
rect 66404 50578 66456 50584
rect 63366 50128 63422 50137
rect 63366 50063 63422 50072
rect 63840 49049 63868 50578
rect 65666 50536 65722 50545
rect 100640 50506 100668 50607
rect 65666 50471 65668 50480
rect 65720 50471 65722 50480
rect 100628 50500 100680 50506
rect 65668 50442 65720 50448
rect 100628 50442 100680 50448
rect 102480 50409 102508 51666
rect 102560 51656 102612 51662
rect 102560 51598 102612 51604
rect 100626 50400 100682 50409
rect 102466 50400 102522 50409
rect 100626 50335 100628 50344
rect 100680 50335 100682 50344
rect 102376 50364 102428 50370
rect 100628 50306 100680 50312
rect 102466 50335 102522 50344
rect 102376 50306 102428 50312
rect 65482 49992 65538 50001
rect 65482 49927 65538 49936
rect 63826 49040 63882 49049
rect 63736 49004 63788 49010
rect 65496 49010 65524 49927
rect 100626 49448 100682 49457
rect 100626 49383 100682 49392
rect 66402 49312 66458 49321
rect 100640 49282 100668 49383
rect 66402 49247 66458 49256
rect 100628 49276 100680 49282
rect 63826 48975 63882 48984
rect 65484 49004 65536 49010
rect 63736 48946 63788 48952
rect 65484 48946 65536 48952
rect 63368 48936 63420 48942
rect 63368 48878 63420 48884
rect 62814 48496 62870 48505
rect 62814 48431 62870 48440
rect 62816 47508 62868 47514
rect 62816 47450 62868 47456
rect 62724 46964 62776 46970
rect 62724 46906 62776 46912
rect 62736 46193 62764 46906
rect 62722 46184 62778 46193
rect 62722 46119 62778 46128
rect 62828 45649 62856 47450
rect 62908 47440 62960 47446
rect 62908 47382 62960 47388
rect 62920 46737 62948 47382
rect 63380 47281 63408 48878
rect 63748 47825 63776 48946
rect 66416 48942 66444 49247
rect 100628 49218 100680 49224
rect 100626 49040 100682 49049
rect 100626 48975 100628 48984
rect 100680 48975 100682 48984
rect 100628 48946 100680 48952
rect 66404 48936 66456 48942
rect 66404 48878 66456 48884
rect 102388 48777 102416 50306
rect 102572 49865 102600 51598
rect 102664 50953 102692 52210
rect 102756 52177 102784 53230
rect 134312 52721 134340 54522
rect 135048 54489 135076 55406
rect 135416 55033 135444 57174
rect 136796 57102 136824 57815
rect 136874 57336 136930 57345
rect 136874 57271 136930 57280
rect 136888 57170 136916 57271
rect 136968 57232 137020 57238
rect 136966 57200 136968 57209
rect 137020 57200 137022 57209
rect 136876 57164 136928 57170
rect 172032 57170 172060 57815
rect 172662 57472 172718 57481
rect 172662 57407 172664 57416
rect 172716 57407 172718 57416
rect 172664 57378 172716 57384
rect 172662 57336 172718 57345
rect 172662 57271 172664 57280
rect 172716 57271 172718 57280
rect 172664 57242 172716 57248
rect 136966 57135 137022 57144
rect 172020 57164 172072 57170
rect 136876 57106 136928 57112
rect 172020 57106 172072 57112
rect 174136 57164 174188 57170
rect 174136 57106 174188 57112
rect 136784 57096 136836 57102
rect 136784 57038 136836 57044
rect 174148 56121 174176 57106
rect 174240 56665 174268 58738
rect 174332 58433 174360 60234
rect 174424 59521 174452 61254
rect 174504 60020 174556 60026
rect 174504 59962 174556 59968
rect 174410 59512 174466 59521
rect 174410 59447 174466 59456
rect 174318 58424 174374 58433
rect 174318 58359 174374 58368
rect 174516 57889 174544 59962
rect 174596 58932 174648 58938
rect 174596 58874 174648 58880
rect 174502 57880 174558 57889
rect 174502 57815 174558 57824
rect 174320 57436 174372 57442
rect 174320 57378 174372 57384
rect 174226 56656 174282 56665
rect 174226 56591 174282 56600
rect 136782 56112 136838 56121
rect 136782 56047 136838 56056
rect 172662 56112 172718 56121
rect 172662 56047 172664 56056
rect 136796 55470 136824 56047
rect 172716 56047 172718 56056
rect 174134 56112 174190 56121
rect 174134 56047 174190 56056
rect 174228 56076 174280 56082
rect 172664 56018 172716 56024
rect 174228 56018 174280 56024
rect 136874 55840 136930 55849
rect 136874 55775 136876 55784
rect 136928 55775 136930 55784
rect 172662 55840 172718 55849
rect 172662 55775 172664 55784
rect 136876 55746 136928 55752
rect 172716 55775 172718 55784
rect 172664 55746 172716 55752
rect 136784 55464 136836 55470
rect 136784 55406 136836 55412
rect 135402 55024 135458 55033
rect 135402 54959 135458 54968
rect 136782 54888 136838 54897
rect 136782 54823 136838 54832
rect 172110 54888 172166 54897
rect 172110 54823 172166 54832
rect 135034 54480 135090 54489
rect 135034 54415 135090 54424
rect 136796 53974 136824 54823
rect 137150 54616 137206 54625
rect 172124 54586 172152 54823
rect 172662 54616 172718 54625
rect 137150 54551 137152 54560
rect 137204 54551 137206 54560
rect 172112 54580 172164 54586
rect 137152 54522 137204 54528
rect 172662 54551 172718 54560
rect 172112 54522 172164 54528
rect 172676 54518 172704 54551
rect 172664 54512 172716 54518
rect 174240 54489 174268 56018
rect 174332 55577 174360 57378
rect 174608 57345 174636 58874
rect 174594 57336 174650 57345
rect 174412 57300 174464 57306
rect 174594 57271 174650 57280
rect 174412 57242 174464 57248
rect 174318 55568 174374 55577
rect 174318 55503 174374 55512
rect 174424 55033 174452 57242
rect 174964 55804 175016 55810
rect 174964 55746 175016 55752
rect 174410 55024 174466 55033
rect 174410 54959 174466 54968
rect 174780 54580 174832 54586
rect 174780 54522 174832 54528
rect 172664 54454 172716 54460
rect 174226 54480 174282 54489
rect 174226 54415 174282 54424
rect 135128 53968 135180 53974
rect 135128 53910 135180 53916
rect 136784 53968 136836 53974
rect 136784 53910 136836 53916
rect 135140 53265 135168 53910
rect 136782 53664 136838 53673
rect 136782 53599 136838 53608
rect 171650 53664 171706 53673
rect 171650 53599 171706 53608
rect 135126 53256 135182 53265
rect 135126 53191 135182 53200
rect 135404 53016 135456 53022
rect 135404 52958 135456 52964
rect 134298 52712 134354 52721
rect 134298 52647 134354 52656
rect 135128 52608 135180 52614
rect 135128 52550 135180 52556
rect 135140 52177 135168 52550
rect 102742 52168 102798 52177
rect 102742 52103 102798 52112
rect 135126 52168 135182 52177
rect 135126 52103 135182 52112
rect 135312 51656 135364 51662
rect 135416 51633 135444 52958
rect 136796 52614 136824 53599
rect 171664 53226 171692 53599
rect 174792 53265 174820 54522
rect 174976 53809 175004 55746
rect 175332 54512 175384 54518
rect 175332 54454 175384 54460
rect 174962 53800 175018 53809
rect 174962 53735 175018 53744
rect 172662 53256 172718 53265
rect 171652 53220 171704 53226
rect 174778 53256 174834 53265
rect 172662 53191 172718 53200
rect 174136 53220 174188 53226
rect 171652 53162 171704 53168
rect 136874 53120 136930 53129
rect 172676 53090 172704 53191
rect 174778 53191 174834 53200
rect 174136 53162 174188 53168
rect 136874 53055 136930 53064
rect 172664 53084 172716 53090
rect 136888 53022 136916 53055
rect 172664 53026 172716 53032
rect 136876 53016 136928 53022
rect 136876 52958 136928 52964
rect 136784 52608 136836 52614
rect 136784 52550 136836 52556
rect 136690 52440 136746 52449
rect 136690 52375 136746 52384
rect 172018 52440 172074 52449
rect 172018 52375 172074 52384
rect 135312 51598 135364 51604
rect 135402 51624 135458 51633
rect 135036 51384 135088 51390
rect 135036 51326 135088 51332
rect 102650 50944 102706 50953
rect 102650 50879 102706 50888
rect 102652 50500 102704 50506
rect 102652 50442 102704 50448
rect 102558 49856 102614 49865
rect 102558 49791 102614 49800
rect 102664 49321 102692 50442
rect 135048 50409 135076 51326
rect 135034 50400 135090 50409
rect 135034 50335 135090 50344
rect 134852 50228 134904 50234
rect 134852 50170 134904 50176
rect 134864 49321 134892 50170
rect 135324 49865 135352 51598
rect 135402 51559 135458 51568
rect 136704 51118 136732 52375
rect 136782 51896 136838 51905
rect 136782 51831 136838 51840
rect 136796 51390 136824 51831
rect 136874 51760 136930 51769
rect 136874 51695 136930 51704
rect 136888 51662 136916 51695
rect 172032 51662 172060 52375
rect 174148 52177 174176 53162
rect 174504 53084 174556 53090
rect 174504 53026 174556 53032
rect 174134 52168 174190 52177
rect 174134 52103 174190 52112
rect 172570 52032 172626 52041
rect 172570 51967 172572 51976
rect 172624 51967 172626 51976
rect 174320 51996 174372 52002
rect 172572 51938 172624 51944
rect 174320 51938 174372 51944
rect 172662 51896 172718 51905
rect 172662 51831 172664 51840
rect 172716 51831 172718 51840
rect 172664 51802 172716 51808
rect 136876 51656 136928 51662
rect 136876 51598 136928 51604
rect 172020 51656 172072 51662
rect 172020 51598 172072 51604
rect 174228 51656 174280 51662
rect 174228 51598 174280 51604
rect 136784 51384 136836 51390
rect 136784 51326 136836 51332
rect 135404 51112 135456 51118
rect 135404 51054 135456 51060
rect 136692 51112 136744 51118
rect 136692 51054 136744 51060
rect 135416 50953 135444 51054
rect 174240 50953 174268 51598
rect 135402 50944 135458 50953
rect 135402 50879 135458 50888
rect 174226 50944 174282 50953
rect 174226 50879 174282 50888
rect 172202 50808 172258 50817
rect 172202 50743 172258 50752
rect 136782 50672 136838 50681
rect 136782 50607 136838 50616
rect 135404 50296 135456 50302
rect 135404 50238 135456 50244
rect 135310 49856 135366 49865
rect 135310 49791 135366 49800
rect 102650 49312 102706 49321
rect 102468 49276 102520 49282
rect 102650 49247 102706 49256
rect 134850 49312 134906 49321
rect 134850 49247 134906 49256
rect 102468 49218 102520 49224
rect 64930 48768 64986 48777
rect 64930 48703 64986 48712
rect 102374 48768 102430 48777
rect 102374 48703 102430 48712
rect 63734 47816 63790 47825
rect 63734 47751 63790 47760
rect 64944 47446 64972 48703
rect 100626 48360 100682 48369
rect 100626 48295 100682 48304
rect 100640 47922 100668 48295
rect 102480 48097 102508 49218
rect 102560 49004 102612 49010
rect 102560 48946 102612 48952
rect 102466 48088 102522 48097
rect 102466 48023 102522 48032
rect 100628 47916 100680 47922
rect 100628 47858 100680 47864
rect 65022 47816 65078 47825
rect 65022 47751 65078 47760
rect 64932 47440 64984 47446
rect 64932 47382 64984 47388
rect 63366 47272 63422 47281
rect 63366 47207 63422 47216
rect 65036 46970 65064 47751
rect 100626 47680 100682 47689
rect 100626 47615 100628 47624
rect 100680 47615 100682 47624
rect 102376 47644 102428 47650
rect 100628 47586 100680 47592
rect 102376 47586 102428 47592
rect 65666 47544 65722 47553
rect 65666 47479 65668 47488
rect 65720 47479 65722 47488
rect 100626 47544 100682 47553
rect 100626 47479 100628 47488
rect 65668 47450 65720 47456
rect 100680 47479 100682 47488
rect 100628 47450 100680 47456
rect 66402 47000 66458 47009
rect 65024 46964 65076 46970
rect 66402 46935 66458 46944
rect 65024 46906 65076 46912
rect 62906 46728 62962 46737
rect 62906 46663 62962 46672
rect 66416 46426 66444 46935
rect 102388 46465 102416 47586
rect 102572 47553 102600 48946
rect 135312 48868 135364 48874
rect 135312 48810 135364 48816
rect 134760 48460 134812 48466
rect 134760 48402 134812 48408
rect 102652 47916 102704 47922
rect 102652 47858 102704 47864
rect 102558 47544 102614 47553
rect 102468 47508 102520 47514
rect 102558 47479 102614 47488
rect 102468 47450 102520 47456
rect 100626 46456 100682 46465
rect 63736 46420 63788 46426
rect 63736 46362 63788 46368
rect 66404 46420 66456 46426
rect 100626 46391 100682 46400
rect 102374 46456 102430 46465
rect 102374 46391 102430 46400
rect 66404 46362 66456 46368
rect 62814 45640 62870 45649
rect 62814 45575 62870 45584
rect 63748 44969 63776 46362
rect 65206 46320 65262 46329
rect 100640 46290 100668 46391
rect 65206 46255 65262 46264
rect 100628 46284 100680 46290
rect 63734 44960 63790 44969
rect 63734 44895 63790 44904
rect 63736 44856 63788 44862
rect 63736 44798 63788 44804
rect 63644 44788 63696 44794
rect 63644 44730 63696 44736
rect 62816 44720 62868 44726
rect 62816 44662 62868 44668
rect 62828 44425 62856 44662
rect 62814 44416 62870 44425
rect 62814 44351 62870 44360
rect 63656 43337 63684 44730
rect 63748 43881 63776 44798
rect 65220 44726 65248 46255
rect 100628 46226 100680 46232
rect 100902 46184 100958 46193
rect 100902 46119 100904 46128
rect 100956 46119 100958 46128
rect 102376 46148 102428 46154
rect 100904 46090 100956 46096
rect 102376 46090 102428 46096
rect 66310 45776 66366 45785
rect 66310 45711 66366 45720
rect 66324 44862 66352 45711
rect 100534 45368 100590 45377
rect 100534 45303 100590 45312
rect 100548 45270 100576 45303
rect 100536 45264 100588 45270
rect 66402 45232 66458 45241
rect 100536 45206 100588 45212
rect 66402 45167 66458 45176
rect 66312 44856 66364 44862
rect 66312 44798 66364 44804
rect 66416 44794 66444 45167
rect 99982 45096 100038 45105
rect 99982 45031 100038 45040
rect 99996 44998 100024 45031
rect 99984 44992 100036 44998
rect 99984 44934 100036 44940
rect 66404 44788 66456 44794
rect 66404 44730 66456 44736
rect 65208 44720 65260 44726
rect 102388 44697 102416 46090
rect 102480 45921 102508 47450
rect 102664 47009 102692 47858
rect 134772 47553 134800 48402
rect 135324 48097 135352 48810
rect 135416 48777 135444 50238
rect 136796 50234 136824 50607
rect 136874 50400 136930 50409
rect 172216 50370 172244 50743
rect 174332 50409 174360 51938
rect 174412 51860 174464 51866
rect 174412 51802 174464 51808
rect 172662 50400 172718 50409
rect 136874 50335 136930 50344
rect 172204 50364 172256 50370
rect 136888 50302 136916 50335
rect 174318 50400 174374 50409
rect 172662 50335 172718 50344
rect 174136 50364 174188 50370
rect 172204 50306 172256 50312
rect 172676 50302 172704 50335
rect 174318 50335 174374 50344
rect 174136 50306 174188 50312
rect 136876 50296 136928 50302
rect 136876 50238 136928 50244
rect 172664 50296 172716 50302
rect 172664 50238 172716 50244
rect 136784 50228 136836 50234
rect 136784 50170 136836 50176
rect 136874 49448 136930 49457
rect 136874 49383 136930 49392
rect 172662 49448 172718 49457
rect 172662 49383 172718 49392
rect 136888 48942 136916 49383
rect 172676 49282 172704 49383
rect 174148 49321 174176 50306
rect 174320 50296 174372 50302
rect 174320 50238 174372 50244
rect 174134 49312 174190 49321
rect 172664 49276 172716 49282
rect 174134 49247 174190 49256
rect 174228 49276 174280 49282
rect 172664 49218 172716 49224
rect 174228 49218 174280 49224
rect 171834 49176 171890 49185
rect 171834 49111 171836 49120
rect 171888 49111 171890 49120
rect 171836 49082 171888 49088
rect 136876 48936 136928 48942
rect 136782 48904 136838 48913
rect 136876 48878 136928 48884
rect 136782 48839 136838 48848
rect 135402 48768 135458 48777
rect 135402 48703 135458 48712
rect 136796 48466 136824 48839
rect 136784 48460 136836 48466
rect 136784 48402 136836 48408
rect 136690 48360 136746 48369
rect 136690 48295 136746 48304
rect 172570 48360 172626 48369
rect 172570 48295 172626 48304
rect 135310 48088 135366 48097
rect 135310 48023 135366 48032
rect 134758 47544 134814 47553
rect 134758 47479 134814 47488
rect 135404 47508 135456 47514
rect 135404 47450 135456 47456
rect 134852 47372 134904 47378
rect 134852 47314 134904 47320
rect 102650 47000 102706 47009
rect 102650 46935 102706 46944
rect 134864 46465 134892 47314
rect 135312 47168 135364 47174
rect 135312 47110 135364 47116
rect 135324 47009 135352 47110
rect 135310 47000 135366 47009
rect 135310 46935 135366 46944
rect 134850 46456 134906 46465
rect 134850 46391 134906 46400
rect 102560 46284 102612 46290
rect 102560 46226 102612 46232
rect 102466 45912 102522 45921
rect 102466 45847 102522 45856
rect 102468 45264 102520 45270
rect 102572 45241 102600 46226
rect 134668 46080 134720 46086
rect 134668 46022 134720 46028
rect 134680 45241 134708 46022
rect 135416 45921 135444 47450
rect 136704 47174 136732 48295
rect 172584 47922 172612 48295
rect 174240 48097 174268 49218
rect 174332 48777 174360 50238
rect 174424 49865 174452 51802
rect 174516 51633 174544 53026
rect 175344 52721 175372 54454
rect 175330 52712 175386 52721
rect 175330 52647 175386 52656
rect 174502 51624 174558 51633
rect 174502 51559 174558 51568
rect 174410 49856 174466 49865
rect 174410 49791 174466 49800
rect 174412 49140 174464 49146
rect 174412 49082 174464 49088
rect 174318 48768 174374 48777
rect 174318 48703 174374 48712
rect 174226 48088 174282 48097
rect 174226 48023 174282 48032
rect 172662 47952 172718 47961
rect 172572 47916 172624 47922
rect 172662 47887 172718 47896
rect 174228 47916 174280 47922
rect 172572 47858 172624 47864
rect 172676 47786 172704 47887
rect 174228 47858 174280 47864
rect 172664 47780 172716 47786
rect 172664 47722 172716 47728
rect 174136 47780 174188 47786
rect 174136 47722 174188 47728
rect 136782 47680 136838 47689
rect 136782 47615 136838 47624
rect 172662 47680 172718 47689
rect 172662 47615 172664 47624
rect 136796 47378 136824 47615
rect 172716 47615 172718 47624
rect 172664 47586 172716 47592
rect 136874 47544 136930 47553
rect 136874 47479 136876 47488
rect 136928 47479 136930 47488
rect 136876 47450 136928 47456
rect 136784 47372 136836 47378
rect 136784 47314 136836 47320
rect 136692 47168 136744 47174
rect 136692 47110 136744 47116
rect 172662 46592 172718 46601
rect 172662 46527 172664 46536
rect 172716 46527 172718 46536
rect 172664 46498 172716 46504
rect 174148 46465 174176 47722
rect 174240 47009 174268 47858
rect 174320 47644 174372 47650
rect 174320 47586 174372 47592
rect 174226 47000 174282 47009
rect 174226 46935 174282 46944
rect 174228 46556 174280 46562
rect 174228 46498 174280 46504
rect 136782 46456 136838 46465
rect 136782 46391 136838 46400
rect 174134 46456 174190 46465
rect 174134 46391 174190 46400
rect 136796 46086 136824 46391
rect 137518 46184 137574 46193
rect 137518 46119 137574 46128
rect 172662 46184 172718 46193
rect 172662 46119 172664 46128
rect 136784 46080 136836 46086
rect 136784 46022 136836 46028
rect 135402 45912 135458 45921
rect 135402 45847 135458 45856
rect 136690 45368 136746 45377
rect 136690 45303 136746 45312
rect 102468 45206 102520 45212
rect 102558 45232 102614 45241
rect 65208 44662 65260 44668
rect 102374 44688 102430 44697
rect 102374 44623 102430 44632
rect 66218 44552 66274 44561
rect 66218 44487 66274 44496
rect 63734 43872 63790 43881
rect 63734 43807 63790 43816
rect 66232 43570 66260 44487
rect 102480 44153 102508 45206
rect 102558 45167 102614 45176
rect 134666 45232 134722 45241
rect 134666 45167 134722 45176
rect 102560 44992 102612 44998
rect 102560 44934 102612 44940
rect 99890 44144 99946 44153
rect 102466 44144 102522 44153
rect 99890 44079 99892 44088
rect 99944 44079 99946 44088
rect 102284 44108 102336 44114
rect 99892 44050 99944 44056
rect 102466 44079 102522 44088
rect 102284 44050 102336 44056
rect 66402 44008 66458 44017
rect 66402 43943 66458 43952
rect 63736 43564 63788 43570
rect 63736 43506 63788 43512
rect 66220 43564 66272 43570
rect 66220 43506 66272 43512
rect 63642 43328 63698 43337
rect 63642 43263 63698 43272
rect 63748 42793 63776 43506
rect 66416 43366 66444 43943
rect 100626 43464 100682 43473
rect 100626 43399 100682 43408
rect 100640 43366 100668 43399
rect 63828 43360 63880 43366
rect 66404 43360 66456 43366
rect 63828 43302 63880 43308
rect 66310 43328 66366 43337
rect 63734 42784 63790 42793
rect 63734 42719 63790 42728
rect 63840 42521 63868 43302
rect 66404 43302 66456 43308
rect 100628 43360 100680 43366
rect 100628 43302 100680 43308
rect 66310 43263 66366 43272
rect 63826 42512 63882 42521
rect 63826 42447 63882 42456
rect 63828 42340 63880 42346
rect 63828 42282 63880 42288
rect 63736 42000 63788 42006
rect 63736 41942 63788 41948
rect 63748 41569 63776 41942
rect 63734 41560 63790 41569
rect 63734 41495 63790 41504
rect 63840 41025 63868 42282
rect 66324 42006 66352 43263
rect 102296 43065 102324 44050
rect 102572 43609 102600 44934
rect 135036 44720 135088 44726
rect 135034 44688 135036 44697
rect 135088 44688 135090 44697
rect 135034 44623 135090 44632
rect 136704 44454 136732 45303
rect 136782 44960 136838 44969
rect 136782 44895 136838 44904
rect 135404 44448 135456 44454
rect 135404 44390 135456 44396
rect 136692 44448 136744 44454
rect 136692 44390 136744 44396
rect 135036 44312 135088 44318
rect 135036 44254 135088 44260
rect 135048 43609 135076 44254
rect 135416 44153 135444 44390
rect 136796 44318 136824 44895
rect 137532 44726 137560 46119
rect 172716 46119 172718 46128
rect 172664 46090 172716 46096
rect 171650 45368 171706 45377
rect 171650 45303 171706 45312
rect 171664 44998 171692 45303
rect 174240 45241 174268 46498
rect 174332 45921 174360 47586
rect 174424 47553 174452 49082
rect 174410 47544 174466 47553
rect 174410 47479 174466 47488
rect 175332 46148 175384 46154
rect 175332 46090 175384 46096
rect 174318 45912 174374 45921
rect 174318 45847 174374 45856
rect 174226 45232 174282 45241
rect 174226 45167 174282 45176
rect 171652 44992 171704 44998
rect 171652 44934 171704 44940
rect 171834 44960 171890 44969
rect 171834 44895 171890 44904
rect 171848 44794 171876 44895
rect 171836 44788 171888 44794
rect 171836 44730 171888 44736
rect 174780 44788 174832 44794
rect 174780 44730 174832 44736
rect 137520 44720 137572 44726
rect 137520 44662 137572 44668
rect 136784 44312 136836 44318
rect 136784 44254 136836 44260
rect 135402 44144 135458 44153
rect 135402 44079 135458 44088
rect 136782 44144 136838 44153
rect 136782 44079 136838 44088
rect 172662 44144 172718 44153
rect 172662 44079 172718 44088
rect 102558 43600 102614 43609
rect 102558 43535 102614 43544
rect 135034 43600 135090 43609
rect 135034 43535 135090 43544
rect 102376 43292 102428 43298
rect 102376 43234 102428 43240
rect 134944 43292 134996 43298
rect 134944 43234 134996 43240
rect 102282 43056 102338 43065
rect 102282 42991 102338 43000
rect 100626 42920 100682 42929
rect 100626 42855 100682 42864
rect 66402 42784 66458 42793
rect 66402 42719 66458 42728
rect 66416 42346 66444 42719
rect 100640 42686 100668 42855
rect 100628 42680 100680 42686
rect 100628 42622 100680 42628
rect 102388 42385 102416 43234
rect 102560 42680 102612 42686
rect 102560 42622 102612 42628
rect 100626 42376 100682 42385
rect 66404 42340 66456 42346
rect 100626 42311 100682 42320
rect 102374 42376 102430 42385
rect 102374 42311 102430 42320
rect 66404 42282 66456 42288
rect 66402 42240 66458 42249
rect 100640 42210 100668 42311
rect 66402 42175 66458 42184
rect 100628 42204 100680 42210
rect 66312 42000 66364 42006
rect 66312 41942 66364 41948
rect 63826 41016 63882 41025
rect 63826 40951 63882 40960
rect 66416 40578 66444 42175
rect 100628 42146 100680 42152
rect 102468 42204 102520 42210
rect 102468 42146 102520 42152
rect 100626 42104 100682 42113
rect 100626 42039 100628 42048
rect 100680 42039 100682 42048
rect 102376 42068 102428 42074
rect 100628 42010 100680 42016
rect 102376 42010 102428 42016
rect 71628 41926 71964 41954
rect 79080 41926 79416 41954
rect 63184 40572 63236 40578
rect 63184 40514 63236 40520
rect 66404 40572 66456 40578
rect 66404 40514 66456 40520
rect 63196 40481 63224 40514
rect 63182 40472 63238 40481
rect 63182 40407 63238 40416
rect 66402 40472 66458 40481
rect 66402 40407 66458 40416
rect 66312 39892 66364 39898
rect 66312 39834 66364 39840
rect 62814 39520 62870 39529
rect 62814 39455 62870 39464
rect 62828 39218 62856 39455
rect 62816 39212 62868 39218
rect 62816 39154 62868 39160
rect 30524 33636 30576 33642
rect 30524 33578 30576 33584
rect 66220 33636 66272 33642
rect 66220 33578 66272 33584
rect 66232 32729 66260 33578
rect 66218 32720 66274 32729
rect 66218 32655 66274 32664
rect 66324 24705 66352 39834
rect 66310 24696 66366 24705
rect 66310 24631 66366 24640
rect 13318 19664 13374 19673
rect 13318 19599 13374 19608
rect 66416 16817 66444 40407
rect 71936 39966 71964 41926
rect 71924 39960 71976 39966
rect 71924 39902 71976 39908
rect 72568 39212 72620 39218
rect 72568 39154 72620 39160
rect 72580 36786 72608 39154
rect 79388 37790 79416 41926
rect 86288 41926 86624 41954
rect 94016 41926 94076 41954
rect 82504 39960 82556 39966
rect 82504 39902 82556 39908
rect 79376 37784 79428 37790
rect 79376 37726 79428 37732
rect 82516 36786 82544 39902
rect 86288 39898 86316 41926
rect 94016 40481 94044 41926
rect 102388 40753 102416 42010
rect 102480 41297 102508 42146
rect 102572 41841 102600 42622
rect 134956 42385 134984 43234
rect 136796 43094 136824 44079
rect 172676 43638 172704 44079
rect 172664 43632 172716 43638
rect 172570 43600 172626 43609
rect 172664 43574 172716 43580
rect 174044 43632 174096 43638
rect 174792 43609 174820 44730
rect 175344 44697 175372 46090
rect 175424 44992 175476 44998
rect 175424 44934 175476 44940
rect 175330 44688 175386 44697
rect 175330 44623 175386 44632
rect 175436 44153 175464 44934
rect 175422 44144 175478 44153
rect 175422 44079 175478 44088
rect 174044 43574 174096 43580
rect 174778 43600 174834 43609
rect 172570 43535 172626 43544
rect 136874 43464 136930 43473
rect 136874 43399 136930 43408
rect 136888 43366 136916 43399
rect 172584 43366 172612 43535
rect 136876 43360 136928 43366
rect 136876 43302 136928 43308
rect 172572 43360 172624 43366
rect 172572 43302 172624 43308
rect 135404 43088 135456 43094
rect 135402 43056 135404 43065
rect 136784 43088 136836 43094
rect 135456 43056 135458 43065
rect 174056 43065 174084 43574
rect 174778 43535 174834 43544
rect 174136 43292 174188 43298
rect 174136 43234 174188 43240
rect 136784 43030 136836 43036
rect 174042 43056 174098 43065
rect 135402 42991 135458 43000
rect 174042 42991 174098 43000
rect 136690 42920 136746 42929
rect 136690 42855 136746 42864
rect 172202 42920 172258 42929
rect 172202 42855 172258 42864
rect 134942 42376 134998 42385
rect 134942 42311 134998 42320
rect 135404 41932 135456 41938
rect 135404 41874 135456 41880
rect 135312 41864 135364 41870
rect 102558 41832 102614 41841
rect 102558 41767 102614 41776
rect 135310 41832 135312 41841
rect 135364 41832 135366 41841
rect 135310 41767 135366 41776
rect 134852 41524 134904 41530
rect 134852 41466 134904 41472
rect 102466 41288 102522 41297
rect 102466 41223 102522 41232
rect 134864 40753 134892 41466
rect 135416 41297 135444 41874
rect 136704 41870 136732 42855
rect 136874 42376 136930 42385
rect 172216 42346 172244 42855
rect 174148 42385 174176 43234
rect 172662 42376 172718 42385
rect 136874 42311 136930 42320
rect 172204 42340 172256 42346
rect 136782 42104 136838 42113
rect 136782 42039 136838 42048
rect 136692 41864 136744 41870
rect 136692 41806 136744 41812
rect 136796 41530 136824 42039
rect 136888 42006 136916 42311
rect 172662 42311 172718 42320
rect 174134 42376 174190 42385
rect 174134 42311 174190 42320
rect 174228 42340 174280 42346
rect 172204 42282 172256 42288
rect 172676 42210 172704 42311
rect 174228 42282 174280 42288
rect 172664 42204 172716 42210
rect 172664 42146 172716 42152
rect 172662 42104 172718 42113
rect 172662 42039 172664 42048
rect 172716 42039 172718 42048
rect 174136 42068 174188 42074
rect 172664 42010 172716 42016
rect 174136 42010 174188 42016
rect 136876 42000 136928 42006
rect 136876 41942 136928 41948
rect 136784 41524 136836 41530
rect 136784 41466 136836 41472
rect 135402 41288 135458 41297
rect 135402 41223 135458 41232
rect 102374 40744 102430 40753
rect 102374 40679 102430 40688
rect 134850 40744 134906 40753
rect 134850 40679 134906 40688
rect 94002 40472 94058 40481
rect 94002 40407 94058 40416
rect 102374 40200 102430 40209
rect 102374 40135 102430 40144
rect 86276 39892 86328 39898
rect 86276 39834 86328 39840
rect 102388 39218 102416 40135
rect 109642 40064 109698 40073
rect 109532 40022 109642 40050
rect 109642 39999 109698 40008
rect 143604 39966 143632 41940
rect 143592 39960 143644 39966
rect 118824 39886 118884 39914
rect 93176 39212 93228 39218
rect 93176 39154 93228 39160
rect 102376 39212 102428 39218
rect 102376 39154 102428 39160
rect 93188 36786 93216 39154
rect 72580 36758 72916 36786
rect 82516 36758 82852 36786
rect 92880 36758 93216 36786
rect 118856 33642 118884 39886
rect 127780 39886 128116 39914
rect 143592 39902 143644 39908
rect 138072 39892 138124 39898
rect 127780 37790 127808 39886
rect 138072 39834 138124 39840
rect 134482 39656 134538 39665
rect 134482 39591 134538 39600
rect 134496 39218 134524 39591
rect 134484 39212 134536 39218
rect 134484 39154 134536 39160
rect 127768 37784 127820 37790
rect 127768 37726 127820 37732
rect 118844 33636 118896 33642
rect 118844 33578 118896 33584
rect 136876 33636 136928 33642
rect 136876 33578 136928 33584
rect 136888 33409 136916 33578
rect 136874 33400 136930 33409
rect 136874 33335 136930 33344
rect 138084 25113 138112 39834
rect 138162 39792 138218 39801
rect 138162 39727 138218 39736
rect 138070 25104 138126 25113
rect 138070 25039 138126 25048
rect 138176 17089 138204 39727
rect 144880 39212 144932 39218
rect 144880 39154 144932 39160
rect 144892 36772 144920 39154
rect 151056 37790 151084 41940
rect 154816 39960 154868 39966
rect 154816 39902 154868 39908
rect 151044 37784 151096 37790
rect 151044 37726 151096 37732
rect 154828 36772 154856 39902
rect 158600 39898 158628 41940
rect 158588 39892 158640 39898
rect 158588 39834 158640 39840
rect 166052 39801 166080 41940
rect 174148 40753 174176 42010
rect 174240 41841 174268 42282
rect 174320 42204 174372 42210
rect 174320 42146 174372 42152
rect 174226 41832 174282 41841
rect 174226 41767 174282 41776
rect 174332 41297 174360 42146
rect 174318 41288 174374 41297
rect 174318 41223 174374 41232
rect 174134 40744 174190 40753
rect 174134 40679 174190 40688
rect 181402 40064 181458 40073
rect 181458 40022 181522 40050
rect 181402 39999 181458 40008
rect 166038 39792 166094 39801
rect 166038 39727 166094 39736
rect 174134 39520 174190 39529
rect 174134 39455 174190 39464
rect 174148 39218 174176 39455
rect 164844 39212 164896 39218
rect 164844 39154 164896 39160
rect 174136 39212 174188 39218
rect 174136 39154 174188 39160
rect 164856 36772 164884 39154
rect 190800 37722 190828 39900
rect 200092 37790 200120 39900
rect 200080 37784 200132 37790
rect 200080 37726 200132 37732
rect 205152 37722 205180 68802
rect 222540 44561 222568 141902
rect 222816 127550 222844 142038
rect 222908 139761 222936 146782
rect 223552 141966 223580 149479
rect 223540 141960 223592 141966
rect 223540 141902 223592 141908
rect 222894 139752 222950 139761
rect 222894 139687 222950 139696
rect 222804 127544 222856 127550
rect 222804 127486 222856 127492
rect 222712 124824 222764 124830
rect 222712 124766 222764 124772
rect 222724 116210 222752 124766
rect 222724 116182 223028 116210
rect 222710 115952 222766 115961
rect 222710 115887 222766 115896
rect 222620 115100 222672 115106
rect 222620 115042 222672 115048
rect 222632 103290 222660 115042
rect 222724 110278 222752 115887
rect 223000 115106 223028 116182
rect 222988 115100 223040 115106
rect 222988 115042 223040 115048
rect 222712 110272 222764 110278
rect 222712 110214 222764 110220
rect 222804 107960 222856 107966
rect 222724 107908 222804 107914
rect 222724 107902 222856 107908
rect 222724 107886 222844 107902
rect 222724 103426 222752 107886
rect 224472 105761 224500 163487
rect 224458 105752 224514 105761
rect 224458 105687 224514 105696
rect 222724 103398 223028 103426
rect 222632 103262 222752 103290
rect 222724 97034 222752 103262
rect 223000 97154 223028 103398
rect 222988 97148 223040 97154
rect 222988 97090 223040 97096
rect 223540 97148 223592 97154
rect 223540 97090 223592 97096
rect 222724 97006 222844 97034
rect 222816 92598 222844 97006
rect 223552 96377 223580 97090
rect 223538 96368 223594 96377
rect 223538 96303 223594 96312
rect 222804 92592 222856 92598
rect 222804 92534 222856 92540
rect 223540 92592 223592 92598
rect 223540 92534 223592 92540
rect 223552 92161 223580 92534
rect 223538 92152 223594 92161
rect 223538 92087 223594 92096
rect 223538 85216 223594 85225
rect 223538 85151 223594 85160
rect 223552 84846 223580 85151
rect 222804 84840 222856 84846
rect 222724 84788 222804 84794
rect 222724 84782 222856 84788
rect 223540 84840 223592 84846
rect 223540 84782 223592 84788
rect 222724 84766 222844 84782
rect 222724 73642 222752 84766
rect 223538 75288 223594 75297
rect 223538 75223 223594 75232
rect 223552 75122 223580 75223
rect 222988 75116 223040 75122
rect 222988 75058 223040 75064
rect 223540 75116 223592 75122
rect 223540 75058 223592 75064
rect 222724 73626 222844 73642
rect 222724 73620 222856 73626
rect 222724 73614 222804 73620
rect 222804 73562 222856 73568
rect 223000 68066 223028 75058
rect 223080 73620 223132 73626
rect 223080 73562 223132 73568
rect 223092 68361 223120 73562
rect 223078 68352 223134 68361
rect 223078 68287 223134 68296
rect 222632 68038 223028 68066
rect 222632 63986 222660 68038
rect 222632 63958 222752 63986
rect 222526 44552 222582 44561
rect 222526 44487 222582 44496
rect 222724 40730 222752 63958
rect 222540 40702 222752 40730
rect 222540 40594 222568 40702
rect 222448 40566 222568 40594
rect 222448 40458 222476 40566
rect 222448 40430 222568 40458
rect 222540 37790 222568 40430
rect 222528 37784 222580 37790
rect 222528 37726 222580 37732
rect 190788 37716 190840 37722
rect 190788 37658 190840 37664
rect 205140 37716 205192 37722
rect 205140 37658 205192 37664
rect 222712 28196 222764 28202
rect 222712 28138 222764 28144
rect 222724 20761 222752 28138
rect 222710 20752 222766 20761
rect 222710 20687 222766 20696
rect 138162 17080 138218 17089
rect 138162 17015 138218 17024
rect 66402 16808 66458 16817
rect 66402 16743 66458 16752
rect 71292 12822 71628 12850
rect 71292 10998 71320 12822
rect 79066 12630 79094 12836
rect 86624 12822 86960 12850
rect 77996 12624 78048 12630
rect 77996 12566 78048 12572
rect 79054 12624 79106 12630
rect 79054 12566 79106 12572
rect 23532 10992 23584 10998
rect 23532 10934 23584 10940
rect 71280 10992 71332 10998
rect 71280 10934 71332 10940
rect 23544 9304 23572 10934
rect 50764 10924 50816 10930
rect 50764 10866 50816 10872
rect 50776 9304 50804 10866
rect 78008 9304 78036 12566
rect 86932 11746 86960 12822
rect 94016 12822 94076 12850
rect 86920 11740 86972 11746
rect 86920 11682 86972 11688
rect 94016 11678 94044 12822
rect 132552 11740 132604 11746
rect 132552 11682 132604 11688
rect 94004 11672 94056 11678
rect 94004 11614 94056 11620
rect 105228 10992 105280 10998
rect 105228 10934 105280 10940
rect 105240 9304 105268 10934
rect 132564 9304 132592 11682
rect 143604 10930 143632 12836
rect 151056 10998 151084 12836
rect 151044 10992 151096 10998
rect 151044 10934 151096 10940
rect 143592 10924 143644 10930
rect 143592 10866 143644 10872
rect 158600 10454 158628 12836
rect 166052 11746 166080 12836
rect 166040 11740 166092 11746
rect 166040 11682 166092 11688
rect 214248 11740 214300 11746
rect 214248 11682 214300 11688
rect 187016 11672 187068 11678
rect 187016 11614 187068 11620
rect 158588 10448 158640 10454
rect 158588 10390 158640 10396
rect 159784 10448 159836 10454
rect 159784 10390 159836 10396
rect 159796 9304 159824 10390
rect 187028 9304 187056 11614
rect 214260 9304 214288 11682
rect 23530 8824 23586 9304
rect 50762 8824 50818 9304
rect 77994 8824 78050 9304
rect 105226 8824 105282 9304
rect 132550 8824 132606 9304
rect 159782 8824 159838 9304
rect 187014 8824 187070 9304
rect 214246 8824 214302 9304
<< via2 >>
rect 98234 238704 98290 238760
rect 169994 238704 170050 238760
rect 12030 235848 12086 235904
rect 11938 214224 11994 214280
rect 55822 217216 55878 217272
rect 62538 215312 62594 215368
rect 62630 214632 62686 214688
rect 63642 213952 63698 214008
rect 62538 213292 62594 213328
rect 62538 213272 62540 213292
rect 62540 213272 62592 213292
rect 62592 213272 62594 213292
rect 98326 230680 98382 230736
rect 168522 230136 168578 230192
rect 98418 222792 98474 222848
rect 135402 215584 135458 215640
rect 102374 215312 102430 215368
rect 102558 214652 102614 214688
rect 102558 214632 102560 214652
rect 102560 214632 102612 214652
rect 102612 214632 102614 214652
rect 135402 214652 135458 214688
rect 135402 214632 135404 214652
rect 135404 214632 135456 214652
rect 135456 214632 135458 214652
rect 103110 213952 103166 214008
rect 135402 213952 135458 214008
rect 100994 213816 101050 213872
rect 65022 213408 65078 213464
rect 62354 212592 62410 212648
rect 62630 211912 62686 211968
rect 66402 212728 66458 212784
rect 102374 213272 102430 213328
rect 135034 213292 135090 213328
rect 135034 213272 135036 213292
rect 135036 213272 135088 213292
rect 135088 213272 135090 213292
rect 136782 213272 136838 213328
rect 151042 215856 151098 215912
rect 223078 234896 223134 234952
rect 170086 222812 170142 222848
rect 170086 222792 170088 222812
rect 170088 222792 170140 222812
rect 170140 222792 170142 222812
rect 174226 215720 174282 215776
rect 174042 214632 174098 214688
rect 174226 213952 174282 214008
rect 172018 213816 172074 213872
rect 174042 213272 174098 213328
rect 100994 212728 101050 212784
rect 136874 212728 136930 212784
rect 102466 212592 102522 212648
rect 135402 212592 135458 212648
rect 100534 212048 100590 212104
rect 102374 211932 102430 211968
rect 102374 211912 102376 211932
rect 102376 211912 102428 211932
rect 102428 211912 102430 211932
rect 65022 211776 65078 211832
rect 62538 211232 62594 211288
rect 62630 210552 62686 210608
rect 65666 211504 65722 211560
rect 100810 211504 100866 211560
rect 65022 210552 65078 210608
rect 64930 210416 64986 210472
rect 62630 209892 62686 209928
rect 62630 209872 62632 209892
rect 62632 209872 62684 209892
rect 62684 209872 62686 209892
rect 135402 211932 135458 211968
rect 135402 211912 135404 211932
rect 135404 211912 135456 211932
rect 135456 211912 135458 211932
rect 172662 213036 172664 213056
rect 172664 213036 172716 213056
rect 172716 213036 172718 213056
rect 172662 213000 172718 213036
rect 174226 212592 174282 212648
rect 172662 212456 172718 212512
rect 137058 212048 137114 212104
rect 174042 211912 174098 211968
rect 172662 211640 172718 211696
rect 136966 211504 137022 211560
rect 172386 211268 172388 211288
rect 172388 211268 172440 211288
rect 172440 211268 172442 211288
rect 172386 211232 172442 211268
rect 174226 211232 174282 211288
rect 100994 210960 101050 211016
rect 136874 210960 136930 211016
rect 103662 210844 103718 210880
rect 103662 210824 103664 210844
rect 103664 210824 103716 210844
rect 103716 210824 103718 210844
rect 65666 210416 65722 210472
rect 102374 210572 102430 210608
rect 102374 210552 102376 210572
rect 102376 210552 102428 210572
rect 102428 210552 102430 210572
rect 134666 210572 134722 210608
rect 172662 210588 172664 210608
rect 172664 210588 172716 210608
rect 172716 210588 172718 210608
rect 134666 210552 134668 210572
rect 134668 210552 134720 210572
rect 134720 210552 134722 210572
rect 172662 210552 172718 210588
rect 174042 210552 174098 210608
rect 65482 210280 65538 210336
rect 100902 210280 100958 210336
rect 65022 209328 65078 209384
rect 62722 209192 62778 209248
rect 172662 210044 172664 210064
rect 172664 210044 172716 210064
rect 172716 210044 172718 210064
rect 172662 210008 172718 210044
rect 174134 209872 174190 209928
rect 100994 209736 101050 209792
rect 136874 209736 136930 209792
rect 171650 209364 171652 209384
rect 171652 209364 171704 209384
rect 171704 209364 171706 209384
rect 171650 209328 171706 209364
rect 135310 209192 135366 209248
rect 174594 209192 174650 209248
rect 66402 209056 66458 209112
rect 62630 208512 62686 208568
rect 63642 207832 63698 207888
rect 172110 208784 172166 208840
rect 65850 208512 65906 208568
rect 137702 208512 137758 208568
rect 66402 207968 66458 208024
rect 135402 207852 135458 207888
rect 135402 207832 135404 207852
rect 135404 207832 135456 207852
rect 135456 207832 135458 207852
rect 65022 207560 65078 207616
rect 65850 207560 65906 207616
rect 65298 207288 65354 207344
rect 136874 207288 136930 207344
rect 62538 207152 62594 207208
rect 174134 207152 174190 207208
rect 65666 206764 65722 206800
rect 65666 206744 65668 206764
rect 65668 206744 65720 206764
rect 65720 206744 65722 206764
rect 171650 206608 171706 206664
rect 62630 206472 62686 206528
rect 135402 206472 135458 206528
rect 174042 206472 174098 206528
rect 62630 205792 62686 205848
rect 136874 206064 136930 206120
rect 171834 205964 171836 205984
rect 171836 205964 171888 205984
rect 171888 205964 171890 205984
rect 171834 205928 171890 205964
rect 66402 205520 66458 205576
rect 64930 205248 64986 205304
rect 62630 204432 62686 204488
rect 65666 204332 65668 204352
rect 65668 204332 65720 204352
rect 65720 204332 65722 204352
rect 65666 204296 65722 204332
rect 62538 203752 62594 203808
rect 65482 203752 65538 203808
rect 100902 200660 100904 200680
rect 100904 200660 100956 200680
rect 100956 200660 100958 200680
rect 100902 200624 100958 200660
rect 136782 200624 136838 200680
rect 65022 200352 65078 200408
rect 66402 200352 66458 200408
rect 102374 200352 102430 200408
rect 135402 200352 135458 200408
rect 65114 200080 65170 200136
rect 66402 199536 66458 199592
rect 136782 199400 136838 199456
rect 172202 199420 172258 199456
rect 172202 199400 172204 199420
rect 172204 199400 172256 199420
rect 172256 199400 172258 199420
rect 65114 199264 65170 199320
rect 100902 199300 100904 199320
rect 100904 199300 100956 199320
rect 100956 199300 100958 199320
rect 100902 199264 100958 199300
rect 62354 198992 62410 199048
rect 102374 198992 102430 199048
rect 134758 198992 134814 199048
rect 175238 198992 175294 199048
rect 172202 198060 172258 198096
rect 172202 198040 172204 198060
rect 172204 198040 172256 198060
rect 172256 198040 172258 198060
rect 65022 197904 65078 197960
rect 100902 197924 100958 197960
rect 100902 197904 100904 197924
rect 100904 197904 100956 197924
rect 100956 197904 100958 197924
rect 136782 197904 136838 197960
rect 62630 197632 62686 197688
rect 102374 197632 102430 197688
rect 135402 197632 135458 197688
rect 174226 197632 174282 197688
rect 65022 196816 65078 196872
rect 172662 196836 172718 196872
rect 172662 196816 172664 196836
rect 172664 196816 172716 196836
rect 172716 196816 172718 196836
rect 62630 196272 62686 196328
rect 63642 195592 63698 195648
rect 100902 196700 100958 196736
rect 100902 196680 100904 196700
rect 100904 196680 100956 196700
rect 100956 196680 100958 196700
rect 136782 196680 136838 196736
rect 172202 196700 172258 196736
rect 172202 196680 172204 196700
rect 172204 196680 172256 196700
rect 172256 196680 172258 196700
rect 66402 196564 66458 196600
rect 66402 196544 66404 196564
rect 66404 196544 66456 196564
rect 66456 196544 66458 196564
rect 100902 196564 100958 196600
rect 100902 196544 100904 196564
rect 100904 196544 100956 196564
rect 100956 196544 100958 196564
rect 136690 196544 136746 196600
rect 102374 196272 102430 196328
rect 135402 196272 135458 196328
rect 174134 196272 174190 196328
rect 174226 196136 174282 196192
rect 134298 196036 134300 196056
rect 134300 196036 134352 196056
rect 134352 196036 134354 196056
rect 134298 196000 134354 196036
rect 65022 195592 65078 195648
rect 102466 195592 102522 195648
rect 171466 195612 171522 195648
rect 171466 195592 171468 195612
rect 171468 195592 171520 195612
rect 171520 195592 171522 195612
rect 100718 195456 100774 195512
rect 136874 195456 136930 195512
rect 66402 195320 66458 195376
rect 100902 195204 100958 195240
rect 100902 195184 100904 195204
rect 100904 195184 100956 195204
rect 100956 195184 100958 195204
rect 62630 194948 62632 194968
rect 62632 194948 62684 194968
rect 62684 194948 62686 194968
rect 62630 194912 62686 194948
rect 65114 194776 65170 194832
rect 65022 194368 65078 194424
rect 62538 194232 62594 194288
rect 136782 195184 136838 195240
rect 102466 194912 102522 194968
rect 135402 194912 135458 194968
rect 172662 195204 172718 195240
rect 172662 195184 172664 195204
rect 172664 195184 172716 195204
rect 172716 195184 172718 195204
rect 174134 194912 174190 194968
rect 135402 194812 135404 194832
rect 135404 194812 135456 194832
rect 135456 194812 135458 194832
rect 135402 194776 135458 194812
rect 174226 194776 174282 194832
rect 100626 194252 100682 194288
rect 100626 194232 100628 194252
rect 100628 194232 100680 194252
rect 100680 194232 100682 194252
rect 102374 194232 102430 194288
rect 136782 194232 136838 194288
rect 171558 194252 171614 194288
rect 171558 194232 171560 194252
rect 171560 194232 171612 194252
rect 171612 194232 171614 194252
rect 65114 193824 65170 193880
rect 100626 193844 100682 193880
rect 100626 193824 100628 193844
rect 100628 193824 100680 193844
rect 100680 193824 100682 193844
rect 66402 193552 66458 193608
rect 62354 192872 62410 192928
rect 12214 192600 12270 192656
rect 65022 192600 65078 192656
rect 12030 179680 12086 179736
rect 12122 170976 12178 171032
rect 12030 149760 12086 149816
rect 11938 105696 11994 105752
rect 11938 75096 11994 75152
rect 64930 192464 64986 192520
rect 62538 192228 62540 192248
rect 62540 192228 62592 192248
rect 62592 192228 62594 192248
rect 62538 192192 62594 192228
rect 99706 193144 99762 193200
rect 136690 193824 136746 193880
rect 102466 193552 102522 193608
rect 135402 193552 135458 193608
rect 172662 193960 172718 194016
rect 174134 193552 174190 193608
rect 135402 193452 135404 193472
rect 135404 193452 135456 193472
rect 135456 193452 135458 193472
rect 135402 193416 135458 193452
rect 174226 193416 174282 193472
rect 136782 193144 136838 193200
rect 171650 193144 171706 193200
rect 102374 192872 102430 192928
rect 66402 192464 66458 192520
rect 100626 192484 100682 192520
rect 100626 192464 100628 192484
rect 100628 192464 100680 192484
rect 100680 192464 100682 192484
rect 66402 192328 66458 192384
rect 66310 191784 66366 191840
rect 62354 191548 62356 191568
rect 62356 191548 62408 191568
rect 62408 191548 62410 191568
rect 62354 191512 62410 191548
rect 65022 191240 65078 191296
rect 65206 191104 65262 191160
rect 62630 190868 62632 190888
rect 62632 190868 62684 190888
rect 62684 190868 62686 190888
rect 62630 190832 62686 190868
rect 62446 190152 62502 190208
rect 62630 189508 62632 189528
rect 62632 189508 62684 189528
rect 62684 189508 62686 189528
rect 62630 189472 62686 189508
rect 62630 188792 62686 188848
rect 65022 189608 65078 189664
rect 99890 191940 99946 191976
rect 99890 191920 99892 191940
rect 99892 191920 99944 191940
rect 99944 191920 99946 191940
rect 66402 191240 66458 191296
rect 100626 191260 100682 191296
rect 100626 191240 100628 191260
rect 100628 191240 100680 191260
rect 100680 191240 100682 191260
rect 100902 191104 100958 191160
rect 66310 190560 66366 190616
rect 136690 192464 136746 192520
rect 102466 192192 102522 192248
rect 172202 192736 172258 192792
rect 135402 192192 135458 192248
rect 223538 211096 223594 211152
rect 207898 201712 207954 201768
rect 207254 192464 207310 192520
rect 207254 192328 207310 192384
rect 174226 192192 174282 192248
rect 134298 192056 134354 192112
rect 174134 192056 174190 192112
rect 136782 191920 136838 191976
rect 172202 191920 172258 191976
rect 102374 191512 102430 191568
rect 136690 191240 136746 191296
rect 102282 190832 102338 190888
rect 100534 190152 100590 190208
rect 102190 190152 102246 190208
rect 66402 190016 66458 190072
rect 99890 189880 99946 189936
rect 66310 189608 66366 189664
rect 172662 191376 172718 191432
rect 136966 191104 137022 191160
rect 172662 191004 172664 191024
rect 172664 191004 172716 191024
rect 172716 191004 172718 191024
rect 172662 190968 172718 191004
rect 135402 190832 135458 190888
rect 174042 190832 174098 190888
rect 134758 190696 134814 190752
rect 173950 190696 174006 190752
rect 136782 190152 136838 190208
rect 172386 190172 172442 190208
rect 172386 190152 172388 190172
rect 172388 190152 172440 190172
rect 172440 190152 172442 190172
rect 102558 189472 102614 189528
rect 134298 189472 134354 189528
rect 172018 189880 172074 189936
rect 137426 189744 137482 189800
rect 134758 189236 134760 189256
rect 134760 189236 134812 189256
rect 134812 189236 134814 189256
rect 134758 189200 134814 189236
rect 102466 188792 102522 188848
rect 174962 189472 175018 189528
rect 174410 189200 174466 189256
rect 63642 188112 63698 188168
rect 102374 188112 102430 188168
rect 135034 188148 135036 188168
rect 135036 188148 135088 188168
rect 135088 188148 135090 188168
rect 135034 188112 135090 188148
rect 175422 188112 175478 188168
rect 37882 184984 37938 185040
rect 40274 184984 40330 185040
rect 37974 184440 38030 184496
rect 39630 184440 39686 184496
rect 54902 184168 54958 184224
rect 60146 184168 60202 184224
rect 31994 178184 32050 178240
rect 37422 178184 37478 178240
rect 59594 178184 59650 178240
rect 12214 170024 12270 170080
rect 105594 184712 105650 184768
rect 105594 182264 105650 182320
rect 105318 178456 105374 178512
rect 105226 177096 105282 177152
rect 105134 175736 105190 175792
rect 57570 174784 57626 174840
rect 106146 183488 106202 183544
rect 117094 185392 117150 185448
rect 116910 184712 116966 184768
rect 117462 185256 117518 185312
rect 118198 185392 118254 185448
rect 118658 185392 118714 185448
rect 118290 185120 118346 185176
rect 117646 184712 117702 184768
rect 118106 184712 118162 184768
rect 118934 185256 118990 185312
rect 119118 184984 119174 185040
rect 120590 185392 120646 185448
rect 120958 185392 121014 185448
rect 120314 185120 120370 185176
rect 120590 185120 120646 185176
rect 119670 184848 119726 184904
rect 119578 184712 119634 184768
rect 121050 185256 121106 185312
rect 121142 184984 121198 185040
rect 121694 184984 121750 185040
rect 121602 184848 121658 184904
rect 122706 184984 122762 185040
rect 122522 184712 122578 184768
rect 123442 185392 123498 185448
rect 123902 185392 123958 185448
rect 123074 185120 123130 185176
rect 123350 185120 123406 185176
rect 124362 185256 124418 185312
rect 124362 184848 124418 184904
rect 125098 185120 125154 185176
rect 124822 184984 124878 185040
rect 124914 184848 124970 184904
rect 125466 184984 125522 185040
rect 125926 185428 125928 185448
rect 125928 185428 125980 185448
rect 125980 185428 125982 185448
rect 125926 185392 125982 185428
rect 125926 185292 125928 185312
rect 125928 185292 125980 185312
rect 125980 185292 125982 185312
rect 125926 185256 125982 185292
rect 126110 185256 126166 185312
rect 126662 185392 126718 185448
rect 125650 184712 125706 184768
rect 126478 184712 126534 184768
rect 127214 185120 127270 185176
rect 127214 185020 127216 185040
rect 127216 185020 127268 185040
rect 127268 185020 127270 185040
rect 127214 184984 127270 185020
rect 127214 184884 127216 184904
rect 127216 184884 127268 184904
rect 127268 184884 127270 184904
rect 127214 184848 127270 184884
rect 120130 184576 120186 184632
rect 122798 184576 122854 184632
rect 124362 184576 124418 184632
rect 127030 184576 127086 184632
rect 131446 185256 131502 185312
rect 131630 184712 131686 184768
rect 123718 184440 123774 184496
rect 127030 184476 127032 184496
rect 127032 184476 127084 184496
rect 127084 184476 127086 184496
rect 127030 184440 127086 184476
rect 108538 183488 108594 183544
rect 108078 181176 108134 181232
rect 106054 181040 106110 181096
rect 105962 179816 106018 179872
rect 107894 178864 107950 178920
rect 106146 174396 106202 174432
rect 106146 174376 106148 174396
rect 106148 174376 106200 174396
rect 106200 174376 106202 174396
rect 105410 173696 105466 173752
rect 107894 176416 107950 176472
rect 106330 172472 106386 172528
rect 108170 174104 108226 174160
rect 107894 171792 107950 171848
rect 106422 171384 106478 171440
rect 106054 170160 106110 170216
rect 107894 169344 107950 169400
rect 105226 168800 105282 168856
rect 105962 167440 106018 167496
rect 107802 167032 107858 167088
rect 106422 166116 106424 166136
rect 106424 166116 106476 166136
rect 106476 166116 106478 166136
rect 106422 166080 106478 166116
rect 32638 164856 32694 164912
rect 37422 164856 37478 164912
rect 12214 159280 12270 159336
rect 12582 149352 12638 149408
rect 31994 151528 32050 151584
rect 12582 142552 12638 142608
rect 59594 164856 59650 164912
rect 106422 163516 106478 163552
rect 106422 163496 106424 163516
rect 106424 163496 106476 163516
rect 106476 163496 106478 163516
rect 107802 162408 107858 162464
rect 106146 162156 106202 162192
rect 106146 162136 106148 162156
rect 106148 162136 106200 162156
rect 106200 162136 106202 162156
rect 105778 160660 105834 160696
rect 105778 160640 105780 160660
rect 105780 160640 105832 160660
rect 105832 160640 105834 160660
rect 106422 159300 106478 159336
rect 106422 159280 106424 159300
rect 106424 159280 106476 159300
rect 106476 159280 106478 159300
rect 105410 158328 105466 158384
rect 105410 156988 105466 157024
rect 105410 156968 105412 156988
rect 105412 156968 105464 156988
rect 105464 156968 105466 156988
rect 105226 155764 105282 155800
rect 105226 155744 105228 155764
rect 105228 155744 105280 155764
rect 105280 155744 105282 155764
rect 57478 154792 57534 154848
rect 105778 154520 105834 154576
rect 105594 153860 105650 153896
rect 105594 153840 105596 153860
rect 105596 153840 105648 153860
rect 105648 153840 105650 153860
rect 106422 152480 106478 152536
rect 59594 151548 59650 151584
rect 59594 151528 59596 151548
rect 59596 151528 59648 151548
rect 59648 151528 59650 151548
rect 105962 149624 106018 149680
rect 105410 148400 105466 148456
rect 105226 147176 105282 147232
rect 31810 141328 31866 141384
rect 62814 142008 62870 142064
rect 62814 140920 62870 140976
rect 62722 140648 62778 140704
rect 62354 139424 62410 139480
rect 62814 139696 62870 139752
rect 62814 138880 62870 138936
rect 62538 137656 62594 137712
rect 30522 137112 30578 137168
rect 30430 127728 30486 127784
rect 12214 106104 12270 106160
rect 12122 95768 12178 95824
rect 62814 137112 62870 137168
rect 90138 141872 90194 141928
rect 91242 141328 91298 141384
rect 66218 139424 66274 139480
rect 66402 138880 66458 138936
rect 102282 142552 102338 142608
rect 100626 139016 100682 139072
rect 100534 138608 100590 138664
rect 63458 138336 63514 138392
rect 66310 138200 66366 138256
rect 100074 137792 100130 137848
rect 66402 137656 66458 137712
rect 99706 137268 99762 137304
rect 99706 137248 99708 137268
rect 99708 137248 99760 137268
rect 99760 137248 99762 137268
rect 105870 145952 105926 146008
rect 106422 144864 106478 144920
rect 106606 150984 106662 151040
rect 108538 159960 108594 160016
rect 107802 157648 107858 157704
rect 107710 155336 107766 155392
rect 107894 152888 107950 152944
rect 107250 150576 107306 150632
rect 107158 148264 107214 148320
rect 108538 145952 108594 146008
rect 132182 185392 132238 185448
rect 132366 151528 132422 151584
rect 176986 181720 177042 181776
rect 177078 180496 177134 180552
rect 177722 184168 177778 184224
rect 177446 182944 177502 183000
rect 197456 184984 197512 185040
rect 202194 184984 202250 185040
rect 198514 184440 198570 184496
rect 198882 184440 198938 184496
rect 203942 184440 203998 184496
rect 203390 184304 203446 184360
rect 180298 183488 180354 183544
rect 179746 181176 179802 181232
rect 177630 179272 177686 179328
rect 179746 178864 179802 178920
rect 177538 178048 177594 178104
rect 176986 176824 177042 176880
rect 179654 176416 179710 176472
rect 176894 175600 176950 175656
rect 177354 174396 177410 174432
rect 177354 174376 177356 174396
rect 177356 174376 177408 174396
rect 177408 174376 177410 174396
rect 176986 173152 177042 173208
rect 177538 172064 177594 172120
rect 179654 174104 179710 174160
rect 225194 187296 225250 187352
rect 207254 182944 207310 183000
rect 225194 179680 225250 179736
rect 201090 178184 201146 178240
rect 204494 178184 204550 178240
rect 179654 171792 179710 171848
rect 177722 170840 177778 170896
rect 177630 169616 177686 169672
rect 179654 169344 179710 169400
rect 178090 168392 178146 168448
rect 177538 167168 177594 167224
rect 179562 167032 179618 167088
rect 223538 169208 223594 169264
rect 177538 165944 177594 166000
rect 200998 164856 201054 164912
rect 204494 164856 204550 164912
rect 177722 163516 177778 163552
rect 177722 163496 177724 163516
rect 177724 163496 177776 163516
rect 177776 163496 177778 163516
rect 179562 162408 179618 162464
rect 176986 162272 177042 162328
rect 176986 161048 177042 161104
rect 177538 159824 177594 159880
rect 177354 158736 177410 158792
rect 177538 157512 177594 157568
rect 177538 156288 177594 156344
rect 179654 159960 179710 160016
rect 179562 157648 179618 157704
rect 179470 155336 179526 155392
rect 177354 155064 177410 155120
rect 178182 153840 178238 153896
rect 179654 152888 179710 152944
rect 178274 152616 178330 152672
rect 177722 148944 177778 149000
rect 177170 147720 177226 147776
rect 134482 142008 134538 142064
rect 103478 141464 103534 141520
rect 102282 140920 102338 140976
rect 102374 140376 102430 140432
rect 102374 139696 102430 139752
rect 102466 139152 102522 139208
rect 102558 138608 102614 138664
rect 102374 137928 102430 137984
rect 65022 136704 65078 136760
rect 62906 136568 62962 136624
rect 62722 135616 62778 135672
rect 62630 135344 62686 135400
rect 62814 134800 62870 134856
rect 62906 134256 62962 134312
rect 100626 136568 100682 136624
rect 66402 136432 66458 136488
rect 65666 135908 65722 135944
rect 65666 135888 65668 135908
rect 65668 135888 65720 135908
rect 65720 135888 65722 135908
rect 100902 136024 100958 136080
rect 100902 135908 100958 135944
rect 100902 135888 100904 135908
rect 100904 135888 100956 135908
rect 100956 135888 100958 135908
rect 65850 135208 65906 135264
rect 99890 134800 99946 134856
rect 66218 134664 66274 134720
rect 100902 134664 100958 134720
rect 65482 134120 65538 134176
rect 62998 133576 63054 133632
rect 100902 133576 100958 133632
rect 66402 133440 66458 133496
rect 62814 132760 62870 132816
rect 62722 132488 62778 132544
rect 62814 130756 62816 130776
rect 62816 130756 62868 130776
rect 62868 130756 62870 130776
rect 62814 130720 62870 130756
rect 62722 128680 62778 128736
rect 100258 133188 100314 133224
rect 100258 133168 100260 133188
rect 100260 133168 100312 133188
rect 100312 133168 100314 133188
rect 63458 131536 63514 131592
rect 65022 132488 65078 132544
rect 63550 131264 63606 131320
rect 100258 132352 100314 132408
rect 66402 132216 66458 132272
rect 65666 131708 65668 131728
rect 65668 131708 65720 131728
rect 65720 131708 65722 131728
rect 65666 131672 65722 131708
rect 100902 131944 100958 132000
rect 100902 131708 100904 131728
rect 100904 131708 100956 131728
rect 100956 131708 100958 131728
rect 100902 131672 100958 131708
rect 66310 131128 66366 131184
rect 100258 130584 100314 130640
rect 66402 130448 66458 130504
rect 100902 130448 100958 130504
rect 102466 137384 102522 137440
rect 102374 136840 102430 136896
rect 102650 136296 102706 136352
rect 102282 135616 102338 135672
rect 102190 135072 102246 135128
rect 102006 133304 102062 133360
rect 102098 132216 102154 132272
rect 102006 131536 102062 131592
rect 101914 131400 101970 131456
rect 63642 130176 63698 130232
rect 65482 129904 65538 129960
rect 63090 129496 63146 129552
rect 100258 129360 100314 129416
rect 66402 129224 66458 129280
rect 100902 128972 100958 129008
rect 100902 128952 100904 128972
rect 100904 128952 100956 128972
rect 100956 128952 100958 128972
rect 62906 128408 62962 128464
rect 100074 128272 100130 128328
rect 66402 128136 66458 128192
rect 65022 127864 65078 127920
rect 62814 127456 62870 127512
rect 62630 127184 62686 127240
rect 62814 126640 62870 126696
rect 102374 134528 102430 134584
rect 102374 133848 102430 133904
rect 102282 132760 102338 132816
rect 102190 130992 102246 131048
rect 102282 130720 102338 130776
rect 102098 129224 102154 129280
rect 102006 128136 102062 128192
rect 100810 127612 100866 127648
rect 100810 127592 100812 127612
rect 100812 127592 100864 127612
rect 100864 127592 100866 127612
rect 100534 127048 100590 127104
rect 66310 126912 66366 126968
rect 65022 126504 65078 126560
rect 62906 125960 62962 126016
rect 66402 126232 66458 126288
rect 100626 126368 100682 126424
rect 100902 126232 100958 126288
rect 66402 125688 66458 125744
rect 62814 125416 62870 125472
rect 65850 125144 65906 125200
rect 65022 124872 65078 124928
rect 62722 124600 62778 124656
rect 62630 124328 62686 124384
rect 62814 123648 62870 123704
rect 100626 125280 100682 125336
rect 66402 124872 66458 124928
rect 100626 124892 100682 124928
rect 100626 124872 100628 124892
rect 100628 124872 100680 124892
rect 100680 124872 100682 124892
rect 102098 127456 102154 127512
rect 102374 129768 102430 129824
rect 102282 128680 102338 128736
rect 102190 126912 102246 126968
rect 135126 138880 135182 138936
rect 134574 138336 134630 138392
rect 135310 140920 135366 140976
rect 135310 140376 135366 140432
rect 135310 139696 135366 139752
rect 163278 142552 163334 142608
rect 162174 141872 162230 141928
rect 135310 139152 135366 139208
rect 136966 139016 137022 139072
rect 136874 138880 136930 138936
rect 135218 137656 135274 137712
rect 174594 142144 174650 142200
rect 177446 145408 177502 145464
rect 178366 151392 178422 151448
rect 178458 150168 178514 150224
rect 178182 146496 178238 146552
rect 200538 151548 200594 151584
rect 200538 151528 200540 151548
rect 200540 151528 200592 151548
rect 200592 151528 200594 151548
rect 180482 150576 180538 150632
rect 180390 148264 180446 148320
rect 180298 145952 180354 146008
rect 224458 163496 224514 163552
rect 207438 163224 207494 163280
rect 223538 159144 223594 159200
rect 207438 153704 207494 153760
rect 207438 152208 207494 152264
rect 204494 151528 204550 151584
rect 207438 142688 207494 142744
rect 207898 142552 207954 142608
rect 174410 140920 174466 140976
rect 174226 140376 174282 140432
rect 174134 139152 174190 139208
rect 172570 139016 172626 139072
rect 172202 138608 172258 138664
rect 136874 137792 136930 137848
rect 136874 137268 136930 137304
rect 136874 137248 136876 137268
rect 136876 137248 136928 137268
rect 136928 137248 136930 137268
rect 174318 139696 174374 139752
rect 174226 138608 174282 138664
rect 174134 137928 174190 137984
rect 172662 137792 172718 137848
rect 172662 137268 172718 137304
rect 172662 137248 172664 137268
rect 172664 137248 172716 137268
rect 172716 137248 172718 137268
rect 135402 136840 135458 136896
rect 135310 136568 135366 136624
rect 136782 136568 136838 136624
rect 172570 136568 172626 136624
rect 135218 135616 135274 135672
rect 135126 135344 135182 135400
rect 135218 134800 135274 134856
rect 134298 133576 134354 133632
rect 136874 136024 136930 136080
rect 136966 135908 137022 135944
rect 136966 135888 136968 135908
rect 136968 135888 137020 135908
rect 137020 135888 137022 135908
rect 172662 136044 172718 136080
rect 172662 136024 172664 136044
rect 172664 136024 172716 136044
rect 172716 136024 172718 136044
rect 172662 135908 172718 135944
rect 172662 135888 172664 135908
rect 172664 135888 172716 135908
rect 172716 135888 172718 135908
rect 174226 137384 174282 137440
rect 136874 134800 136930 134856
rect 172662 134800 172718 134856
rect 136966 134664 137022 134720
rect 172570 134528 172626 134584
rect 135310 134256 135366 134312
rect 135126 132488 135182 132544
rect 134298 130756 134300 130776
rect 134300 130756 134352 130776
rect 134352 130756 134354 130776
rect 134298 130720 134354 130756
rect 135218 131536 135274 131592
rect 136966 133576 137022 133632
rect 171650 133576 171706 133632
rect 173766 133304 173822 133360
rect 136874 133052 136930 133088
rect 136874 133032 136876 133052
rect 136876 133032 136928 133052
rect 136928 133032 136930 133052
rect 172662 133032 172718 133088
rect 135402 132760 135458 132816
rect 136782 132352 136838 132408
rect 172018 132352 172074 132408
rect 135310 131264 135366 131320
rect 135034 129496 135090 129552
rect 102282 126368 102338 126424
rect 102006 125688 102062 125744
rect 100626 124056 100682 124112
rect 66402 123920 66458 123976
rect 65022 123512 65078 123568
rect 62906 123104 62962 123160
rect 62814 122596 62816 122616
rect 62816 122596 62868 122616
rect 62868 122596 62870 122616
rect 62814 122560 62870 122596
rect 62814 121336 62870 121392
rect 99890 123396 99946 123432
rect 99890 123376 99892 123396
rect 99892 123376 99944 123396
rect 99944 123376 99946 123396
rect 102374 125144 102430 125200
rect 102282 124600 102338 124656
rect 102374 123920 102430 123976
rect 102098 123376 102154 123432
rect 100166 122832 100222 122888
rect 102006 122832 102062 122888
rect 66310 122696 66366 122752
rect 65022 122424 65078 122480
rect 63550 121608 63606 121664
rect 63458 120520 63514 120576
rect 100994 122288 101050 122344
rect 66402 122152 66458 122208
rect 100902 122152 100958 122208
rect 100626 121064 100682 121120
rect 66218 120928 66274 120984
rect 65022 120656 65078 120712
rect 63642 120248 63698 120304
rect 62814 119568 62870 119624
rect 65022 119432 65078 119488
rect 62722 118752 62778 118808
rect 62814 118480 62870 118536
rect 100626 120676 100682 120712
rect 100626 120656 100628 120676
rect 100628 120656 100680 120676
rect 100680 120656 100682 120676
rect 102282 122288 102338 122344
rect 102190 121608 102246 121664
rect 102282 121064 102338 121120
rect 100626 119840 100682 119896
rect 102098 119840 102154 119896
rect 66402 119704 66458 119760
rect 100902 119296 100958 119352
rect 66402 119160 66458 119216
rect 64930 118480 64986 118536
rect 62906 117800 62962 117856
rect 62814 117292 62816 117312
rect 62816 117292 62868 117312
rect 62868 117292 62870 117312
rect 62814 117256 62870 117292
rect 100626 118616 100682 118672
rect 65022 118208 65078 118264
rect 66402 118208 66458 118264
rect 100626 118072 100682 118128
rect 66402 117936 66458 117992
rect 100718 117936 100774 117992
rect 100534 116848 100590 116904
rect 62814 116712 62870 116768
rect 66402 116712 66458 116768
rect 65022 116440 65078 116496
rect 62722 116168 62778 116224
rect 62814 115488 62870 115544
rect 65022 115080 65078 115136
rect 62814 114672 62870 114728
rect 100626 116712 100682 116768
rect 102374 120556 102376 120576
rect 102376 120556 102428 120576
rect 102428 120556 102430 120576
rect 102374 120520 102430 120556
rect 102282 119568 102338 119624
rect 102190 118752 102246 118808
rect 135126 128408 135182 128464
rect 134298 127184 134354 127240
rect 134666 126640 134722 126696
rect 136874 131944 136930 132000
rect 171650 131944 171706 132000
rect 136966 131708 136968 131728
rect 136968 131708 137020 131728
rect 137020 131708 137022 131728
rect 136966 131672 137022 131708
rect 172662 131808 172718 131864
rect 136874 130584 136930 130640
rect 172386 130604 172442 130640
rect 172386 130584 172388 130604
rect 172388 130584 172440 130604
rect 172440 130584 172442 130604
rect 136966 130448 137022 130504
rect 172662 130312 172718 130368
rect 135402 130176 135458 130232
rect 136874 129360 136930 129416
rect 172662 129360 172718 129416
rect 136966 128988 136968 129008
rect 136968 128988 137020 129008
rect 137020 128988 137022 129008
rect 136966 128952 137022 128988
rect 172662 128972 172718 129008
rect 172662 128952 172664 128972
rect 172664 128952 172716 128972
rect 172716 128952 172718 128972
rect 174134 136840 174190 136896
rect 204770 136568 204826 136624
rect 174226 136296 174282 136352
rect 174134 135652 174136 135672
rect 174136 135652 174188 135672
rect 174188 135652 174190 135672
rect 174134 135616 174190 135652
rect 174042 135072 174098 135128
rect 174226 134528 174282 134584
rect 173950 133848 174006 133904
rect 174042 132760 174098 132816
rect 173858 132216 173914 132272
rect 174134 131572 174136 131592
rect 174136 131572 174188 131592
rect 174188 131572 174190 131592
rect 174134 131536 174190 131572
rect 135310 128680 135366 128736
rect 136782 128272 136838 128328
rect 171650 128272 171706 128328
rect 135218 127456 135274 127512
rect 136874 127612 136930 127648
rect 136874 127592 136876 127612
rect 136876 127592 136928 127612
rect 136928 127592 136930 127612
rect 172662 127592 172718 127648
rect 136782 127048 136838 127104
rect 172018 127048 172074 127104
rect 135126 125960 135182 126016
rect 134850 125416 134906 125472
rect 135310 124600 135366 124656
rect 136874 126368 136930 126424
rect 136966 126252 137022 126288
rect 136966 126232 136968 126252
rect 136968 126232 137020 126252
rect 137020 126232 137022 126252
rect 172386 126388 172442 126424
rect 172386 126368 172388 126388
rect 172388 126368 172440 126388
rect 172440 126368 172442 126388
rect 172662 126096 172718 126152
rect 175054 130992 175110 131048
rect 174134 130448 174190 130504
rect 174134 129768 174190 129824
rect 174502 129224 174558 129280
rect 174042 128680 174098 128736
rect 174134 128136 174190 128192
rect 173950 127456 174006 127512
rect 173858 126912 173914 126968
rect 174226 126368 174282 126424
rect 136782 125280 136838 125336
rect 172018 125280 172074 125336
rect 136874 124872 136930 124928
rect 172662 124892 172718 124928
rect 172662 124872 172664 124892
rect 172664 124872 172716 124892
rect 172716 124872 172718 124892
rect 135402 124328 135458 124384
rect 136782 124056 136838 124112
rect 172386 124056 172442 124112
rect 135218 123648 135274 123704
rect 135126 123104 135182 123160
rect 135310 122560 135366 122616
rect 136874 123396 136930 123432
rect 173858 123920 173914 123976
rect 136874 123376 136876 123396
rect 136876 123376 136928 123396
rect 136928 123376 136930 123396
rect 172662 123376 172718 123432
rect 136874 122832 136930 122888
rect 171558 122832 171614 122888
rect 136966 122424 137022 122480
rect 137058 122172 137114 122208
rect 137058 122152 137060 122172
rect 137060 122152 137112 122172
rect 137112 122152 137114 122172
rect 172662 122016 172718 122072
rect 135402 121880 135458 121936
rect 135310 121336 135366 121392
rect 136782 121064 136838 121120
rect 171742 121064 171798 121120
rect 135218 120520 135274 120576
rect 135126 120248 135182 120304
rect 136874 120656 136930 120712
rect 172662 120676 172718 120712
rect 172662 120656 172664 120676
rect 172664 120656 172716 120676
rect 172716 120656 172718 120676
rect 136782 119840 136838 119896
rect 134850 119568 134906 119624
rect 135034 118480 135090 118536
rect 102282 118208 102338 118264
rect 102190 116984 102246 117040
rect 62814 114400 62870 114456
rect 56926 113176 56982 113232
rect 31994 104200 32050 104256
rect 37422 104200 37478 104256
rect 32638 90872 32694 90928
rect 36410 90872 36466 90928
rect 72842 113584 72898 113640
rect 73210 113176 73266 113232
rect 100626 115488 100682 115544
rect 102374 117528 102430 117584
rect 102282 116440 102338 116496
rect 102466 115760 102522 115816
rect 102374 115216 102430 115272
rect 102190 114672 102246 114728
rect 135310 119060 135312 119080
rect 135312 119060 135364 119080
rect 135364 119060 135366 119080
rect 135310 119024 135366 119060
rect 174226 125688 174282 125744
rect 174134 125144 174190 125200
rect 174042 124600 174098 124656
rect 174226 123376 174282 123432
rect 173950 122832 174006 122888
rect 172938 122288 172994 122344
rect 174042 122288 174098 122344
rect 174318 121608 174374 121664
rect 174134 121064 174190 121120
rect 172662 119840 172718 119896
rect 136966 119316 137022 119352
rect 136966 119296 136968 119316
rect 136968 119296 137020 119316
rect 137020 119296 137022 119316
rect 172662 119296 172718 119352
rect 136966 118616 137022 118672
rect 172018 118616 172074 118672
rect 136782 118072 136838 118128
rect 135218 117528 135274 117584
rect 134114 117256 134170 117312
rect 134666 116712 134722 116768
rect 136874 117956 136930 117992
rect 136874 117936 136876 117956
rect 136876 117936 136928 117956
rect 136928 117936 136930 117956
rect 172662 118092 172718 118128
rect 172662 118072 172664 118092
rect 172664 118072 172716 118092
rect 172716 118072 172718 118092
rect 172478 117936 172534 117992
rect 136782 116848 136838 116904
rect 135310 116168 135366 116224
rect 136874 116440 136930 116496
rect 134482 115488 134538 115544
rect 136782 115488 136838 115544
rect 135310 114980 135312 115000
rect 135312 114980 135364 115000
rect 135364 114980 135366 115000
rect 135310 114944 135366 114980
rect 174134 120556 174136 120576
rect 174136 120556 174188 120576
rect 174188 120556 174190 120576
rect 174134 120520 174190 120556
rect 173950 118752 174006 118808
rect 174318 119840 174374 119896
rect 174134 119296 174190 119352
rect 174042 118208 174098 118264
rect 172662 116848 172718 116904
rect 172570 116440 172626 116496
rect 134850 114436 134852 114456
rect 134852 114436 134904 114456
rect 134904 114436 134906 114456
rect 134850 114400 134906 114436
rect 102282 114128 102338 114184
rect 92806 112632 92862 112688
rect 60514 104200 60570 104256
rect 105502 106512 105558 106568
rect 105226 105288 105282 105344
rect 105962 110184 106018 110240
rect 105778 108960 105834 109016
rect 105686 107736 105742 107792
rect 108630 109504 108686 109560
rect 108538 107192 108594 107248
rect 107894 104880 107950 104936
rect 106146 104064 106202 104120
rect 105594 102840 105650 102896
rect 105134 101616 105190 101672
rect 57570 100800 57626 100856
rect 105594 99168 105650 99224
rect 107894 102432 107950 102488
rect 105962 100392 106018 100448
rect 105686 98080 105742 98136
rect 107894 100120 107950 100176
rect 106330 96856 106386 96912
rect 107894 97808 107950 97864
rect 106422 95632 106478 95688
rect 107802 95360 107858 95416
rect 105778 94408 105834 94464
rect 105778 93184 105834 93240
rect 107802 93048 107858 93104
rect 105226 91960 105282 92016
rect 59594 90872 59650 90928
rect 105778 89260 105834 89296
rect 105778 89240 105780 89260
rect 105780 89240 105832 89260
rect 105832 89240 105834 89260
rect 107802 88424 107858 88480
rect 105410 87900 105466 87936
rect 105410 87880 105412 87900
rect 105412 87880 105464 87900
rect 105464 87880 105466 87900
rect 106422 86520 106478 86576
rect 107894 85976 107950 86032
rect 105134 85296 105190 85352
rect 105686 84772 105742 84808
rect 105686 84752 105688 84772
rect 105688 84752 105740 84772
rect 105740 84752 105742 84772
rect 105226 83412 105282 83448
rect 105226 83392 105228 83412
rect 105228 83392 105280 83412
rect 105280 83392 105282 83412
rect 106422 82188 106478 82224
rect 106422 82168 106424 82188
rect 106424 82168 106476 82188
rect 106476 82168 106478 82188
rect 56926 81896 56982 81952
rect 57478 81896 57534 81952
rect 57478 80808 57534 80864
rect 105962 80828 106018 80864
rect 105962 80808 105964 80828
rect 105964 80808 106016 80828
rect 106016 80808 106018 80828
rect 105410 79584 105466 79640
rect 107618 78904 107674 78960
rect 105226 77952 105282 78008
rect 31994 77544 32050 77600
rect 37422 77544 37478 77600
rect 59594 77580 59596 77600
rect 59596 77580 59648 77600
rect 59648 77580 59650 77600
rect 31902 69420 31904 69440
rect 31904 69420 31956 69440
rect 31956 69420 31958 69440
rect 31902 69384 31958 69420
rect 59594 77544 59650 77580
rect 106974 76728 107030 76784
rect 105962 75504 106018 75560
rect 105410 74280 105466 74336
rect 105226 73736 105282 73792
rect 62814 66700 62816 66720
rect 62816 66700 62868 66720
rect 62868 66700 62870 66720
rect 62814 66664 62870 66700
rect 62722 66120 62778 66176
rect 62906 65576 62962 65632
rect 62814 64896 62870 64952
rect 62722 64352 62778 64408
rect 63366 67208 63422 67264
rect 62998 63808 63054 63864
rect 62354 63264 62410 63320
rect 12030 62856 12086 62912
rect 29234 62856 29290 62912
rect 66402 65440 66458 65496
rect 66402 64896 66458 64952
rect 63366 62720 63422 62776
rect 11938 41232 11994 41288
rect 65666 64236 65722 64272
rect 65666 64216 65668 64236
rect 65668 64216 65720 64236
rect 65720 64216 65722 64236
rect 101362 71152 101418 71208
rect 101914 71016 101970 71072
rect 102374 66392 102430 66448
rect 102466 65848 102522 65904
rect 100902 65460 100958 65496
rect 100902 65440 100904 65460
rect 100904 65440 100956 65460
rect 100956 65440 100958 65460
rect 100626 64508 100682 64544
rect 100626 64488 100628 64508
rect 100628 64488 100680 64508
rect 100680 64488 100682 64508
rect 100902 64100 100958 64136
rect 100902 64080 100904 64100
rect 100904 64080 100956 64100
rect 100956 64080 100958 64100
rect 66402 63672 66458 63728
rect 65666 63128 65722 63184
rect 100626 63264 100682 63320
rect 105870 72512 105926 72568
rect 106514 71016 106570 71072
rect 107986 83664 108042 83720
rect 107802 81352 107858 81408
rect 107710 76592 107766 76648
rect 107894 74280 107950 74336
rect 108538 71968 108594 72024
rect 117830 69112 117886 69168
rect 119394 69112 119450 69168
rect 119118 68976 119174 69032
rect 121142 68976 121198 69032
rect 144878 113584 144934 113640
rect 172662 115644 172718 115680
rect 172662 115624 172664 115644
rect 172664 115624 172716 115644
rect 172716 115624 172718 115644
rect 204770 117936 204826 117992
rect 174134 117528 174190 117584
rect 174042 116984 174098 117040
rect 173950 116440 174006 116496
rect 174134 115760 174190 115816
rect 173858 114672 173914 114728
rect 174226 115216 174282 115272
rect 174042 114128 174098 114184
rect 164842 113584 164898 113640
rect 176986 107736 177042 107792
rect 176894 106512 176950 106568
rect 177078 105288 177134 105344
rect 177354 108996 177356 109016
rect 177356 108996 177408 109016
rect 177408 108996 177410 109016
rect 177354 108960 177410 108996
rect 177262 104064 177318 104120
rect 177722 110184 177778 110240
rect 180298 109504 180354 109560
rect 179654 104880 179710 104936
rect 177538 102840 177594 102896
rect 176894 101616 176950 101672
rect 176986 100392 177042 100448
rect 177354 99168 177410 99224
rect 132366 95768 132422 95824
rect 132550 95768 132606 95824
rect 177630 96856 177686 96912
rect 179654 102432 179710 102488
rect 180390 107192 180446 107248
rect 179654 100120 179710 100176
rect 223538 149488 223594 149544
rect 207990 127728 208046 127784
rect 207898 118480 207954 118536
rect 201090 104200 201146 104256
rect 204678 104200 204734 104256
rect 178182 98080 178238 98136
rect 179654 97808 179710 97864
rect 177722 95632 177778 95688
rect 179562 95360 179618 95416
rect 177538 94408 177594 94464
rect 177354 93184 177410 93240
rect 179562 93048 179618 93104
rect 176986 91996 176988 92016
rect 176988 91996 177040 92016
rect 177040 91996 177042 92016
rect 176986 91960 177042 91996
rect 200998 90872 201054 90928
rect 204494 90872 204550 90928
rect 177354 88288 177410 88344
rect 177538 87064 177594 87120
rect 179654 85976 179710 86032
rect 176986 85840 177042 85896
rect 178182 84772 178238 84808
rect 178182 84752 178184 84772
rect 178184 84752 178236 84772
rect 178236 84752 178238 84772
rect 178090 83528 178146 83584
rect 177722 82324 177778 82360
rect 177722 82304 177724 82324
rect 177724 82304 177776 82324
rect 177776 82304 177778 82324
rect 178090 81080 178146 81136
rect 177630 79856 177686 79912
rect 176986 78632 177042 78688
rect 178826 77408 178882 77464
rect 178274 76184 178330 76240
rect 177722 74960 177778 75016
rect 177170 73736 177226 73792
rect 103478 67480 103534 67536
rect 102926 66936 102982 66992
rect 102742 65168 102798 65224
rect 102650 64624 102706 64680
rect 102558 64080 102614 64136
rect 102374 62992 102430 63048
rect 100626 62740 100682 62776
rect 100626 62720 100628 62740
rect 100628 62720 100680 62740
rect 100680 62720 100682 62740
rect 66402 62448 66458 62504
rect 63550 62040 63606 62096
rect 65666 61904 65722 61960
rect 63458 61496 63514 61552
rect 62814 60952 62870 61008
rect 62722 60408 62778 60464
rect 100626 62040 100682 62096
rect 100534 61360 100590 61416
rect 65482 61224 65538 61280
rect 102558 63536 102614 63592
rect 102466 61768 102522 61824
rect 102374 61224 102430 61280
rect 100626 60816 100682 60872
rect 66310 60680 66366 60736
rect 63734 59864 63790 59920
rect 62906 59184 62962 59240
rect 100626 60292 100682 60328
rect 100626 60272 100628 60292
rect 100628 60272 100680 60292
rect 100680 60272 100682 60292
rect 66402 60156 66458 60192
rect 66402 60136 66404 60156
rect 66404 60136 66456 60156
rect 66456 60136 66458 60156
rect 100626 60020 100682 60056
rect 100626 60000 100628 60020
rect 100628 60000 100680 60020
rect 100680 60000 100682 60020
rect 66310 59456 66366 59512
rect 63826 58640 63882 58696
rect 100626 59048 100682 59104
rect 66402 58912 66458 58968
rect 62722 58096 62778 58152
rect 62630 57552 62686 57608
rect 62538 55784 62594 55840
rect 100626 58660 100682 58696
rect 100626 58640 100628 58660
rect 100628 58640 100680 58660
rect 100680 58640 100682 58660
rect 62814 57008 62870 57064
rect 135310 67480 135366 67536
rect 135034 66936 135090 66992
rect 135310 66428 135312 66448
rect 135312 66428 135364 66448
rect 135364 66428 135366 66448
rect 135310 66392 135366 66428
rect 134666 65848 134722 65904
rect 134482 64080 134538 64136
rect 135310 65204 135312 65224
rect 135312 65204 135364 65224
rect 135364 65204 135366 65224
rect 135310 65168 135366 65204
rect 134850 64624 134906 64680
rect 134666 62992 134722 63048
rect 102742 62312 102798 62368
rect 102558 60680 102614 60736
rect 102466 60136 102522 60192
rect 102374 58368 102430 58424
rect 65022 58232 65078 58288
rect 100626 57824 100682 57880
rect 66402 57688 66458 57744
rect 100626 57280 100682 57336
rect 66402 57164 66458 57200
rect 66402 57144 66404 57164
rect 66404 57144 66456 57164
rect 66456 57144 66458 57164
rect 100534 57164 100590 57200
rect 100534 57144 100536 57164
rect 100536 57144 100588 57164
rect 100588 57144 100590 57164
rect 66402 56464 66458 56520
rect 62906 56328 62962 56384
rect 62722 55240 62778 55296
rect 62630 54696 62686 54752
rect 30522 53472 30578 53528
rect 63274 53472 63330 53528
rect 134850 62312 134906 62368
rect 135402 63536 135458 63592
rect 136874 65460 136930 65496
rect 136874 65440 136876 65460
rect 136876 65440 136928 65460
rect 136928 65440 136930 65460
rect 136874 64488 136930 64544
rect 136966 64116 136968 64136
rect 136968 64116 137020 64136
rect 137020 64116 137022 64136
rect 136966 64080 137022 64116
rect 174042 66936 174098 66992
rect 173950 66392 174006 66448
rect 173858 65848 173914 65904
rect 172662 65596 172718 65632
rect 172662 65576 172664 65596
rect 172664 65576 172716 65596
rect 172716 65576 172718 65596
rect 174134 65168 174190 65224
rect 174226 64624 174282 64680
rect 172662 64488 172718 64544
rect 171834 64100 171890 64136
rect 171834 64080 171836 64100
rect 171836 64080 171888 64100
rect 171888 64080 171890 64100
rect 174134 63536 174190 63592
rect 136874 63264 136930 63320
rect 172662 63264 172718 63320
rect 172662 62856 172718 62912
rect 136966 62740 137022 62776
rect 136966 62720 136968 62740
rect 136968 62720 137020 62740
rect 137020 62720 137022 62740
rect 135310 61768 135366 61824
rect 136782 62040 136838 62096
rect 172662 62040 172718 62096
rect 134482 60680 134538 60736
rect 135034 60136 135090 60192
rect 102742 59456 102798 59512
rect 102650 58912 102706 58968
rect 102558 57824 102614 57880
rect 102466 57280 102522 57336
rect 100626 56056 100682 56112
rect 102374 56056 102430 56112
rect 66402 55940 66458 55976
rect 66402 55920 66404 55940
rect 66404 55920 66456 55940
rect 66456 55920 66458 55940
rect 100902 55804 100958 55840
rect 100902 55784 100904 55804
rect 100904 55784 100956 55804
rect 100956 55784 100958 55804
rect 66310 55240 66366 55296
rect 100626 54852 100682 54888
rect 100626 54832 100628 54852
rect 100628 54832 100680 54852
rect 100680 54832 100682 54852
rect 66402 54716 66458 54752
rect 66402 54696 66404 54716
rect 66404 54696 66456 54716
rect 66456 54696 66458 54716
rect 100810 54580 100866 54616
rect 100810 54560 100812 54580
rect 100812 54560 100864 54580
rect 100864 54560 100866 54580
rect 102466 55512 102522 55568
rect 135402 61224 135458 61280
rect 171834 61632 171890 61688
rect 136874 61360 136930 61416
rect 177630 72512 177686 72568
rect 177354 71424 177410 71480
rect 179562 81352 179618 81408
rect 179746 83664 179802 83720
rect 179654 78904 179710 78960
rect 179470 76592 179526 76648
rect 179746 74280 179802 74336
rect 180298 71968 180354 72024
rect 189314 69112 189370 69168
rect 190234 69112 190290 69168
rect 191338 69112 191394 69168
rect 193086 69112 193142 69168
rect 201090 77544 201146 77600
rect 204494 77544 204550 77600
rect 201090 69284 201092 69304
rect 201092 69284 201144 69304
rect 201144 69284 201146 69304
rect 201090 69248 201146 69284
rect 175054 67480 175110 67536
rect 174410 64080 174466 64136
rect 174226 62312 174282 62368
rect 174134 61224 174190 61280
rect 136782 60816 136838 60872
rect 172202 60816 172258 60872
rect 135310 59456 135366 59512
rect 135034 58912 135090 58968
rect 134482 58368 134538 58424
rect 135034 57280 135090 57336
rect 102650 56600 102706 56656
rect 102558 54968 102614 55024
rect 102374 54424 102430 54480
rect 63642 54152 63698 54208
rect 66402 54152 66458 54208
rect 65298 53472 65354 53528
rect 100626 53608 100682 53664
rect 102466 53200 102522 53256
rect 100626 53084 100682 53120
rect 100626 53064 100628 53084
rect 100628 53064 100680 53084
rect 100680 53064 100682 53084
rect 63550 52928 63606 52984
rect 63366 52384 63422 52440
rect 62814 51296 62870 51352
rect 62722 49528 62778 49584
rect 66310 52928 66366 52984
rect 65298 52248 65354 52304
rect 63734 51840 63790 51896
rect 65666 51724 65722 51760
rect 65666 51704 65668 51724
rect 65668 51704 65720 51724
rect 65720 51704 65722 51724
rect 100626 52384 100682 52440
rect 100626 51840 100682 51896
rect 100534 51704 100590 51760
rect 136966 60272 137022 60328
rect 172662 60292 172718 60328
rect 172662 60272 172664 60292
rect 172664 60272 172716 60292
rect 172716 60272 172718 60292
rect 175330 62992 175386 63048
rect 175238 61768 175294 61824
rect 174318 60680 174374 60736
rect 174226 60136 174282 60192
rect 136874 60000 136930 60056
rect 172662 60020 172718 60056
rect 172662 60000 172664 60020
rect 172664 60000 172716 60020
rect 172716 60000 172718 60020
rect 136782 59048 136838 59104
rect 172202 59048 172258 59104
rect 174134 58912 174190 58968
rect 171834 58796 171890 58832
rect 171834 58776 171836 58796
rect 171836 58776 171888 58796
rect 171888 58776 171890 58796
rect 136874 58640 136930 58696
rect 135402 57824 135458 57880
rect 136782 57824 136838 57880
rect 172018 57824 172074 57880
rect 135310 56600 135366 56656
rect 135034 56056 135090 56112
rect 134758 55512 134814 55568
rect 102650 53744 102706 53800
rect 134206 53744 134262 53800
rect 102558 52656 102614 52712
rect 102374 51568 102430 51624
rect 66402 51160 66458 51216
rect 63734 50616 63790 50672
rect 100626 50616 100682 50672
rect 63366 50072 63422 50128
rect 65666 50500 65722 50536
rect 65666 50480 65668 50500
rect 65668 50480 65720 50500
rect 65720 50480 65722 50500
rect 100626 50364 100682 50400
rect 100626 50344 100628 50364
rect 100628 50344 100680 50364
rect 100680 50344 100682 50364
rect 102466 50344 102522 50400
rect 65482 49936 65538 49992
rect 63826 48984 63882 49040
rect 100626 49392 100682 49448
rect 66402 49256 66458 49312
rect 62814 48440 62870 48496
rect 62722 46128 62778 46184
rect 100626 49004 100682 49040
rect 100626 48984 100628 49004
rect 100628 48984 100680 49004
rect 100680 48984 100682 49004
rect 136874 57280 136930 57336
rect 136966 57180 136968 57200
rect 136968 57180 137020 57200
rect 137020 57180 137022 57200
rect 136966 57144 137022 57180
rect 172662 57436 172718 57472
rect 172662 57416 172664 57436
rect 172664 57416 172716 57436
rect 172716 57416 172718 57436
rect 172662 57300 172718 57336
rect 172662 57280 172664 57300
rect 172664 57280 172716 57300
rect 172716 57280 172718 57300
rect 174410 59456 174466 59512
rect 174318 58368 174374 58424
rect 174502 57824 174558 57880
rect 174226 56600 174282 56656
rect 136782 56056 136838 56112
rect 172662 56076 172718 56112
rect 172662 56056 172664 56076
rect 172664 56056 172716 56076
rect 172716 56056 172718 56076
rect 174134 56056 174190 56112
rect 136874 55804 136930 55840
rect 136874 55784 136876 55804
rect 136876 55784 136928 55804
rect 136928 55784 136930 55804
rect 172662 55804 172718 55840
rect 172662 55784 172664 55804
rect 172664 55784 172716 55804
rect 172716 55784 172718 55804
rect 135402 54968 135458 55024
rect 136782 54832 136838 54888
rect 172110 54832 172166 54888
rect 135034 54424 135090 54480
rect 137150 54580 137206 54616
rect 137150 54560 137152 54580
rect 137152 54560 137204 54580
rect 137204 54560 137206 54580
rect 172662 54560 172718 54616
rect 174594 57280 174650 57336
rect 174318 55512 174374 55568
rect 174410 54968 174466 55024
rect 174226 54424 174282 54480
rect 136782 53608 136838 53664
rect 171650 53608 171706 53664
rect 135126 53200 135182 53256
rect 134298 52656 134354 52712
rect 102742 52112 102798 52168
rect 135126 52112 135182 52168
rect 174962 53744 175018 53800
rect 172662 53200 172718 53256
rect 136874 53064 136930 53120
rect 174778 53200 174834 53256
rect 136690 52384 136746 52440
rect 172018 52384 172074 52440
rect 102650 50888 102706 50944
rect 102558 49800 102614 49856
rect 135034 50344 135090 50400
rect 135402 51568 135458 51624
rect 136782 51840 136838 51896
rect 136874 51704 136930 51760
rect 174134 52112 174190 52168
rect 172570 51996 172626 52032
rect 172570 51976 172572 51996
rect 172572 51976 172624 51996
rect 172624 51976 172626 51996
rect 172662 51860 172718 51896
rect 172662 51840 172664 51860
rect 172664 51840 172716 51860
rect 172716 51840 172718 51860
rect 135402 50888 135458 50944
rect 174226 50888 174282 50944
rect 172202 50752 172258 50808
rect 136782 50616 136838 50672
rect 135310 49800 135366 49856
rect 102650 49256 102706 49312
rect 134850 49256 134906 49312
rect 64930 48712 64986 48768
rect 102374 48712 102430 48768
rect 63734 47760 63790 47816
rect 100626 48304 100682 48360
rect 102466 48032 102522 48088
rect 65022 47760 65078 47816
rect 63366 47216 63422 47272
rect 100626 47644 100682 47680
rect 100626 47624 100628 47644
rect 100628 47624 100680 47644
rect 100680 47624 100682 47644
rect 65666 47508 65722 47544
rect 65666 47488 65668 47508
rect 65668 47488 65720 47508
rect 65720 47488 65722 47508
rect 100626 47508 100682 47544
rect 100626 47488 100628 47508
rect 100628 47488 100680 47508
rect 100680 47488 100682 47508
rect 66402 46944 66458 47000
rect 62906 46672 62962 46728
rect 102558 47488 102614 47544
rect 100626 46400 100682 46456
rect 102374 46400 102430 46456
rect 62814 45584 62870 45640
rect 65206 46264 65262 46320
rect 63734 44904 63790 44960
rect 62814 44360 62870 44416
rect 100902 46148 100958 46184
rect 100902 46128 100904 46148
rect 100904 46128 100956 46148
rect 100956 46128 100958 46148
rect 66310 45720 66366 45776
rect 100534 45312 100590 45368
rect 66402 45176 66458 45232
rect 99982 45040 100038 45096
rect 136874 50344 136930 50400
rect 172662 50344 172718 50400
rect 174318 50344 174374 50400
rect 136874 49392 136930 49448
rect 172662 49392 172718 49448
rect 174134 49256 174190 49312
rect 171834 49140 171890 49176
rect 171834 49120 171836 49140
rect 171836 49120 171888 49140
rect 171888 49120 171890 49140
rect 136782 48848 136838 48904
rect 135402 48712 135458 48768
rect 136690 48304 136746 48360
rect 172570 48304 172626 48360
rect 135310 48032 135366 48088
rect 134758 47488 134814 47544
rect 102650 46944 102706 47000
rect 135310 46944 135366 47000
rect 134850 46400 134906 46456
rect 102466 45856 102522 45912
rect 175330 52656 175386 52712
rect 174502 51568 174558 51624
rect 174410 49800 174466 49856
rect 174318 48712 174374 48768
rect 174226 48032 174282 48088
rect 172662 47896 172718 47952
rect 136782 47624 136838 47680
rect 172662 47644 172718 47680
rect 172662 47624 172664 47644
rect 172664 47624 172716 47644
rect 172716 47624 172718 47644
rect 136874 47508 136930 47544
rect 136874 47488 136876 47508
rect 136876 47488 136928 47508
rect 136928 47488 136930 47508
rect 172662 46556 172718 46592
rect 172662 46536 172664 46556
rect 172664 46536 172716 46556
rect 172716 46536 172718 46556
rect 174226 46944 174282 47000
rect 136782 46400 136838 46456
rect 174134 46400 174190 46456
rect 137518 46128 137574 46184
rect 172662 46148 172718 46184
rect 172662 46128 172664 46148
rect 172664 46128 172716 46148
rect 172716 46128 172718 46148
rect 135402 45856 135458 45912
rect 136690 45312 136746 45368
rect 102374 44632 102430 44688
rect 66218 44496 66274 44552
rect 63734 43816 63790 43872
rect 102558 45176 102614 45232
rect 134666 45176 134722 45232
rect 99890 44108 99946 44144
rect 99890 44088 99892 44108
rect 99892 44088 99944 44108
rect 99944 44088 99946 44108
rect 102466 44088 102522 44144
rect 66402 43952 66458 44008
rect 63642 43272 63698 43328
rect 100626 43408 100682 43464
rect 63734 42728 63790 42784
rect 66310 43272 66366 43328
rect 63826 42456 63882 42512
rect 63734 41504 63790 41560
rect 135034 44668 135036 44688
rect 135036 44668 135088 44688
rect 135088 44668 135090 44688
rect 135034 44632 135090 44668
rect 136782 44904 136838 44960
rect 171650 45312 171706 45368
rect 174410 47488 174466 47544
rect 174318 45856 174374 45912
rect 174226 45176 174282 45232
rect 171834 44904 171890 44960
rect 135402 44088 135458 44144
rect 136782 44088 136838 44144
rect 172662 44088 172718 44144
rect 102558 43544 102614 43600
rect 135034 43544 135090 43600
rect 102282 43000 102338 43056
rect 100626 42864 100682 42920
rect 66402 42728 66458 42784
rect 100626 42320 100682 42376
rect 102374 42320 102430 42376
rect 66402 42184 66458 42240
rect 63826 40960 63882 41016
rect 100626 42068 100682 42104
rect 100626 42048 100628 42068
rect 100628 42048 100680 42068
rect 100680 42048 100682 42068
rect 63182 40416 63238 40472
rect 66402 40416 66458 40472
rect 62814 39464 62870 39520
rect 66218 32664 66274 32720
rect 66310 24640 66366 24696
rect 13318 19608 13374 19664
rect 172570 43544 172626 43600
rect 175330 44632 175386 44688
rect 175422 44088 175478 44144
rect 136874 43408 136930 43464
rect 135402 43036 135404 43056
rect 135404 43036 135456 43056
rect 135456 43036 135458 43056
rect 135402 43000 135458 43036
rect 174778 43544 174834 43600
rect 174042 43000 174098 43056
rect 136690 42864 136746 42920
rect 172202 42864 172258 42920
rect 134942 42320 134998 42376
rect 102558 41776 102614 41832
rect 135310 41812 135312 41832
rect 135312 41812 135364 41832
rect 135364 41812 135366 41832
rect 135310 41776 135366 41812
rect 102466 41232 102522 41288
rect 136874 42320 136930 42376
rect 136782 42048 136838 42104
rect 172662 42320 172718 42376
rect 174134 42320 174190 42376
rect 172662 42068 172718 42104
rect 172662 42048 172664 42068
rect 172664 42048 172716 42068
rect 172716 42048 172718 42068
rect 135402 41232 135458 41288
rect 102374 40688 102430 40744
rect 134850 40688 134906 40744
rect 94002 40416 94058 40472
rect 102374 40144 102430 40200
rect 109642 40008 109698 40064
rect 134482 39600 134538 39656
rect 136874 33344 136930 33400
rect 138162 39736 138218 39792
rect 138070 25048 138126 25104
rect 174226 41776 174282 41832
rect 174318 41232 174374 41288
rect 174134 40688 174190 40744
rect 181402 40008 181458 40064
rect 166038 39736 166094 39792
rect 174134 39464 174190 39520
rect 222894 139696 222950 139752
rect 222710 115896 222766 115952
rect 224458 105696 224514 105752
rect 223538 96312 223594 96368
rect 223538 92096 223594 92152
rect 223538 85160 223594 85216
rect 223538 75232 223594 75288
rect 223078 68296 223134 68352
rect 222526 44496 222582 44552
rect 222710 20696 222766 20752
rect 138162 17024 138218 17080
rect 66402 16752 66458 16808
<< metal3 >>
rect 98229 238762 98295 238765
rect 169989 238762 170055 238765
rect 96652 238760 98295 238762
rect 96652 238704 98234 238760
rect 98290 238704 98295 238760
rect 96652 238702 98295 238704
rect 168780 238760 170055 238762
rect 168780 238704 169994 238760
rect 170050 238704 170055 238760
rect 168780 238702 170055 238704
rect 98229 238699 98295 238702
rect 169989 238699 170055 238702
rect 9896 235906 10376 235936
rect 12025 235906 12091 235909
rect 9896 235904 12091 235906
rect 9896 235848 12030 235904
rect 12086 235848 12091 235904
rect 9896 235846 12091 235848
rect 9896 235816 10376 235846
rect 12025 235843 12091 235846
rect 223073 234954 223139 234957
rect 227416 234954 227896 234984
rect 223073 234952 227896 234954
rect 223073 234896 223078 234952
rect 223134 234896 227896 234952
rect 223073 234894 227896 234896
rect 223073 234891 223139 234894
rect 227416 234864 227896 234894
rect 98321 230738 98387 230741
rect 96652 230736 98387 230738
rect 96652 230680 98326 230736
rect 98382 230680 98387 230736
rect 96652 230678 98387 230680
rect 98321 230675 98387 230678
rect 168566 230197 168626 230708
rect 168517 230192 168626 230197
rect 168517 230136 168522 230192
rect 168578 230136 168626 230192
rect 168517 230134 168626 230136
rect 168517 230131 168583 230134
rect 98413 222850 98479 222853
rect 170081 222850 170147 222853
rect 96652 222848 98479 222850
rect 96652 222792 98418 222848
rect 98474 222792 98479 222848
rect 96652 222790 98479 222792
rect 168780 222848 170147 222850
rect 168780 222792 170086 222848
rect 170142 222792 170147 222848
rect 168780 222790 170147 222792
rect 98413 222787 98479 222790
rect 170081 222787 170147 222790
rect 37918 217212 37924 217276
rect 37988 217274 37994 217276
rect 55817 217274 55883 217277
rect 37988 217272 55883 217274
rect 37988 217216 55822 217272
rect 55878 217216 55883 217272
rect 37988 217214 55883 217216
rect 37988 217212 37994 217214
rect 55817 217211 55883 217214
rect 151037 215914 151103 215917
rect 204254 215914 204260 215916
rect 151037 215912 204260 215914
rect 151037 215856 151042 215912
rect 151098 215856 204260 215912
rect 151037 215854 204260 215856
rect 151037 215851 151103 215854
rect 204254 215852 204260 215854
rect 204324 215852 204330 215916
rect 174221 215778 174287 215781
rect 174221 215776 177090 215778
rect 174221 215720 174226 215776
rect 174282 215720 177090 215776
rect 174221 215718 177090 215720
rect 174221 215715 174287 215718
rect 135397 215642 135463 215645
rect 132686 215640 135463 215642
rect 132686 215584 135402 215640
rect 135458 215584 135463 215640
rect 132686 215582 135463 215584
rect 132686 215408 132746 215582
rect 135397 215579 135463 215582
rect 177030 215408 177090 215718
rect 62533 215370 62599 215373
rect 60588 215368 62599 215370
rect 60588 215312 62538 215368
rect 62594 215312 62599 215368
rect 60588 215310 62599 215312
rect 62533 215307 62599 215310
rect 102369 215370 102435 215373
rect 102369 215368 104932 215370
rect 102369 215312 102374 215368
rect 102430 215312 104932 215368
rect 102369 215310 104932 215312
rect 102369 215307 102435 215310
rect 62625 214690 62691 214693
rect 60588 214688 62691 214690
rect 60588 214632 62630 214688
rect 62686 214632 62691 214688
rect 60588 214630 62691 214632
rect 62625 214627 62691 214630
rect 102553 214690 102619 214693
rect 135397 214690 135463 214693
rect 102553 214688 104932 214690
rect 102553 214632 102558 214688
rect 102614 214632 104932 214688
rect 102553 214630 104932 214632
rect 132716 214688 135463 214690
rect 132716 214632 135402 214688
rect 135458 214632 135463 214688
rect 132716 214630 135463 214632
rect 102553 214627 102619 214630
rect 135397 214627 135463 214630
rect 174037 214690 174103 214693
rect 174037 214688 177060 214690
rect 174037 214632 174042 214688
rect 174098 214632 177060 214688
rect 174037 214630 177060 214632
rect 174037 214627 174103 214630
rect 9896 214282 10376 214312
rect 11933 214282 11999 214285
rect 9896 214280 11999 214282
rect 9896 214224 11938 214280
rect 11994 214224 11999 214280
rect 9896 214222 11999 214224
rect 9896 214192 10376 214222
rect 11933 214219 11999 214222
rect 63637 214010 63703 214013
rect 60588 214008 63703 214010
rect 60588 213952 63642 214008
rect 63698 213952 63703 214008
rect 60588 213950 63703 213952
rect 63637 213947 63703 213950
rect 103105 214010 103171 214013
rect 135397 214010 135463 214013
rect 103105 214008 104932 214010
rect 103105 213952 103110 214008
rect 103166 213952 104932 214008
rect 103105 213950 104932 213952
rect 132716 214008 135463 214010
rect 132716 213952 135402 214008
rect 135458 213952 135463 214008
rect 132716 213950 135463 213952
rect 103105 213947 103171 213950
rect 135397 213947 135463 213950
rect 174221 214010 174287 214013
rect 174221 214008 177060 214010
rect 174221 213952 174226 214008
rect 174282 213952 177060 214008
rect 174221 213950 177060 213952
rect 174221 213947 174287 213950
rect 100989 213874 101055 213877
rect 172013 213874 172079 213877
rect 97726 213872 101055 213874
rect 97726 213816 100994 213872
rect 101050 213816 101055 213872
rect 97726 213814 101055 213816
rect 65017 213466 65083 213469
rect 65017 213464 67978 213466
rect 65017 213408 65022 213464
rect 65078 213408 67978 213464
rect 65017 213406 67978 213408
rect 65017 213403 65083 213406
rect 62533 213330 62599 213333
rect 60588 213328 62599 213330
rect 60588 213272 62538 213328
rect 62594 213272 62599 213328
rect 67918 213300 67978 213406
rect 97726 213300 97786 213814
rect 100989 213811 101055 213814
rect 169670 213872 172079 213874
rect 169670 213816 172018 213872
rect 172074 213816 172079 213872
rect 169670 213814 172079 213816
rect 102369 213330 102435 213333
rect 135029 213330 135095 213333
rect 102369 213328 104932 213330
rect 60588 213270 62599 213272
rect 62533 213267 62599 213270
rect 102369 213272 102374 213328
rect 102430 213272 104932 213328
rect 102369 213270 104932 213272
rect 132716 213328 135095 213330
rect 132716 213272 135034 213328
rect 135090 213272 135095 213328
rect 132716 213270 135095 213272
rect 102369 213267 102435 213270
rect 135029 213267 135095 213270
rect 136777 213330 136843 213333
rect 136777 213328 140076 213330
rect 136777 213272 136782 213328
rect 136838 213272 140076 213328
rect 169670 213300 169730 213814
rect 172013 213811 172079 213814
rect 174037 213330 174103 213333
rect 174037 213328 177060 213330
rect 136777 213270 140076 213272
rect 174037 213272 174042 213328
rect 174098 213272 177060 213328
rect 174037 213270 177060 213272
rect 136777 213267 136843 213270
rect 174037 213267 174103 213270
rect 172657 213058 172723 213061
rect 169670 213056 172723 213058
rect 169670 213000 172662 213056
rect 172718 213000 172723 213056
rect 169670 212998 172723 213000
rect 66397 212786 66463 212789
rect 100989 212786 101055 212789
rect 66397 212784 67948 212786
rect 66397 212728 66402 212784
rect 66458 212728 67948 212784
rect 66397 212726 67948 212728
rect 97756 212784 101055 212786
rect 97756 212728 100994 212784
rect 101050 212728 101055 212784
rect 97756 212726 101055 212728
rect 66397 212723 66463 212726
rect 100989 212723 101055 212726
rect 136869 212786 136935 212789
rect 136869 212784 140076 212786
rect 136869 212728 136874 212784
rect 136930 212728 140076 212784
rect 169670 212756 169730 212998
rect 172657 212995 172723 212998
rect 136869 212726 140076 212728
rect 136869 212723 136935 212726
rect 62349 212650 62415 212653
rect 60588 212648 62415 212650
rect 60588 212592 62354 212648
rect 62410 212592 62415 212648
rect 60588 212590 62415 212592
rect 62349 212587 62415 212590
rect 102461 212650 102527 212653
rect 135397 212650 135463 212653
rect 102461 212648 104932 212650
rect 102461 212592 102466 212648
rect 102522 212592 104932 212648
rect 102461 212590 104932 212592
rect 132716 212648 135463 212650
rect 132716 212592 135402 212648
rect 135458 212592 135463 212648
rect 132716 212590 135463 212592
rect 102461 212587 102527 212590
rect 135397 212587 135463 212590
rect 174221 212650 174287 212653
rect 174221 212648 177060 212650
rect 174221 212592 174226 212648
rect 174282 212592 177060 212648
rect 174221 212590 177060 212592
rect 174221 212587 174287 212590
rect 172657 212514 172723 212517
rect 169670 212512 172723 212514
rect 169670 212456 172662 212512
rect 172718 212456 172723 212512
rect 169670 212454 172723 212456
rect 100529 212106 100595 212109
rect 97756 212104 100595 212106
rect 62625 211970 62691 211973
rect 60588 211968 62691 211970
rect 60588 211912 62630 211968
rect 62686 211912 62691 211968
rect 60588 211910 62691 211912
rect 62625 211907 62691 211910
rect 65017 211834 65083 211837
rect 67918 211834 67978 212076
rect 97756 212048 100534 212104
rect 100590 212048 100595 212104
rect 97756 212046 100595 212048
rect 100529 212043 100595 212046
rect 137053 212106 137119 212109
rect 137053 212104 140076 212106
rect 137053 212048 137058 212104
rect 137114 212048 140076 212104
rect 169670 212076 169730 212454
rect 172657 212451 172723 212454
rect 137053 212046 140076 212048
rect 137053 212043 137119 212046
rect 102369 211970 102435 211973
rect 135397 211970 135463 211973
rect 102369 211968 104932 211970
rect 102369 211912 102374 211968
rect 102430 211912 104932 211968
rect 102369 211910 104932 211912
rect 132716 211968 135463 211970
rect 132716 211912 135402 211968
rect 135458 211912 135463 211968
rect 132716 211910 135463 211912
rect 102369 211907 102435 211910
rect 135397 211907 135463 211910
rect 174037 211970 174103 211973
rect 174037 211968 177060 211970
rect 174037 211912 174042 211968
rect 174098 211912 177060 211968
rect 174037 211910 177060 211912
rect 174037 211907 174103 211910
rect 65017 211832 67978 211834
rect 65017 211776 65022 211832
rect 65078 211776 67978 211832
rect 65017 211774 67978 211776
rect 65017 211771 65083 211774
rect 172657 211698 172723 211701
rect 169670 211696 172723 211698
rect 169670 211640 172662 211696
rect 172718 211640 172723 211696
rect 169670 211638 172723 211640
rect 65661 211562 65727 211565
rect 100805 211562 100871 211565
rect 65661 211560 67948 211562
rect 65661 211504 65666 211560
rect 65722 211504 67948 211560
rect 65661 211502 67948 211504
rect 97756 211560 100871 211562
rect 97756 211504 100810 211560
rect 100866 211504 100871 211560
rect 97756 211502 100871 211504
rect 65661 211499 65727 211502
rect 100805 211499 100871 211502
rect 136961 211562 137027 211565
rect 136961 211560 140076 211562
rect 136961 211504 136966 211560
rect 137022 211504 140076 211560
rect 169670 211532 169730 211638
rect 172657 211635 172723 211638
rect 204806 211636 204812 211700
rect 204876 211636 204882 211700
rect 136961 211502 140076 211504
rect 136961 211499 137027 211502
rect 62533 211290 62599 211293
rect 172381 211290 172447 211293
rect 60588 211288 62599 211290
rect 60588 211232 62538 211288
rect 62594 211232 62599 211288
rect 169670 211288 172447 211290
rect 60588 211230 62599 211232
rect 62533 211227 62599 211230
rect 100989 211018 101055 211021
rect 97756 211016 101055 211018
rect 62625 210610 62691 210613
rect 60588 210608 62691 210610
rect 60588 210552 62630 210608
rect 62686 210552 62691 210608
rect 60588 210550 62691 210552
rect 62625 210547 62691 210550
rect 65017 210610 65083 210613
rect 67918 210610 67978 210988
rect 97756 210960 100994 211016
rect 101050 210960 101055 211016
rect 97756 210958 101055 210960
rect 100989 210955 101055 210958
rect 103657 210882 103723 210885
rect 104902 210882 104962 211260
rect 103657 210880 104962 210882
rect 103657 210824 103662 210880
rect 103718 210824 104962 210880
rect 103657 210822 104962 210824
rect 132686 210882 132746 211260
rect 169670 211232 172386 211288
rect 172442 211232 172447 211288
rect 169670 211230 172447 211232
rect 136869 211018 136935 211021
rect 136869 211016 140076 211018
rect 136869 210960 136874 211016
rect 136930 210960 140076 211016
rect 169670 210988 169730 211230
rect 172381 211227 172447 211230
rect 174221 211290 174287 211293
rect 174221 211288 177060 211290
rect 174221 211232 174226 211288
rect 174282 211232 177060 211288
rect 174221 211230 177060 211232
rect 174221 211227 174287 211230
rect 204814 211124 204874 211636
rect 223533 211154 223599 211157
rect 227416 211154 227896 211184
rect 223533 211152 227896 211154
rect 223533 211096 223538 211152
rect 223594 211096 227896 211152
rect 223533 211094 227896 211096
rect 223533 211091 223599 211094
rect 227416 211064 227896 211094
rect 136869 210958 140076 210960
rect 136869 210955 136935 210958
rect 132686 210822 133114 210882
rect 103657 210819 103723 210822
rect 133054 210746 133114 210822
rect 133054 210686 140106 210746
rect 65017 210608 67978 210610
rect 65017 210552 65022 210608
rect 65078 210552 67978 210608
rect 65017 210550 67978 210552
rect 102369 210610 102435 210613
rect 134661 210610 134727 210613
rect 102369 210608 104932 210610
rect 102369 210552 102374 210608
rect 102430 210552 104932 210608
rect 102369 210550 104932 210552
rect 132716 210608 134727 210610
rect 132716 210552 134666 210608
rect 134722 210552 134727 210608
rect 132716 210550 134727 210552
rect 65017 210547 65083 210550
rect 102369 210547 102435 210550
rect 134661 210547 134727 210550
rect 64925 210474 64991 210477
rect 65661 210474 65727 210477
rect 64925 210472 65727 210474
rect 64925 210416 64930 210472
rect 64986 210416 65666 210472
rect 65722 210416 65727 210472
rect 64925 210414 65727 210416
rect 64925 210411 64991 210414
rect 65661 210411 65727 210414
rect 65477 210338 65543 210341
rect 100897 210338 100963 210341
rect 65477 210336 67948 210338
rect 65477 210280 65482 210336
rect 65538 210280 67948 210336
rect 65477 210278 67948 210280
rect 97756 210336 100963 210338
rect 97756 210280 100902 210336
rect 100958 210280 100963 210336
rect 140046 210308 140106 210686
rect 172657 210610 172723 210613
rect 169670 210608 172723 210610
rect 169670 210552 172662 210608
rect 172718 210552 172723 210608
rect 169670 210550 172723 210552
rect 169670 210308 169730 210550
rect 172657 210547 172723 210550
rect 174037 210610 174103 210613
rect 174037 210608 177060 210610
rect 174037 210552 174042 210608
rect 174098 210552 177060 210608
rect 174037 210550 177060 210552
rect 174037 210547 174103 210550
rect 97756 210278 100963 210280
rect 65477 210275 65543 210278
rect 100897 210275 100963 210278
rect 172657 210066 172723 210069
rect 169670 210064 172723 210066
rect 169670 210008 172662 210064
rect 172718 210008 172723 210064
rect 169670 210006 172723 210008
rect 62625 209930 62691 209933
rect 60588 209928 62691 209930
rect 60588 209872 62630 209928
rect 62686 209872 62691 209928
rect 60588 209870 62691 209872
rect 62625 209867 62691 209870
rect 100989 209794 101055 209797
rect 97756 209792 101055 209794
rect 65017 209386 65083 209389
rect 67918 209386 67978 209764
rect 97756 209736 100994 209792
rect 101050 209736 101055 209792
rect 97756 209734 101055 209736
rect 100989 209731 101055 209734
rect 104902 209522 104962 209900
rect 65017 209384 67978 209386
rect 65017 209328 65022 209384
rect 65078 209328 67978 209384
rect 65017 209326 67978 209328
rect 97726 209462 104962 209522
rect 132686 209522 132746 209900
rect 136869 209794 136935 209797
rect 136869 209792 140076 209794
rect 136869 209736 136874 209792
rect 136930 209736 140076 209792
rect 169670 209764 169730 210006
rect 172657 210003 172723 210006
rect 174129 209930 174195 209933
rect 174129 209928 177060 209930
rect 174129 209872 174134 209928
rect 174190 209872 177060 209928
rect 174129 209870 177060 209872
rect 174129 209867 174195 209870
rect 136869 209734 140076 209736
rect 136869 209731 136935 209734
rect 132686 209462 140106 209522
rect 65017 209323 65083 209326
rect 62717 209250 62783 209253
rect 60588 209248 62783 209250
rect 60588 209192 62722 209248
rect 62778 209192 62783 209248
rect 60588 209190 62783 209192
rect 62717 209187 62783 209190
rect 66397 209114 66463 209117
rect 66397 209112 67948 209114
rect 66397 209056 66402 209112
rect 66458 209056 67948 209112
rect 97726 209084 97786 209462
rect 135305 209250 135371 209253
rect 132716 209248 135371 209250
rect 66397 209054 67948 209056
rect 66397 209051 66463 209054
rect 104902 208978 104962 209220
rect 132716 209192 135310 209248
rect 135366 209192 135371 209248
rect 132716 209190 135371 209192
rect 135305 209187 135371 209190
rect 140046 209084 140106 209462
rect 171645 209386 171711 209389
rect 169670 209384 171711 209386
rect 169670 209328 171650 209384
rect 171706 209328 171711 209384
rect 169670 209326 171711 209328
rect 169670 209084 169730 209326
rect 171645 209323 171711 209326
rect 174589 209250 174655 209253
rect 174589 209248 177060 209250
rect 174589 209192 174594 209248
rect 174650 209192 177060 209248
rect 174589 209190 177060 209192
rect 174589 209187 174655 209190
rect 101038 208918 104962 208978
rect 101038 208842 101098 208918
rect 172105 208842 172171 208845
rect 97726 208782 101098 208842
rect 169670 208840 172171 208842
rect 169670 208784 172110 208840
rect 172166 208784 172171 208840
rect 169670 208782 172171 208784
rect 62625 208570 62691 208573
rect 60588 208568 62691 208570
rect 60588 208512 62630 208568
rect 62686 208512 62691 208568
rect 60588 208510 62691 208512
rect 62625 208507 62691 208510
rect 65845 208570 65911 208573
rect 65845 208568 67948 208570
rect 65845 208512 65850 208568
rect 65906 208512 67948 208568
rect 97726 208540 97786 208782
rect 137697 208570 137763 208573
rect 137697 208568 140076 208570
rect 65845 208510 67948 208512
rect 65845 208507 65911 208510
rect 104902 208298 104962 208540
rect 97726 208238 104962 208298
rect 132686 208298 132746 208540
rect 137697 208512 137702 208568
rect 137758 208512 140076 208568
rect 169670 208540 169730 208782
rect 172105 208779 172171 208782
rect 137697 208510 140076 208512
rect 137697 208507 137763 208510
rect 132686 208238 140106 208298
rect 66397 208026 66463 208029
rect 66397 208024 67948 208026
rect 66397 207968 66402 208024
rect 66458 207968 67948 208024
rect 97726 207996 97786 208238
rect 140046 207996 140106 208238
rect 177030 208162 177090 208540
rect 169670 208102 177090 208162
rect 169670 207996 169730 208102
rect 66397 207966 67948 207968
rect 66397 207963 66463 207966
rect 63637 207890 63703 207893
rect 135397 207890 135463 207893
rect 60588 207888 63703 207890
rect 60588 207832 63642 207888
rect 63698 207832 63703 207888
rect 132716 207888 135463 207890
rect 60588 207830 63703 207832
rect 63637 207827 63703 207830
rect 65017 207618 65083 207621
rect 65845 207618 65911 207621
rect 104902 207618 104962 207860
rect 132716 207832 135402 207888
rect 135458 207832 135463 207888
rect 132716 207830 135463 207832
rect 135397 207827 135463 207830
rect 177030 207618 177090 207860
rect 65017 207616 65911 207618
rect 65017 207560 65022 207616
rect 65078 207560 65850 207616
rect 65906 207560 65911 207616
rect 65017 207558 65911 207560
rect 65017 207555 65083 207558
rect 65845 207555 65911 207558
rect 102326 207558 104962 207618
rect 174086 207558 177090 207618
rect 102326 207482 102386 207558
rect 174086 207482 174146 207558
rect 97726 207422 102386 207482
rect 169670 207422 174146 207482
rect 65293 207346 65359 207349
rect 65293 207344 67948 207346
rect 65293 207288 65298 207344
rect 65354 207288 67948 207344
rect 97726 207316 97786 207422
rect 136869 207346 136935 207349
rect 136869 207344 140076 207346
rect 65293 207286 67948 207288
rect 136869 207288 136874 207344
rect 136930 207288 140076 207344
rect 169670 207316 169730 207422
rect 136869 207286 140076 207288
rect 65293 207283 65359 207286
rect 136869 207283 136935 207286
rect 62533 207210 62599 207213
rect 60588 207208 62599 207210
rect 60588 207152 62538 207208
rect 62594 207152 62599 207208
rect 174129 207210 174195 207213
rect 174129 207208 177060 207210
rect 60588 207150 62599 207152
rect 62533 207147 62599 207150
rect 65661 206802 65727 206805
rect 104902 206802 104962 207180
rect 65661 206800 67948 206802
rect 65661 206744 65666 206800
rect 65722 206744 67948 206800
rect 65661 206742 67948 206744
rect 97756 206742 104962 206802
rect 132686 206802 132746 207180
rect 174129 207152 174134 207208
rect 174190 207152 177060 207208
rect 174129 207150 177060 207152
rect 174129 207147 174195 207150
rect 132686 206742 140076 206802
rect 65661 206739 65727 206742
rect 169854 206666 169914 206772
rect 171645 206666 171711 206669
rect 169854 206664 171711 206666
rect 169854 206608 171650 206664
rect 171706 206608 171711 206664
rect 169854 206606 171711 206608
rect 171645 206603 171711 206606
rect 62625 206530 62691 206533
rect 135397 206530 135463 206533
rect 60588 206528 62691 206530
rect 60588 206472 62630 206528
rect 62686 206472 62691 206528
rect 132716 206528 135463 206530
rect 60588 206470 62691 206472
rect 62625 206467 62691 206470
rect 104902 206258 104962 206500
rect 132716 206472 135402 206528
rect 135458 206472 135463 206528
rect 132716 206470 135463 206472
rect 135397 206467 135463 206470
rect 174037 206530 174103 206533
rect 174037 206528 177060 206530
rect 174037 206472 174042 206528
rect 174098 206472 177060 206528
rect 174037 206470 177060 206472
rect 174037 206467 174103 206470
rect 102326 206198 104962 206258
rect 102326 206122 102386 206198
rect 62625 205850 62691 205853
rect 60588 205848 62691 205850
rect 60588 205792 62630 205848
rect 62686 205792 62691 205848
rect 60588 205790 62691 205792
rect 62625 205787 62691 205790
rect 67918 205714 67978 206092
rect 97756 206062 102386 206122
rect 136869 206122 136935 206125
rect 136869 206120 140076 206122
rect 136869 206064 136874 206120
rect 136930 206064 140076 206120
rect 136869 206062 140076 206064
rect 136869 206059 136935 206062
rect 169854 205986 169914 206092
rect 171829 205986 171895 205989
rect 169854 205984 171895 205986
rect 169854 205928 171834 205984
rect 171890 205928 171895 205984
rect 169854 205926 171895 205928
rect 171829 205923 171895 205926
rect 65158 205654 67978 205714
rect 65158 205578 65218 205654
rect 65112 205518 65218 205578
rect 66397 205578 66463 205581
rect 104902 205578 104962 205820
rect 132716 205790 140106 205850
rect 66397 205576 67948 205578
rect 66397 205520 66402 205576
rect 66458 205520 67948 205576
rect 66397 205518 67948 205520
rect 97756 205518 104962 205578
rect 140046 205548 140106 205790
rect 64925 205306 64991 205309
rect 65112 205306 65172 205518
rect 66397 205515 66463 205518
rect 169854 205442 169914 205548
rect 177030 205442 177090 205820
rect 169854 205382 177090 205442
rect 64925 205304 65172 205306
rect 64925 205248 64930 205304
rect 64986 205248 65172 205304
rect 64925 205246 65172 205248
rect 169670 205246 176538 205306
rect 64925 205243 64991 205246
rect 60558 204898 60618 205140
rect 104902 205034 104962 205140
rect 132716 205110 140106 205170
rect 67918 204898 67978 205004
rect 97756 204974 104962 205034
rect 140046 205004 140106 205110
rect 169670 205004 169730 205246
rect 176478 205238 176538 205246
rect 176478 205178 177060 205238
rect 60558 204838 67978 204898
rect 62625 204490 62691 204493
rect 60588 204488 62691 204490
rect 60588 204432 62630 204488
rect 62686 204432 62691 204488
rect 60588 204430 62691 204432
rect 62625 204427 62691 204430
rect 65661 204354 65727 204357
rect 104902 204354 104962 204460
rect 132716 204430 140106 204490
rect 65661 204352 67948 204354
rect 65661 204296 65666 204352
rect 65722 204296 67948 204352
rect 65661 204294 67948 204296
rect 97756 204294 104962 204354
rect 140046 204324 140106 204430
rect 65661 204291 65727 204294
rect 169854 204218 169914 204324
rect 177030 204218 177090 204460
rect 169854 204158 177090 204218
rect 169670 203886 176538 203946
rect 62533 203810 62599 203813
rect 60588 203808 62599 203810
rect 60588 203752 62538 203808
rect 62594 203752 62599 203808
rect 60588 203750 62599 203752
rect 62533 203747 62599 203750
rect 65477 203810 65543 203813
rect 65477 203808 67948 203810
rect 65477 203752 65482 203808
rect 65538 203752 67948 203808
rect 65477 203750 67948 203752
rect 97756 203750 104932 203810
rect 132716 203750 140076 203810
rect 169670 203780 169730 203886
rect 176478 203878 176538 203886
rect 176478 203818 177060 203878
rect 65477 203747 65543 203750
rect 60558 203342 67978 203402
rect 60558 203100 60618 203342
rect 67918 203100 67978 203342
rect 97756 203070 104932 203130
rect 132716 203070 140076 203130
rect 169854 202994 169914 203100
rect 177030 202994 177090 203100
rect 169854 202934 177090 202994
rect 169670 202662 177090 202722
rect 169670 202556 169730 202662
rect 60558 202178 60618 202420
rect 67918 202178 67978 202556
rect 177030 202488 177090 202662
rect 97726 202450 97786 202488
rect 140046 202450 140106 202488
rect 97726 202390 104932 202450
rect 132716 202390 140106 202450
rect 60558 202118 67978 202178
rect 60558 201634 60618 201740
rect 67918 201634 67978 202012
rect 97726 201770 97786 201944
rect 140046 201770 140106 201944
rect 97726 201710 104932 201770
rect 132716 201710 140106 201770
rect 169854 201770 169914 202012
rect 207893 201770 207959 201773
rect 169854 201710 177060 201770
rect 204844 201768 207959 201770
rect 204844 201712 207898 201768
rect 207954 201712 207959 201768
rect 204844 201710 207959 201712
rect 207893 201707 207959 201710
rect 60558 201574 67978 201634
rect 60558 200954 60618 201060
rect 67918 200954 67978 201332
rect 97726 201090 97786 201264
rect 140046 201090 140106 201264
rect 169854 201226 169914 201332
rect 169854 201166 176538 201226
rect 176478 201158 176538 201166
rect 176478 201098 177060 201158
rect 97726 201030 104932 201090
rect 132716 201030 140106 201090
rect 60558 200894 67978 200954
rect 67918 200682 67978 200788
rect 63640 200622 67978 200682
rect 97726 200682 97786 200720
rect 100897 200682 100963 200685
rect 97726 200680 100963 200682
rect 97726 200624 100902 200680
rect 100958 200624 100963 200680
rect 97726 200622 100963 200624
rect 63640 200546 63700 200622
rect 100897 200619 100963 200622
rect 136777 200682 136843 200685
rect 140046 200682 140106 200720
rect 136777 200680 140106 200682
rect 136777 200624 136782 200680
rect 136838 200624 140106 200680
rect 136777 200622 140106 200624
rect 169854 200682 169914 200788
rect 169854 200622 174146 200682
rect 136777 200619 136843 200622
rect 60558 200486 63700 200546
rect 174086 200546 174146 200622
rect 174086 200486 176538 200546
rect 60558 200380 60618 200486
rect 176478 200478 176538 200486
rect 176478 200418 177060 200478
rect 65017 200410 65083 200413
rect 66397 200410 66463 200413
rect 65017 200408 66463 200410
rect 65017 200352 65022 200408
rect 65078 200352 66402 200408
rect 66458 200352 66463 200408
rect 65017 200350 66463 200352
rect 65017 200347 65083 200350
rect 66397 200347 66463 200350
rect 102369 200410 102435 200413
rect 135397 200410 135463 200413
rect 102369 200408 104932 200410
rect 102369 200352 102374 200408
rect 102430 200352 104932 200408
rect 102369 200350 104932 200352
rect 132716 200408 135463 200410
rect 132716 200352 135402 200408
rect 135458 200352 135463 200408
rect 132716 200350 135463 200352
rect 102369 200347 102435 200350
rect 135397 200347 135463 200350
rect 65109 200138 65175 200141
rect 65109 200136 67948 200138
rect 65109 200080 65114 200136
rect 65170 200080 67948 200136
rect 65109 200078 67948 200080
rect 65109 200075 65175 200078
rect 97726 199730 97786 200040
rect 140046 199730 140106 200040
rect 169854 200002 169914 200108
rect 169854 199942 177090 200002
rect 177030 199768 177090 199942
rect 60558 199322 60618 199700
rect 97726 199670 104932 199730
rect 132716 199670 140106 199730
rect 66397 199594 66463 199597
rect 66397 199592 67948 199594
rect 66397 199536 66402 199592
rect 66458 199536 67948 199592
rect 66397 199534 67948 199536
rect 66397 199531 66463 199534
rect 65109 199322 65175 199325
rect 60558 199320 65175 199322
rect 60558 199264 65114 199320
rect 65170 199264 65175 199320
rect 60558 199262 65175 199264
rect 97726 199322 97786 199496
rect 136777 199458 136843 199461
rect 140046 199458 140106 199496
rect 136777 199456 140106 199458
rect 136777 199400 136782 199456
rect 136838 199400 140106 199456
rect 136777 199398 140106 199400
rect 169854 199458 169914 199564
rect 172197 199458 172263 199461
rect 169854 199456 172263 199458
rect 169854 199400 172202 199456
rect 172258 199400 172263 199456
rect 169854 199398 172263 199400
rect 136777 199395 136843 199398
rect 172197 199395 172263 199398
rect 100897 199322 100963 199325
rect 97726 199320 100963 199322
rect 97726 199264 100902 199320
rect 100958 199264 100963 199320
rect 97726 199262 100963 199264
rect 65109 199259 65175 199262
rect 100897 199259 100963 199262
rect 62349 199050 62415 199053
rect 60588 199048 62415 199050
rect 60588 198992 62354 199048
rect 62410 198992 62415 199048
rect 102369 199050 102435 199053
rect 134753 199050 134819 199053
rect 102369 199048 104932 199050
rect 60588 198990 62415 198992
rect 62349 198987 62415 198990
rect 67918 198642 67978 199020
rect 102369 198992 102374 199048
rect 102430 198992 104932 199048
rect 102369 198990 104932 198992
rect 132716 199048 134819 199050
rect 132716 198992 134758 199048
rect 134814 198992 134819 199048
rect 175233 199050 175299 199053
rect 175233 199048 177060 199050
rect 132716 198990 134819 198992
rect 102369 198987 102435 198990
rect 134753 198987 134819 198990
rect 97726 198778 97786 198952
rect 97726 198718 104962 198778
rect 60558 198582 67978 198642
rect 60558 198340 60618 198582
rect 104902 198340 104962 198718
rect 140046 198642 140106 198952
rect 169854 198778 169914 199020
rect 175233 198992 175238 199048
rect 175294 198992 177060 199048
rect 175233 198990 177060 198992
rect 175233 198987 175299 198990
rect 169854 198718 177090 198778
rect 132686 198582 140106 198642
rect 132686 198408 132746 198582
rect 177030 198408 177090 198718
rect 65017 197962 65083 197965
rect 67918 197962 67978 198340
rect 65017 197960 67978 197962
rect 65017 197904 65022 197960
rect 65078 197904 67978 197960
rect 65017 197902 67978 197904
rect 97726 197962 97786 198272
rect 100897 197962 100963 197965
rect 97726 197960 100963 197962
rect 97726 197904 100902 197960
rect 100958 197904 100963 197960
rect 97726 197902 100963 197904
rect 65017 197899 65083 197902
rect 100897 197899 100963 197902
rect 136777 197962 136843 197965
rect 140046 197962 140106 198272
rect 169854 198098 169914 198340
rect 172197 198098 172263 198101
rect 169854 198096 172263 198098
rect 169854 198040 172202 198096
rect 172258 198040 172263 198096
rect 169854 198038 172263 198040
rect 172197 198035 172263 198038
rect 136777 197960 140106 197962
rect 136777 197904 136782 197960
rect 136838 197904 140106 197960
rect 136777 197902 140106 197904
rect 136777 197899 136843 197902
rect 62625 197690 62691 197693
rect 60588 197688 62691 197690
rect 60588 197632 62630 197688
rect 62686 197632 62691 197688
rect 60588 197630 62691 197632
rect 62625 197627 62691 197630
rect 67918 197418 67978 197796
rect 60558 197358 67978 197418
rect 97726 197418 97786 197728
rect 102369 197690 102435 197693
rect 135397 197690 135463 197693
rect 102369 197688 104932 197690
rect 102369 197632 102374 197688
rect 102430 197632 104932 197688
rect 102369 197630 104932 197632
rect 132716 197688 135463 197690
rect 132716 197632 135402 197688
rect 135458 197632 135463 197688
rect 132716 197630 135463 197632
rect 102369 197627 102435 197630
rect 135397 197627 135463 197630
rect 140046 197418 140106 197728
rect 169854 197554 169914 197796
rect 174221 197690 174287 197693
rect 174221 197688 177060 197690
rect 174221 197632 174226 197688
rect 174282 197632 177060 197688
rect 174221 197630 177060 197632
rect 174221 197627 174287 197630
rect 169854 197494 177090 197554
rect 97726 197358 104962 197418
rect 60558 196980 60618 197358
rect 65017 196874 65083 196877
rect 67918 196874 67978 197116
rect 65017 196872 67978 196874
rect 65017 196816 65022 196872
rect 65078 196816 67978 196872
rect 65017 196814 67978 196816
rect 65017 196811 65083 196814
rect 97726 196738 97786 197048
rect 104902 196980 104962 197358
rect 132686 197358 140106 197418
rect 132686 197048 132746 197358
rect 100897 196738 100963 196741
rect 97726 196736 100963 196738
rect 97726 196680 100902 196736
rect 100958 196680 100963 196736
rect 97726 196678 100963 196680
rect 100897 196675 100963 196678
rect 136777 196738 136843 196741
rect 140046 196738 140106 197048
rect 169854 196874 169914 197116
rect 177030 197048 177090 197494
rect 172657 196874 172723 196877
rect 169854 196872 172723 196874
rect 169854 196816 172662 196872
rect 172718 196816 172723 196872
rect 169854 196814 172723 196816
rect 172657 196811 172723 196814
rect 172197 196738 172263 196741
rect 136777 196736 140106 196738
rect 136777 196680 136782 196736
rect 136838 196680 140106 196736
rect 136777 196678 140106 196680
rect 169670 196736 172263 196738
rect 169670 196680 172202 196736
rect 172258 196680 172263 196736
rect 169670 196678 172263 196680
rect 136777 196675 136843 196678
rect 66397 196602 66463 196605
rect 100897 196602 100963 196605
rect 66397 196600 67948 196602
rect 66397 196544 66402 196600
rect 66458 196544 67948 196600
rect 66397 196542 67948 196544
rect 97756 196600 100963 196602
rect 97756 196544 100902 196600
rect 100958 196544 100963 196600
rect 97756 196542 100963 196544
rect 66397 196539 66463 196542
rect 100897 196539 100963 196542
rect 136685 196602 136751 196605
rect 136685 196600 140076 196602
rect 136685 196544 136690 196600
rect 136746 196544 140076 196600
rect 169670 196572 169730 196678
rect 172197 196675 172263 196678
rect 136685 196542 140076 196544
rect 136685 196539 136751 196542
rect 62625 196330 62691 196333
rect 60588 196328 62691 196330
rect 60588 196272 62630 196328
rect 62686 196272 62691 196328
rect 60588 196270 62691 196272
rect 62625 196267 62691 196270
rect 102369 196330 102435 196333
rect 135397 196330 135463 196333
rect 102369 196328 104932 196330
rect 102369 196272 102374 196328
rect 102430 196272 104932 196328
rect 102369 196270 104932 196272
rect 132716 196328 135463 196330
rect 132716 196272 135402 196328
rect 135458 196272 135463 196328
rect 132716 196270 135463 196272
rect 102369 196267 102435 196270
rect 135397 196267 135463 196270
rect 174129 196330 174195 196333
rect 174129 196328 177060 196330
rect 174129 196272 174134 196328
rect 174190 196272 177060 196328
rect 174129 196270 177060 196272
rect 174129 196267 174195 196270
rect 174221 196194 174287 196197
rect 174221 196192 177090 196194
rect 174221 196136 174226 196192
rect 174282 196136 177090 196192
rect 174221 196134 177090 196136
rect 174221 196131 174287 196134
rect 134293 196058 134359 196061
rect 132686 196056 134359 196058
rect 63637 195650 63703 195653
rect 60588 195648 63703 195650
rect 60588 195592 63642 195648
rect 63698 195592 63703 195648
rect 60588 195590 63703 195592
rect 63637 195587 63703 195590
rect 65017 195650 65083 195653
rect 67918 195650 67978 196028
rect 132686 196000 134298 196056
rect 134354 196000 134359 196056
rect 132686 195998 134359 196000
rect 65017 195648 67978 195650
rect 65017 195592 65022 195648
rect 65078 195592 67978 195648
rect 65017 195590 67978 195592
rect 65017 195587 65083 195590
rect 97726 195514 97786 195960
rect 132686 195688 132746 195998
rect 134293 195995 134359 195998
rect 102461 195650 102527 195653
rect 102461 195648 104932 195650
rect 102461 195592 102466 195648
rect 102522 195592 104932 195648
rect 102461 195590 104932 195592
rect 102461 195587 102527 195590
rect 100713 195514 100779 195517
rect 97726 195512 100779 195514
rect 97726 195456 100718 195512
rect 100774 195456 100779 195512
rect 97726 195454 100779 195456
rect 100713 195451 100779 195454
rect 136869 195514 136935 195517
rect 140046 195514 140106 195960
rect 169854 195650 169914 196028
rect 177030 195688 177090 196134
rect 171461 195650 171527 195653
rect 169854 195648 171527 195650
rect 169854 195592 171466 195648
rect 171522 195592 171527 195648
rect 169854 195590 171527 195592
rect 171461 195587 171527 195590
rect 136869 195512 140106 195514
rect 136869 195456 136874 195512
rect 136930 195456 140106 195512
rect 136869 195454 140106 195456
rect 136869 195451 136935 195454
rect 66397 195378 66463 195381
rect 66397 195376 67948 195378
rect 66397 195320 66402 195376
rect 66458 195320 67948 195376
rect 66397 195318 67948 195320
rect 66397 195315 66463 195318
rect 97726 195242 97786 195280
rect 100897 195242 100963 195245
rect 97726 195240 100963 195242
rect 97726 195184 100902 195240
rect 100958 195184 100963 195240
rect 97726 195182 100963 195184
rect 100897 195179 100963 195182
rect 136777 195242 136843 195245
rect 140046 195242 140106 195280
rect 136777 195240 140106 195242
rect 136777 195184 136782 195240
rect 136838 195184 140106 195240
rect 136777 195182 140106 195184
rect 169854 195242 169914 195348
rect 172657 195242 172723 195245
rect 169854 195240 172723 195242
rect 169854 195184 172662 195240
rect 172718 195184 172723 195240
rect 169854 195182 172723 195184
rect 136777 195179 136843 195182
rect 172657 195179 172723 195182
rect 62625 194970 62691 194973
rect 60588 194968 62691 194970
rect 60588 194912 62630 194968
rect 62686 194912 62691 194968
rect 60588 194910 62691 194912
rect 62625 194907 62691 194910
rect 102461 194970 102527 194973
rect 135397 194970 135463 194973
rect 102461 194968 104932 194970
rect 102461 194912 102466 194968
rect 102522 194912 104932 194968
rect 102461 194910 104932 194912
rect 132716 194968 135463 194970
rect 132716 194912 135402 194968
rect 135458 194912 135463 194968
rect 132716 194910 135463 194912
rect 102461 194907 102527 194910
rect 135397 194907 135463 194910
rect 174129 194970 174195 194973
rect 174129 194968 177060 194970
rect 174129 194912 174134 194968
rect 174190 194912 177060 194968
rect 174129 194910 177060 194912
rect 174129 194907 174195 194910
rect 65109 194834 65175 194837
rect 135397 194834 135463 194837
rect 65109 194832 67948 194834
rect 65109 194776 65114 194832
rect 65170 194776 67948 194832
rect 65109 194774 67948 194776
rect 132686 194832 135463 194834
rect 132686 194776 135402 194832
rect 135458 194776 135463 194832
rect 174221 194834 174287 194837
rect 174221 194832 177090 194834
rect 132686 194774 135463 194776
rect 65109 194771 65175 194774
rect 65017 194426 65083 194429
rect 65017 194424 67978 194426
rect 65017 194368 65022 194424
rect 65078 194368 67978 194424
rect 65017 194366 67978 194368
rect 65017 194363 65083 194366
rect 62533 194290 62599 194293
rect 60588 194288 62599 194290
rect 60588 194232 62538 194288
rect 62594 194232 62599 194288
rect 60588 194230 62599 194232
rect 62533 194227 62599 194230
rect 67918 194124 67978 194366
rect 97726 194290 97786 194736
rect 132686 194328 132746 194774
rect 135397 194771 135463 194774
rect 100621 194290 100687 194293
rect 97726 194288 100687 194290
rect 97726 194232 100626 194288
rect 100682 194232 100687 194288
rect 97726 194230 100687 194232
rect 100621 194227 100687 194230
rect 102369 194290 102435 194293
rect 136777 194290 136843 194293
rect 140046 194290 140106 194736
rect 102369 194288 104932 194290
rect 102369 194232 102374 194288
rect 102430 194232 104932 194288
rect 102369 194230 104932 194232
rect 136777 194288 140106 194290
rect 136777 194232 136782 194288
rect 136838 194232 140106 194288
rect 136777 194230 140106 194232
rect 169854 194290 169914 194804
rect 174221 194776 174226 194832
rect 174282 194776 177090 194832
rect 174221 194774 177090 194776
rect 174221 194771 174287 194774
rect 177030 194328 177090 194774
rect 171553 194290 171619 194293
rect 169854 194288 171619 194290
rect 169854 194232 171558 194288
rect 171614 194232 171619 194288
rect 169854 194230 171619 194232
rect 102369 194227 102435 194230
rect 136777 194227 136843 194230
rect 171553 194227 171619 194230
rect 65109 193880 65175 193885
rect 65109 193824 65114 193880
rect 65170 193824 65175 193880
rect 65109 193819 65175 193824
rect 97726 193882 97786 194056
rect 100621 193882 100687 193885
rect 97726 193880 100687 193882
rect 97726 193824 100626 193880
rect 100682 193824 100687 193880
rect 97726 193822 100687 193824
rect 100621 193819 100687 193822
rect 136685 193882 136751 193885
rect 140046 193882 140106 194056
rect 169854 194018 169914 194124
rect 172657 194018 172723 194021
rect 169854 194016 172723 194018
rect 169854 193960 172662 194016
rect 172718 193960 172723 194016
rect 169854 193958 172723 193960
rect 172657 193955 172723 193958
rect 136685 193880 140106 193882
rect 136685 193824 136690 193880
rect 136746 193824 140106 193880
rect 136685 193822 140106 193824
rect 136685 193819 136751 193822
rect 65112 193746 65172 193819
rect 60558 193686 65172 193746
rect 60558 193580 60618 193686
rect 66397 193610 66463 193613
rect 102461 193610 102527 193613
rect 135397 193610 135463 193613
rect 66397 193608 67948 193610
rect 66397 193552 66402 193608
rect 66458 193552 67948 193608
rect 66397 193550 67948 193552
rect 102461 193608 104932 193610
rect 102461 193552 102466 193608
rect 102522 193552 104932 193608
rect 102461 193550 104932 193552
rect 132716 193608 135463 193610
rect 132716 193552 135402 193608
rect 135458 193552 135463 193608
rect 174129 193610 174195 193613
rect 174129 193608 177060 193610
rect 132716 193550 135463 193552
rect 66397 193547 66463 193550
rect 102461 193547 102527 193550
rect 135397 193547 135463 193550
rect 97726 193202 97786 193512
rect 135397 193474 135463 193477
rect 132686 193472 135463 193474
rect 132686 193416 135402 193472
rect 135458 193416 135463 193472
rect 132686 193414 135463 193416
rect 99701 193202 99767 193205
rect 97726 193200 99767 193202
rect 97726 193144 99706 193200
rect 99762 193144 99767 193200
rect 97726 193142 99767 193144
rect 99701 193139 99767 193142
rect 62349 192930 62415 192933
rect 60588 192928 62415 192930
rect 60588 192872 62354 192928
rect 62410 192872 62415 192928
rect 60588 192870 62415 192872
rect 62349 192867 62415 192870
rect 9896 192658 10376 192688
rect 12209 192658 12275 192661
rect 9896 192656 12275 192658
rect 9896 192600 12214 192656
rect 12270 192600 12275 192656
rect 9896 192598 12275 192600
rect 9896 192568 10376 192598
rect 12209 192595 12275 192598
rect 65017 192658 65083 192661
rect 67918 192658 67978 193036
rect 132686 192968 132746 193414
rect 135397 193411 135463 193414
rect 136777 193202 136843 193205
rect 140046 193202 140106 193512
rect 136777 193200 140106 193202
rect 136777 193144 136782 193200
rect 136838 193144 140106 193200
rect 136777 193142 140106 193144
rect 169854 193202 169914 193580
rect 174129 193552 174134 193608
rect 174190 193552 177060 193608
rect 174129 193550 177060 193552
rect 174129 193547 174195 193550
rect 174221 193474 174287 193477
rect 174221 193472 177090 193474
rect 174221 193416 174226 193472
rect 174282 193416 177090 193472
rect 174221 193414 177090 193416
rect 174221 193411 174287 193414
rect 171645 193202 171711 193205
rect 169854 193200 171711 193202
rect 169854 193144 171650 193200
rect 171706 193144 171711 193200
rect 169854 193142 171711 193144
rect 136777 193139 136843 193142
rect 171645 193139 171711 193142
rect 65017 192656 67978 192658
rect 65017 192600 65022 192656
rect 65078 192600 67978 192656
rect 65017 192598 67978 192600
rect 65017 192595 65083 192598
rect 64925 192522 64991 192525
rect 66397 192522 66463 192525
rect 64925 192520 66463 192522
rect 64925 192464 64930 192520
rect 64986 192464 66402 192520
rect 66458 192464 66463 192520
rect 64925 192462 66463 192464
rect 97726 192522 97786 192968
rect 102369 192930 102435 192933
rect 102369 192928 104932 192930
rect 102369 192872 102374 192928
rect 102430 192872 104932 192928
rect 102369 192870 104932 192872
rect 102369 192867 102435 192870
rect 100621 192522 100687 192525
rect 97726 192520 100687 192522
rect 97726 192464 100626 192520
rect 100682 192464 100687 192520
rect 97726 192462 100687 192464
rect 64925 192459 64991 192462
rect 66397 192459 66463 192462
rect 100621 192459 100687 192462
rect 136685 192522 136751 192525
rect 140046 192522 140106 192968
rect 169854 192794 169914 193036
rect 177030 192968 177090 193414
rect 172197 192794 172263 192797
rect 169854 192792 172263 192794
rect 169854 192736 172202 192792
rect 172258 192736 172263 192792
rect 169854 192734 172263 192736
rect 172197 192731 172263 192734
rect 207249 192522 207315 192525
rect 207566 192522 207572 192524
rect 136685 192520 140106 192522
rect 136685 192464 136690 192520
rect 136746 192464 140106 192520
rect 136685 192462 140106 192464
rect 204844 192520 207572 192522
rect 204844 192464 207254 192520
rect 207310 192464 207572 192520
rect 204844 192462 207572 192464
rect 136685 192459 136751 192462
rect 207249 192459 207315 192462
rect 207566 192460 207572 192462
rect 207636 192460 207642 192524
rect 66397 192386 66463 192389
rect 207249 192386 207315 192389
rect 207566 192386 207572 192388
rect 66397 192384 67948 192386
rect 66397 192328 66402 192384
rect 66458 192328 67948 192384
rect 207249 192384 207572 192386
rect 66397 192326 67948 192328
rect 66397 192323 66463 192326
rect 62533 192250 62599 192253
rect 60588 192248 62599 192250
rect 60588 192192 62538 192248
rect 62594 192192 62599 192248
rect 60588 192190 62599 192192
rect 62533 192187 62599 192190
rect 97726 191978 97786 192288
rect 102461 192250 102527 192253
rect 135397 192250 135463 192253
rect 102461 192248 104932 192250
rect 102461 192192 102466 192248
rect 102522 192192 104932 192248
rect 102461 192190 104932 192192
rect 132716 192248 135463 192250
rect 132716 192192 135402 192248
rect 135458 192192 135463 192248
rect 132716 192190 135463 192192
rect 102461 192187 102527 192190
rect 135397 192187 135463 192190
rect 134293 192114 134359 192117
rect 132686 192112 134359 192114
rect 132686 192056 134298 192112
rect 134354 192056 134359 192112
rect 132686 192054 134359 192056
rect 99885 191978 99951 191981
rect 97726 191976 99951 191978
rect 97726 191920 99890 191976
rect 99946 191920 99951 191976
rect 97726 191918 99951 191920
rect 99885 191915 99951 191918
rect 66305 191842 66371 191845
rect 66305 191840 67948 191842
rect 66305 191784 66310 191840
rect 66366 191784 67948 191840
rect 66305 191782 67948 191784
rect 66305 191779 66371 191782
rect 62349 191570 62415 191573
rect 60588 191568 62415 191570
rect 60588 191512 62354 191568
rect 62410 191512 62415 191568
rect 60588 191510 62415 191512
rect 62349 191507 62415 191510
rect 65017 191298 65083 191301
rect 66397 191298 66463 191301
rect 65017 191296 66463 191298
rect 65017 191240 65022 191296
rect 65078 191240 66402 191296
rect 66458 191240 66463 191296
rect 65017 191238 66463 191240
rect 97726 191298 97786 191744
rect 132686 191608 132746 192054
rect 134293 192051 134359 192054
rect 136777 191978 136843 191981
rect 140046 191978 140106 192288
rect 136777 191976 140106 191978
rect 136777 191920 136782 191976
rect 136838 191920 140106 191976
rect 136777 191918 140106 191920
rect 169854 191978 169914 192356
rect 207249 192328 207254 192384
rect 207310 192328 207572 192384
rect 207249 192326 207572 192328
rect 207249 192323 207315 192326
rect 207566 192324 207572 192326
rect 207636 192324 207642 192388
rect 174221 192250 174287 192253
rect 174221 192248 177060 192250
rect 174221 192192 174226 192248
rect 174282 192192 177060 192248
rect 174221 192190 177060 192192
rect 174221 192187 174287 192190
rect 174129 192114 174195 192117
rect 174129 192112 177090 192114
rect 174129 192056 174134 192112
rect 174190 192056 177090 192112
rect 174129 192054 177090 192056
rect 174129 192051 174195 192054
rect 172197 191978 172263 191981
rect 169854 191976 172263 191978
rect 169854 191920 172202 191976
rect 172258 191920 172263 191976
rect 169854 191918 172263 191920
rect 136777 191915 136843 191918
rect 172197 191915 172263 191918
rect 102369 191570 102435 191573
rect 102369 191568 104932 191570
rect 102369 191512 102374 191568
rect 102430 191512 104932 191568
rect 102369 191510 104932 191512
rect 102369 191507 102435 191510
rect 100621 191298 100687 191301
rect 97726 191296 100687 191298
rect 97726 191240 100626 191296
rect 100682 191240 100687 191296
rect 97726 191238 100687 191240
rect 65017 191235 65083 191238
rect 66397 191235 66463 191238
rect 100621 191235 100687 191238
rect 136685 191298 136751 191301
rect 140046 191298 140106 191744
rect 169854 191434 169914 191812
rect 177030 191608 177090 192054
rect 172657 191434 172723 191437
rect 169854 191432 172723 191434
rect 169854 191376 172662 191432
rect 172718 191376 172723 191432
rect 169854 191374 172723 191376
rect 172657 191371 172723 191374
rect 136685 191296 140106 191298
rect 136685 191240 136690 191296
rect 136746 191240 140106 191296
rect 136685 191238 140106 191240
rect 136685 191235 136751 191238
rect 65201 191162 65267 191165
rect 100897 191162 100963 191165
rect 65201 191160 67948 191162
rect 65201 191104 65206 191160
rect 65262 191104 67948 191160
rect 65201 191102 67948 191104
rect 97756 191160 100963 191162
rect 97756 191104 100902 191160
rect 100958 191104 100963 191160
rect 97756 191102 100963 191104
rect 65201 191099 65267 191102
rect 100897 191099 100963 191102
rect 136961 191162 137027 191165
rect 136961 191160 140076 191162
rect 136961 191104 136966 191160
rect 137022 191104 140076 191160
rect 136961 191102 140076 191104
rect 136961 191099 137027 191102
rect 169854 191026 169914 191132
rect 172657 191026 172723 191029
rect 169854 191024 172723 191026
rect 169854 190968 172662 191024
rect 172718 190968 172723 191024
rect 169854 190966 172723 190968
rect 172657 190963 172723 190966
rect 62625 190890 62691 190893
rect 60588 190888 62691 190890
rect 60588 190832 62630 190888
rect 62686 190832 62691 190888
rect 60588 190830 62691 190832
rect 62625 190827 62691 190830
rect 102277 190890 102343 190893
rect 135397 190890 135463 190893
rect 102277 190888 104932 190890
rect 102277 190832 102282 190888
rect 102338 190832 104932 190888
rect 102277 190830 104932 190832
rect 132716 190888 135463 190890
rect 132716 190832 135402 190888
rect 135458 190832 135463 190888
rect 132716 190830 135463 190832
rect 102277 190827 102343 190830
rect 135397 190827 135463 190830
rect 174037 190890 174103 190893
rect 174037 190888 177060 190890
rect 174037 190832 174042 190888
rect 174098 190832 177060 190888
rect 174037 190830 177060 190832
rect 174037 190827 174103 190830
rect 134753 190754 134819 190757
rect 132686 190752 134819 190754
rect 132686 190696 134758 190752
rect 134814 190696 134819 190752
rect 132686 190694 134819 190696
rect 66305 190618 66371 190621
rect 66305 190616 67948 190618
rect 66305 190560 66310 190616
rect 66366 190560 67948 190616
rect 66305 190558 67948 190560
rect 66305 190555 66371 190558
rect 62441 190210 62507 190213
rect 60588 190208 62507 190210
rect 60588 190152 62446 190208
rect 62502 190152 62507 190208
rect 60588 190150 62507 190152
rect 97726 190210 97786 190520
rect 132686 190248 132746 190694
rect 134753 190691 134819 190694
rect 173945 190754 174011 190757
rect 173945 190752 177090 190754
rect 173945 190696 173950 190752
rect 174006 190696 177090 190752
rect 173945 190694 177090 190696
rect 173945 190691 174011 190694
rect 100529 190210 100595 190213
rect 97726 190208 100595 190210
rect 97726 190152 100534 190208
rect 100590 190152 100595 190208
rect 97726 190150 100595 190152
rect 62441 190147 62507 190150
rect 100529 190147 100595 190150
rect 102185 190210 102251 190213
rect 136777 190210 136843 190213
rect 140046 190210 140106 190520
rect 102185 190208 104932 190210
rect 102185 190152 102190 190208
rect 102246 190152 104932 190208
rect 102185 190150 104932 190152
rect 136777 190208 140106 190210
rect 136777 190152 136782 190208
rect 136838 190152 140106 190208
rect 136777 190150 140106 190152
rect 169854 190210 169914 190588
rect 177030 190248 177090 190694
rect 172381 190210 172447 190213
rect 169854 190208 172447 190210
rect 169854 190152 172386 190208
rect 172442 190152 172447 190208
rect 169854 190150 172447 190152
rect 102185 190147 102251 190150
rect 136777 190147 136843 190150
rect 172381 190147 172447 190150
rect 66397 190074 66463 190077
rect 66397 190072 67948 190074
rect 66397 190016 66402 190072
rect 66458 190016 67948 190072
rect 66397 190014 67948 190016
rect 66397 190011 66463 190014
rect 97726 189938 97786 189976
rect 99885 189938 99951 189941
rect 97726 189936 99951 189938
rect 97726 189880 99890 189936
rect 99946 189880 99951 189936
rect 97726 189878 99951 189880
rect 99885 189875 99951 189878
rect 137421 189802 137487 189805
rect 140046 189802 140106 189976
rect 169854 189938 169914 190044
rect 172013 189938 172079 189941
rect 169854 189936 172079 189938
rect 169854 189880 172018 189936
rect 172074 189880 172079 189936
rect 169854 189878 172079 189880
rect 172013 189875 172079 189878
rect 137421 189800 140106 189802
rect 137421 189744 137426 189800
rect 137482 189744 140106 189800
rect 137421 189742 140106 189744
rect 137421 189739 137487 189742
rect 65017 189666 65083 189669
rect 66305 189666 66371 189669
rect 65017 189664 66371 189666
rect 65017 189608 65022 189664
rect 65078 189608 66310 189664
rect 66366 189608 66371 189664
rect 65017 189606 66371 189608
rect 65017 189603 65083 189606
rect 66305 189603 66371 189606
rect 62625 189530 62691 189533
rect 60588 189528 62691 189530
rect 60588 189472 62630 189528
rect 62686 189472 62691 189528
rect 60588 189470 62691 189472
rect 62625 189467 62691 189470
rect 102553 189530 102619 189533
rect 134293 189530 134359 189533
rect 102553 189528 104932 189530
rect 102553 189472 102558 189528
rect 102614 189472 104932 189528
rect 102553 189470 104932 189472
rect 132716 189528 134359 189530
rect 132716 189472 134298 189528
rect 134354 189472 134359 189528
rect 132716 189470 134359 189472
rect 102553 189467 102619 189470
rect 134293 189467 134359 189470
rect 174957 189530 175023 189533
rect 174957 189528 177060 189530
rect 174957 189472 174962 189528
rect 175018 189472 177060 189528
rect 174957 189470 177060 189472
rect 174957 189467 175023 189470
rect 134753 189258 134819 189261
rect 132686 189256 134819 189258
rect 132686 189200 134758 189256
rect 134814 189200 134819 189256
rect 132686 189198 134819 189200
rect 132686 188888 132746 189198
rect 134753 189195 134819 189198
rect 174405 189258 174471 189261
rect 174405 189256 177090 189258
rect 174405 189200 174410 189256
rect 174466 189200 177090 189256
rect 174405 189198 177090 189200
rect 174405 189195 174471 189198
rect 177030 188888 177090 189198
rect 62625 188850 62691 188853
rect 60588 188848 62691 188850
rect 60588 188792 62630 188848
rect 62686 188792 62691 188848
rect 60588 188790 62691 188792
rect 62625 188787 62691 188790
rect 102461 188850 102527 188853
rect 102461 188848 104932 188850
rect 102461 188792 102466 188848
rect 102522 188792 104932 188848
rect 102461 188790 104932 188792
rect 102461 188787 102527 188790
rect 63637 188170 63703 188173
rect 60588 188168 63703 188170
rect 60588 188112 63642 188168
rect 63698 188112 63703 188168
rect 60588 188110 63703 188112
rect 63637 188107 63703 188110
rect 102369 188170 102435 188173
rect 135029 188170 135095 188173
rect 102369 188168 104932 188170
rect 102369 188112 102374 188168
rect 102430 188112 104932 188168
rect 102369 188110 104932 188112
rect 132716 188168 135095 188170
rect 132716 188112 135034 188168
rect 135090 188112 135095 188168
rect 132716 188110 135095 188112
rect 102369 188107 102435 188110
rect 135029 188107 135095 188110
rect 175417 188170 175483 188173
rect 175417 188168 177060 188170
rect 175417 188112 175422 188168
rect 175478 188112 177060 188168
rect 175417 188110 177060 188112
rect 175417 188107 175483 188110
rect 225189 187354 225255 187357
rect 227416 187354 227896 187384
rect 225189 187352 227896 187354
rect 225189 187296 225194 187352
rect 225250 187296 227896 187352
rect 225189 187294 227896 187296
rect 225189 187291 225255 187294
rect 227416 187264 227896 187294
rect 117089 185450 117155 185453
rect 118193 185450 118259 185453
rect 117089 185448 118259 185450
rect 117089 185392 117094 185448
rect 117150 185392 118198 185448
rect 118254 185392 118259 185448
rect 117089 185390 118259 185392
rect 117089 185387 117155 185390
rect 118193 185387 118259 185390
rect 118653 185450 118719 185453
rect 120585 185450 120651 185453
rect 118653 185448 120651 185450
rect 118653 185392 118658 185448
rect 118714 185392 120590 185448
rect 120646 185392 120651 185448
rect 118653 185390 120651 185392
rect 118653 185387 118719 185390
rect 120585 185387 120651 185390
rect 120953 185450 121019 185453
rect 123437 185450 123503 185453
rect 120953 185448 123503 185450
rect 120953 185392 120958 185448
rect 121014 185392 123442 185448
rect 123498 185392 123503 185448
rect 120953 185390 123503 185392
rect 120953 185387 121019 185390
rect 123437 185387 123503 185390
rect 123897 185450 123963 185453
rect 125921 185450 125987 185453
rect 123897 185448 125987 185450
rect 123897 185392 123902 185448
rect 123958 185392 125926 185448
rect 125982 185392 125987 185448
rect 123897 185390 125987 185392
rect 123897 185387 123963 185390
rect 125921 185387 125987 185390
rect 126657 185450 126723 185453
rect 132177 185450 132243 185453
rect 126657 185448 132243 185450
rect 126657 185392 126662 185448
rect 126718 185392 132182 185448
rect 132238 185392 132243 185448
rect 126657 185390 132243 185392
rect 126657 185387 126723 185390
rect 132177 185387 132243 185390
rect 117457 185314 117523 185317
rect 118929 185314 118995 185317
rect 117457 185312 118995 185314
rect 117457 185256 117462 185312
rect 117518 185256 118934 185312
rect 118990 185256 118995 185312
rect 117457 185254 118995 185256
rect 117457 185251 117523 185254
rect 118929 185251 118995 185254
rect 121045 185314 121111 185317
rect 124357 185314 124423 185317
rect 125921 185314 125987 185317
rect 121045 185312 124423 185314
rect 121045 185256 121050 185312
rect 121106 185256 124362 185312
rect 124418 185256 124423 185312
rect 121045 185254 124423 185256
rect 121045 185251 121111 185254
rect 124357 185251 124423 185254
rect 124590 185312 125987 185314
rect 124590 185256 125926 185312
rect 125982 185256 125987 185312
rect 124590 185254 125987 185256
rect 118285 185178 118351 185181
rect 120309 185178 120375 185181
rect 118285 185176 120375 185178
rect 118285 185120 118290 185176
rect 118346 185120 120314 185176
rect 120370 185120 120375 185176
rect 118285 185118 120375 185120
rect 118285 185115 118351 185118
rect 120309 185115 120375 185118
rect 120585 185178 120651 185181
rect 123069 185178 123135 185181
rect 120585 185176 123135 185178
rect 120585 185120 120590 185176
rect 120646 185120 123074 185176
rect 123130 185120 123135 185176
rect 120585 185118 123135 185120
rect 120585 185115 120651 185118
rect 123069 185115 123135 185118
rect 123345 185178 123411 185181
rect 124590 185178 124650 185254
rect 125921 185251 125987 185254
rect 126105 185314 126171 185317
rect 131441 185314 131507 185317
rect 126105 185312 131507 185314
rect 126105 185256 126110 185312
rect 126166 185256 131446 185312
rect 131502 185256 131507 185312
rect 126105 185254 131507 185256
rect 126105 185251 126171 185254
rect 131441 185251 131507 185254
rect 123345 185176 124650 185178
rect 123345 185120 123350 185176
rect 123406 185120 124650 185176
rect 123345 185118 124650 185120
rect 125093 185178 125159 185181
rect 127209 185178 127275 185181
rect 125093 185176 127275 185178
rect 125093 185120 125098 185176
rect 125154 185120 127214 185176
rect 127270 185120 127275 185176
rect 125093 185118 127275 185120
rect 123345 185115 123411 185118
rect 125093 185115 125159 185118
rect 127209 185115 127275 185118
rect 37877 185042 37943 185045
rect 40269 185042 40335 185045
rect 37877 185040 40335 185042
rect 37877 184984 37882 185040
rect 37938 184984 40274 185040
rect 40330 184984 40335 185040
rect 37877 184982 40335 184984
rect 37877 184979 37943 184982
rect 40269 184979 40335 184982
rect 119113 185042 119179 185045
rect 121137 185042 121203 185045
rect 121689 185042 121755 185045
rect 119113 185040 121203 185042
rect 119113 184984 119118 185040
rect 119174 184984 121142 185040
rect 121198 184984 121203 185040
rect 119113 184982 121203 184984
rect 119113 184979 119179 184982
rect 121137 184979 121203 184982
rect 121278 185040 121755 185042
rect 121278 184984 121694 185040
rect 121750 184984 121755 185040
rect 121278 184982 121755 184984
rect 119665 184906 119731 184909
rect 121278 184906 121338 184982
rect 121689 184979 121755 184982
rect 122701 185042 122767 185045
rect 124817 185042 124883 185045
rect 122701 185040 124883 185042
rect 122701 184984 122706 185040
rect 122762 184984 124822 185040
rect 124878 184984 124883 185040
rect 122701 184982 124883 184984
rect 122701 184979 122767 184982
rect 124817 184979 124883 184982
rect 125461 185042 125527 185045
rect 127209 185042 127275 185045
rect 125461 185040 127275 185042
rect 125461 184984 125466 185040
rect 125522 184984 127214 185040
rect 127270 184984 127275 185040
rect 125461 184982 127275 184984
rect 125461 184979 125527 184982
rect 127209 184979 127275 184982
rect 197451 185042 197517 185045
rect 202189 185042 202255 185045
rect 197451 185040 202255 185042
rect 197451 184984 197456 185040
rect 197512 184984 202194 185040
rect 202250 184984 202255 185040
rect 197451 184982 202255 184984
rect 197451 184979 197517 184982
rect 202189 184979 202255 184982
rect 119665 184904 121338 184906
rect 119665 184848 119670 184904
rect 119726 184848 121338 184904
rect 119665 184846 121338 184848
rect 121597 184906 121663 184909
rect 124357 184906 124423 184909
rect 121597 184904 124423 184906
rect 121597 184848 121602 184904
rect 121658 184848 124362 184904
rect 124418 184848 124423 184904
rect 121597 184846 124423 184848
rect 119665 184843 119731 184846
rect 121597 184843 121663 184846
rect 124357 184843 124423 184846
rect 124909 184906 124975 184909
rect 127209 184906 127275 184909
rect 124909 184904 127275 184906
rect 124909 184848 124914 184904
rect 124970 184848 127214 184904
rect 127270 184848 127275 184904
rect 124909 184846 127275 184848
rect 124909 184843 124975 184846
rect 127209 184843 127275 184846
rect 105589 184770 105655 184773
rect 102694 184768 105655 184770
rect 102694 184712 105594 184768
rect 105650 184712 105655 184768
rect 102694 184710 105655 184712
rect 37969 184498 38035 184501
rect 39625 184498 39691 184501
rect 37969 184496 39691 184498
rect 37969 184440 37974 184496
rect 38030 184440 39630 184496
rect 39686 184440 39691 184496
rect 37969 184438 39691 184440
rect 37969 184435 38035 184438
rect 39625 184435 39691 184438
rect 54897 184226 54963 184229
rect 60141 184226 60207 184229
rect 54897 184224 60207 184226
rect 102694 184224 102754 184710
rect 105589 184707 105655 184710
rect 116905 184770 116971 184773
rect 117641 184770 117707 184773
rect 116905 184768 117707 184770
rect 116905 184712 116910 184768
rect 116966 184712 117646 184768
rect 117702 184712 117707 184768
rect 116905 184710 117707 184712
rect 116905 184707 116971 184710
rect 117641 184707 117707 184710
rect 118101 184770 118167 184773
rect 119573 184770 119639 184773
rect 118101 184768 119639 184770
rect 118101 184712 118106 184768
rect 118162 184712 119578 184768
rect 119634 184712 119639 184768
rect 118101 184710 119639 184712
rect 118101 184707 118167 184710
rect 119573 184707 119639 184710
rect 122517 184770 122583 184773
rect 125645 184770 125711 184773
rect 122517 184768 125711 184770
rect 122517 184712 122522 184768
rect 122578 184712 125650 184768
rect 125706 184712 125711 184768
rect 122517 184710 125711 184712
rect 122517 184707 122583 184710
rect 125645 184707 125711 184710
rect 126473 184770 126539 184773
rect 131625 184770 131691 184773
rect 126473 184768 131691 184770
rect 126473 184712 126478 184768
rect 126534 184712 131630 184768
rect 131686 184712 131691 184768
rect 126473 184710 131691 184712
rect 126473 184707 126539 184710
rect 131625 184707 131691 184710
rect 120125 184634 120191 184637
rect 122793 184634 122859 184637
rect 120125 184632 122859 184634
rect 120125 184576 120130 184632
rect 120186 184576 122798 184632
rect 122854 184576 122859 184632
rect 120125 184574 122859 184576
rect 120125 184571 120191 184574
rect 122793 184571 122859 184574
rect 124357 184634 124423 184637
rect 127025 184634 127091 184637
rect 124357 184632 127091 184634
rect 124357 184576 124362 184632
rect 124418 184576 127030 184632
rect 127086 184576 127091 184632
rect 124357 184574 127091 184576
rect 124357 184571 124423 184574
rect 127025 184571 127091 184574
rect 123713 184498 123779 184501
rect 127025 184498 127091 184501
rect 123713 184496 127091 184498
rect 123713 184440 123718 184496
rect 123774 184440 127030 184496
rect 127086 184440 127091 184496
rect 123713 184438 127091 184440
rect 123713 184435 123779 184438
rect 127025 184435 127091 184438
rect 198509 184498 198575 184501
rect 198877 184498 198943 184501
rect 203937 184498 204003 184501
rect 198509 184496 198802 184498
rect 198509 184440 198514 184496
rect 198570 184440 198802 184496
rect 198509 184438 198802 184440
rect 198509 184435 198575 184438
rect 198742 184362 198802 184438
rect 198877 184496 204003 184498
rect 198877 184440 198882 184496
rect 198938 184440 203942 184496
rect 203998 184440 204003 184496
rect 198877 184438 204003 184440
rect 198877 184435 198943 184438
rect 203937 184435 204003 184438
rect 203385 184362 203451 184365
rect 198742 184360 203451 184362
rect 198742 184304 203390 184360
rect 203446 184304 203451 184360
rect 198742 184302 203451 184304
rect 203385 184299 203451 184302
rect 177717 184226 177783 184229
rect 174852 184224 177783 184226
rect 54897 184168 54902 184224
rect 54958 184168 60146 184224
rect 60202 184168 60207 184224
rect 54897 184166 60207 184168
rect 174852 184168 177722 184224
rect 177778 184168 177783 184224
rect 174852 184166 177783 184168
rect 54897 184163 54963 184166
rect 60141 184163 60207 184166
rect 177717 184163 177783 184166
rect 106141 183546 106207 183549
rect 102694 183544 106207 183546
rect 102694 183488 106146 183544
rect 106202 183488 106207 183544
rect 102694 183486 106207 183488
rect 102694 183000 102754 183486
rect 106141 183483 106207 183486
rect 108533 183546 108599 183549
rect 180293 183546 180359 183549
rect 108533 183544 111004 183546
rect 108533 183488 108538 183544
rect 108594 183488 111004 183544
rect 108533 183486 111004 183488
rect 180293 183544 182948 183546
rect 180293 183488 180298 183544
rect 180354 183488 182948 183544
rect 180293 183486 182948 183488
rect 108533 183483 108599 183486
rect 180293 183483 180359 183486
rect 177441 183002 177507 183005
rect 207249 183002 207315 183005
rect 174852 183000 177507 183002
rect 174852 182944 177446 183000
rect 177502 182944 177507 183000
rect 174852 182942 177507 182944
rect 177441 182939 177507 182942
rect 207206 183000 207315 183002
rect 207206 182944 207254 183000
rect 207310 182944 207315 183000
rect 207206 182939 207315 182944
rect 207206 182868 207266 182939
rect 207198 182804 207204 182868
rect 207268 182804 207274 182868
rect 105589 182322 105655 182325
rect 102694 182320 105655 182322
rect 102694 182264 105594 182320
rect 105650 182264 105655 182320
rect 102694 182262 105655 182264
rect 102694 181776 102754 182262
rect 105589 182259 105655 182262
rect 176981 181778 177047 181781
rect 174852 181776 177047 181778
rect 174852 181720 176986 181776
rect 177042 181720 177047 181776
rect 174852 181718 177047 181720
rect 176981 181715 177047 181718
rect 108073 181234 108139 181237
rect 179741 181234 179807 181237
rect 108073 181232 111004 181234
rect 108073 181176 108078 181232
rect 108134 181176 111004 181232
rect 108073 181174 111004 181176
rect 179741 181232 182948 181234
rect 179741 181176 179746 181232
rect 179802 181176 182948 181232
rect 179741 181174 182948 181176
rect 108073 181171 108139 181174
rect 179741 181171 179807 181174
rect 106049 181098 106115 181101
rect 102694 181096 106115 181098
rect 102694 181040 106054 181096
rect 106110 181040 106115 181096
rect 102694 181038 106115 181040
rect 102694 180552 102754 181038
rect 106049 181035 106115 181038
rect 177073 180554 177139 180557
rect 174852 180552 177139 180554
rect 174852 180496 177078 180552
rect 177134 180496 177139 180552
rect 174852 180494 177139 180496
rect 177073 180491 177139 180494
rect 105957 179874 106023 179877
rect 102694 179872 106023 179874
rect 102694 179816 105962 179872
rect 106018 179816 106023 179872
rect 102694 179814 106023 179816
rect 12025 179738 12091 179741
rect 12025 179736 14036 179738
rect 12025 179680 12030 179736
rect 12086 179680 14036 179736
rect 12025 179678 14036 179680
rect 12025 179675 12091 179678
rect 102694 179328 102754 179814
rect 105957 179811 106023 179814
rect 225189 179738 225255 179741
rect 223796 179736 225255 179738
rect 223796 179680 225194 179736
rect 225250 179680 225255 179736
rect 223796 179678 225255 179680
rect 225189 179675 225255 179678
rect 177625 179330 177691 179333
rect 174852 179328 177691 179330
rect 174852 179272 177630 179328
rect 177686 179272 177691 179328
rect 174852 179270 177691 179272
rect 177625 179267 177691 179270
rect 107889 178922 107955 178925
rect 179741 178922 179807 178925
rect 107889 178920 111004 178922
rect 107889 178864 107894 178920
rect 107950 178864 111004 178920
rect 107889 178862 111004 178864
rect 179741 178920 182948 178922
rect 179741 178864 179746 178920
rect 179802 178864 182948 178920
rect 179741 178862 182948 178864
rect 107889 178859 107955 178862
rect 179741 178859 179807 178862
rect 105313 178514 105379 178517
rect 102694 178512 105379 178514
rect 102694 178456 105318 178512
rect 105374 178456 105379 178512
rect 102694 178454 105379 178456
rect 31989 178242 32055 178245
rect 29860 178240 32055 178242
rect 29860 178184 31994 178240
rect 32050 178184 32055 178240
rect 29860 178182 32055 178184
rect 31989 178179 32055 178182
rect 37417 178242 37483 178245
rect 59589 178242 59655 178245
rect 37417 178240 39060 178242
rect 37417 178184 37422 178240
rect 37478 178184 39060 178240
rect 37417 178182 39060 178184
rect 59589 178240 62980 178242
rect 59589 178184 59594 178240
rect 59650 178184 62980 178240
rect 59589 178182 62980 178184
rect 37417 178179 37483 178182
rect 59589 178179 59655 178182
rect 102694 178104 102754 178454
rect 105313 178451 105379 178454
rect 201085 178242 201151 178245
rect 126828 178182 134924 178242
rect 198772 178240 201151 178242
rect 198772 178184 201090 178240
rect 201146 178184 201151 178240
rect 198772 178182 201151 178184
rect 201085 178179 201151 178182
rect 204489 178242 204555 178245
rect 204489 178240 207972 178242
rect 204489 178184 204494 178240
rect 204550 178184 207972 178240
rect 204489 178182 207972 178184
rect 204489 178179 204555 178182
rect 177533 178106 177599 178109
rect 174852 178104 177599 178106
rect 174852 178048 177538 178104
rect 177594 178048 177599 178104
rect 174852 178046 177599 178048
rect 177533 178043 177599 178046
rect 105221 177154 105287 177157
rect 102694 177152 105287 177154
rect 102694 177096 105226 177152
rect 105282 177096 105287 177152
rect 102694 177094 105287 177096
rect 102694 176880 102754 177094
rect 105221 177091 105287 177094
rect 176981 176882 177047 176885
rect 174852 176880 177047 176882
rect 174852 176824 176986 176880
rect 177042 176824 177047 176880
rect 174852 176822 177047 176824
rect 176981 176819 177047 176822
rect 107889 176474 107955 176477
rect 179649 176474 179715 176477
rect 107889 176472 111004 176474
rect 107889 176416 107894 176472
rect 107950 176416 111004 176472
rect 107889 176414 111004 176416
rect 179649 176472 182948 176474
rect 179649 176416 179654 176472
rect 179710 176416 182948 176472
rect 179649 176414 182948 176416
rect 107889 176411 107955 176414
rect 179649 176411 179715 176414
rect 105129 175794 105195 175797
rect 103062 175792 105195 175794
rect 103062 175736 105134 175792
rect 105190 175736 105195 175792
rect 103062 175734 105195 175736
rect 103062 175686 103122 175734
rect 105129 175731 105195 175734
rect 102724 175626 103122 175686
rect 176889 175658 176955 175661
rect 174852 175656 176955 175658
rect 174852 175600 176894 175656
rect 176950 175600 176955 175656
rect 174852 175598 176955 175600
rect 176889 175595 176955 175598
rect 57565 174842 57631 174845
rect 54884 174840 57631 174842
rect 54884 174784 57570 174840
rect 57626 174784 57631 174840
rect 54884 174782 57631 174784
rect 57565 174779 57631 174782
rect 106141 174434 106207 174437
rect 177349 174434 177415 174437
rect 102724 174432 106207 174434
rect 102724 174376 106146 174432
rect 106202 174376 106207 174432
rect 102724 174374 106207 174376
rect 174852 174432 177415 174434
rect 174852 174376 177354 174432
rect 177410 174376 177415 174432
rect 174852 174374 177415 174376
rect 106141 174371 106207 174374
rect 177349 174371 177415 174374
rect 108165 174162 108231 174165
rect 179649 174162 179715 174165
rect 108165 174160 111004 174162
rect 108165 174104 108170 174160
rect 108226 174104 111004 174160
rect 108165 174102 111004 174104
rect 179649 174160 182948 174162
rect 179649 174104 179654 174160
rect 179710 174104 182948 174160
rect 179649 174102 182948 174104
rect 108165 174099 108231 174102
rect 179649 174099 179715 174102
rect 105405 173754 105471 173757
rect 102694 173752 105471 173754
rect 102694 173696 105410 173752
rect 105466 173696 105471 173752
rect 102694 173694 105471 173696
rect 102694 173208 102754 173694
rect 105405 173691 105471 173694
rect 176981 173210 177047 173213
rect 174852 173208 177047 173210
rect 174852 173152 176986 173208
rect 177042 173152 177047 173208
rect 174852 173150 177047 173152
rect 176981 173147 177047 173150
rect 207382 172876 207388 172940
rect 207452 172938 207458 172940
rect 207566 172938 207572 172940
rect 207452 172878 207572 172938
rect 207452 172876 207458 172878
rect 207566 172876 207572 172878
rect 207636 172876 207642 172940
rect 106325 172530 106391 172533
rect 102694 172528 106391 172530
rect 102694 172472 106330 172528
rect 106386 172472 106391 172528
rect 102694 172470 106391 172472
rect 102694 172120 102754 172470
rect 106325 172467 106391 172470
rect 177533 172122 177599 172125
rect 174852 172120 177599 172122
rect 174852 172064 177538 172120
rect 177594 172064 177599 172120
rect 174852 172062 177599 172064
rect 177533 172059 177599 172062
rect 107889 171850 107955 171853
rect 179649 171850 179715 171853
rect 107889 171848 111004 171850
rect 107889 171792 107894 171848
rect 107950 171792 111004 171848
rect 107889 171790 111004 171792
rect 179649 171848 182948 171850
rect 179649 171792 179654 171848
rect 179710 171792 182948 171848
rect 179649 171790 182948 171792
rect 107889 171787 107955 171790
rect 179649 171787 179715 171790
rect 106417 171442 106483 171445
rect 102694 171440 106483 171442
rect 102694 171384 106422 171440
rect 106478 171384 106483 171440
rect 102694 171382 106483 171384
rect 9896 171034 10376 171064
rect 12117 171034 12183 171037
rect 9896 171032 12183 171034
rect 9896 170976 12122 171032
rect 12178 170976 12183 171032
rect 9896 170974 12183 170976
rect 9896 170944 10376 170974
rect 12117 170971 12183 170974
rect 102694 170896 102754 171382
rect 106417 171379 106483 171382
rect 177717 170898 177783 170901
rect 174852 170896 177783 170898
rect 174852 170840 177722 170896
rect 177778 170840 177783 170896
rect 174852 170838 177783 170840
rect 177717 170835 177783 170838
rect 106049 170218 106115 170221
rect 102694 170216 106115 170218
rect 102694 170160 106054 170216
rect 106110 170160 106115 170216
rect 102694 170158 106115 170160
rect 12209 170082 12275 170085
rect 12209 170080 14066 170082
rect 12209 170024 12214 170080
rect 12270 170024 14066 170080
rect 12209 170022 14066 170024
rect 12209 170019 12275 170022
rect 14006 169808 14066 170022
rect 102694 169672 102754 170158
rect 106049 170155 106115 170158
rect 177625 169674 177691 169677
rect 174852 169672 177691 169674
rect 174852 169616 177630 169672
rect 177686 169616 177691 169672
rect 174852 169614 177691 169616
rect 177625 169611 177691 169614
rect 107889 169402 107955 169405
rect 179649 169402 179715 169405
rect 107889 169400 111004 169402
rect 107889 169344 107894 169400
rect 107950 169344 111004 169400
rect 107889 169342 111004 169344
rect 179649 169400 182948 169402
rect 179649 169344 179654 169400
rect 179710 169344 182948 169400
rect 179649 169342 182948 169344
rect 107889 169339 107955 169342
rect 179649 169339 179715 169342
rect 223582 169269 223642 169780
rect 223533 169264 223642 169269
rect 223533 169208 223538 169264
rect 223594 169208 223642 169264
rect 223533 169206 223642 169208
rect 223533 169203 223599 169206
rect 105221 168858 105287 168861
rect 102694 168856 105287 168858
rect 102694 168800 105226 168856
rect 105282 168800 105287 168856
rect 102694 168798 105287 168800
rect 102694 168448 102754 168798
rect 105221 168795 105287 168798
rect 178085 168450 178151 168453
rect 174852 168448 178151 168450
rect 174852 168392 178090 168448
rect 178146 168392 178151 168448
rect 174852 168390 178151 168392
rect 178085 168387 178151 168390
rect 105957 167498 106023 167501
rect 102694 167496 106023 167498
rect 102694 167440 105962 167496
rect 106018 167440 106023 167496
rect 102694 167438 106023 167440
rect 102694 167224 102754 167438
rect 105957 167435 106023 167438
rect 177533 167226 177599 167229
rect 174852 167224 177599 167226
rect 174852 167168 177538 167224
rect 177594 167168 177599 167224
rect 174852 167166 177599 167168
rect 177533 167163 177599 167166
rect 107797 167090 107863 167093
rect 179557 167090 179623 167093
rect 107797 167088 111004 167090
rect 107797 167032 107802 167088
rect 107858 167032 111004 167088
rect 107797 167030 111004 167032
rect 179557 167088 182948 167090
rect 179557 167032 179562 167088
rect 179618 167032 182948 167088
rect 179557 167030 182948 167032
rect 107797 167027 107863 167030
rect 179557 167027 179623 167030
rect 106417 166138 106483 166141
rect 103062 166136 106483 166138
rect 103062 166080 106422 166136
rect 106478 166080 106483 166136
rect 103062 166078 106483 166080
rect 103062 166030 103122 166078
rect 106417 166075 106483 166078
rect 102724 165970 103122 166030
rect 177533 166002 177599 166005
rect 174852 166000 177599 166002
rect 174852 165944 177538 166000
rect 177594 165944 177599 166000
rect 174852 165942 177599 165944
rect 177533 165939 177599 165942
rect 32633 164914 32699 164917
rect 29860 164912 32699 164914
rect 29860 164856 32638 164912
rect 32694 164856 32699 164912
rect 29860 164854 32699 164856
rect 32633 164851 32699 164854
rect 37417 164914 37483 164917
rect 59589 164914 59655 164917
rect 200993 164914 201059 164917
rect 37417 164912 39060 164914
rect 37417 164856 37422 164912
rect 37478 164856 39060 164912
rect 37417 164854 39060 164856
rect 59589 164912 62980 164914
rect 59589 164856 59594 164912
rect 59650 164856 62980 164912
rect 59589 164854 62980 164856
rect 126828 164854 134924 164914
rect 198772 164912 201059 164914
rect 198772 164856 200998 164912
rect 201054 164856 201059 164912
rect 198772 164854 201059 164856
rect 37417 164851 37483 164854
rect 59589 164851 59655 164854
rect 200993 164851 201059 164854
rect 204489 164914 204555 164917
rect 204489 164912 207972 164914
rect 204489 164856 204494 164912
rect 204550 164856 207972 164912
rect 204489 164854 207972 164856
rect 204489 164851 204555 164854
rect 102694 164234 102754 164720
rect 110974 164234 111034 164748
rect 174852 164718 182948 164778
rect 102694 164174 111034 164234
rect 106417 163554 106483 163557
rect 177717 163554 177783 163557
rect 102724 163552 106483 163554
rect 102724 163496 106422 163552
rect 106478 163496 106483 163552
rect 102724 163494 106483 163496
rect 174852 163552 177783 163554
rect 174852 163496 177722 163552
rect 177778 163496 177783 163552
rect 174852 163494 177783 163496
rect 106417 163491 106483 163494
rect 177717 163491 177783 163494
rect 224453 163554 224519 163557
rect 227416 163554 227896 163584
rect 224453 163552 227896 163554
rect 224453 163496 224458 163552
rect 224514 163496 227896 163552
rect 224453 163494 227896 163496
rect 224453 163491 224519 163494
rect 227416 163464 227896 163494
rect 207433 163282 207499 163285
rect 207566 163282 207572 163284
rect 207433 163280 207572 163282
rect 207433 163224 207438 163280
rect 207494 163224 207572 163280
rect 207433 163222 207572 163224
rect 207433 163219 207499 163222
rect 207566 163220 207572 163222
rect 207636 163220 207642 163284
rect 107797 162466 107863 162469
rect 179557 162466 179623 162469
rect 107797 162464 111004 162466
rect 107797 162408 107802 162464
rect 107858 162408 111004 162464
rect 107797 162406 111004 162408
rect 179557 162464 182948 162466
rect 179557 162408 179562 162464
rect 179618 162408 182948 162464
rect 179557 162406 182948 162408
rect 107797 162403 107863 162406
rect 179557 162403 179623 162406
rect 176981 162330 177047 162333
rect 174852 162328 177047 162330
rect 102724 162242 103122 162302
rect 174852 162272 176986 162328
rect 177042 162272 177047 162328
rect 174852 162270 177047 162272
rect 176981 162267 177047 162270
rect 103062 162194 103122 162242
rect 106141 162194 106207 162197
rect 103062 162192 106207 162194
rect 103062 162136 106146 162192
rect 106202 162136 106207 162192
rect 103062 162134 106207 162136
rect 106141 162131 106207 162134
rect 176981 161106 177047 161109
rect 174852 161104 177047 161106
rect 174852 161048 176986 161104
rect 177042 161048 177047 161104
rect 102694 160698 102754 161048
rect 174852 161046 177047 161048
rect 176981 161043 177047 161046
rect 105773 160698 105839 160701
rect 102694 160696 105839 160698
rect 102694 160640 105778 160696
rect 105834 160640 105839 160696
rect 102694 160638 105839 160640
rect 105773 160635 105839 160638
rect 108533 160018 108599 160021
rect 179649 160018 179715 160021
rect 108533 160016 111004 160018
rect 108533 159960 108538 160016
rect 108594 159960 111004 160016
rect 108533 159958 111004 159960
rect 179649 160016 182948 160018
rect 179649 159960 179654 160016
rect 179710 159960 182948 160016
rect 179649 159958 182948 159960
rect 108533 159955 108599 159958
rect 179649 159955 179715 159958
rect 177533 159882 177599 159885
rect 174852 159880 177599 159882
rect 174852 159824 177538 159880
rect 177594 159824 177599 159880
rect 12209 159338 12275 159341
rect 14006 159338 14066 159688
rect 12209 159336 14066 159338
rect 12209 159280 12214 159336
rect 12270 159280 14066 159336
rect 12209 159278 14066 159280
rect 102694 159338 102754 159824
rect 174852 159822 177599 159824
rect 177533 159819 177599 159822
rect 106417 159338 106483 159341
rect 102694 159336 106483 159338
rect 102694 159280 106422 159336
rect 106478 159280 106483 159336
rect 102694 159278 106483 159280
rect 12209 159275 12275 159278
rect 106417 159275 106483 159278
rect 223582 159205 223642 159716
rect 223533 159200 223642 159205
rect 223533 159144 223538 159200
rect 223594 159144 223642 159200
rect 223533 159142 223642 159144
rect 223533 159139 223599 159142
rect 177349 158794 177415 158797
rect 174852 158792 177415 158794
rect 174852 158736 177354 158792
rect 177410 158736 177415 158792
rect 102694 158386 102754 158736
rect 174852 158734 177415 158736
rect 177349 158731 177415 158734
rect 105405 158386 105471 158389
rect 102694 158384 105471 158386
rect 102694 158328 105410 158384
rect 105466 158328 105471 158384
rect 102694 158326 105471 158328
rect 105405 158323 105471 158326
rect 107797 157706 107863 157709
rect 179557 157706 179623 157709
rect 107797 157704 111004 157706
rect 107797 157648 107802 157704
rect 107858 157648 111004 157704
rect 107797 157646 111004 157648
rect 179557 157704 182948 157706
rect 179557 157648 179562 157704
rect 179618 157648 182948 157704
rect 179557 157646 182948 157648
rect 107797 157643 107863 157646
rect 179557 157643 179623 157646
rect 177533 157570 177599 157573
rect 174852 157568 177599 157570
rect 174852 157512 177538 157568
rect 177594 157512 177599 157568
rect 102694 157026 102754 157512
rect 174852 157510 177599 157512
rect 177533 157507 177599 157510
rect 105405 157026 105471 157029
rect 102694 157024 105471 157026
rect 102694 156968 105410 157024
rect 105466 156968 105471 157024
rect 102694 156966 105471 156968
rect 105405 156963 105471 156966
rect 177533 156346 177599 156349
rect 174852 156344 177599 156346
rect 174852 156288 177538 156344
rect 177594 156288 177599 156344
rect 102694 155802 102754 156288
rect 174852 156286 177599 156288
rect 177533 156283 177599 156286
rect 105221 155802 105287 155805
rect 102694 155800 105287 155802
rect 102694 155744 105226 155800
rect 105282 155744 105287 155800
rect 102694 155742 105287 155744
rect 105221 155739 105287 155742
rect 107705 155394 107771 155397
rect 179465 155394 179531 155397
rect 107705 155392 111004 155394
rect 107705 155336 107710 155392
rect 107766 155336 111004 155392
rect 107705 155334 111004 155336
rect 179465 155392 182948 155394
rect 179465 155336 179470 155392
rect 179526 155336 182948 155392
rect 179465 155334 182948 155336
rect 107705 155331 107771 155334
rect 179465 155331 179531 155334
rect 177349 155122 177415 155125
rect 174852 155120 177415 155122
rect 174852 155064 177354 155120
rect 177410 155064 177415 155120
rect 57473 154850 57539 154853
rect 54884 154848 57539 154850
rect 54884 154792 57478 154848
rect 57534 154792 57539 154848
rect 54884 154790 57539 154792
rect 57473 154787 57539 154790
rect 102694 154578 102754 155064
rect 174852 155062 177415 155064
rect 177349 155059 177415 155062
rect 105773 154578 105839 154581
rect 102694 154576 105839 154578
rect 102694 154520 105778 154576
rect 105834 154520 105839 154576
rect 102694 154518 105839 154520
rect 105773 154515 105839 154518
rect 105589 153898 105655 153901
rect 178177 153898 178243 153901
rect 102724 153896 105655 153898
rect 102724 153840 105594 153896
rect 105650 153840 105655 153896
rect 102724 153838 105655 153840
rect 174852 153896 178243 153898
rect 174852 153840 178182 153896
rect 178238 153840 178243 153896
rect 174852 153838 178243 153840
rect 105589 153835 105655 153838
rect 178177 153835 178243 153838
rect 207433 153764 207499 153765
rect 207382 153762 207388 153764
rect 207342 153702 207388 153762
rect 207452 153760 207499 153764
rect 207494 153704 207499 153760
rect 207382 153700 207388 153702
rect 207452 153700 207499 153704
rect 207433 153699 207499 153700
rect 107889 152946 107955 152949
rect 179649 152946 179715 152949
rect 107889 152944 111004 152946
rect 107889 152888 107894 152944
rect 107950 152888 111004 152944
rect 107889 152886 111004 152888
rect 179649 152944 182948 152946
rect 179649 152888 179654 152944
rect 179710 152888 182948 152944
rect 179649 152886 182948 152888
rect 107889 152883 107955 152886
rect 179649 152883 179715 152886
rect 178269 152674 178335 152677
rect 174852 152672 178335 152674
rect 102724 152586 103122 152646
rect 174852 152616 178274 152672
rect 178330 152616 178335 152672
rect 174852 152614 178335 152616
rect 178269 152611 178335 152614
rect 103062 152538 103122 152586
rect 106417 152538 106483 152541
rect 103062 152536 106483 152538
rect 103062 152480 106422 152536
rect 106478 152480 106483 152536
rect 103062 152478 106483 152480
rect 106417 152475 106483 152478
rect 207433 152268 207499 152269
rect 207382 152266 207388 152268
rect 207342 152206 207388 152266
rect 207452 152264 207499 152268
rect 207494 152208 207499 152264
rect 207382 152204 207388 152206
rect 207452 152204 207499 152208
rect 207433 152203 207499 152204
rect 31989 151586 32055 151589
rect 29860 151584 32055 151586
rect 29860 151528 31994 151584
rect 32050 151528 32055 151584
rect 29860 151526 32055 151528
rect 31989 151523 32055 151526
rect 37918 151524 37924 151588
rect 37988 151586 37994 151588
rect 59589 151586 59655 151589
rect 132361 151586 132427 151589
rect 200533 151586 200599 151589
rect 37988 151526 39060 151586
rect 59589 151584 62980 151586
rect 59589 151528 59594 151584
rect 59650 151528 62980 151584
rect 59589 151526 62980 151528
rect 126828 151584 134924 151586
rect 126828 151528 132366 151584
rect 132422 151528 134924 151584
rect 126828 151526 134924 151528
rect 198772 151584 200599 151586
rect 198772 151528 200538 151584
rect 200594 151528 200599 151584
rect 198772 151526 200599 151528
rect 37988 151524 37994 151526
rect 59589 151523 59655 151526
rect 132361 151523 132427 151526
rect 200533 151523 200599 151526
rect 204489 151586 204555 151589
rect 204489 151584 207972 151586
rect 204489 151528 204494 151584
rect 204550 151528 207972 151584
rect 204489 151526 207972 151528
rect 204489 151523 204555 151526
rect 178361 151450 178427 151453
rect 174852 151448 178427 151450
rect 174852 151392 178366 151448
rect 178422 151392 178427 151448
rect 102694 151042 102754 151392
rect 174852 151390 178427 151392
rect 178361 151387 178427 151390
rect 106601 151042 106667 151045
rect 102694 151040 106667 151042
rect 102694 150984 106606 151040
rect 106662 150984 106667 151040
rect 102694 150982 106667 150984
rect 106601 150979 106667 150982
rect 107245 150634 107311 150637
rect 180477 150634 180543 150637
rect 107245 150632 111004 150634
rect 107245 150576 107250 150632
rect 107306 150576 111004 150632
rect 107245 150574 111004 150576
rect 180477 150632 182948 150634
rect 180477 150576 180482 150632
rect 180538 150576 182948 150632
rect 180477 150574 182948 150576
rect 107245 150571 107311 150574
rect 180477 150571 180543 150574
rect 178453 150226 178519 150229
rect 174852 150224 178519 150226
rect 174852 150168 178458 150224
rect 178514 150168 178519 150224
rect 12025 149818 12091 149821
rect 12025 149816 14036 149818
rect 12025 149760 12030 149816
rect 12086 149760 14036 149816
rect 12025 149758 14036 149760
rect 12025 149755 12091 149758
rect 102694 149682 102754 150168
rect 174852 150166 178519 150168
rect 178453 150163 178519 150166
rect 105957 149682 106023 149685
rect 102694 149680 106023 149682
rect 102694 149624 105962 149680
rect 106018 149624 106023 149680
rect 102694 149622 106023 149624
rect 105957 149619 106023 149622
rect 223582 149549 223642 149788
rect 223533 149544 223642 149549
rect 223533 149488 223538 149544
rect 223594 149488 223642 149544
rect 223533 149486 223642 149488
rect 223533 149483 223599 149486
rect 9896 149410 10376 149440
rect 12577 149410 12643 149413
rect 9896 149408 12643 149410
rect 9896 149352 12582 149408
rect 12638 149352 12643 149408
rect 9896 149350 12643 149352
rect 9896 149320 10376 149350
rect 12577 149347 12643 149350
rect 177717 149002 177783 149005
rect 174852 149000 177783 149002
rect 174852 148944 177722 149000
rect 177778 148944 177783 149000
rect 102694 148458 102754 148944
rect 174852 148942 177783 148944
rect 177717 148939 177783 148942
rect 105405 148458 105471 148461
rect 102694 148456 105471 148458
rect 102694 148400 105410 148456
rect 105466 148400 105471 148456
rect 102694 148398 105471 148400
rect 105405 148395 105471 148398
rect 107153 148322 107219 148325
rect 180385 148322 180451 148325
rect 107153 148320 111004 148322
rect 107153 148264 107158 148320
rect 107214 148264 111004 148320
rect 107153 148262 111004 148264
rect 180385 148320 182948 148322
rect 180385 148264 180390 148320
rect 180446 148264 182948 148320
rect 180385 148262 182948 148264
rect 107153 148259 107219 148262
rect 180385 148259 180451 148262
rect 177165 147778 177231 147781
rect 174852 147776 177231 147778
rect 174852 147720 177170 147776
rect 177226 147720 177231 147776
rect 102694 147234 102754 147720
rect 174852 147718 177231 147720
rect 177165 147715 177231 147718
rect 105221 147234 105287 147237
rect 102694 147232 105287 147234
rect 102694 147176 105226 147232
rect 105282 147176 105287 147232
rect 102694 147174 105287 147176
rect 105221 147171 105287 147174
rect 178177 146554 178243 146557
rect 174852 146552 178243 146554
rect 174852 146496 178182 146552
rect 178238 146496 178243 146552
rect 102694 146010 102754 146496
rect 174852 146494 178243 146496
rect 178177 146491 178243 146494
rect 105865 146010 105931 146013
rect 102694 146008 105931 146010
rect 102694 145952 105870 146008
rect 105926 145952 105931 146008
rect 102694 145950 105931 145952
rect 105865 145947 105931 145950
rect 108533 146010 108599 146013
rect 180293 146010 180359 146013
rect 108533 146008 111004 146010
rect 108533 145952 108538 146008
rect 108594 145952 111004 146008
rect 108533 145950 111004 145952
rect 180293 146008 182948 146010
rect 180293 145952 180298 146008
rect 180354 145952 182948 146008
rect 180293 145950 182948 145952
rect 108533 145947 108599 145950
rect 180293 145947 180359 145950
rect 177441 145466 177507 145469
rect 174852 145464 177507 145466
rect 174852 145408 177446 145464
rect 177502 145408 177507 145464
rect 102694 144922 102754 145408
rect 174852 145406 177507 145408
rect 177441 145403 177507 145406
rect 106417 144922 106483 144925
rect 102694 144920 106483 144922
rect 102694 144864 106422 144920
rect 106478 144864 106483 144920
rect 102694 144862 106483 144864
rect 106417 144859 106483 144862
rect 207433 142746 207499 142749
rect 207750 142746 207756 142748
rect 207433 142744 207756 142746
rect 207433 142688 207438 142744
rect 207494 142688 207756 142744
rect 207433 142686 207756 142688
rect 207433 142683 207499 142686
rect 207750 142684 207756 142686
rect 207820 142684 207826 142748
rect 12577 142610 12643 142613
rect 101030 142610 101036 142612
rect 12577 142608 101036 142610
rect 12577 142552 12582 142608
rect 12638 142552 101036 142608
rect 12577 142550 101036 142552
rect 12577 142547 12643 142550
rect 101030 142548 101036 142550
rect 101100 142610 101106 142612
rect 102277 142610 102343 142613
rect 101100 142608 102343 142610
rect 101100 142552 102282 142608
rect 102338 142552 102343 142608
rect 101100 142550 102343 142552
rect 101100 142548 101106 142550
rect 102277 142547 102343 142550
rect 163273 142610 163339 142613
rect 167270 142610 167276 142612
rect 163273 142608 167276 142610
rect 163273 142552 163278 142608
rect 163334 142552 167276 142608
rect 163273 142550 167276 142552
rect 163273 142547 163339 142550
rect 167270 142548 167276 142550
rect 167340 142548 167346 142612
rect 207750 142548 207756 142612
rect 207820 142610 207826 142612
rect 207893 142610 207959 142613
rect 207820 142608 207959 142610
rect 207820 142552 207898 142608
rect 207954 142552 207959 142608
rect 207820 142550 207959 142552
rect 207820 142548 207826 142550
rect 207893 142547 207959 142550
rect 174589 142202 174655 142205
rect 174589 142200 177090 142202
rect 174589 142144 174594 142200
rect 174650 142144 177090 142200
rect 174589 142142 177090 142144
rect 174589 142139 174655 142142
rect 62809 142066 62875 142069
rect 134477 142066 134543 142069
rect 60742 142064 62875 142066
rect 60742 142008 62814 142064
rect 62870 142008 62875 142064
rect 60742 142006 62875 142008
rect 60742 141560 60802 142006
rect 62809 142003 62875 142006
rect 132686 142064 134543 142066
rect 132686 142008 134482 142064
rect 134538 142008 134543 142064
rect 132686 142006 134543 142008
rect 71038 141868 71044 141932
rect 71108 141930 71114 141932
rect 90133 141930 90199 141933
rect 71108 141928 90199 141930
rect 71108 141872 90138 141928
rect 90194 141872 90199 141928
rect 71108 141870 90199 141872
rect 71108 141868 71114 141870
rect 90133 141867 90199 141870
rect 132686 141560 132746 142006
rect 134477 142003 134543 142006
rect 146294 141868 146300 141932
rect 146364 141930 146370 141932
rect 162169 141930 162235 141933
rect 146364 141928 162235 141930
rect 146364 141872 162174 141928
rect 162230 141872 162235 141928
rect 146364 141870 162235 141872
rect 146364 141868 146370 141870
rect 162169 141867 162235 141870
rect 177030 141560 177090 142142
rect 103473 141522 103539 141525
rect 103473 141520 104932 141522
rect 103473 141464 103478 141520
rect 103534 141464 104932 141520
rect 103473 141462 104932 141464
rect 103473 141459 103539 141462
rect 31805 141388 31871 141389
rect 31805 141384 31852 141388
rect 31916 141386 31922 141388
rect 91237 141386 91303 141389
rect 94222 141386 94228 141388
rect 31805 141328 31810 141384
rect 31805 141324 31852 141328
rect 31916 141326 31962 141386
rect 91237 141384 94228 141386
rect 91237 141328 91242 141384
rect 91298 141328 94228 141384
rect 91237 141326 94228 141328
rect 31916 141324 31922 141326
rect 31805 141323 31871 141324
rect 91237 141323 91303 141326
rect 94222 141324 94228 141326
rect 94292 141324 94298 141388
rect 62809 140978 62875 140981
rect 60772 140976 62875 140978
rect 60772 140920 62814 140976
rect 62870 140920 62875 140976
rect 60772 140918 62875 140920
rect 62809 140915 62875 140918
rect 102277 140978 102343 140981
rect 135305 140978 135371 140981
rect 102277 140976 104932 140978
rect 102277 140920 102282 140976
rect 102338 140920 104932 140976
rect 102277 140918 104932 140920
rect 132716 140976 135371 140978
rect 132716 140920 135310 140976
rect 135366 140920 135371 140976
rect 132716 140918 135371 140920
rect 102277 140915 102343 140918
rect 135305 140915 135371 140918
rect 174405 140978 174471 140981
rect 174405 140976 177060 140978
rect 174405 140920 174410 140976
rect 174466 140920 177060 140976
rect 174405 140918 177060 140920
rect 174405 140915 174471 140918
rect 62717 140706 62783 140709
rect 60742 140704 62783 140706
rect 60742 140648 62722 140704
rect 62778 140648 62783 140704
rect 60742 140646 62783 140648
rect 60742 140472 60802 140646
rect 62717 140643 62783 140646
rect 102369 140434 102435 140437
rect 135305 140434 135371 140437
rect 102369 140432 104932 140434
rect 102369 140376 102374 140432
rect 102430 140376 104932 140432
rect 102369 140374 104932 140376
rect 132716 140432 135371 140434
rect 132716 140376 135310 140432
rect 135366 140376 135371 140432
rect 132716 140374 135371 140376
rect 102369 140371 102435 140374
rect 135305 140371 135371 140374
rect 174221 140434 174287 140437
rect 174221 140432 177060 140434
rect 174221 140376 174226 140432
rect 174282 140376 177060 140432
rect 174221 140374 177060 140376
rect 174221 140371 174287 140374
rect 62809 139754 62875 139757
rect 60772 139752 62875 139754
rect 60772 139696 62814 139752
rect 62870 139696 62875 139752
rect 60772 139694 62875 139696
rect 62809 139691 62875 139694
rect 102369 139754 102435 139757
rect 135305 139754 135371 139757
rect 102369 139752 104932 139754
rect 102369 139696 102374 139752
rect 102430 139696 104932 139752
rect 102369 139694 104932 139696
rect 132716 139752 135371 139754
rect 132716 139696 135310 139752
rect 135366 139696 135371 139752
rect 132716 139694 135371 139696
rect 102369 139691 102435 139694
rect 135305 139691 135371 139694
rect 174313 139754 174379 139757
rect 222889 139754 222955 139757
rect 227416 139754 227896 139784
rect 174313 139752 177060 139754
rect 174313 139696 174318 139752
rect 174374 139696 177060 139752
rect 174313 139694 177060 139696
rect 222889 139752 227896 139754
rect 222889 139696 222894 139752
rect 222950 139696 227896 139752
rect 222889 139694 227896 139696
rect 174313 139691 174379 139694
rect 222889 139691 222955 139694
rect 227416 139664 227896 139694
rect 62349 139482 62415 139485
rect 60742 139480 62415 139482
rect 60742 139424 62354 139480
rect 62410 139424 62415 139480
rect 60742 139422 62415 139424
rect 60742 139248 60802 139422
rect 62349 139419 62415 139422
rect 66213 139482 66279 139485
rect 66213 139480 67948 139482
rect 66213 139424 66218 139480
rect 66274 139424 67948 139480
rect 66213 139422 67948 139424
rect 66213 139419 66279 139422
rect 97726 139074 97786 139384
rect 102461 139210 102527 139213
rect 135305 139210 135371 139213
rect 102461 139208 104932 139210
rect 102461 139152 102466 139208
rect 102522 139152 104932 139208
rect 102461 139150 104932 139152
rect 132716 139208 135371 139210
rect 132716 139152 135310 139208
rect 135366 139152 135371 139208
rect 132716 139150 135371 139152
rect 102461 139147 102527 139150
rect 135305 139147 135371 139150
rect 100621 139074 100687 139077
rect 97726 139072 100687 139074
rect 97726 139016 100626 139072
rect 100682 139016 100687 139072
rect 97726 139014 100687 139016
rect 100621 139011 100687 139014
rect 136961 139074 137027 139077
rect 140046 139074 140106 139384
rect 136961 139072 140106 139074
rect 136961 139016 136966 139072
rect 137022 139016 140106 139072
rect 136961 139014 140106 139016
rect 169854 139074 169914 139452
rect 174129 139210 174195 139213
rect 174129 139208 177060 139210
rect 174129 139152 174134 139208
rect 174190 139152 177060 139208
rect 174129 139150 177060 139152
rect 174129 139147 174195 139150
rect 172565 139074 172631 139077
rect 169854 139072 172631 139074
rect 169854 139016 172570 139072
rect 172626 139016 172631 139072
rect 169854 139014 172631 139016
rect 136961 139011 137027 139014
rect 172565 139011 172631 139014
rect 62809 138938 62875 138941
rect 60742 138936 62875 138938
rect 60742 138880 62814 138936
rect 62870 138880 62875 138936
rect 60742 138878 62875 138880
rect 60742 138704 60802 138878
rect 62809 138875 62875 138878
rect 66397 138938 66463 138941
rect 135121 138938 135187 138941
rect 66397 138936 67948 138938
rect 66397 138880 66402 138936
rect 66458 138880 67948 138936
rect 66397 138878 67948 138880
rect 132686 138936 135187 138938
rect 132686 138880 135126 138936
rect 135182 138880 135187 138936
rect 132686 138878 135187 138880
rect 66397 138875 66463 138878
rect 97726 138666 97786 138840
rect 132686 138704 132746 138878
rect 135121 138875 135187 138878
rect 136869 138938 136935 138941
rect 136869 138936 140076 138938
rect 136869 138880 136874 138936
rect 136930 138880 140076 138936
rect 136869 138878 140076 138880
rect 136869 138875 136935 138878
rect 100529 138666 100595 138669
rect 97726 138664 100595 138666
rect 97726 138608 100534 138664
rect 100590 138608 100595 138664
rect 97726 138606 100595 138608
rect 100529 138603 100595 138606
rect 102553 138666 102619 138669
rect 169854 138666 169914 138908
rect 172197 138666 172263 138669
rect 102553 138664 104932 138666
rect 102553 138608 102558 138664
rect 102614 138608 104932 138664
rect 102553 138606 104932 138608
rect 169854 138664 172263 138666
rect 169854 138608 172202 138664
rect 172258 138608 172263 138664
rect 169854 138606 172263 138608
rect 102553 138603 102619 138606
rect 172197 138603 172263 138606
rect 174221 138666 174287 138669
rect 174221 138664 177060 138666
rect 174221 138608 174226 138664
rect 174282 138608 177060 138664
rect 174221 138606 177060 138608
rect 174221 138603 174287 138606
rect 63453 138394 63519 138397
rect 134569 138394 134635 138397
rect 60742 138392 63519 138394
rect 60742 138336 63458 138392
rect 63514 138336 63519 138392
rect 60742 138334 63519 138336
rect 60742 138024 60802 138334
rect 63453 138331 63519 138334
rect 132686 138392 134635 138394
rect 132686 138336 134574 138392
rect 134630 138336 134635 138392
rect 132686 138334 134635 138336
rect 66305 138258 66371 138261
rect 66305 138256 67948 138258
rect 66305 138200 66310 138256
rect 66366 138200 67948 138256
rect 66305 138198 67948 138200
rect 66305 138195 66371 138198
rect 97726 137850 97786 138160
rect 132686 138024 132746 138334
rect 134569 138331 134635 138334
rect 102369 137986 102435 137989
rect 102369 137984 104932 137986
rect 102369 137928 102374 137984
rect 102430 137928 104932 137984
rect 102369 137926 104932 137928
rect 102369 137923 102435 137926
rect 100069 137850 100135 137853
rect 97726 137848 100135 137850
rect 97726 137792 100074 137848
rect 100130 137792 100135 137848
rect 97726 137790 100135 137792
rect 100069 137787 100135 137790
rect 136869 137850 136935 137853
rect 140046 137850 140106 138160
rect 136869 137848 140106 137850
rect 136869 137792 136874 137848
rect 136930 137792 140106 137848
rect 136869 137790 140106 137792
rect 169854 137850 169914 138228
rect 174129 137986 174195 137989
rect 174129 137984 177060 137986
rect 174129 137928 174134 137984
rect 174190 137928 177060 137984
rect 174129 137926 177060 137928
rect 174129 137923 174195 137926
rect 172657 137850 172723 137853
rect 169854 137848 172723 137850
rect 169854 137792 172662 137848
rect 172718 137792 172723 137848
rect 169854 137790 172723 137792
rect 136869 137787 136935 137790
rect 172657 137787 172723 137790
rect 62533 137714 62599 137717
rect 60742 137712 62599 137714
rect 60742 137656 62538 137712
rect 62594 137656 62599 137712
rect 60742 137654 62599 137656
rect 60742 137480 60802 137654
rect 62533 137651 62599 137654
rect 66397 137714 66463 137717
rect 135213 137714 135279 137717
rect 66397 137712 67948 137714
rect 66397 137656 66402 137712
rect 66458 137656 67948 137712
rect 66397 137654 67948 137656
rect 132686 137712 135279 137714
rect 132686 137656 135218 137712
rect 135274 137656 135279 137712
rect 132686 137654 135279 137656
rect 66397 137651 66463 137654
rect 97726 137306 97786 137616
rect 132686 137480 132746 137654
rect 135213 137651 135279 137654
rect 102461 137442 102527 137445
rect 102461 137440 104932 137442
rect 102461 137384 102466 137440
rect 102522 137384 104932 137440
rect 102461 137382 104932 137384
rect 102461 137379 102527 137382
rect 99701 137306 99767 137309
rect 97726 137304 99767 137306
rect 97726 137248 99706 137304
rect 99762 137248 99767 137304
rect 97726 137246 99767 137248
rect 99701 137243 99767 137246
rect 136869 137306 136935 137309
rect 140046 137306 140106 137616
rect 136869 137304 140106 137306
rect 136869 137248 136874 137304
rect 136930 137248 140106 137304
rect 136869 137246 140106 137248
rect 169854 137306 169914 137684
rect 174221 137442 174287 137445
rect 174221 137440 177060 137442
rect 174221 137384 174226 137440
rect 174282 137384 177060 137440
rect 174221 137382 177060 137384
rect 174221 137379 174287 137382
rect 172657 137306 172723 137309
rect 169854 137304 172723 137306
rect 169854 137248 172662 137304
rect 172718 137248 172723 137304
rect 169854 137246 172723 137248
rect 136869 137243 136935 137246
rect 172657 137243 172723 137246
rect 30517 137170 30583 137173
rect 62809 137170 62875 137173
rect 30517 137168 32988 137170
rect 30517 137112 30522 137168
rect 30578 137112 32988 137168
rect 30517 137110 32988 137112
rect 60742 137168 62875 137170
rect 60742 137112 62814 137168
rect 62870 137112 62875 137168
rect 60742 137110 62875 137112
rect 30517 137107 30583 137110
rect 60742 136936 60802 137110
rect 62809 137107 62875 137110
rect 65017 136762 65083 136765
rect 67918 136762 67978 137140
rect 65017 136760 67978 136762
rect 65017 136704 65022 136760
rect 65078 136704 67978 136760
rect 65017 136702 67978 136704
rect 65017 136699 65083 136702
rect 62901 136626 62967 136629
rect 60742 136624 62967 136626
rect 60742 136568 62906 136624
rect 62962 136568 62967 136624
rect 60742 136566 62967 136568
rect 97726 136626 97786 137072
rect 102369 136898 102435 136901
rect 135397 136898 135463 136901
rect 102369 136896 104932 136898
rect 102369 136840 102374 136896
rect 102430 136840 104932 136896
rect 102369 136838 104932 136840
rect 132716 136896 135463 136898
rect 132716 136840 135402 136896
rect 135458 136840 135463 136896
rect 132716 136838 135463 136840
rect 102369 136835 102435 136838
rect 135397 136835 135463 136838
rect 100621 136626 100687 136629
rect 135305 136626 135371 136629
rect 97726 136624 100687 136626
rect 97726 136568 100626 136624
rect 100682 136568 100687 136624
rect 97726 136566 100687 136568
rect 60742 136392 60802 136566
rect 62901 136563 62967 136566
rect 100621 136563 100687 136566
rect 132686 136624 135371 136626
rect 132686 136568 135310 136624
rect 135366 136568 135371 136624
rect 132686 136566 135371 136568
rect 66397 136490 66463 136493
rect 66397 136488 67948 136490
rect 66397 136432 66402 136488
rect 66458 136432 67948 136488
rect 66397 136430 67948 136432
rect 66397 136427 66463 136430
rect 132686 136392 132746 136566
rect 135305 136563 135371 136566
rect 136777 136626 136843 136629
rect 140046 136626 140106 137072
rect 136777 136624 140106 136626
rect 136777 136568 136782 136624
rect 136838 136568 140106 136624
rect 136777 136566 140106 136568
rect 169854 136626 169914 137140
rect 174129 136898 174195 136901
rect 174129 136896 177060 136898
rect 174129 136840 174134 136896
rect 174190 136840 177060 136896
rect 174129 136838 177060 136840
rect 174129 136835 174195 136838
rect 204814 136629 204874 137140
rect 172565 136626 172631 136629
rect 169854 136624 172631 136626
rect 169854 136568 172570 136624
rect 172626 136568 172631 136624
rect 169854 136566 172631 136568
rect 136777 136563 136843 136566
rect 172565 136563 172631 136566
rect 204765 136624 204874 136629
rect 204765 136568 204770 136624
rect 204826 136568 204874 136624
rect 204765 136566 204874 136568
rect 204765 136563 204831 136566
rect 97726 136082 97786 136392
rect 102645 136354 102711 136357
rect 102645 136352 104932 136354
rect 102645 136296 102650 136352
rect 102706 136296 104932 136352
rect 102645 136294 104932 136296
rect 102645 136291 102711 136294
rect 100897 136082 100963 136085
rect 97726 136080 100963 136082
rect 97726 136024 100902 136080
rect 100958 136024 100963 136080
rect 97726 136022 100963 136024
rect 100897 136019 100963 136022
rect 136869 136082 136935 136085
rect 140046 136082 140106 136392
rect 169854 136218 169914 136460
rect 174221 136354 174287 136357
rect 174221 136352 177060 136354
rect 174221 136296 174226 136352
rect 174282 136296 177060 136352
rect 174221 136294 177060 136296
rect 174221 136291 174287 136294
rect 169854 136158 170282 136218
rect 170222 136082 170282 136158
rect 172657 136082 172723 136085
rect 136869 136080 140106 136082
rect 136869 136024 136874 136080
rect 136930 136024 140106 136080
rect 136869 136022 140106 136024
rect 169670 136022 170098 136082
rect 170222 136080 172723 136082
rect 170222 136024 172662 136080
rect 172718 136024 172723 136080
rect 170222 136022 172723 136024
rect 136869 136019 136935 136022
rect 65661 135946 65727 135949
rect 100897 135946 100963 135949
rect 65661 135944 67948 135946
rect 65661 135888 65666 135944
rect 65722 135888 67948 135944
rect 65661 135886 67948 135888
rect 97756 135944 100963 135946
rect 97756 135888 100902 135944
rect 100958 135888 100963 135944
rect 97756 135886 100963 135888
rect 65661 135883 65727 135886
rect 100897 135883 100963 135886
rect 136961 135946 137027 135949
rect 136961 135944 140076 135946
rect 136961 135888 136966 135944
rect 137022 135888 140076 135944
rect 169670 135916 169730 136022
rect 170038 135946 170098 136022
rect 172657 136019 172723 136022
rect 172657 135946 172723 135949
rect 170038 135944 172723 135946
rect 136961 135886 140076 135888
rect 170038 135888 172662 135944
rect 172718 135888 172723 135944
rect 170038 135886 172723 135888
rect 136961 135883 137027 135886
rect 172657 135883 172723 135886
rect 62717 135674 62783 135677
rect 60772 135672 62783 135674
rect 60772 135616 62722 135672
rect 62778 135616 62783 135672
rect 60772 135614 62783 135616
rect 62717 135611 62783 135614
rect 102277 135674 102343 135677
rect 135213 135674 135279 135677
rect 102277 135672 104932 135674
rect 102277 135616 102282 135672
rect 102338 135616 104932 135672
rect 102277 135614 104932 135616
rect 132716 135672 135279 135674
rect 132716 135616 135218 135672
rect 135274 135616 135279 135672
rect 132716 135614 135279 135616
rect 102277 135611 102343 135614
rect 135213 135611 135279 135614
rect 174129 135674 174195 135677
rect 174129 135672 177060 135674
rect 174129 135616 174134 135672
rect 174190 135616 177060 135672
rect 174129 135614 177060 135616
rect 174129 135611 174195 135614
rect 62625 135402 62691 135405
rect 135121 135402 135187 135405
rect 60742 135400 62691 135402
rect 60742 135344 62630 135400
rect 62686 135344 62691 135400
rect 60742 135342 62691 135344
rect 60742 135168 60802 135342
rect 62625 135339 62691 135342
rect 132686 135400 135187 135402
rect 132686 135344 135126 135400
rect 135182 135344 135187 135400
rect 132686 135342 135187 135344
rect 65845 135266 65911 135269
rect 65845 135264 67948 135266
rect 65845 135208 65850 135264
rect 65906 135208 67948 135264
rect 65845 135206 67948 135208
rect 65845 135203 65911 135206
rect 132686 135168 132746 135342
rect 135121 135339 135187 135342
rect 62809 134858 62875 134861
rect 60742 134856 62875 134858
rect 60742 134800 62814 134856
rect 62870 134800 62875 134856
rect 60742 134798 62875 134800
rect 97726 134858 97786 135168
rect 102185 135130 102251 135133
rect 102185 135128 104932 135130
rect 102185 135072 102190 135128
rect 102246 135072 104932 135128
rect 102185 135070 104932 135072
rect 102185 135067 102251 135070
rect 99885 134858 99951 134861
rect 135213 134858 135279 134861
rect 97726 134856 99951 134858
rect 97726 134800 99890 134856
rect 99946 134800 99951 134856
rect 97726 134798 99951 134800
rect 60742 134624 60802 134798
rect 62809 134795 62875 134798
rect 99885 134795 99951 134798
rect 132686 134856 135279 134858
rect 132686 134800 135218 134856
rect 135274 134800 135279 134856
rect 132686 134798 135279 134800
rect 66213 134722 66279 134725
rect 100897 134722 100963 134725
rect 66213 134720 67948 134722
rect 66213 134664 66218 134720
rect 66274 134664 67948 134720
rect 66213 134662 67948 134664
rect 97756 134720 100963 134722
rect 97756 134664 100902 134720
rect 100958 134664 100963 134720
rect 97756 134662 100963 134664
rect 66213 134659 66279 134662
rect 100897 134659 100963 134662
rect 132686 134624 132746 134798
rect 135213 134795 135279 134798
rect 136869 134858 136935 134861
rect 140046 134858 140106 135168
rect 136869 134856 140106 134858
rect 136869 134800 136874 134856
rect 136930 134800 140106 134856
rect 136869 134798 140106 134800
rect 169854 134858 169914 135236
rect 174037 135130 174103 135133
rect 174037 135128 177060 135130
rect 174037 135072 174042 135128
rect 174098 135072 177060 135128
rect 174037 135070 177060 135072
rect 174037 135067 174103 135070
rect 172657 134858 172723 134861
rect 169854 134856 172723 134858
rect 169854 134800 172662 134856
rect 172718 134800 172723 134856
rect 169854 134798 172723 134800
rect 136869 134795 136935 134798
rect 172657 134795 172723 134798
rect 136961 134722 137027 134725
rect 136961 134720 140076 134722
rect 136961 134664 136966 134720
rect 137022 134664 140076 134720
rect 136961 134662 140076 134664
rect 136961 134659 137027 134662
rect 102369 134586 102435 134589
rect 169854 134586 169914 134692
rect 172565 134586 172631 134589
rect 102369 134584 104932 134586
rect 102369 134528 102374 134584
rect 102430 134528 104932 134584
rect 102369 134526 104932 134528
rect 169854 134584 172631 134586
rect 169854 134528 172570 134584
rect 172626 134528 172631 134584
rect 169854 134526 172631 134528
rect 102369 134523 102435 134526
rect 172565 134523 172631 134526
rect 174221 134586 174287 134589
rect 174221 134584 177060 134586
rect 174221 134528 174226 134584
rect 174282 134528 177060 134584
rect 174221 134526 177060 134528
rect 174221 134523 174287 134526
rect 62901 134314 62967 134317
rect 135305 134314 135371 134317
rect 60742 134312 62967 134314
rect 60742 134256 62906 134312
rect 62962 134256 62967 134312
rect 60742 134254 62967 134256
rect 60742 133944 60802 134254
rect 62901 134251 62967 134254
rect 132686 134312 135371 134314
rect 132686 134256 135310 134312
rect 135366 134256 135371 134312
rect 132686 134254 135371 134256
rect 65477 134178 65543 134181
rect 65477 134176 67948 134178
rect 65477 134120 65482 134176
rect 65538 134120 67948 134176
rect 65477 134118 67948 134120
rect 65477 134115 65543 134118
rect 62993 133634 63059 133637
rect 60742 133632 63059 133634
rect 60742 133576 62998 133632
rect 63054 133576 63059 133632
rect 60742 133574 63059 133576
rect 97726 133634 97786 134080
rect 132686 133944 132746 134254
rect 135305 134251 135371 134254
rect 102369 133906 102435 133909
rect 102369 133904 104932 133906
rect 102369 133848 102374 133904
rect 102430 133848 104932 133904
rect 102369 133846 104932 133848
rect 102369 133843 102435 133846
rect 100897 133634 100963 133637
rect 134293 133634 134359 133637
rect 97726 133632 100963 133634
rect 97726 133576 100902 133632
rect 100958 133576 100963 133632
rect 97726 133574 100963 133576
rect 60742 133400 60802 133574
rect 62993 133571 63059 133574
rect 100897 133571 100963 133574
rect 132686 133632 134359 133634
rect 132686 133576 134298 133632
rect 134354 133576 134359 133632
rect 132686 133574 134359 133576
rect 66397 133498 66463 133501
rect 66397 133496 67948 133498
rect 66397 133440 66402 133496
rect 66458 133440 67948 133496
rect 66397 133438 67948 133440
rect 66397 133435 66463 133438
rect 132686 133400 132746 133574
rect 134293 133571 134359 133574
rect 136961 133634 137027 133637
rect 140046 133634 140106 134080
rect 136961 133632 140106 133634
rect 136961 133576 136966 133632
rect 137022 133576 140106 133632
rect 136961 133574 140106 133576
rect 169854 133634 169914 134148
rect 173945 133906 174011 133909
rect 173945 133904 177060 133906
rect 173945 133848 173950 133904
rect 174006 133848 177060 133904
rect 173945 133846 177060 133848
rect 173945 133843 174011 133846
rect 171645 133634 171711 133637
rect 169854 133632 171711 133634
rect 169854 133576 171650 133632
rect 171706 133576 171711 133632
rect 169854 133574 171711 133576
rect 136961 133571 137027 133574
rect 171645 133571 171711 133574
rect 97726 133226 97786 133400
rect 102001 133362 102067 133365
rect 102001 133360 104932 133362
rect 102001 133304 102006 133360
rect 102062 133304 104932 133360
rect 102001 133302 104932 133304
rect 102001 133299 102067 133302
rect 100253 133226 100319 133229
rect 97726 133224 100319 133226
rect 97726 133168 100258 133224
rect 100314 133168 100319 133224
rect 97726 133166 100319 133168
rect 100253 133163 100319 133166
rect 136869 133090 136935 133093
rect 140046 133090 140106 133400
rect 136869 133088 140106 133090
rect 136869 133032 136874 133088
rect 136930 133032 140106 133088
rect 136869 133030 140106 133032
rect 169854 133090 169914 133468
rect 173761 133362 173827 133365
rect 173761 133360 177060 133362
rect 173761 133304 173766 133360
rect 173822 133304 177060 133360
rect 173761 133302 177060 133304
rect 173761 133299 173827 133302
rect 172657 133090 172723 133093
rect 169854 133088 172723 133090
rect 169854 133032 172662 133088
rect 172718 133032 172723 133088
rect 169854 133030 172723 133032
rect 136869 133027 136935 133030
rect 172657 133027 172723 133030
rect 62809 132818 62875 132821
rect 60772 132816 62875 132818
rect 60772 132760 62814 132816
rect 62870 132760 62875 132816
rect 60772 132758 62875 132760
rect 62809 132755 62875 132758
rect 62717 132546 62783 132549
rect 60742 132544 62783 132546
rect 60742 132488 62722 132544
rect 62778 132488 62783 132544
rect 60742 132486 62783 132488
rect 60742 132312 60802 132486
rect 62717 132483 62783 132486
rect 65017 132546 65083 132549
rect 67918 132546 67978 132924
rect 65017 132544 67978 132546
rect 65017 132488 65022 132544
rect 65078 132488 67978 132544
rect 65017 132486 67978 132488
rect 65017 132483 65083 132486
rect 97726 132410 97786 132856
rect 102277 132818 102343 132821
rect 135397 132818 135463 132821
rect 102277 132816 104932 132818
rect 102277 132760 102282 132816
rect 102338 132760 104932 132816
rect 102277 132758 104932 132760
rect 132716 132816 135463 132818
rect 132716 132760 135402 132816
rect 135458 132760 135463 132816
rect 132716 132758 135463 132760
rect 102277 132755 102343 132758
rect 135397 132755 135463 132758
rect 135121 132546 135187 132549
rect 132686 132544 135187 132546
rect 132686 132488 135126 132544
rect 135182 132488 135187 132544
rect 132686 132486 135187 132488
rect 100253 132410 100319 132413
rect 97726 132408 100319 132410
rect 97726 132352 100258 132408
rect 100314 132352 100319 132408
rect 97726 132350 100319 132352
rect 100253 132347 100319 132350
rect 132686 132312 132746 132486
rect 135121 132483 135187 132486
rect 136777 132410 136843 132413
rect 140046 132410 140106 132856
rect 136777 132408 140106 132410
rect 136777 132352 136782 132408
rect 136838 132352 140106 132408
rect 136777 132350 140106 132352
rect 169854 132410 169914 132924
rect 174037 132818 174103 132821
rect 174037 132816 177060 132818
rect 174037 132760 174042 132816
rect 174098 132760 177060 132816
rect 174037 132758 177060 132760
rect 174037 132755 174103 132758
rect 172013 132410 172079 132413
rect 169854 132408 172079 132410
rect 169854 132352 172018 132408
rect 172074 132352 172079 132408
rect 169854 132350 172079 132352
rect 136777 132347 136843 132350
rect 172013 132347 172079 132350
rect 66397 132274 66463 132277
rect 102093 132274 102159 132277
rect 173853 132274 173919 132277
rect 66397 132272 67948 132274
rect 66397 132216 66402 132272
rect 66458 132216 67948 132272
rect 66397 132214 67948 132216
rect 102093 132272 104932 132274
rect 102093 132216 102098 132272
rect 102154 132216 104932 132272
rect 173853 132272 177060 132274
rect 102093 132214 104932 132216
rect 66397 132211 66463 132214
rect 102093 132211 102159 132214
rect 97726 132002 97786 132176
rect 100897 132002 100963 132005
rect 97726 132000 100963 132002
rect 97726 131944 100902 132000
rect 100958 131944 100963 132000
rect 97726 131942 100963 131944
rect 100897 131939 100963 131942
rect 136869 132002 136935 132005
rect 140046 132002 140106 132176
rect 136869 132000 140106 132002
rect 136869 131944 136874 132000
rect 136930 131944 140106 132000
rect 136869 131942 140106 131944
rect 169854 132002 169914 132244
rect 173853 132216 173858 132272
rect 173914 132216 177060 132272
rect 173853 132214 177060 132216
rect 173853 132211 173919 132214
rect 171645 132002 171711 132005
rect 169854 132000 171711 132002
rect 169854 131944 171650 132000
rect 171706 131944 171711 132000
rect 169854 131942 171711 131944
rect 136869 131939 136935 131942
rect 171645 131939 171711 131942
rect 172657 131866 172723 131869
rect 169670 131864 172723 131866
rect 169670 131808 172662 131864
rect 172718 131808 172723 131864
rect 169670 131806 172723 131808
rect 65661 131730 65727 131733
rect 100897 131730 100963 131733
rect 65661 131728 67948 131730
rect 65661 131672 65666 131728
rect 65722 131672 67948 131728
rect 65661 131670 67948 131672
rect 97756 131728 100963 131730
rect 97756 131672 100902 131728
rect 100958 131672 100963 131728
rect 97756 131670 100963 131672
rect 65661 131667 65727 131670
rect 100897 131667 100963 131670
rect 136961 131730 137027 131733
rect 136961 131728 140076 131730
rect 136961 131672 136966 131728
rect 137022 131672 140076 131728
rect 169670 131700 169730 131806
rect 172657 131803 172723 131806
rect 136961 131670 140076 131672
rect 136961 131667 137027 131670
rect 63453 131594 63519 131597
rect 60772 131592 63519 131594
rect 60772 131536 63458 131592
rect 63514 131536 63519 131592
rect 60772 131534 63519 131536
rect 63453 131531 63519 131534
rect 102001 131594 102067 131597
rect 135213 131594 135279 131597
rect 102001 131592 104932 131594
rect 102001 131536 102006 131592
rect 102062 131536 104932 131592
rect 102001 131534 104932 131536
rect 132716 131592 135279 131594
rect 132716 131536 135218 131592
rect 135274 131536 135279 131592
rect 132716 131534 135279 131536
rect 102001 131531 102067 131534
rect 135213 131531 135279 131534
rect 174129 131594 174195 131597
rect 174129 131592 177060 131594
rect 174129 131536 174134 131592
rect 174190 131536 177060 131592
rect 174129 131534 177060 131536
rect 174129 131531 174195 131534
rect 101398 131396 101404 131460
rect 101468 131458 101474 131460
rect 101909 131458 101975 131461
rect 101468 131456 101975 131458
rect 101468 131400 101914 131456
rect 101970 131400 101975 131456
rect 101468 131398 101975 131400
rect 101468 131396 101474 131398
rect 101909 131395 101975 131398
rect 63545 131322 63611 131325
rect 135305 131322 135371 131325
rect 60742 131320 63611 131322
rect 60742 131264 63550 131320
rect 63606 131264 63611 131320
rect 60742 131262 63611 131264
rect 60742 131088 60802 131262
rect 63545 131259 63611 131262
rect 132686 131320 135371 131322
rect 132686 131264 135310 131320
rect 135366 131264 135371 131320
rect 132686 131262 135371 131264
rect 66305 131186 66371 131189
rect 66305 131184 67948 131186
rect 66305 131128 66310 131184
rect 66366 131128 67948 131184
rect 66305 131126 67948 131128
rect 66305 131123 66371 131126
rect 132686 131088 132746 131262
rect 135305 131259 135371 131262
rect 62809 130778 62875 130781
rect 60742 130776 62875 130778
rect 60742 130720 62814 130776
rect 62870 130720 62875 130776
rect 60742 130718 62875 130720
rect 60742 130544 60802 130718
rect 62809 130715 62875 130718
rect 97726 130642 97786 131088
rect 102185 131050 102251 131053
rect 102185 131048 104932 131050
rect 102185 130992 102190 131048
rect 102246 130992 104932 131048
rect 102185 130990 104932 130992
rect 102185 130987 102251 130990
rect 102277 130778 102343 130781
rect 134293 130778 134359 130781
rect 102277 130776 104962 130778
rect 102277 130720 102282 130776
rect 102338 130720 104962 130776
rect 102277 130718 104962 130720
rect 102277 130715 102343 130718
rect 100253 130642 100319 130645
rect 97726 130640 100319 130642
rect 97726 130584 100258 130640
rect 100314 130584 100319 130640
rect 97726 130582 100319 130584
rect 100253 130579 100319 130582
rect 66397 130506 66463 130509
rect 100897 130506 100963 130509
rect 66397 130504 67948 130506
rect 66397 130448 66402 130504
rect 66458 130448 67948 130504
rect 66397 130446 67948 130448
rect 97756 130504 100963 130506
rect 97756 130448 100902 130504
rect 100958 130448 100963 130504
rect 104902 130476 104962 130718
rect 132686 130776 134359 130778
rect 132686 130720 134298 130776
rect 134354 130720 134359 130776
rect 132686 130718 134359 130720
rect 132686 130544 132746 130718
rect 134293 130715 134359 130718
rect 136869 130642 136935 130645
rect 140046 130642 140106 131088
rect 136869 130640 140106 130642
rect 136869 130584 136874 130640
rect 136930 130584 140106 130640
rect 136869 130582 140106 130584
rect 169854 130642 169914 131156
rect 175049 131050 175115 131053
rect 175049 131048 177060 131050
rect 175049 130992 175054 131048
rect 175110 130992 177060 131048
rect 175049 130990 177060 130992
rect 175049 130987 175115 130990
rect 172381 130642 172447 130645
rect 169854 130640 172447 130642
rect 169854 130584 172386 130640
rect 172442 130584 172447 130640
rect 169854 130582 172447 130584
rect 136869 130579 136935 130582
rect 172381 130579 172447 130582
rect 136961 130506 137027 130509
rect 174129 130506 174195 130509
rect 136961 130504 140076 130506
rect 97756 130446 100963 130448
rect 66397 130443 66463 130446
rect 100897 130443 100963 130446
rect 136961 130448 136966 130504
rect 137022 130448 140076 130504
rect 174129 130504 177060 130506
rect 136961 130446 140076 130448
rect 136961 130443 137027 130446
rect 169854 130370 169914 130476
rect 174129 130448 174134 130504
rect 174190 130448 177060 130504
rect 174129 130446 177060 130448
rect 174129 130443 174195 130446
rect 172657 130370 172723 130373
rect 169854 130368 172723 130370
rect 169854 130312 172662 130368
rect 172718 130312 172723 130368
rect 169854 130310 172723 130312
rect 172657 130307 172723 130310
rect 63637 130234 63703 130237
rect 135397 130234 135463 130237
rect 60742 130232 63703 130234
rect 60742 130176 63642 130232
rect 63698 130176 63703 130232
rect 60742 130174 63703 130176
rect 60742 129864 60802 130174
rect 63637 130171 63703 130174
rect 132686 130232 135463 130234
rect 132686 130176 135402 130232
rect 135458 130176 135463 130232
rect 132686 130174 135463 130176
rect 65477 129962 65543 129965
rect 65477 129960 67948 129962
rect 65477 129904 65482 129960
rect 65538 129904 67948 129960
rect 65477 129902 67948 129904
rect 65477 129899 65543 129902
rect 132686 129864 132746 130174
rect 135397 130171 135463 130174
rect 63085 129554 63151 129557
rect 60742 129552 63151 129554
rect 60742 129496 63090 129552
rect 63146 129496 63151 129552
rect 60742 129494 63151 129496
rect 60742 129320 60802 129494
rect 63085 129491 63151 129494
rect 97726 129418 97786 129864
rect 102369 129826 102435 129829
rect 102369 129824 104932 129826
rect 102369 129768 102374 129824
rect 102430 129768 104932 129824
rect 102369 129766 104932 129768
rect 102369 129763 102435 129766
rect 135029 129554 135095 129557
rect 132686 129552 135095 129554
rect 132686 129496 135034 129552
rect 135090 129496 135095 129552
rect 132686 129494 135095 129496
rect 100253 129418 100319 129421
rect 97726 129416 100319 129418
rect 97726 129360 100258 129416
rect 100314 129360 100319 129416
rect 97726 129358 100319 129360
rect 100253 129355 100319 129358
rect 132686 129320 132746 129494
rect 135029 129491 135095 129494
rect 136869 129418 136935 129421
rect 140046 129418 140106 129864
rect 136869 129416 140106 129418
rect 136869 129360 136874 129416
rect 136930 129360 140106 129416
rect 136869 129358 140106 129360
rect 169854 129418 169914 129932
rect 174129 129826 174195 129829
rect 174129 129824 177060 129826
rect 174129 129768 174134 129824
rect 174190 129768 177060 129824
rect 174129 129766 177060 129768
rect 174129 129763 174195 129766
rect 172657 129418 172723 129421
rect 169854 129416 172723 129418
rect 169854 129360 172662 129416
rect 172718 129360 172723 129416
rect 169854 129358 172723 129360
rect 136869 129355 136935 129358
rect 172657 129355 172723 129358
rect 66397 129282 66463 129285
rect 102093 129282 102159 129285
rect 174497 129282 174563 129285
rect 66397 129280 67948 129282
rect 66397 129224 66402 129280
rect 66458 129224 67948 129280
rect 66397 129222 67948 129224
rect 102093 129280 104932 129282
rect 102093 129224 102098 129280
rect 102154 129224 104932 129280
rect 174497 129280 177060 129282
rect 102093 129222 104932 129224
rect 66397 129219 66463 129222
rect 102093 129219 102159 129222
rect 97726 129010 97786 129184
rect 100897 129010 100963 129013
rect 97726 129008 100963 129010
rect 97726 128952 100902 129008
rect 100958 128952 100963 129008
rect 97726 128950 100963 128952
rect 100897 128947 100963 128950
rect 136961 129010 137027 129013
rect 140046 129010 140106 129184
rect 136961 129008 140106 129010
rect 136961 128952 136966 129008
rect 137022 128952 140106 129008
rect 136961 128950 140106 128952
rect 169854 129010 169914 129252
rect 174497 129224 174502 129280
rect 174558 129224 177060 129280
rect 174497 129222 177060 129224
rect 174497 129219 174563 129222
rect 172657 129010 172723 129013
rect 169854 129008 172723 129010
rect 169854 128952 172662 129008
rect 172718 128952 172723 129008
rect 169854 128950 172723 128952
rect 136961 128947 137027 128950
rect 172657 128947 172723 128950
rect 62717 128738 62783 128741
rect 60772 128736 62783 128738
rect 60772 128680 62722 128736
rect 62778 128680 62783 128736
rect 102277 128738 102343 128741
rect 135305 128738 135371 128741
rect 102277 128736 104932 128738
rect 60772 128678 62783 128680
rect 62717 128675 62783 128678
rect 62901 128466 62967 128469
rect 60742 128464 62967 128466
rect 60742 128408 62906 128464
rect 62962 128408 62967 128464
rect 60742 128406 62967 128408
rect 60742 128232 60802 128406
rect 62901 128403 62967 128406
rect 67918 128330 67978 128708
rect 102277 128680 102282 128736
rect 102338 128680 104932 128736
rect 102277 128678 104932 128680
rect 132716 128736 135371 128738
rect 132716 128680 135310 128736
rect 135366 128680 135371 128736
rect 174037 128738 174103 128741
rect 174037 128736 177060 128738
rect 132716 128678 135371 128680
rect 102277 128675 102343 128678
rect 135305 128675 135371 128678
rect 66262 128270 67978 128330
rect 97726 128330 97786 128640
rect 135121 128466 135187 128469
rect 132686 128464 135187 128466
rect 132686 128408 135126 128464
rect 135182 128408 135187 128464
rect 132686 128406 135187 128408
rect 100069 128330 100135 128333
rect 97726 128328 100135 128330
rect 97726 128272 100074 128328
rect 100130 128272 100135 128328
rect 97726 128270 100135 128272
rect 65017 127922 65083 127925
rect 66262 127922 66322 128270
rect 100069 128267 100135 128270
rect 132686 128232 132746 128406
rect 135121 128403 135187 128406
rect 136777 128330 136843 128333
rect 140046 128330 140106 128640
rect 136777 128328 140106 128330
rect 136777 128272 136782 128328
rect 136838 128272 140106 128328
rect 136777 128270 140106 128272
rect 169854 128330 169914 128708
rect 174037 128680 174042 128736
rect 174098 128680 177060 128736
rect 174037 128678 177060 128680
rect 174037 128675 174103 128678
rect 171645 128330 171711 128333
rect 169854 128328 171711 128330
rect 169854 128272 171650 128328
rect 171706 128272 171711 128328
rect 169854 128270 171711 128272
rect 136777 128267 136843 128270
rect 171645 128267 171711 128270
rect 66397 128194 66463 128197
rect 102001 128194 102067 128197
rect 174129 128194 174195 128197
rect 66397 128192 67948 128194
rect 66397 128136 66402 128192
rect 66458 128136 67948 128192
rect 66397 128134 67948 128136
rect 102001 128192 104932 128194
rect 102001 128136 102006 128192
rect 102062 128136 104932 128192
rect 174129 128192 177060 128194
rect 102001 128134 104932 128136
rect 66397 128131 66463 128134
rect 102001 128131 102067 128134
rect 65017 127920 66322 127922
rect 65017 127864 65022 127920
rect 65078 127864 66322 127920
rect 65017 127862 66322 127864
rect 65017 127859 65083 127862
rect 9896 127786 10376 127816
rect 30425 127786 30491 127789
rect 9896 127726 10570 127786
rect 9896 127696 10376 127726
rect 10510 127650 10570 127726
rect 30425 127784 32988 127786
rect 30425 127728 30430 127784
rect 30486 127728 32988 127784
rect 30425 127726 32988 127728
rect 30425 127723 30491 127726
rect 21542 127650 21548 127652
rect 10510 127590 21548 127650
rect 21542 127588 21548 127590
rect 21612 127588 21618 127652
rect 97726 127650 97786 128096
rect 100805 127650 100871 127653
rect 97726 127648 100871 127650
rect 97726 127592 100810 127648
rect 100866 127592 100871 127648
rect 97726 127590 100871 127592
rect 100805 127587 100871 127590
rect 136869 127650 136935 127653
rect 140046 127650 140106 128096
rect 136869 127648 140106 127650
rect 136869 127592 136874 127648
rect 136930 127592 140106 127648
rect 136869 127590 140106 127592
rect 169854 127650 169914 128164
rect 174129 128136 174134 128192
rect 174190 128136 177060 128192
rect 174129 128134 177060 128136
rect 174129 128131 174195 128134
rect 207985 127786 208051 127789
rect 204844 127784 208051 127786
rect 204844 127728 207990 127784
rect 208046 127728 208051 127784
rect 204844 127726 208051 127728
rect 207985 127723 208051 127726
rect 172657 127650 172723 127653
rect 169854 127648 172723 127650
rect 169854 127592 172662 127648
rect 172718 127592 172723 127648
rect 169854 127590 172723 127592
rect 136869 127587 136935 127590
rect 172657 127587 172723 127590
rect 62809 127514 62875 127517
rect 60772 127512 62875 127514
rect 60772 127456 62814 127512
rect 62870 127456 62875 127512
rect 102093 127514 102159 127517
rect 135213 127514 135279 127517
rect 102093 127512 104932 127514
rect 60772 127454 62875 127456
rect 62809 127451 62875 127454
rect 62625 127242 62691 127245
rect 60742 127240 62691 127242
rect 60742 127184 62630 127240
rect 62686 127184 62691 127240
rect 60742 127182 62691 127184
rect 60742 127008 60802 127182
rect 62625 127179 62691 127182
rect 67918 127106 67978 127484
rect 102093 127456 102098 127512
rect 102154 127456 104932 127512
rect 102093 127454 104932 127456
rect 132716 127512 135279 127514
rect 132716 127456 135218 127512
rect 135274 127456 135279 127512
rect 173945 127514 174011 127517
rect 173945 127512 177060 127514
rect 132716 127454 135279 127456
rect 102093 127451 102159 127454
rect 135213 127451 135279 127454
rect 66078 127046 67978 127106
rect 97726 127106 97786 127416
rect 134293 127242 134359 127245
rect 132686 127240 134359 127242
rect 132686 127184 134298 127240
rect 134354 127184 134359 127240
rect 132686 127182 134359 127184
rect 100529 127106 100595 127109
rect 97726 127104 100595 127106
rect 97726 127048 100534 127104
rect 100590 127048 100595 127104
rect 97726 127046 100595 127048
rect 62809 126698 62875 126701
rect 60742 126696 62875 126698
rect 60742 126640 62814 126696
rect 62870 126640 62875 126696
rect 60742 126638 62875 126640
rect 60742 126464 60802 126638
rect 62809 126635 62875 126638
rect 65017 126562 65083 126565
rect 66078 126562 66138 127046
rect 100529 127043 100595 127046
rect 132686 127008 132746 127182
rect 134293 127179 134359 127182
rect 136777 127106 136843 127109
rect 140046 127106 140106 127416
rect 136777 127104 140106 127106
rect 136777 127048 136782 127104
rect 136838 127048 140106 127104
rect 136777 127046 140106 127048
rect 169854 127106 169914 127484
rect 173945 127456 173950 127512
rect 174006 127456 177060 127512
rect 173945 127454 177060 127456
rect 173945 127451 174011 127454
rect 172013 127106 172079 127109
rect 169854 127104 172079 127106
rect 169854 127048 172018 127104
rect 172074 127048 172079 127104
rect 169854 127046 172079 127048
rect 136777 127043 136843 127046
rect 172013 127043 172079 127046
rect 66305 126970 66371 126973
rect 102185 126970 102251 126973
rect 173853 126970 173919 126973
rect 66305 126968 67948 126970
rect 66305 126912 66310 126968
rect 66366 126912 67948 126968
rect 66305 126910 67948 126912
rect 102185 126968 104932 126970
rect 102185 126912 102190 126968
rect 102246 126912 104932 126968
rect 173853 126968 177060 126970
rect 102185 126910 104932 126912
rect 66305 126907 66371 126910
rect 102185 126907 102251 126910
rect 65017 126560 66138 126562
rect 65017 126504 65022 126560
rect 65078 126504 66138 126560
rect 65017 126502 66138 126504
rect 65017 126499 65083 126502
rect 97726 126426 97786 126872
rect 134661 126698 134727 126701
rect 132686 126696 134727 126698
rect 132686 126640 134666 126696
rect 134722 126640 134727 126696
rect 132686 126638 134727 126640
rect 132686 126464 132746 126638
rect 134661 126635 134727 126638
rect 100621 126426 100687 126429
rect 97726 126424 100687 126426
rect 97726 126368 100626 126424
rect 100682 126368 100687 126424
rect 97726 126366 100687 126368
rect 100621 126363 100687 126366
rect 102277 126426 102343 126429
rect 136869 126426 136935 126429
rect 140046 126426 140106 126872
rect 102277 126424 104932 126426
rect 102277 126368 102282 126424
rect 102338 126368 104932 126424
rect 102277 126366 104932 126368
rect 136869 126424 140106 126426
rect 136869 126368 136874 126424
rect 136930 126368 140106 126424
rect 136869 126366 140106 126368
rect 169854 126426 169914 126940
rect 173853 126912 173858 126968
rect 173914 126912 177060 126968
rect 173853 126910 177060 126912
rect 173853 126907 173919 126910
rect 172381 126426 172447 126429
rect 169854 126424 172447 126426
rect 169854 126368 172386 126424
rect 172442 126368 172447 126424
rect 169854 126366 172447 126368
rect 102277 126363 102343 126366
rect 136869 126363 136935 126366
rect 172381 126363 172447 126366
rect 174221 126426 174287 126429
rect 174221 126424 177060 126426
rect 174221 126368 174226 126424
rect 174282 126368 177060 126424
rect 174221 126366 177060 126368
rect 174221 126363 174287 126366
rect 66397 126290 66463 126293
rect 100897 126290 100963 126293
rect 66397 126288 67948 126290
rect 66397 126232 66402 126288
rect 66458 126232 67948 126288
rect 66397 126230 67948 126232
rect 97756 126288 100963 126290
rect 97756 126232 100902 126288
rect 100958 126232 100963 126288
rect 97756 126230 100963 126232
rect 66397 126227 66463 126230
rect 100897 126227 100963 126230
rect 136961 126290 137027 126293
rect 136961 126288 140076 126290
rect 136961 126232 136966 126288
rect 137022 126232 140076 126288
rect 136961 126230 140076 126232
rect 136961 126227 137027 126230
rect 169854 126154 169914 126260
rect 172657 126154 172723 126157
rect 169854 126152 172723 126154
rect 169854 126096 172662 126152
rect 172718 126096 172723 126152
rect 169854 126094 172723 126096
rect 172657 126091 172723 126094
rect 62901 126018 62967 126021
rect 135121 126018 135187 126021
rect 60742 126016 62967 126018
rect 60742 125960 62906 126016
rect 62962 125960 62967 126016
rect 60742 125958 62967 125960
rect 60742 125784 60802 125958
rect 62901 125955 62967 125958
rect 132686 126016 135187 126018
rect 132686 125960 135126 126016
rect 135182 125960 135187 126016
rect 132686 125958 135187 125960
rect 132686 125784 132746 125958
rect 135121 125955 135187 125958
rect 66397 125746 66463 125749
rect 102001 125746 102067 125749
rect 174221 125746 174287 125749
rect 66397 125744 67948 125746
rect 66397 125688 66402 125744
rect 66458 125688 67948 125744
rect 66397 125686 67948 125688
rect 102001 125744 104932 125746
rect 102001 125688 102006 125744
rect 102062 125688 104932 125744
rect 174221 125744 177060 125746
rect 102001 125686 104932 125688
rect 66397 125683 66463 125686
rect 102001 125683 102067 125686
rect 62809 125474 62875 125477
rect 60742 125472 62875 125474
rect 60742 125416 62814 125472
rect 62870 125416 62875 125472
rect 60742 125414 62875 125416
rect 60742 125240 60802 125414
rect 62809 125411 62875 125414
rect 97726 125338 97786 125648
rect 134845 125474 134911 125477
rect 132686 125472 134911 125474
rect 132686 125416 134850 125472
rect 134906 125416 134911 125472
rect 132686 125414 134911 125416
rect 100621 125338 100687 125341
rect 97726 125336 100687 125338
rect 97726 125280 100626 125336
rect 100682 125280 100687 125336
rect 97726 125278 100687 125280
rect 100621 125275 100687 125278
rect 132686 125240 132746 125414
rect 134845 125411 134911 125414
rect 136777 125338 136843 125341
rect 140046 125338 140106 125648
rect 136777 125336 140106 125338
rect 136777 125280 136782 125336
rect 136838 125280 140106 125336
rect 136777 125278 140106 125280
rect 169854 125338 169914 125716
rect 174221 125688 174226 125744
rect 174282 125688 177060 125744
rect 174221 125686 177060 125688
rect 174221 125683 174287 125686
rect 172013 125338 172079 125341
rect 169854 125336 172079 125338
rect 169854 125280 172018 125336
rect 172074 125280 172079 125336
rect 169854 125278 172079 125280
rect 136777 125275 136843 125278
rect 172013 125275 172079 125278
rect 65845 125202 65911 125205
rect 102369 125202 102435 125205
rect 174129 125202 174195 125205
rect 65845 125200 67948 125202
rect 65845 125144 65850 125200
rect 65906 125144 67948 125200
rect 65845 125142 67948 125144
rect 102369 125200 104932 125202
rect 102369 125144 102374 125200
rect 102430 125144 104932 125200
rect 174129 125200 177060 125202
rect 102369 125142 104932 125144
rect 65845 125139 65911 125142
rect 102369 125139 102435 125142
rect 65017 124930 65083 124933
rect 66397 124930 66463 124933
rect 65017 124928 66463 124930
rect 65017 124872 65022 124928
rect 65078 124872 66402 124928
rect 66458 124872 66463 124928
rect 65017 124870 66463 124872
rect 97726 124930 97786 125104
rect 100621 124930 100687 124933
rect 97726 124928 100687 124930
rect 97726 124872 100626 124928
rect 100682 124872 100687 124928
rect 97726 124870 100687 124872
rect 65017 124867 65083 124870
rect 66397 124867 66463 124870
rect 100621 124867 100687 124870
rect 136869 124930 136935 124933
rect 140046 124930 140106 125104
rect 136869 124928 140106 124930
rect 136869 124872 136874 124928
rect 136930 124872 140106 124928
rect 136869 124870 140106 124872
rect 169854 124930 169914 125172
rect 174129 125144 174134 125200
rect 174190 125144 177060 125200
rect 174129 125142 177060 125144
rect 174129 125139 174195 125142
rect 172657 124930 172723 124933
rect 169854 124928 172723 124930
rect 169854 124872 172662 124928
rect 172718 124872 172723 124928
rect 169854 124870 172723 124872
rect 136869 124867 136935 124870
rect 172657 124867 172723 124870
rect 62717 124658 62783 124661
rect 60772 124656 62783 124658
rect 60772 124600 62722 124656
rect 62778 124600 62783 124656
rect 60772 124598 62783 124600
rect 62717 124595 62783 124598
rect 102277 124658 102343 124661
rect 135305 124658 135371 124661
rect 102277 124656 104932 124658
rect 102277 124600 102282 124656
rect 102338 124600 104932 124656
rect 102277 124598 104932 124600
rect 132716 124656 135371 124658
rect 132716 124600 135310 124656
rect 135366 124600 135371 124656
rect 132716 124598 135371 124600
rect 102277 124595 102343 124598
rect 135305 124595 135371 124598
rect 174037 124658 174103 124661
rect 174037 124656 177060 124658
rect 174037 124600 174042 124656
rect 174098 124600 177060 124656
rect 174037 124598 177060 124600
rect 174037 124595 174103 124598
rect 62625 124386 62691 124389
rect 60742 124384 62691 124386
rect 60742 124328 62630 124384
rect 62686 124328 62691 124384
rect 60742 124326 62691 124328
rect 60742 124016 60802 124326
rect 62625 124323 62691 124326
rect 67918 124114 67978 124492
rect 66262 124054 67978 124114
rect 97726 124114 97786 124424
rect 135397 124386 135463 124389
rect 132686 124384 135463 124386
rect 132686 124328 135402 124384
rect 135458 124328 135463 124384
rect 132686 124326 135463 124328
rect 100621 124114 100687 124117
rect 97726 124112 100687 124114
rect 97726 124056 100626 124112
rect 100682 124056 100687 124112
rect 97726 124054 100687 124056
rect 62809 123706 62875 123709
rect 60742 123704 62875 123706
rect 60742 123648 62814 123704
rect 62870 123648 62875 123704
rect 60742 123646 62875 123648
rect 60742 123472 60802 123646
rect 62809 123643 62875 123646
rect 65017 123570 65083 123573
rect 66262 123570 66322 124054
rect 100621 124051 100687 124054
rect 132686 124016 132746 124326
rect 135397 124323 135463 124326
rect 136777 124114 136843 124117
rect 140046 124114 140106 124424
rect 136777 124112 140106 124114
rect 136777 124056 136782 124112
rect 136838 124056 140106 124112
rect 136777 124054 140106 124056
rect 169854 124114 169914 124492
rect 172381 124114 172447 124117
rect 169854 124112 172447 124114
rect 169854 124056 172386 124112
rect 172442 124056 172447 124112
rect 169854 124054 172447 124056
rect 136777 124051 136843 124054
rect 172381 124051 172447 124054
rect 66397 123978 66463 123981
rect 102369 123978 102435 123981
rect 173853 123978 173919 123981
rect 66397 123976 67948 123978
rect 66397 123920 66402 123976
rect 66458 123920 67948 123976
rect 66397 123918 67948 123920
rect 102369 123976 104932 123978
rect 102369 123920 102374 123976
rect 102430 123920 104932 123976
rect 173853 123976 177060 123978
rect 102369 123918 104932 123920
rect 66397 123915 66463 123918
rect 102369 123915 102435 123918
rect 65017 123568 66322 123570
rect 65017 123512 65022 123568
rect 65078 123512 66322 123568
rect 65017 123510 66322 123512
rect 65017 123507 65083 123510
rect 97726 123434 97786 123880
rect 135213 123706 135279 123709
rect 132686 123704 135279 123706
rect 132686 123648 135218 123704
rect 135274 123648 135279 123704
rect 132686 123646 135279 123648
rect 132686 123472 132746 123646
rect 135213 123643 135279 123646
rect 99885 123434 99951 123437
rect 97726 123432 99951 123434
rect 97726 123376 99890 123432
rect 99946 123376 99951 123432
rect 97726 123374 99951 123376
rect 99885 123371 99951 123374
rect 102093 123434 102159 123437
rect 136869 123434 136935 123437
rect 140046 123434 140106 123880
rect 102093 123432 104932 123434
rect 102093 123376 102098 123432
rect 102154 123376 104932 123432
rect 102093 123374 104932 123376
rect 136869 123432 140106 123434
rect 136869 123376 136874 123432
rect 136930 123376 140106 123432
rect 136869 123374 140106 123376
rect 169854 123434 169914 123948
rect 173853 123920 173858 123976
rect 173914 123920 177060 123976
rect 173853 123918 177060 123920
rect 173853 123915 173919 123918
rect 172657 123434 172723 123437
rect 169854 123432 172723 123434
rect 169854 123376 172662 123432
rect 172718 123376 172723 123432
rect 169854 123374 172723 123376
rect 102093 123371 102159 123374
rect 136869 123371 136935 123374
rect 172657 123371 172723 123374
rect 174221 123434 174287 123437
rect 174221 123432 177060 123434
rect 174221 123376 174226 123432
rect 174282 123376 177060 123432
rect 174221 123374 177060 123376
rect 174221 123371 174287 123374
rect 62901 123162 62967 123165
rect 60742 123160 62967 123162
rect 60742 123104 62906 123160
rect 62962 123104 62967 123160
rect 60742 123102 62967 123104
rect 60742 122928 60802 123102
rect 62901 123099 62967 123102
rect 67918 122890 67978 123268
rect 66078 122830 67978 122890
rect 97726 122890 97786 123200
rect 135121 123162 135187 123165
rect 132686 123160 135187 123162
rect 132686 123104 135126 123160
rect 135182 123104 135187 123160
rect 132686 123102 135187 123104
rect 132686 122928 132746 123102
rect 135121 123099 135187 123102
rect 100161 122890 100227 122893
rect 97726 122888 100227 122890
rect 97726 122832 100166 122888
rect 100222 122832 100227 122888
rect 97726 122830 100227 122832
rect 62809 122618 62875 122621
rect 60742 122616 62875 122618
rect 60742 122560 62814 122616
rect 62870 122560 62875 122616
rect 60742 122558 62875 122560
rect 60742 122384 60802 122558
rect 62809 122555 62875 122558
rect 65017 122482 65083 122485
rect 66078 122482 66138 122830
rect 100161 122827 100227 122830
rect 102001 122890 102067 122893
rect 136869 122890 136935 122893
rect 140046 122890 140106 123200
rect 102001 122888 104932 122890
rect 102001 122832 102006 122888
rect 102062 122832 104932 122888
rect 102001 122830 104932 122832
rect 136869 122888 140106 122890
rect 136869 122832 136874 122888
rect 136930 122832 140106 122888
rect 136869 122830 140106 122832
rect 169854 122890 169914 123268
rect 171553 122890 171619 122893
rect 169854 122888 171619 122890
rect 169854 122832 171558 122888
rect 171614 122832 171619 122888
rect 169854 122830 171619 122832
rect 102001 122827 102067 122830
rect 136869 122827 136935 122830
rect 171553 122827 171619 122830
rect 173945 122890 174011 122893
rect 173945 122888 177060 122890
rect 173945 122832 173950 122888
rect 174006 122832 177060 122888
rect 173945 122830 177060 122832
rect 173945 122827 174011 122830
rect 66305 122754 66371 122757
rect 66305 122752 67948 122754
rect 66305 122696 66310 122752
rect 66366 122696 67948 122752
rect 66305 122694 67948 122696
rect 66305 122691 66371 122694
rect 65017 122480 66138 122482
rect 65017 122424 65022 122480
rect 65078 122424 66138 122480
rect 65017 122422 66138 122424
rect 65017 122419 65083 122422
rect 97726 122346 97786 122656
rect 135305 122618 135371 122621
rect 132686 122616 135371 122618
rect 132686 122560 135310 122616
rect 135366 122560 135371 122616
rect 132686 122558 135371 122560
rect 132686 122384 132746 122558
rect 135305 122555 135371 122558
rect 136961 122482 137027 122485
rect 140046 122482 140106 122656
rect 136961 122480 140106 122482
rect 136961 122424 136966 122480
rect 137022 122424 140106 122480
rect 136961 122422 140106 122424
rect 136961 122419 137027 122422
rect 100989 122346 101055 122349
rect 97726 122344 101055 122346
rect 97726 122288 100994 122344
rect 101050 122288 101055 122344
rect 97726 122286 101055 122288
rect 100989 122283 101055 122286
rect 102277 122346 102343 122349
rect 169854 122346 169914 122724
rect 172933 122346 172999 122349
rect 102277 122344 104932 122346
rect 102277 122288 102282 122344
rect 102338 122288 104932 122344
rect 102277 122286 104932 122288
rect 169854 122344 172999 122346
rect 169854 122288 172938 122344
rect 172994 122288 172999 122344
rect 169854 122286 172999 122288
rect 102277 122283 102343 122286
rect 172933 122283 172999 122286
rect 174037 122346 174103 122349
rect 174037 122344 177060 122346
rect 174037 122288 174042 122344
rect 174098 122288 177060 122344
rect 174037 122286 177060 122288
rect 174037 122283 174103 122286
rect 66397 122210 66463 122213
rect 100897 122210 100963 122213
rect 66397 122208 67948 122210
rect 66397 122152 66402 122208
rect 66458 122152 67948 122208
rect 66397 122150 67948 122152
rect 97756 122208 100963 122210
rect 97756 122152 100902 122208
rect 100958 122152 100963 122208
rect 97756 122150 100963 122152
rect 66397 122147 66463 122150
rect 100897 122147 100963 122150
rect 137053 122210 137119 122213
rect 137053 122208 140076 122210
rect 137053 122152 137058 122208
rect 137114 122152 140076 122208
rect 137053 122150 140076 122152
rect 137053 122147 137119 122150
rect 169854 122074 169914 122180
rect 172657 122074 172723 122077
rect 169854 122072 172723 122074
rect 169854 122016 172662 122072
rect 172718 122016 172723 122072
rect 169854 122014 172723 122016
rect 172657 122011 172723 122014
rect 135397 121938 135463 121941
rect 132686 121936 135463 121938
rect 132686 121880 135402 121936
rect 135458 121880 135463 121936
rect 132686 121878 135463 121880
rect 132686 121704 132746 121878
rect 135397 121875 135463 121878
rect 63545 121666 63611 121669
rect 60772 121664 63611 121666
rect 60772 121608 63550 121664
rect 63606 121608 63611 121664
rect 60772 121606 63611 121608
rect 63545 121603 63611 121606
rect 102185 121666 102251 121669
rect 174313 121666 174379 121669
rect 102185 121664 104932 121666
rect 102185 121608 102190 121664
rect 102246 121608 104932 121664
rect 102185 121606 104932 121608
rect 174313 121664 177060 121666
rect 174313 121608 174318 121664
rect 174374 121608 177060 121664
rect 174313 121606 177060 121608
rect 102185 121603 102251 121606
rect 174313 121603 174379 121606
rect 62809 121394 62875 121397
rect 60742 121392 62875 121394
rect 60742 121336 62814 121392
rect 62870 121336 62875 121392
rect 60742 121334 62875 121336
rect 60742 121160 60802 121334
rect 62809 121331 62875 121334
rect 67918 121122 67978 121500
rect 66078 121062 67978 121122
rect 97726 121122 97786 121432
rect 135305 121394 135371 121397
rect 132686 121392 135371 121394
rect 132686 121336 135310 121392
rect 135366 121336 135371 121392
rect 132686 121334 135371 121336
rect 132686 121160 132746 121334
rect 135305 121331 135371 121334
rect 100621 121122 100687 121125
rect 97726 121120 100687 121122
rect 97726 121064 100626 121120
rect 100682 121064 100687 121120
rect 97726 121062 100687 121064
rect 65017 120714 65083 120717
rect 66078 120714 66138 121062
rect 100621 121059 100687 121062
rect 102277 121122 102343 121125
rect 136777 121122 136843 121125
rect 140046 121122 140106 121432
rect 102277 121120 104932 121122
rect 102277 121064 102282 121120
rect 102338 121064 104932 121120
rect 102277 121062 104932 121064
rect 136777 121120 140106 121122
rect 136777 121064 136782 121120
rect 136838 121064 140106 121120
rect 136777 121062 140106 121064
rect 169854 121122 169914 121500
rect 171737 121122 171803 121125
rect 169854 121120 171803 121122
rect 169854 121064 171742 121120
rect 171798 121064 171803 121120
rect 169854 121062 171803 121064
rect 102277 121059 102343 121062
rect 136777 121059 136843 121062
rect 171737 121059 171803 121062
rect 174129 121122 174195 121125
rect 174129 121120 177060 121122
rect 174129 121064 174134 121120
rect 174190 121064 177060 121120
rect 174129 121062 177060 121064
rect 174129 121059 174195 121062
rect 66213 120986 66279 120989
rect 66213 120984 67948 120986
rect 66213 120928 66218 120984
rect 66274 120928 67948 120984
rect 66213 120926 67948 120928
rect 66213 120923 66279 120926
rect 65017 120712 66138 120714
rect 65017 120656 65022 120712
rect 65078 120656 66138 120712
rect 65017 120654 66138 120656
rect 97726 120714 97786 120888
rect 100621 120714 100687 120717
rect 97726 120712 100687 120714
rect 97726 120656 100626 120712
rect 100682 120656 100687 120712
rect 97726 120654 100687 120656
rect 65017 120651 65083 120654
rect 100621 120651 100687 120654
rect 136869 120714 136935 120717
rect 140046 120714 140106 120888
rect 136869 120712 140106 120714
rect 136869 120656 136874 120712
rect 136930 120656 140106 120712
rect 136869 120654 140106 120656
rect 169854 120714 169914 120956
rect 172657 120714 172723 120717
rect 169854 120712 172723 120714
rect 169854 120656 172662 120712
rect 172718 120656 172723 120712
rect 169854 120654 172723 120656
rect 136869 120651 136935 120654
rect 172657 120651 172723 120654
rect 63453 120578 63519 120581
rect 60772 120576 63519 120578
rect 60772 120520 63458 120576
rect 63514 120520 63519 120576
rect 60772 120518 63519 120520
rect 63453 120515 63519 120518
rect 102369 120578 102435 120581
rect 135213 120578 135279 120581
rect 102369 120576 104932 120578
rect 102369 120520 102374 120576
rect 102430 120520 104932 120576
rect 102369 120518 104932 120520
rect 132716 120576 135279 120578
rect 132716 120520 135218 120576
rect 135274 120520 135279 120576
rect 132716 120518 135279 120520
rect 102369 120515 102435 120518
rect 135213 120515 135279 120518
rect 174129 120578 174195 120581
rect 174129 120576 177060 120578
rect 174129 120520 174134 120576
rect 174190 120520 177060 120576
rect 174129 120518 177060 120520
rect 174129 120515 174195 120518
rect 63637 120306 63703 120309
rect 135121 120306 135187 120309
rect 60742 120304 63703 120306
rect 60742 120248 63642 120304
rect 63698 120248 63703 120304
rect 132686 120304 135187 120306
rect 60742 120246 63703 120248
rect 60742 119936 60802 120246
rect 63637 120243 63703 120246
rect 67918 119898 67978 120276
rect 132686 120248 135126 120304
rect 135182 120248 135187 120304
rect 132686 120246 135187 120248
rect 66262 119838 67978 119898
rect 97726 119898 97786 120208
rect 132686 119936 132746 120246
rect 135121 120243 135187 120246
rect 100621 119898 100687 119901
rect 97726 119896 100687 119898
rect 97726 119840 100626 119896
rect 100682 119840 100687 119896
rect 97726 119838 100687 119840
rect 62809 119626 62875 119629
rect 60742 119624 62875 119626
rect 60742 119568 62814 119624
rect 62870 119568 62875 119624
rect 60742 119566 62875 119568
rect 60742 119392 60802 119566
rect 62809 119563 62875 119566
rect 65017 119490 65083 119493
rect 66262 119490 66322 119838
rect 100621 119835 100687 119838
rect 102093 119898 102159 119901
rect 136777 119898 136843 119901
rect 140046 119898 140106 120208
rect 102093 119896 104932 119898
rect 102093 119840 102098 119896
rect 102154 119840 104932 119896
rect 102093 119838 104932 119840
rect 136777 119896 140106 119898
rect 136777 119840 136782 119896
rect 136838 119840 140106 119896
rect 136777 119838 140106 119840
rect 169854 119898 169914 120276
rect 172657 119898 172723 119901
rect 169854 119896 172723 119898
rect 169854 119840 172662 119896
rect 172718 119840 172723 119896
rect 169854 119838 172723 119840
rect 102093 119835 102159 119838
rect 136777 119835 136843 119838
rect 172657 119835 172723 119838
rect 174313 119898 174379 119901
rect 174313 119896 177060 119898
rect 174313 119840 174318 119896
rect 174374 119840 177060 119896
rect 174313 119838 177060 119840
rect 174313 119835 174379 119838
rect 66397 119762 66463 119765
rect 66397 119760 67948 119762
rect 66397 119704 66402 119760
rect 66458 119704 67948 119760
rect 66397 119702 67948 119704
rect 66397 119699 66463 119702
rect 65017 119488 66322 119490
rect 65017 119432 65022 119488
rect 65078 119432 66322 119488
rect 65017 119430 66322 119432
rect 65017 119427 65083 119430
rect 97726 119354 97786 119664
rect 102277 119626 102343 119629
rect 134845 119626 134911 119629
rect 102277 119624 104962 119626
rect 102277 119568 102282 119624
rect 102338 119568 104962 119624
rect 102277 119566 104962 119568
rect 102277 119563 102343 119566
rect 100897 119354 100963 119357
rect 97726 119352 100963 119354
rect 97726 119296 100902 119352
rect 100958 119296 100963 119352
rect 104902 119324 104962 119566
rect 132686 119624 134911 119626
rect 132686 119568 134850 119624
rect 134906 119568 134911 119624
rect 132686 119566 134911 119568
rect 132686 119392 132746 119566
rect 134845 119563 134911 119566
rect 136961 119354 137027 119357
rect 140046 119354 140106 119664
rect 136961 119352 140106 119354
rect 97726 119294 100963 119296
rect 100897 119291 100963 119294
rect 136961 119296 136966 119352
rect 137022 119296 140106 119352
rect 136961 119294 140106 119296
rect 169854 119354 169914 119732
rect 172657 119354 172723 119357
rect 169854 119352 172723 119354
rect 169854 119296 172662 119352
rect 172718 119296 172723 119352
rect 169854 119294 172723 119296
rect 136961 119291 137027 119294
rect 172657 119291 172723 119294
rect 174129 119354 174195 119357
rect 174129 119352 177060 119354
rect 174129 119296 174134 119352
rect 174190 119296 177060 119352
rect 174129 119294 177060 119296
rect 174129 119291 174195 119294
rect 66397 119218 66463 119221
rect 66397 119216 67948 119218
rect 66397 119160 66402 119216
rect 66458 119160 67948 119216
rect 66397 119158 67948 119160
rect 66397 119155 66463 119158
rect 62717 118810 62783 118813
rect 60772 118808 62783 118810
rect 60772 118752 62722 118808
rect 62778 118752 62783 118808
rect 60772 118750 62783 118752
rect 62717 118747 62783 118750
rect 97726 118674 97786 119120
rect 135305 119082 135371 119085
rect 132686 119080 135371 119082
rect 132686 119024 135310 119080
rect 135366 119024 135371 119080
rect 132686 119022 135371 119024
rect 132686 118848 132746 119022
rect 135305 119019 135371 119022
rect 102185 118810 102251 118813
rect 102185 118808 104932 118810
rect 102185 118752 102190 118808
rect 102246 118752 104932 118808
rect 102185 118750 104932 118752
rect 102185 118747 102251 118750
rect 100621 118674 100687 118677
rect 97726 118672 100687 118674
rect 97726 118616 100626 118672
rect 100682 118616 100687 118672
rect 97726 118614 100687 118616
rect 100621 118611 100687 118614
rect 136961 118674 137027 118677
rect 140046 118674 140106 119120
rect 136961 118672 140106 118674
rect 136961 118616 136966 118672
rect 137022 118616 140106 118672
rect 136961 118614 140106 118616
rect 169854 118674 169914 119188
rect 173945 118810 174011 118813
rect 173945 118808 177060 118810
rect 173945 118752 173950 118808
rect 174006 118752 177060 118808
rect 173945 118750 177060 118752
rect 173945 118747 174011 118750
rect 172013 118674 172079 118677
rect 169854 118672 172079 118674
rect 169854 118616 172018 118672
rect 172074 118616 172079 118672
rect 169854 118614 172079 118616
rect 136961 118611 137027 118614
rect 172013 118611 172079 118614
rect 31846 118476 31852 118540
rect 31916 118538 31922 118540
rect 62809 118538 62875 118541
rect 31916 118478 32988 118538
rect 60742 118536 62875 118538
rect 60742 118480 62814 118536
rect 62870 118480 62875 118536
rect 60742 118478 62875 118480
rect 31916 118476 31922 118478
rect 60742 118304 60802 118478
rect 62809 118475 62875 118478
rect 64925 118538 64991 118541
rect 135029 118538 135095 118541
rect 207893 118538 207959 118541
rect 64925 118536 67948 118538
rect 64925 118480 64930 118536
rect 64986 118480 67948 118536
rect 64925 118478 67948 118480
rect 132686 118536 135095 118538
rect 132686 118480 135034 118536
rect 135090 118480 135095 118536
rect 204844 118536 207959 118538
rect 204844 118508 207898 118536
rect 132686 118478 135095 118480
rect 64925 118475 64991 118478
rect 65017 118266 65083 118269
rect 66397 118266 66463 118269
rect 65017 118264 66463 118266
rect 65017 118208 65022 118264
rect 65078 118208 66402 118264
rect 66458 118208 66463 118264
rect 65017 118206 66463 118208
rect 65017 118203 65083 118206
rect 66397 118203 66463 118206
rect 97726 118130 97786 118440
rect 132686 118304 132746 118478
rect 135029 118475 135095 118478
rect 102277 118266 102343 118269
rect 102277 118264 104932 118266
rect 102277 118208 102282 118264
rect 102338 118208 104932 118264
rect 102277 118206 104932 118208
rect 102277 118203 102343 118206
rect 100621 118130 100687 118133
rect 97726 118128 100687 118130
rect 97726 118072 100626 118128
rect 100682 118072 100687 118128
rect 97726 118070 100687 118072
rect 100621 118067 100687 118070
rect 136777 118130 136843 118133
rect 140046 118130 140106 118440
rect 169854 118402 169914 118508
rect 204814 118480 207898 118508
rect 207954 118480 207959 118536
rect 204814 118478 207959 118480
rect 169854 118342 170282 118402
rect 170222 118130 170282 118342
rect 174037 118266 174103 118269
rect 174037 118264 177060 118266
rect 174037 118208 174042 118264
rect 174098 118208 177060 118264
rect 174037 118206 177060 118208
rect 174037 118203 174103 118206
rect 172657 118130 172723 118133
rect 136777 118128 140106 118130
rect 136777 118072 136782 118128
rect 136838 118072 140106 118128
rect 136777 118070 140106 118072
rect 169670 118070 170098 118130
rect 170222 118128 172723 118130
rect 170222 118072 172662 118128
rect 172718 118072 172723 118128
rect 170222 118070 172723 118072
rect 136777 118067 136843 118070
rect 66397 117994 66463 117997
rect 100713 117994 100779 117997
rect 66397 117992 67948 117994
rect 66397 117936 66402 117992
rect 66458 117936 67948 117992
rect 66397 117934 67948 117936
rect 97756 117992 100779 117994
rect 97756 117936 100718 117992
rect 100774 117936 100779 117992
rect 97756 117934 100779 117936
rect 66397 117931 66463 117934
rect 100713 117931 100779 117934
rect 136869 117994 136935 117997
rect 136869 117992 140076 117994
rect 136869 117936 136874 117992
rect 136930 117936 140076 117992
rect 169670 117964 169730 118070
rect 170038 117994 170098 118070
rect 172657 118067 172723 118070
rect 204814 117997 204874 118478
rect 207893 118475 207959 118478
rect 172473 117994 172539 117997
rect 170038 117992 172539 117994
rect 136869 117934 140076 117936
rect 170038 117936 172478 117992
rect 172534 117936 172539 117992
rect 170038 117934 172539 117936
rect 136869 117931 136935 117934
rect 172473 117931 172539 117934
rect 204765 117992 204874 117997
rect 204765 117936 204770 117992
rect 204826 117936 204874 117992
rect 204765 117934 204874 117936
rect 204765 117931 204831 117934
rect 62901 117858 62967 117861
rect 60742 117856 62967 117858
rect 60742 117800 62906 117856
rect 62962 117800 62967 117856
rect 60742 117798 62967 117800
rect 60742 117624 60802 117798
rect 62901 117795 62967 117798
rect 102369 117586 102435 117589
rect 135213 117586 135279 117589
rect 102369 117584 104932 117586
rect 102369 117528 102374 117584
rect 102430 117528 104932 117584
rect 102369 117526 104932 117528
rect 132716 117584 135279 117586
rect 132716 117528 135218 117584
rect 135274 117528 135279 117584
rect 132716 117526 135279 117528
rect 102369 117523 102435 117526
rect 135213 117523 135279 117526
rect 174129 117586 174195 117589
rect 174129 117584 177060 117586
rect 174129 117528 174134 117584
rect 174190 117528 177060 117584
rect 174129 117526 177060 117528
rect 174129 117523 174195 117526
rect 62809 117314 62875 117317
rect 134109 117314 134175 117317
rect 60742 117312 62875 117314
rect 60742 117256 62814 117312
rect 62870 117256 62875 117312
rect 132686 117312 134175 117314
rect 60742 117254 62875 117256
rect 60742 117080 60802 117254
rect 62809 117251 62875 117254
rect 67918 116906 67978 117284
rect 132686 117256 134114 117312
rect 134170 117256 134175 117312
rect 132686 117254 134175 117256
rect 66262 116846 67978 116906
rect 97726 116906 97786 117216
rect 132686 117080 132746 117254
rect 134109 117251 134175 117254
rect 102185 117042 102251 117045
rect 102185 117040 104932 117042
rect 102185 116984 102190 117040
rect 102246 116984 104932 117040
rect 102185 116982 104932 116984
rect 102185 116979 102251 116982
rect 100529 116906 100595 116909
rect 97726 116904 100595 116906
rect 97726 116848 100534 116904
rect 100590 116848 100595 116904
rect 97726 116846 100595 116848
rect 62809 116770 62875 116773
rect 60742 116768 62875 116770
rect 60742 116712 62814 116768
rect 62870 116712 62875 116768
rect 60742 116710 62875 116712
rect 60742 116536 60802 116710
rect 62809 116707 62875 116710
rect 65017 116498 65083 116501
rect 66262 116498 66322 116846
rect 100529 116843 100595 116846
rect 136777 116906 136843 116909
rect 140046 116906 140106 117216
rect 136777 116904 140106 116906
rect 136777 116848 136782 116904
rect 136838 116848 140106 116904
rect 136777 116846 140106 116848
rect 169854 116906 169914 117284
rect 174037 117042 174103 117045
rect 174037 117040 177060 117042
rect 174037 116984 174042 117040
rect 174098 116984 177060 117040
rect 174037 116982 177060 116984
rect 174037 116979 174103 116982
rect 172657 116906 172723 116909
rect 169854 116904 172723 116906
rect 169854 116848 172662 116904
rect 172718 116848 172723 116904
rect 169854 116846 172723 116848
rect 136777 116843 136843 116846
rect 172657 116843 172723 116846
rect 66397 116770 66463 116773
rect 100621 116770 100687 116773
rect 134661 116770 134727 116773
rect 66397 116768 67948 116770
rect 66397 116712 66402 116768
rect 66458 116712 67948 116768
rect 66397 116710 67948 116712
rect 97756 116768 100687 116770
rect 97756 116712 100626 116768
rect 100682 116712 100687 116768
rect 97756 116710 100687 116712
rect 66397 116707 66463 116710
rect 100621 116707 100687 116710
rect 132686 116768 134727 116770
rect 132686 116712 134666 116768
rect 134722 116712 134727 116768
rect 132686 116710 134727 116712
rect 132686 116536 132746 116710
rect 134661 116707 134727 116710
rect 65017 116496 66322 116498
rect 65017 116440 65022 116496
rect 65078 116440 66322 116496
rect 65017 116438 66322 116440
rect 102277 116498 102343 116501
rect 136869 116498 136935 116501
rect 140046 116498 140106 116672
rect 102277 116496 104932 116498
rect 102277 116440 102282 116496
rect 102338 116440 104932 116496
rect 102277 116438 104932 116440
rect 136869 116496 140106 116498
rect 136869 116440 136874 116496
rect 136930 116440 140106 116496
rect 136869 116438 140106 116440
rect 169854 116498 169914 116740
rect 172565 116498 172631 116501
rect 169854 116496 172631 116498
rect 169854 116440 172570 116496
rect 172626 116440 172631 116496
rect 169854 116438 172631 116440
rect 65017 116435 65083 116438
rect 102277 116435 102343 116438
rect 136869 116435 136935 116438
rect 172565 116435 172631 116438
rect 173945 116498 174011 116501
rect 173945 116496 177060 116498
rect 173945 116440 173950 116496
rect 174006 116440 177060 116496
rect 173945 116438 177060 116440
rect 173945 116435 174011 116438
rect 62717 116226 62783 116229
rect 135305 116226 135371 116229
rect 60742 116224 62783 116226
rect 60742 116168 62722 116224
rect 62778 116168 62783 116224
rect 132686 116224 135371 116226
rect 60742 116166 62783 116168
rect 60742 115856 60802 116166
rect 62717 116163 62783 116166
rect 62809 115546 62875 115549
rect 60742 115544 62875 115546
rect 60742 115488 62814 115544
rect 62870 115488 62875 115544
rect 60742 115486 62875 115488
rect 60742 115312 60802 115486
rect 62809 115483 62875 115486
rect 65017 115138 65083 115141
rect 67918 115138 67978 116196
rect 132686 116168 135310 116224
rect 135366 116168 135371 116224
rect 132686 116166 135371 116168
rect 97726 115546 97786 116128
rect 132686 115856 132746 116166
rect 135305 116163 135371 116166
rect 102461 115818 102527 115821
rect 102461 115816 104932 115818
rect 102461 115760 102466 115816
rect 102522 115760 104932 115816
rect 102461 115758 104932 115760
rect 102461 115755 102527 115758
rect 100621 115546 100687 115549
rect 134477 115546 134543 115549
rect 97726 115544 100687 115546
rect 97726 115488 100626 115544
rect 100682 115488 100687 115544
rect 97726 115486 100687 115488
rect 100621 115483 100687 115486
rect 132686 115544 134543 115546
rect 132686 115488 134482 115544
rect 134538 115488 134543 115544
rect 132686 115486 134543 115488
rect 132686 115312 132746 115486
rect 134477 115483 134543 115486
rect 136777 115546 136843 115549
rect 140046 115546 140106 116128
rect 169854 115682 169914 116196
rect 222705 115954 222771 115957
rect 227416 115954 227896 115984
rect 222705 115952 227896 115954
rect 222705 115896 222710 115952
rect 222766 115896 227896 115952
rect 222705 115894 227896 115896
rect 222705 115891 222771 115894
rect 227416 115864 227896 115894
rect 174129 115818 174195 115821
rect 174129 115816 177060 115818
rect 174129 115760 174134 115816
rect 174190 115760 177060 115816
rect 174129 115758 177060 115760
rect 174129 115755 174195 115758
rect 172657 115682 172723 115685
rect 169854 115680 172723 115682
rect 169854 115624 172662 115680
rect 172718 115624 172723 115680
rect 169854 115622 172723 115624
rect 172657 115619 172723 115622
rect 136777 115544 140106 115546
rect 136777 115488 136782 115544
rect 136838 115488 140106 115544
rect 136777 115486 140106 115488
rect 136777 115483 136843 115486
rect 102369 115274 102435 115277
rect 174221 115274 174287 115277
rect 102369 115272 104932 115274
rect 102369 115216 102374 115272
rect 102430 115216 104932 115272
rect 102369 115214 104932 115216
rect 174221 115272 177060 115274
rect 174221 115216 174226 115272
rect 174282 115216 177060 115272
rect 174221 115214 177060 115216
rect 102369 115211 102435 115214
rect 174221 115211 174287 115214
rect 65017 115136 67978 115138
rect 65017 115080 65022 115136
rect 65078 115080 67978 115136
rect 65017 115078 67978 115080
rect 65017 115075 65083 115078
rect 135305 115002 135371 115005
rect 132686 115000 135371 115002
rect 132686 114944 135310 115000
rect 135366 114944 135371 115000
rect 132686 114942 135371 114944
rect 132686 114768 132746 114942
rect 135305 114939 135371 114942
rect 62809 114730 62875 114733
rect 60772 114728 62875 114730
rect 60772 114672 62814 114728
rect 62870 114672 62875 114728
rect 60772 114670 62875 114672
rect 62809 114667 62875 114670
rect 102185 114730 102251 114733
rect 173853 114730 173919 114733
rect 102185 114728 104932 114730
rect 102185 114672 102190 114728
rect 102246 114672 104932 114728
rect 102185 114670 104932 114672
rect 173853 114728 177060 114730
rect 173853 114672 173858 114728
rect 173914 114672 177060 114728
rect 173853 114670 177060 114672
rect 102185 114667 102251 114670
rect 173853 114667 173919 114670
rect 62809 114458 62875 114461
rect 134845 114458 134911 114461
rect 60742 114456 62875 114458
rect 60742 114400 62814 114456
rect 62870 114400 62875 114456
rect 60742 114398 62875 114400
rect 60742 114224 60802 114398
rect 62809 114395 62875 114398
rect 132686 114456 134911 114458
rect 132686 114400 134850 114456
rect 134906 114400 134911 114456
rect 132686 114398 134911 114400
rect 132686 114224 132746 114398
rect 134845 114395 134911 114398
rect 102277 114186 102343 114189
rect 174037 114186 174103 114189
rect 102277 114184 104932 114186
rect 102277 114128 102282 114184
rect 102338 114128 104932 114184
rect 102277 114126 104932 114128
rect 174037 114184 177060 114186
rect 174037 114128 174042 114184
rect 174098 114128 177060 114184
rect 174037 114126 177060 114128
rect 102277 114123 102343 114126
rect 174037 114123 174103 114126
rect 71038 113580 71044 113644
rect 71108 113642 71114 113644
rect 72837 113642 72903 113645
rect 71108 113640 72903 113642
rect 71108 113584 72842 113640
rect 72898 113584 72903 113640
rect 71108 113582 72903 113584
rect 71108 113580 71114 113582
rect 72837 113579 72903 113582
rect 142982 113580 142988 113644
rect 143052 113642 143058 113644
rect 144873 113642 144939 113645
rect 143052 113640 144939 113642
rect 143052 113584 144878 113640
rect 144934 113584 144939 113640
rect 143052 113582 144939 113584
rect 143052 113580 143058 113582
rect 144873 113579 144939 113582
rect 164837 113642 164903 113645
rect 167270 113642 167276 113644
rect 164837 113640 167276 113642
rect 164837 113584 164842 113640
rect 164898 113584 167276 113640
rect 164837 113582 167276 113584
rect 164837 113579 164903 113582
rect 167270 113580 167276 113582
rect 167340 113580 167346 113644
rect 56921 113236 56987 113237
rect 56870 113172 56876 113236
rect 56940 113234 56987 113236
rect 56940 113232 57032 113234
rect 56982 113176 57032 113232
rect 56940 113174 57032 113176
rect 56940 113172 56987 113174
rect 73062 113172 73068 113236
rect 73132 113234 73138 113236
rect 73205 113234 73271 113237
rect 73132 113232 73271 113234
rect 73132 113176 73210 113232
rect 73266 113176 73271 113232
rect 73132 113174 73271 113176
rect 73132 113172 73138 113174
rect 56921 113171 56987 113172
rect 73205 113171 73271 113174
rect 92801 112690 92867 112693
rect 94222 112690 94228 112692
rect 92801 112688 94228 112690
rect 92801 112632 92806 112688
rect 92862 112632 94228 112688
rect 92801 112630 94228 112632
rect 92801 112627 92867 112630
rect 94222 112628 94228 112630
rect 94292 112628 94298 112692
rect 105957 110242 106023 110245
rect 177717 110242 177783 110245
rect 102724 110240 106023 110242
rect 102724 110184 105962 110240
rect 106018 110184 106023 110240
rect 102724 110182 106023 110184
rect 174852 110240 177783 110242
rect 174852 110184 177722 110240
rect 177778 110184 177783 110240
rect 174852 110182 177783 110184
rect 105957 110179 106023 110182
rect 177717 110179 177783 110182
rect 108625 109562 108691 109565
rect 180293 109562 180359 109565
rect 108625 109560 111004 109562
rect 108625 109504 108630 109560
rect 108686 109504 111004 109560
rect 108625 109502 111004 109504
rect 180293 109560 182948 109562
rect 180293 109504 180298 109560
rect 180354 109504 182948 109560
rect 180293 109502 182948 109504
rect 108625 109499 108691 109502
rect 180293 109499 180359 109502
rect 105773 109018 105839 109021
rect 177349 109018 177415 109021
rect 102724 109016 105839 109018
rect 102724 108960 105778 109016
rect 105834 108960 105839 109016
rect 102724 108958 105839 108960
rect 174852 109016 177415 109018
rect 174852 108960 177354 109016
rect 177410 108960 177415 109016
rect 174852 108958 177415 108960
rect 105773 108955 105839 108958
rect 177349 108955 177415 108958
rect 105681 107794 105747 107797
rect 176981 107794 177047 107797
rect 102724 107792 105747 107794
rect 102724 107736 105686 107792
rect 105742 107736 105747 107792
rect 102724 107734 105747 107736
rect 174852 107792 177047 107794
rect 174852 107736 176986 107792
rect 177042 107736 177047 107792
rect 174852 107734 177047 107736
rect 105681 107731 105747 107734
rect 176981 107731 177047 107734
rect 108533 107250 108599 107253
rect 180385 107250 180451 107253
rect 108533 107248 111004 107250
rect 108533 107192 108538 107248
rect 108594 107192 111004 107248
rect 108533 107190 111004 107192
rect 180385 107248 182948 107250
rect 180385 107192 180390 107248
rect 180446 107192 182948 107248
rect 180385 107190 182948 107192
rect 108533 107187 108599 107190
rect 180385 107187 180451 107190
rect 105497 106570 105563 106573
rect 176889 106570 176955 106573
rect 102724 106568 105563 106570
rect 102724 106512 105502 106568
rect 105558 106512 105563 106568
rect 102724 106510 105563 106512
rect 174852 106568 176955 106570
rect 174852 106512 176894 106568
rect 176950 106512 176955 106568
rect 174852 106510 176955 106512
rect 105497 106507 105563 106510
rect 176889 106507 176955 106510
rect 9896 106162 10376 106192
rect 12209 106162 12275 106165
rect 9896 106160 12275 106162
rect 9896 106104 12214 106160
rect 12270 106104 12275 106160
rect 9896 106102 12275 106104
rect 9896 106072 10376 106102
rect 12209 106099 12275 106102
rect 11933 105754 11999 105757
rect 224453 105754 224519 105757
rect 11933 105752 14036 105754
rect 11933 105696 11938 105752
rect 11994 105696 14036 105752
rect 11933 105694 14036 105696
rect 223796 105752 224519 105754
rect 223796 105696 224458 105752
rect 224514 105696 224519 105752
rect 223796 105694 224519 105696
rect 11933 105691 11999 105694
rect 224453 105691 224519 105694
rect 105221 105346 105287 105349
rect 177073 105346 177139 105349
rect 102724 105344 105287 105346
rect 102724 105288 105226 105344
rect 105282 105288 105287 105344
rect 102724 105286 105287 105288
rect 174852 105344 177139 105346
rect 174852 105288 177078 105344
rect 177134 105288 177139 105344
rect 174852 105286 177139 105288
rect 105221 105283 105287 105286
rect 177073 105283 177139 105286
rect 107889 104938 107955 104941
rect 179649 104938 179715 104941
rect 107889 104936 111004 104938
rect 107889 104880 107894 104936
rect 107950 104880 111004 104936
rect 107889 104878 111004 104880
rect 179649 104936 182948 104938
rect 179649 104880 179654 104936
rect 179710 104880 182948 104936
rect 179649 104878 182948 104880
rect 107889 104875 107955 104878
rect 179649 104875 179715 104878
rect 31989 104258 32055 104261
rect 29860 104256 32055 104258
rect 29860 104200 31994 104256
rect 32050 104200 32055 104256
rect 29860 104198 32055 104200
rect 31989 104195 32055 104198
rect 37417 104258 37483 104261
rect 60509 104258 60575 104261
rect 201085 104258 201151 104261
rect 37417 104256 39060 104258
rect 37417 104200 37422 104256
rect 37478 104200 39060 104256
rect 37417 104198 39060 104200
rect 60509 104256 62980 104258
rect 60509 104200 60514 104256
rect 60570 104200 62980 104256
rect 60509 104198 62980 104200
rect 126828 104198 134924 104258
rect 198772 104256 201151 104258
rect 198772 104200 201090 104256
rect 201146 104200 201151 104256
rect 198772 104198 201151 104200
rect 37417 104195 37483 104198
rect 60509 104195 60575 104198
rect 201085 104195 201151 104198
rect 204673 104258 204739 104261
rect 204673 104256 207972 104258
rect 204673 104200 204678 104256
rect 204734 104200 207972 104256
rect 204673 104198 207972 104200
rect 204673 104195 204739 104198
rect 106141 104122 106207 104125
rect 177257 104122 177323 104125
rect 102724 104120 106207 104122
rect 102724 104064 106146 104120
rect 106202 104064 106207 104120
rect 102724 104062 106207 104064
rect 174852 104120 177323 104122
rect 174852 104064 177262 104120
rect 177318 104064 177323 104120
rect 174852 104062 177323 104064
rect 106141 104059 106207 104062
rect 177257 104059 177323 104062
rect 105589 102898 105655 102901
rect 177533 102898 177599 102901
rect 102724 102896 105655 102898
rect 102724 102840 105594 102896
rect 105650 102840 105655 102896
rect 102724 102838 105655 102840
rect 174852 102896 177599 102898
rect 174852 102840 177538 102896
rect 177594 102840 177599 102896
rect 174852 102838 177599 102840
rect 105589 102835 105655 102838
rect 177533 102835 177599 102838
rect 107889 102490 107955 102493
rect 179649 102490 179715 102493
rect 107889 102488 111004 102490
rect 107889 102432 107894 102488
rect 107950 102432 111004 102488
rect 107889 102430 111004 102432
rect 179649 102488 182948 102490
rect 179649 102432 179654 102488
rect 179710 102432 182948 102488
rect 179649 102430 182948 102432
rect 107889 102427 107955 102430
rect 179649 102427 179715 102430
rect 105129 101674 105195 101677
rect 176889 101674 176955 101677
rect 102724 101672 105195 101674
rect 102724 101616 105134 101672
rect 105190 101616 105195 101672
rect 102724 101614 105195 101616
rect 174852 101672 176955 101674
rect 174852 101616 176894 101672
rect 176950 101616 176955 101672
rect 174852 101614 176955 101616
rect 105129 101611 105195 101614
rect 176889 101611 176955 101614
rect 57565 100858 57631 100861
rect 54884 100856 57631 100858
rect 54884 100800 57570 100856
rect 57626 100800 57631 100856
rect 54884 100798 57631 100800
rect 57565 100795 57631 100798
rect 105957 100450 106023 100453
rect 176981 100450 177047 100453
rect 102724 100448 106023 100450
rect 102724 100392 105962 100448
rect 106018 100392 106023 100448
rect 102724 100390 106023 100392
rect 174852 100448 177047 100450
rect 174852 100392 176986 100448
rect 177042 100392 177047 100448
rect 174852 100390 177047 100392
rect 105957 100387 106023 100390
rect 176981 100387 177047 100390
rect 107889 100178 107955 100181
rect 179649 100178 179715 100181
rect 107889 100176 111004 100178
rect 107889 100120 107894 100176
rect 107950 100120 111004 100176
rect 107889 100118 111004 100120
rect 179649 100176 182948 100178
rect 179649 100120 179654 100176
rect 179710 100120 182948 100176
rect 179649 100118 182948 100120
rect 107889 100115 107955 100118
rect 179649 100115 179715 100118
rect 105589 99226 105655 99229
rect 177349 99226 177415 99229
rect 102724 99224 105655 99226
rect 102724 99168 105594 99224
rect 105650 99168 105655 99224
rect 102724 99166 105655 99168
rect 174852 99224 177415 99226
rect 174852 99168 177354 99224
rect 177410 99168 177415 99224
rect 174852 99166 177415 99168
rect 105589 99163 105655 99166
rect 177349 99163 177415 99166
rect 105681 98138 105747 98141
rect 178177 98138 178243 98141
rect 102724 98136 105747 98138
rect 102724 98080 105686 98136
rect 105742 98080 105747 98136
rect 102724 98078 105747 98080
rect 174852 98136 178243 98138
rect 174852 98080 178182 98136
rect 178238 98080 178243 98136
rect 174852 98078 178243 98080
rect 105681 98075 105747 98078
rect 178177 98075 178243 98078
rect 107889 97866 107955 97869
rect 179649 97866 179715 97869
rect 107889 97864 111004 97866
rect 107889 97808 107894 97864
rect 107950 97808 111004 97864
rect 107889 97806 111004 97808
rect 179649 97864 182948 97866
rect 179649 97808 179654 97864
rect 179710 97808 182948 97864
rect 179649 97806 182948 97808
rect 107889 97803 107955 97806
rect 179649 97803 179715 97806
rect 106325 96914 106391 96917
rect 177625 96914 177691 96917
rect 102724 96912 106391 96914
rect 102724 96856 106330 96912
rect 106386 96856 106391 96912
rect 102724 96854 106391 96856
rect 174852 96912 177691 96914
rect 174852 96856 177630 96912
rect 177686 96856 177691 96912
rect 174852 96854 177691 96856
rect 106325 96851 106391 96854
rect 177625 96851 177691 96854
rect 223533 96370 223599 96373
rect 223533 96368 223642 96370
rect 223533 96312 223538 96368
rect 223594 96312 223642 96368
rect 223533 96307 223642 96312
rect 12117 95826 12183 95829
rect 132361 95826 132427 95829
rect 132545 95826 132611 95829
rect 12117 95824 14036 95826
rect 12117 95768 12122 95824
rect 12178 95768 14036 95824
rect 12117 95766 14036 95768
rect 132361 95824 132611 95826
rect 132361 95768 132366 95824
rect 132422 95768 132550 95824
rect 132606 95768 132611 95824
rect 223582 95796 223642 96307
rect 132361 95766 132611 95768
rect 12117 95763 12183 95766
rect 132361 95763 132427 95766
rect 132545 95763 132611 95766
rect 106417 95690 106483 95693
rect 177717 95690 177783 95693
rect 102724 95688 106483 95690
rect 102724 95632 106422 95688
rect 106478 95632 106483 95688
rect 102724 95630 106483 95632
rect 174852 95688 177783 95690
rect 174852 95632 177722 95688
rect 177778 95632 177783 95688
rect 174852 95630 177783 95632
rect 106417 95627 106483 95630
rect 177717 95627 177783 95630
rect 107797 95418 107863 95421
rect 179557 95418 179623 95421
rect 107797 95416 111004 95418
rect 107797 95360 107802 95416
rect 107858 95360 111004 95416
rect 107797 95358 111004 95360
rect 179557 95416 182948 95418
rect 179557 95360 179562 95416
rect 179618 95360 182948 95416
rect 179557 95358 182948 95360
rect 107797 95355 107863 95358
rect 179557 95355 179623 95358
rect 105773 94466 105839 94469
rect 177533 94466 177599 94469
rect 102724 94464 105839 94466
rect 102724 94408 105778 94464
rect 105834 94408 105839 94464
rect 102724 94406 105839 94408
rect 174852 94464 177599 94466
rect 174852 94408 177538 94464
rect 177594 94408 177599 94464
rect 174852 94406 177599 94408
rect 105773 94403 105839 94406
rect 177533 94403 177599 94406
rect 105773 93242 105839 93245
rect 177349 93242 177415 93245
rect 102724 93240 105839 93242
rect 102724 93184 105778 93240
rect 105834 93184 105839 93240
rect 102724 93182 105839 93184
rect 174852 93240 177415 93242
rect 174852 93184 177354 93240
rect 177410 93184 177415 93240
rect 174852 93182 177415 93184
rect 105773 93179 105839 93182
rect 177349 93179 177415 93182
rect 107797 93106 107863 93109
rect 179557 93106 179623 93109
rect 107797 93104 111004 93106
rect 107797 93048 107802 93104
rect 107858 93048 111004 93104
rect 107797 93046 111004 93048
rect 179557 93104 182948 93106
rect 179557 93048 179562 93104
rect 179618 93048 182948 93104
rect 179557 93046 182948 93048
rect 107797 93043 107863 93046
rect 179557 93043 179623 93046
rect 223533 92154 223599 92157
rect 227416 92154 227896 92184
rect 223533 92152 227896 92154
rect 223533 92096 223538 92152
rect 223594 92096 227896 92152
rect 223533 92094 227896 92096
rect 223533 92091 223599 92094
rect 227416 92064 227896 92094
rect 105221 92018 105287 92021
rect 176981 92018 177047 92021
rect 102724 92016 105287 92018
rect 102724 91960 105226 92016
rect 105282 91960 105287 92016
rect 102724 91958 105287 91960
rect 174852 92016 177047 92018
rect 174852 91960 176986 92016
rect 177042 91960 177047 92016
rect 174852 91958 177047 91960
rect 105221 91955 105287 91958
rect 176981 91955 177047 91958
rect 32633 90930 32699 90933
rect 29860 90928 32699 90930
rect 29860 90872 32638 90928
rect 32694 90872 32699 90928
rect 29860 90870 32699 90872
rect 32633 90867 32699 90870
rect 36405 90930 36471 90933
rect 59589 90930 59655 90933
rect 200993 90930 201059 90933
rect 36405 90928 39060 90930
rect 36405 90872 36410 90928
rect 36466 90872 39060 90928
rect 36405 90870 39060 90872
rect 59589 90928 62980 90930
rect 59589 90872 59594 90928
rect 59650 90872 62980 90928
rect 59589 90870 62980 90872
rect 126828 90870 134924 90930
rect 198772 90928 201059 90930
rect 198772 90872 200998 90928
rect 201054 90872 201059 90928
rect 198772 90870 201059 90872
rect 36405 90867 36471 90870
rect 59589 90867 59655 90870
rect 200993 90867 201059 90870
rect 204489 90930 204555 90933
rect 204489 90928 207972 90930
rect 204489 90872 204494 90928
rect 204550 90872 207972 90928
rect 204489 90870 207972 90872
rect 204489 90867 204555 90870
rect 102724 90734 111004 90794
rect 174852 90734 182948 90794
rect 102694 89298 102754 89472
rect 105773 89298 105839 89301
rect 102694 89296 105839 89298
rect 102694 89240 105778 89296
rect 105834 89240 105839 89296
rect 102694 89238 105839 89240
rect 105773 89235 105839 89238
rect 174822 89026 174882 89540
rect 174822 88966 178378 89026
rect 178318 88890 178378 88966
rect 178318 88830 182978 88890
rect 107797 88482 107863 88485
rect 107797 88480 111004 88482
rect 107797 88424 107802 88480
rect 107858 88424 111004 88480
rect 182918 88452 182978 88830
rect 107797 88422 111004 88424
rect 107797 88419 107863 88422
rect 177349 88346 177415 88349
rect 174852 88344 177415 88346
rect 174852 88288 177354 88344
rect 177410 88288 177415 88344
rect 174852 88286 177415 88288
rect 177349 88283 177415 88286
rect 102694 87938 102754 88248
rect 105405 87938 105471 87941
rect 102694 87936 105471 87938
rect 102694 87880 105410 87936
rect 105466 87880 105471 87936
rect 102694 87878 105471 87880
rect 105405 87875 105471 87878
rect 177533 87122 177599 87125
rect 174852 87120 177599 87122
rect 174852 87064 177538 87120
rect 177594 87064 177599 87120
rect 174852 87062 177599 87064
rect 177533 87059 177599 87062
rect 102694 86578 102754 87024
rect 106417 86578 106483 86581
rect 102694 86576 106483 86578
rect 102694 86520 106422 86576
rect 106478 86520 106483 86576
rect 102694 86518 106483 86520
rect 106417 86515 106483 86518
rect 107889 86034 107955 86037
rect 179649 86034 179715 86037
rect 107889 86032 111004 86034
rect 107889 85976 107894 86032
rect 107950 85976 111004 86032
rect 107889 85974 111004 85976
rect 179649 86032 182948 86034
rect 179649 85976 179654 86032
rect 179710 85976 182948 86032
rect 179649 85974 182948 85976
rect 107889 85971 107955 85974
rect 179649 85971 179715 85974
rect 176981 85898 177047 85901
rect 174852 85896 177047 85898
rect 174852 85840 176986 85896
rect 177042 85840 177047 85896
rect 174852 85838 177047 85840
rect 176981 85835 177047 85838
rect 14006 84810 14066 85664
rect 102694 85354 102754 85800
rect 105129 85354 105195 85357
rect 102694 85352 105195 85354
rect 102694 85296 105134 85352
rect 105190 85296 105195 85352
rect 102694 85294 105195 85296
rect 105129 85291 105195 85294
rect 223582 85221 223642 85732
rect 223533 85216 223642 85221
rect 223533 85160 223538 85216
rect 223594 85160 223642 85216
rect 223533 85158 223642 85160
rect 223533 85155 223599 85158
rect 105681 84810 105747 84813
rect 178177 84810 178243 84813
rect 11982 84750 14066 84810
rect 102724 84808 105747 84810
rect 102724 84752 105686 84808
rect 105742 84752 105747 84808
rect 102724 84750 105747 84752
rect 174852 84808 178243 84810
rect 174852 84752 178182 84808
rect 178238 84752 178243 84808
rect 174852 84750 178243 84752
rect 9896 84538 10376 84568
rect 11982 84538 12042 84750
rect 105681 84747 105747 84750
rect 178177 84747 178243 84750
rect 9896 84478 12042 84538
rect 9896 84448 10376 84478
rect 107981 83722 108047 83725
rect 179741 83722 179807 83725
rect 107981 83720 111004 83722
rect 107981 83664 107986 83720
rect 108042 83664 111004 83720
rect 107981 83662 111004 83664
rect 179741 83720 182948 83722
rect 179741 83664 179746 83720
rect 179802 83664 182948 83720
rect 179741 83662 182948 83664
rect 107981 83659 108047 83662
rect 179741 83659 179807 83662
rect 178085 83586 178151 83589
rect 174852 83584 178151 83586
rect 174852 83528 178090 83584
rect 178146 83528 178151 83584
rect 174852 83526 178151 83528
rect 178085 83523 178151 83526
rect 102724 83458 103122 83518
rect 103062 83450 103122 83458
rect 105221 83450 105287 83453
rect 103062 83448 105287 83450
rect 103062 83392 105226 83448
rect 105282 83392 105287 83448
rect 103062 83390 105287 83392
rect 105221 83387 105287 83390
rect 177717 82362 177783 82365
rect 174852 82360 177783 82362
rect 174852 82304 177722 82360
rect 177778 82304 177783 82360
rect 174852 82302 177783 82304
rect 177717 82299 177783 82302
rect 102724 82234 103122 82294
rect 103062 82226 103122 82234
rect 106417 82226 106483 82229
rect 103062 82224 106483 82226
rect 103062 82168 106422 82224
rect 106478 82168 106483 82224
rect 103062 82166 106483 82168
rect 106417 82163 106483 82166
rect 56921 81954 56987 81957
rect 57473 81954 57539 81957
rect 56921 81952 57539 81954
rect 56921 81896 56926 81952
rect 56982 81896 57478 81952
rect 57534 81896 57539 81952
rect 56921 81894 57539 81896
rect 56921 81891 56987 81894
rect 57473 81891 57539 81894
rect 107797 81410 107863 81413
rect 179557 81410 179623 81413
rect 107797 81408 111004 81410
rect 107797 81352 107802 81408
rect 107858 81352 111004 81408
rect 107797 81350 111004 81352
rect 179557 81408 182948 81410
rect 179557 81352 179562 81408
rect 179618 81352 182948 81408
rect 179557 81350 182948 81352
rect 107797 81347 107863 81350
rect 179557 81347 179623 81350
rect 178085 81138 178151 81141
rect 174852 81136 178151 81138
rect 174852 81080 178090 81136
rect 178146 81080 178151 81136
rect 174852 81078 178151 81080
rect 178085 81075 178151 81078
rect 57473 80866 57539 80869
rect 54884 80864 57539 80866
rect 54884 80808 57478 80864
rect 57534 80808 57539 80864
rect 54884 80806 57539 80808
rect 102694 80866 102754 81040
rect 105957 80866 106023 80869
rect 102694 80864 106023 80866
rect 102694 80808 105962 80864
rect 106018 80808 106023 80864
rect 102694 80806 106023 80808
rect 57473 80803 57539 80806
rect 105957 80803 106023 80806
rect 177625 79914 177691 79917
rect 174852 79912 177691 79914
rect 174852 79856 177630 79912
rect 177686 79856 177691 79912
rect 174852 79854 177691 79856
rect 177625 79851 177691 79854
rect 102694 79642 102754 79816
rect 105405 79642 105471 79645
rect 102694 79640 105471 79642
rect 102694 79584 105410 79640
rect 105466 79584 105471 79640
rect 102694 79582 105471 79584
rect 105405 79579 105471 79582
rect 107613 78962 107679 78965
rect 179649 78962 179715 78965
rect 107613 78960 111004 78962
rect 107613 78904 107618 78960
rect 107674 78904 111004 78960
rect 107613 78902 111004 78904
rect 179649 78960 182948 78962
rect 179649 78904 179654 78960
rect 179710 78904 182948 78960
rect 179649 78902 182948 78904
rect 107613 78899 107679 78902
rect 179649 78899 179715 78902
rect 176981 78690 177047 78693
rect 174852 78688 177047 78690
rect 174852 78632 176986 78688
rect 177042 78632 177047 78688
rect 174852 78630 177047 78632
rect 176981 78627 177047 78630
rect 102694 78010 102754 78592
rect 105221 78010 105287 78013
rect 102694 78008 105287 78010
rect 102694 77952 105226 78008
rect 105282 77952 105287 78008
rect 102694 77950 105287 77952
rect 105221 77947 105287 77950
rect 31989 77602 32055 77605
rect 29860 77600 32055 77602
rect 29860 77544 31994 77600
rect 32050 77544 32055 77600
rect 29860 77542 32055 77544
rect 31989 77539 32055 77542
rect 37417 77602 37483 77605
rect 59589 77602 59655 77605
rect 129734 77602 129740 77604
rect 37417 77600 39060 77602
rect 37417 77544 37422 77600
rect 37478 77544 39060 77600
rect 37417 77542 39060 77544
rect 59589 77600 62980 77602
rect 59589 77544 59594 77600
rect 59650 77544 62980 77600
rect 59589 77542 62980 77544
rect 126828 77542 129740 77602
rect 37417 77539 37483 77542
rect 59589 77539 59655 77542
rect 129734 77540 129740 77542
rect 129804 77602 129810 77604
rect 201085 77602 201151 77605
rect 129804 77542 134924 77602
rect 198772 77600 201151 77602
rect 198772 77544 201090 77600
rect 201146 77544 201151 77600
rect 198772 77542 201151 77544
rect 129804 77540 129810 77542
rect 201085 77539 201151 77542
rect 204489 77602 204555 77605
rect 204489 77600 207972 77602
rect 204489 77544 204494 77600
rect 204550 77544 207972 77600
rect 204489 77542 207972 77544
rect 204489 77539 204555 77542
rect 178821 77466 178887 77469
rect 174852 77464 178887 77466
rect 174852 77408 178826 77464
rect 178882 77408 178887 77464
rect 174852 77406 178887 77408
rect 178821 77403 178887 77406
rect 102694 76786 102754 77368
rect 106969 76786 107035 76789
rect 102694 76784 107035 76786
rect 102694 76728 106974 76784
rect 107030 76728 107035 76784
rect 102694 76726 107035 76728
rect 106969 76723 107035 76726
rect 107705 76650 107771 76653
rect 179465 76650 179531 76653
rect 107705 76648 111004 76650
rect 107705 76592 107710 76648
rect 107766 76592 111004 76648
rect 107705 76590 111004 76592
rect 179465 76648 182948 76650
rect 179465 76592 179470 76648
rect 179526 76592 182948 76648
rect 179465 76590 182948 76592
rect 107705 76587 107771 76590
rect 179465 76587 179531 76590
rect 178269 76242 178335 76245
rect 174852 76240 178335 76242
rect 174852 76184 178274 76240
rect 178330 76184 178335 76240
rect 174852 76182 178335 76184
rect 178269 76179 178335 76182
rect 11933 75154 11999 75157
rect 14006 75154 14066 75736
rect 102694 75562 102754 76144
rect 105957 75562 106023 75565
rect 102694 75560 106023 75562
rect 102694 75504 105962 75560
rect 106018 75504 106023 75560
rect 102694 75502 106023 75504
rect 105957 75499 106023 75502
rect 223582 75293 223642 75804
rect 223533 75288 223642 75293
rect 223533 75232 223538 75288
rect 223594 75232 223642 75288
rect 223533 75230 223642 75232
rect 223533 75227 223599 75230
rect 11933 75152 14066 75154
rect 11933 75096 11938 75152
rect 11994 75096 14066 75152
rect 11933 75094 14066 75096
rect 11933 75091 11999 75094
rect 177717 75018 177783 75021
rect 174852 75016 177783 75018
rect 174852 74960 177722 75016
rect 177778 74960 177783 75016
rect 174852 74958 177783 74960
rect 177717 74955 177783 74958
rect 102694 74338 102754 74920
rect 105405 74338 105471 74341
rect 102694 74336 105471 74338
rect 102694 74280 105410 74336
rect 105466 74280 105471 74336
rect 102694 74278 105471 74280
rect 105405 74275 105471 74278
rect 107889 74338 107955 74341
rect 179741 74338 179807 74341
rect 107889 74336 111004 74338
rect 107889 74280 107894 74336
rect 107950 74280 111004 74336
rect 107889 74278 111004 74280
rect 179741 74336 182948 74338
rect 179741 74280 179746 74336
rect 179802 74280 182948 74336
rect 179741 74278 182948 74280
rect 107889 74275 107955 74278
rect 179741 74275 179807 74278
rect 105221 73794 105287 73797
rect 177165 73794 177231 73797
rect 102724 73792 105287 73794
rect 102724 73736 105226 73792
rect 105282 73736 105287 73792
rect 102724 73734 105287 73736
rect 174852 73792 177231 73794
rect 174852 73736 177170 73792
rect 177226 73736 177231 73792
rect 174852 73734 177231 73736
rect 105221 73731 105287 73734
rect 177165 73731 177231 73734
rect 105865 72570 105931 72573
rect 177625 72570 177691 72573
rect 102724 72568 105931 72570
rect 102724 72512 105870 72568
rect 105926 72512 105931 72568
rect 102724 72510 105931 72512
rect 174852 72568 177691 72570
rect 174852 72512 177630 72568
rect 177686 72512 177691 72568
rect 174852 72510 177691 72512
rect 105865 72507 105931 72510
rect 177625 72507 177691 72510
rect 108533 72026 108599 72029
rect 180293 72026 180359 72029
rect 108533 72024 111004 72026
rect 108533 71968 108538 72024
rect 108594 71968 111004 72024
rect 108533 71966 111004 71968
rect 180293 72024 182948 72026
rect 180293 71968 180298 72024
rect 180354 71968 182948 72024
rect 180293 71966 182948 71968
rect 108533 71963 108599 71966
rect 180293 71963 180359 71966
rect 177349 71482 177415 71485
rect 174852 71480 177415 71482
rect 174852 71424 177354 71480
rect 177410 71424 177415 71480
rect 174852 71422 177415 71424
rect 177349 71419 177415 71422
rect 101357 71212 101423 71213
rect 101357 71210 101404 71212
rect 101312 71208 101404 71210
rect 101312 71152 101362 71208
rect 101312 71150 101404 71152
rect 101357 71148 101404 71150
rect 101468 71148 101474 71212
rect 101357 71147 101423 71148
rect 101030 71012 101036 71076
rect 101100 71074 101106 71076
rect 101909 71074 101975 71077
rect 101100 71072 101975 71074
rect 101100 71016 101914 71072
rect 101970 71016 101975 71072
rect 101100 71014 101975 71016
rect 102694 71074 102754 71384
rect 106509 71074 106575 71077
rect 102694 71072 106575 71074
rect 102694 71016 106514 71072
rect 106570 71016 106575 71072
rect 102694 71014 106575 71016
rect 101100 71012 101106 71014
rect 101909 71011 101975 71014
rect 106509 71011 106575 71014
rect 31897 69444 31963 69445
rect 31846 69442 31852 69444
rect 31806 69382 31852 69442
rect 31916 69440 31963 69444
rect 31958 69384 31963 69440
rect 31846 69380 31852 69382
rect 31916 69380 31963 69384
rect 31897 69379 31963 69380
rect 201085 69306 201151 69309
rect 201494 69306 201500 69308
rect 201085 69304 201500 69306
rect 201085 69248 201090 69304
rect 201146 69248 201500 69304
rect 201085 69246 201500 69248
rect 201085 69243 201151 69246
rect 201494 69244 201500 69246
rect 201564 69244 201570 69308
rect 117825 69170 117891 69173
rect 119389 69170 119455 69173
rect 117825 69168 119455 69170
rect 117825 69112 117830 69168
rect 117886 69112 119394 69168
rect 119450 69112 119455 69168
rect 117825 69110 119455 69112
rect 117825 69107 117891 69110
rect 119389 69107 119455 69110
rect 189309 69170 189375 69173
rect 190229 69170 190295 69173
rect 189309 69168 190295 69170
rect 189309 69112 189314 69168
rect 189370 69112 190234 69168
rect 190290 69112 190295 69168
rect 189309 69110 190295 69112
rect 189309 69107 189375 69110
rect 190229 69107 190295 69110
rect 191333 69170 191399 69173
rect 193081 69170 193147 69173
rect 191333 69168 193147 69170
rect 191333 69112 191338 69168
rect 191394 69112 193086 69168
rect 193142 69112 193147 69168
rect 191333 69110 193147 69112
rect 191333 69107 191399 69110
rect 193081 69107 193147 69110
rect 119113 69034 119179 69037
rect 121137 69034 121203 69037
rect 119113 69032 121203 69034
rect 119113 68976 119118 69032
rect 119174 68976 121142 69032
rect 121198 68976 121203 69032
rect 119113 68974 121203 68976
rect 119113 68971 119179 68974
rect 121137 68971 121203 68974
rect 223073 68354 223139 68357
rect 227416 68354 227896 68384
rect 223073 68352 227896 68354
rect 223073 68296 223078 68352
rect 223134 68296 227896 68352
rect 223073 68294 227896 68296
rect 223073 68291 223139 68294
rect 227416 68264 227896 68294
rect 103473 67538 103539 67541
rect 135305 67538 135371 67541
rect 103473 67536 104932 67538
rect 103473 67480 103478 67536
rect 103534 67480 104932 67536
rect 103473 67478 104932 67480
rect 132716 67536 135371 67538
rect 132716 67480 135310 67536
rect 135366 67480 135371 67536
rect 132716 67478 135371 67480
rect 103473 67475 103539 67478
rect 135305 67475 135371 67478
rect 175049 67538 175115 67541
rect 175049 67536 177060 67538
rect 175049 67480 175054 67536
rect 175110 67480 177060 67536
rect 175049 67478 177060 67480
rect 175049 67475 175115 67478
rect 63361 67266 63427 67269
rect 60772 67264 63427 67266
rect 60772 67208 63366 67264
rect 63422 67208 63427 67264
rect 60772 67206 63427 67208
rect 63361 67203 63427 67206
rect 102921 66994 102987 66997
rect 135029 66994 135095 66997
rect 102921 66992 104932 66994
rect 102921 66936 102926 66992
rect 102982 66936 104932 66992
rect 102921 66934 104932 66936
rect 132716 66992 135095 66994
rect 132716 66936 135034 66992
rect 135090 66936 135095 66992
rect 132716 66934 135095 66936
rect 102921 66931 102987 66934
rect 135029 66931 135095 66934
rect 174037 66994 174103 66997
rect 174037 66992 177060 66994
rect 174037 66936 174042 66992
rect 174098 66936 177060 66992
rect 174037 66934 177060 66936
rect 174037 66931 174103 66934
rect 62809 66722 62875 66725
rect 60772 66720 62875 66722
rect 60772 66664 62814 66720
rect 62870 66664 62875 66720
rect 60772 66662 62875 66664
rect 62809 66659 62875 66662
rect 102369 66450 102435 66453
rect 135305 66450 135371 66453
rect 102369 66448 104932 66450
rect 102369 66392 102374 66448
rect 102430 66392 104932 66448
rect 102369 66390 104932 66392
rect 132716 66448 135371 66450
rect 132716 66392 135310 66448
rect 135366 66392 135371 66448
rect 132716 66390 135371 66392
rect 102369 66387 102435 66390
rect 135305 66387 135371 66390
rect 173945 66450 174011 66453
rect 173945 66448 177060 66450
rect 173945 66392 173950 66448
rect 174006 66392 177060 66448
rect 173945 66390 177060 66392
rect 173945 66387 174011 66390
rect 62717 66178 62783 66181
rect 60772 66176 62783 66178
rect 60772 66120 62722 66176
rect 62778 66120 62783 66176
rect 60772 66118 62783 66120
rect 62717 66115 62783 66118
rect 102461 65906 102527 65909
rect 134661 65906 134727 65909
rect 102461 65904 104932 65906
rect 102461 65848 102466 65904
rect 102522 65848 104932 65904
rect 102461 65846 104932 65848
rect 132716 65904 134727 65906
rect 132716 65848 134666 65904
rect 134722 65848 134727 65904
rect 132716 65846 134727 65848
rect 102461 65843 102527 65846
rect 134661 65843 134727 65846
rect 173853 65906 173919 65909
rect 173853 65904 177060 65906
rect 173853 65848 173858 65904
rect 173914 65848 177060 65904
rect 173853 65846 177060 65848
rect 173853 65843 173919 65846
rect 62901 65634 62967 65637
rect 172657 65634 172723 65637
rect 60772 65632 62967 65634
rect 60772 65576 62906 65632
rect 62962 65576 62967 65632
rect 60772 65574 62967 65576
rect 62901 65571 62967 65574
rect 169670 65632 172723 65634
rect 169670 65576 172662 65632
rect 172718 65576 172723 65632
rect 169670 65574 172723 65576
rect 66397 65498 66463 65501
rect 100897 65498 100963 65501
rect 66397 65496 67948 65498
rect 66397 65440 66402 65496
rect 66458 65440 67948 65496
rect 66397 65438 67948 65440
rect 97756 65496 100963 65498
rect 97756 65440 100902 65496
rect 100958 65440 100963 65496
rect 97756 65438 100963 65440
rect 66397 65435 66463 65438
rect 100897 65435 100963 65438
rect 136869 65498 136935 65501
rect 136869 65496 140076 65498
rect 136869 65440 136874 65496
rect 136930 65440 140076 65496
rect 169670 65468 169730 65574
rect 172657 65571 172723 65574
rect 136869 65438 140076 65440
rect 136869 65435 136935 65438
rect 102737 65226 102803 65229
rect 135305 65226 135371 65229
rect 102737 65224 104932 65226
rect 102737 65168 102742 65224
rect 102798 65168 104932 65224
rect 102737 65166 104932 65168
rect 132716 65224 135371 65226
rect 132716 65168 135310 65224
rect 135366 65168 135371 65224
rect 132716 65166 135371 65168
rect 102737 65163 102803 65166
rect 135305 65163 135371 65166
rect 174129 65226 174195 65229
rect 174129 65224 177060 65226
rect 174129 65168 174134 65224
rect 174190 65168 177060 65224
rect 174129 65166 177060 65168
rect 174129 65163 174195 65166
rect 62809 64954 62875 64957
rect 60772 64952 62875 64954
rect 60772 64896 62814 64952
rect 62870 64896 62875 64952
rect 60772 64894 62875 64896
rect 62809 64891 62875 64894
rect 66397 64954 66463 64957
rect 66397 64952 67948 64954
rect 66397 64896 66402 64952
rect 66458 64896 67948 64952
rect 66397 64894 67948 64896
rect 66397 64891 66463 64894
rect 97726 64546 97786 64856
rect 102645 64682 102711 64685
rect 134845 64682 134911 64685
rect 102645 64680 104932 64682
rect 102645 64624 102650 64680
rect 102706 64624 104932 64680
rect 102645 64622 104932 64624
rect 132716 64680 134911 64682
rect 132716 64624 134850 64680
rect 134906 64624 134911 64680
rect 132716 64622 134911 64624
rect 102645 64619 102711 64622
rect 134845 64619 134911 64622
rect 100621 64546 100687 64549
rect 97726 64544 100687 64546
rect 97726 64488 100626 64544
rect 100682 64488 100687 64544
rect 97726 64486 100687 64488
rect 100621 64483 100687 64486
rect 136869 64546 136935 64549
rect 140046 64546 140106 64856
rect 136869 64544 140106 64546
rect 136869 64488 136874 64544
rect 136930 64488 140106 64544
rect 136869 64486 140106 64488
rect 169854 64546 169914 64924
rect 174221 64682 174287 64685
rect 174221 64680 177060 64682
rect 174221 64624 174226 64680
rect 174282 64624 177060 64680
rect 174221 64622 177060 64624
rect 174221 64619 174287 64622
rect 172657 64546 172723 64549
rect 169854 64544 172723 64546
rect 169854 64488 172662 64544
rect 172718 64488 172723 64544
rect 169854 64486 172723 64488
rect 136869 64483 136935 64486
rect 172657 64483 172723 64486
rect 62717 64410 62783 64413
rect 60772 64408 62783 64410
rect 60772 64352 62722 64408
rect 62778 64352 62783 64408
rect 60772 64350 62783 64352
rect 62717 64347 62783 64350
rect 65661 64274 65727 64277
rect 65661 64272 67948 64274
rect 65661 64216 65666 64272
rect 65722 64216 67948 64272
rect 65661 64214 67948 64216
rect 65661 64211 65727 64214
rect 97726 64138 97786 64176
rect 100897 64138 100963 64141
rect 97726 64136 100963 64138
rect 97726 64080 100902 64136
rect 100958 64080 100963 64136
rect 97726 64078 100963 64080
rect 100897 64075 100963 64078
rect 102553 64138 102619 64141
rect 134477 64138 134543 64141
rect 102553 64136 104932 64138
rect 102553 64080 102558 64136
rect 102614 64080 104932 64136
rect 102553 64078 104932 64080
rect 132716 64136 134543 64138
rect 132716 64080 134482 64136
rect 134538 64080 134543 64136
rect 132716 64078 134543 64080
rect 102553 64075 102619 64078
rect 134477 64075 134543 64078
rect 136961 64138 137027 64141
rect 140046 64138 140106 64176
rect 136961 64136 140106 64138
rect 136961 64080 136966 64136
rect 137022 64080 140106 64136
rect 136961 64078 140106 64080
rect 169854 64138 169914 64244
rect 171829 64138 171895 64141
rect 169854 64136 171895 64138
rect 169854 64080 171834 64136
rect 171890 64080 171895 64136
rect 169854 64078 171895 64080
rect 136961 64075 137027 64078
rect 171829 64075 171895 64078
rect 174405 64138 174471 64141
rect 174405 64136 177060 64138
rect 174405 64080 174410 64136
rect 174466 64080 177060 64136
rect 174405 64078 177060 64080
rect 174405 64075 174471 64078
rect 62993 63866 63059 63869
rect 60772 63864 63059 63866
rect 60772 63808 62998 63864
rect 63054 63808 63059 63864
rect 60772 63806 63059 63808
rect 62993 63803 63059 63806
rect 66397 63730 66463 63733
rect 66397 63728 67948 63730
rect 66397 63672 66402 63728
rect 66458 63672 67948 63728
rect 66397 63670 67948 63672
rect 66397 63667 66463 63670
rect 62349 63322 62415 63325
rect 60772 63320 62415 63322
rect 60772 63264 62354 63320
rect 62410 63264 62415 63320
rect 60772 63262 62415 63264
rect 97726 63322 97786 63632
rect 102553 63594 102619 63597
rect 135397 63594 135463 63597
rect 102553 63592 104932 63594
rect 102553 63536 102558 63592
rect 102614 63536 104932 63592
rect 102553 63534 104932 63536
rect 132716 63592 135463 63594
rect 132716 63536 135402 63592
rect 135458 63536 135463 63592
rect 132716 63534 135463 63536
rect 102553 63531 102619 63534
rect 135397 63531 135463 63534
rect 100621 63322 100687 63325
rect 97726 63320 100687 63322
rect 97726 63264 100626 63320
rect 100682 63264 100687 63320
rect 97726 63262 100687 63264
rect 62349 63259 62415 63262
rect 100621 63259 100687 63262
rect 136869 63322 136935 63325
rect 140046 63322 140106 63632
rect 136869 63320 140106 63322
rect 136869 63264 136874 63320
rect 136930 63264 140106 63320
rect 136869 63262 140106 63264
rect 169854 63322 169914 63700
rect 174129 63594 174195 63597
rect 174129 63592 177060 63594
rect 174129 63536 174134 63592
rect 174190 63536 177060 63592
rect 174129 63534 177060 63536
rect 174129 63531 174195 63534
rect 172657 63322 172723 63325
rect 169854 63320 172723 63322
rect 169854 63264 172662 63320
rect 172718 63264 172723 63320
rect 169854 63262 172723 63264
rect 136869 63259 136935 63262
rect 172657 63259 172723 63262
rect 65661 63186 65727 63189
rect 65661 63184 67948 63186
rect 65661 63128 65666 63184
rect 65722 63128 67948 63184
rect 65661 63126 67948 63128
rect 65661 63123 65727 63126
rect 9896 62914 10376 62944
rect 12025 62914 12091 62917
rect 9896 62912 12091 62914
rect 9896 62856 12030 62912
rect 12086 62856 12091 62912
rect 9896 62854 12091 62856
rect 9896 62824 10376 62854
rect 12025 62851 12091 62854
rect 29229 62914 29295 62917
rect 29229 62912 32988 62914
rect 29229 62856 29234 62912
rect 29290 62856 32988 62912
rect 29229 62854 32988 62856
rect 29229 62851 29295 62854
rect 63361 62778 63427 62781
rect 60772 62776 63427 62778
rect 60772 62720 63366 62776
rect 63422 62720 63427 62776
rect 60772 62718 63427 62720
rect 97726 62778 97786 63088
rect 102369 63050 102435 63053
rect 134661 63050 134727 63053
rect 102369 63048 104932 63050
rect 102369 62992 102374 63048
rect 102430 62992 104932 63048
rect 102369 62990 104932 62992
rect 132716 63048 134727 63050
rect 132716 62992 134666 63048
rect 134722 62992 134727 63048
rect 132716 62990 134727 62992
rect 102369 62987 102435 62990
rect 134661 62987 134727 62990
rect 100621 62778 100687 62781
rect 97726 62776 100687 62778
rect 97726 62720 100626 62776
rect 100682 62720 100687 62776
rect 97726 62718 100687 62720
rect 63361 62715 63427 62718
rect 100621 62715 100687 62718
rect 136961 62778 137027 62781
rect 140046 62778 140106 63088
rect 169854 62914 169914 63156
rect 175325 63050 175391 63053
rect 175325 63048 177060 63050
rect 175325 62992 175330 63048
rect 175386 62992 177060 63048
rect 175325 62990 177060 62992
rect 175325 62987 175391 62990
rect 172657 62914 172723 62917
rect 169854 62912 172723 62914
rect 169854 62856 172662 62912
rect 172718 62856 172723 62912
rect 169854 62854 172723 62856
rect 172657 62851 172723 62854
rect 136961 62776 140106 62778
rect 136961 62720 136966 62776
rect 137022 62720 140106 62776
rect 136961 62718 140106 62720
rect 136961 62715 137027 62718
rect 66397 62506 66463 62509
rect 66397 62504 67948 62506
rect 66397 62448 66402 62504
rect 66458 62448 67948 62504
rect 66397 62446 67948 62448
rect 66397 62443 66463 62446
rect 63545 62098 63611 62101
rect 60772 62096 63611 62098
rect 60772 62040 63550 62096
rect 63606 62040 63611 62096
rect 60772 62038 63611 62040
rect 97726 62098 97786 62408
rect 102737 62370 102803 62373
rect 134845 62370 134911 62373
rect 102737 62368 104932 62370
rect 102737 62312 102742 62368
rect 102798 62312 104932 62368
rect 102737 62310 104932 62312
rect 132716 62368 134911 62370
rect 132716 62312 134850 62368
rect 134906 62312 134911 62368
rect 132716 62310 134911 62312
rect 102737 62307 102803 62310
rect 134845 62307 134911 62310
rect 100621 62098 100687 62101
rect 97726 62096 100687 62098
rect 97726 62040 100626 62096
rect 100682 62040 100687 62096
rect 97726 62038 100687 62040
rect 63545 62035 63611 62038
rect 100621 62035 100687 62038
rect 136777 62098 136843 62101
rect 140046 62098 140106 62408
rect 136777 62096 140106 62098
rect 136777 62040 136782 62096
rect 136838 62040 140106 62096
rect 136777 62038 140106 62040
rect 169854 62098 169914 62476
rect 174221 62370 174287 62373
rect 174221 62368 177060 62370
rect 174221 62312 174226 62368
rect 174282 62312 177060 62368
rect 174221 62310 177060 62312
rect 174221 62307 174287 62310
rect 172657 62098 172723 62101
rect 169854 62096 172723 62098
rect 169854 62040 172662 62096
rect 172718 62040 172723 62096
rect 169854 62038 172723 62040
rect 136777 62035 136843 62038
rect 172657 62035 172723 62038
rect 65661 61962 65727 61965
rect 65661 61960 67948 61962
rect 65661 61904 65666 61960
rect 65722 61904 67948 61960
rect 65661 61902 67948 61904
rect 65661 61899 65727 61902
rect 63453 61554 63519 61557
rect 60772 61552 63519 61554
rect 60772 61496 63458 61552
rect 63514 61496 63519 61552
rect 60772 61494 63519 61496
rect 63453 61491 63519 61494
rect 97726 61418 97786 61864
rect 102461 61826 102527 61829
rect 135305 61826 135371 61829
rect 102461 61824 104932 61826
rect 102461 61768 102466 61824
rect 102522 61768 104932 61824
rect 102461 61766 104932 61768
rect 132716 61824 135371 61826
rect 132716 61768 135310 61824
rect 135366 61768 135371 61824
rect 132716 61766 135371 61768
rect 102461 61763 102527 61766
rect 135305 61763 135371 61766
rect 100529 61418 100595 61421
rect 97726 61416 100595 61418
rect 97726 61360 100534 61416
rect 100590 61360 100595 61416
rect 97726 61358 100595 61360
rect 100529 61355 100595 61358
rect 136869 61418 136935 61421
rect 140046 61418 140106 61864
rect 169854 61690 169914 61932
rect 175233 61826 175299 61829
rect 175233 61824 177060 61826
rect 175233 61768 175238 61824
rect 175294 61768 177060 61824
rect 175233 61766 177060 61768
rect 175233 61763 175299 61766
rect 171829 61690 171895 61693
rect 169854 61688 171895 61690
rect 169854 61632 171834 61688
rect 171890 61632 171895 61688
rect 169854 61630 171895 61632
rect 171829 61627 171895 61630
rect 136869 61416 140106 61418
rect 136869 61360 136874 61416
rect 136930 61360 140106 61416
rect 136869 61358 140106 61360
rect 136869 61355 136935 61358
rect 65477 61282 65543 61285
rect 102369 61282 102435 61285
rect 135397 61282 135463 61285
rect 65477 61280 67948 61282
rect 65477 61224 65482 61280
rect 65538 61224 67948 61280
rect 65477 61222 67948 61224
rect 102369 61280 104932 61282
rect 102369 61224 102374 61280
rect 102430 61224 104932 61280
rect 102369 61222 104932 61224
rect 132716 61280 135463 61282
rect 132716 61224 135402 61280
rect 135458 61224 135463 61280
rect 174129 61282 174195 61285
rect 174129 61280 177060 61282
rect 132716 61222 135463 61224
rect 65477 61219 65543 61222
rect 102369 61219 102435 61222
rect 135397 61219 135463 61222
rect 62809 61010 62875 61013
rect 60772 61008 62875 61010
rect 60772 60952 62814 61008
rect 62870 60952 62875 61008
rect 60772 60950 62875 60952
rect 62809 60947 62875 60950
rect 97726 60874 97786 61184
rect 100621 60874 100687 60877
rect 97726 60872 100687 60874
rect 97726 60816 100626 60872
rect 100682 60816 100687 60872
rect 97726 60814 100687 60816
rect 100621 60811 100687 60814
rect 136777 60874 136843 60877
rect 140046 60874 140106 61184
rect 136777 60872 140106 60874
rect 136777 60816 136782 60872
rect 136838 60816 140106 60872
rect 136777 60814 140106 60816
rect 169854 60874 169914 61252
rect 174129 61224 174134 61280
rect 174190 61224 177060 61280
rect 174129 61222 177060 61224
rect 174129 61219 174195 61222
rect 172197 60874 172263 60877
rect 169854 60872 172263 60874
rect 169854 60816 172202 60872
rect 172258 60816 172263 60872
rect 169854 60814 172263 60816
rect 136777 60811 136843 60814
rect 172197 60811 172263 60814
rect 66305 60738 66371 60741
rect 102553 60738 102619 60741
rect 134477 60738 134543 60741
rect 66305 60736 67948 60738
rect 66305 60680 66310 60736
rect 66366 60680 67948 60736
rect 66305 60678 67948 60680
rect 102553 60736 104932 60738
rect 102553 60680 102558 60736
rect 102614 60680 104932 60736
rect 102553 60678 104932 60680
rect 132716 60736 134543 60738
rect 132716 60680 134482 60736
rect 134538 60680 134543 60736
rect 174313 60738 174379 60741
rect 174313 60736 177060 60738
rect 132716 60678 134543 60680
rect 66305 60675 66371 60678
rect 102553 60675 102619 60678
rect 134477 60675 134543 60678
rect 62717 60466 62783 60469
rect 60772 60464 62783 60466
rect 60772 60408 62722 60464
rect 62778 60408 62783 60464
rect 60772 60406 62783 60408
rect 62717 60403 62783 60406
rect 97726 60330 97786 60640
rect 100621 60330 100687 60333
rect 97726 60328 100687 60330
rect 97726 60272 100626 60328
rect 100682 60272 100687 60328
rect 97726 60270 100687 60272
rect 100621 60267 100687 60270
rect 136961 60330 137027 60333
rect 140046 60330 140106 60640
rect 136961 60328 140106 60330
rect 136961 60272 136966 60328
rect 137022 60272 140106 60328
rect 136961 60270 140106 60272
rect 169854 60330 169914 60708
rect 174313 60680 174318 60736
rect 174374 60680 177060 60736
rect 174313 60678 177060 60680
rect 174313 60675 174379 60678
rect 172657 60330 172723 60333
rect 169854 60328 172723 60330
rect 169854 60272 172662 60328
rect 172718 60272 172723 60328
rect 169854 60270 172723 60272
rect 136961 60267 137027 60270
rect 172657 60267 172723 60270
rect 66397 60194 66463 60197
rect 102461 60194 102527 60197
rect 135029 60194 135095 60197
rect 66397 60192 67948 60194
rect 66397 60136 66402 60192
rect 66458 60136 67948 60192
rect 66397 60134 67948 60136
rect 102461 60192 104932 60194
rect 102461 60136 102466 60192
rect 102522 60136 104932 60192
rect 102461 60134 104932 60136
rect 132716 60192 135095 60194
rect 132716 60136 135034 60192
rect 135090 60136 135095 60192
rect 174221 60194 174287 60197
rect 174221 60192 177060 60194
rect 132716 60134 135095 60136
rect 66397 60131 66463 60134
rect 102461 60131 102527 60134
rect 135029 60131 135095 60134
rect 97726 60058 97786 60096
rect 100621 60058 100687 60061
rect 97726 60056 100687 60058
rect 97726 60000 100626 60056
rect 100682 60000 100687 60056
rect 97726 59998 100687 60000
rect 100621 59995 100687 59998
rect 136869 60058 136935 60061
rect 140046 60058 140106 60096
rect 136869 60056 140106 60058
rect 136869 60000 136874 60056
rect 136930 60000 140106 60056
rect 136869 59998 140106 60000
rect 169854 60058 169914 60164
rect 174221 60136 174226 60192
rect 174282 60136 177060 60192
rect 174221 60134 177060 60136
rect 174221 60131 174287 60134
rect 172657 60058 172723 60061
rect 169854 60056 172723 60058
rect 169854 60000 172662 60056
rect 172718 60000 172723 60056
rect 169854 59998 172723 60000
rect 136869 59995 136935 59998
rect 172657 59995 172723 59998
rect 63729 59922 63795 59925
rect 60772 59920 63795 59922
rect 60772 59864 63734 59920
rect 63790 59864 63795 59920
rect 60772 59862 63795 59864
rect 63729 59859 63795 59862
rect 66305 59514 66371 59517
rect 102737 59514 102803 59517
rect 135305 59514 135371 59517
rect 66305 59512 67948 59514
rect 66305 59456 66310 59512
rect 66366 59456 67948 59512
rect 66305 59454 67948 59456
rect 102737 59512 104932 59514
rect 102737 59456 102742 59512
rect 102798 59456 104932 59512
rect 102737 59454 104932 59456
rect 132716 59512 135371 59514
rect 132716 59456 135310 59512
rect 135366 59456 135371 59512
rect 174405 59514 174471 59517
rect 174405 59512 177060 59514
rect 132716 59454 135371 59456
rect 66305 59451 66371 59454
rect 102737 59451 102803 59454
rect 135305 59451 135371 59454
rect 62901 59242 62967 59245
rect 60772 59240 62967 59242
rect 60772 59184 62906 59240
rect 62962 59184 62967 59240
rect 60772 59182 62967 59184
rect 62901 59179 62967 59182
rect 97726 59106 97786 59416
rect 100621 59106 100687 59109
rect 97726 59104 100687 59106
rect 97726 59048 100626 59104
rect 100682 59048 100687 59104
rect 97726 59046 100687 59048
rect 100621 59043 100687 59046
rect 136777 59106 136843 59109
rect 140046 59106 140106 59416
rect 136777 59104 140106 59106
rect 136777 59048 136782 59104
rect 136838 59048 140106 59104
rect 136777 59046 140106 59048
rect 169854 59106 169914 59484
rect 174405 59456 174410 59512
rect 174466 59456 177060 59512
rect 174405 59454 177060 59456
rect 174405 59451 174471 59454
rect 172197 59106 172263 59109
rect 169854 59104 172263 59106
rect 169854 59048 172202 59104
rect 172258 59048 172263 59104
rect 169854 59046 172263 59048
rect 136777 59043 136843 59046
rect 172197 59043 172263 59046
rect 66397 58970 66463 58973
rect 102645 58970 102711 58973
rect 135029 58970 135095 58973
rect 66397 58968 67948 58970
rect 66397 58912 66402 58968
rect 66458 58912 67948 58968
rect 66397 58910 67948 58912
rect 102645 58968 104932 58970
rect 102645 58912 102650 58968
rect 102706 58912 104932 58968
rect 102645 58910 104932 58912
rect 132716 58968 135095 58970
rect 132716 58912 135034 58968
rect 135090 58912 135095 58968
rect 174129 58970 174195 58973
rect 174129 58968 177060 58970
rect 132716 58910 135095 58912
rect 66397 58907 66463 58910
rect 102645 58907 102711 58910
rect 135029 58907 135095 58910
rect 63821 58698 63887 58701
rect 60772 58696 63887 58698
rect 60772 58640 63826 58696
rect 63882 58640 63887 58696
rect 60772 58638 63887 58640
rect 97726 58698 97786 58872
rect 100621 58698 100687 58701
rect 97726 58696 100687 58698
rect 97726 58640 100626 58696
rect 100682 58640 100687 58696
rect 97726 58638 100687 58640
rect 63821 58635 63887 58638
rect 100621 58635 100687 58638
rect 136869 58698 136935 58701
rect 140046 58698 140106 58872
rect 169854 58834 169914 58940
rect 174129 58912 174134 58968
rect 174190 58912 177060 58968
rect 174129 58910 177060 58912
rect 174129 58907 174195 58910
rect 171829 58834 171895 58837
rect 169854 58832 171895 58834
rect 169854 58776 171834 58832
rect 171890 58776 171895 58832
rect 169854 58774 171895 58776
rect 171829 58771 171895 58774
rect 136869 58696 140106 58698
rect 136869 58640 136874 58696
rect 136930 58640 140106 58696
rect 136869 58638 140106 58640
rect 136869 58635 136935 58638
rect 102369 58426 102435 58429
rect 134477 58426 134543 58429
rect 102369 58424 104932 58426
rect 102369 58368 102374 58424
rect 102430 58368 104932 58424
rect 102369 58366 104932 58368
rect 132716 58424 134543 58426
rect 132716 58368 134482 58424
rect 134538 58368 134543 58424
rect 132716 58366 134543 58368
rect 102369 58363 102435 58366
rect 134477 58363 134543 58366
rect 174313 58426 174379 58429
rect 174313 58424 177060 58426
rect 174313 58368 174318 58424
rect 174374 58368 177060 58424
rect 174313 58366 177060 58368
rect 174313 58363 174379 58366
rect 65017 58290 65083 58293
rect 65017 58288 67948 58290
rect 65017 58232 65022 58288
rect 65078 58232 67948 58288
rect 65017 58230 67948 58232
rect 65017 58227 65083 58230
rect 62717 58154 62783 58157
rect 60772 58152 62783 58154
rect 60772 58096 62722 58152
rect 62778 58096 62783 58152
rect 60772 58094 62783 58096
rect 62717 58091 62783 58094
rect 97726 57882 97786 58192
rect 100621 57882 100687 57885
rect 97726 57880 100687 57882
rect 97726 57824 100626 57880
rect 100682 57824 100687 57880
rect 97726 57822 100687 57824
rect 100621 57819 100687 57822
rect 102553 57882 102619 57885
rect 135397 57882 135463 57885
rect 102553 57880 104932 57882
rect 102553 57824 102558 57880
rect 102614 57824 104932 57880
rect 102553 57822 104932 57824
rect 132716 57880 135463 57882
rect 132716 57824 135402 57880
rect 135458 57824 135463 57880
rect 132716 57822 135463 57824
rect 102553 57819 102619 57822
rect 135397 57819 135463 57822
rect 136777 57882 136843 57885
rect 140046 57882 140106 58192
rect 136777 57880 140106 57882
rect 136777 57824 136782 57880
rect 136838 57824 140106 57880
rect 136777 57822 140106 57824
rect 169854 57882 169914 58260
rect 172013 57882 172079 57885
rect 169854 57880 172079 57882
rect 169854 57824 172018 57880
rect 172074 57824 172079 57880
rect 169854 57822 172079 57824
rect 136777 57819 136843 57822
rect 172013 57819 172079 57822
rect 174497 57882 174563 57885
rect 174497 57880 177060 57882
rect 174497 57824 174502 57880
rect 174558 57824 177060 57880
rect 174497 57822 177060 57824
rect 174497 57819 174563 57822
rect 66397 57746 66463 57749
rect 66397 57744 67948 57746
rect 66397 57688 66402 57744
rect 66458 57688 67948 57744
rect 66397 57686 67948 57688
rect 66397 57683 66463 57686
rect 62625 57610 62691 57613
rect 60772 57608 62691 57610
rect 60772 57552 62630 57608
rect 62686 57552 62691 57608
rect 60772 57550 62691 57552
rect 62625 57547 62691 57550
rect 97726 57338 97786 57648
rect 100621 57338 100687 57341
rect 97726 57336 100687 57338
rect 97726 57280 100626 57336
rect 100682 57280 100687 57336
rect 97726 57278 100687 57280
rect 100621 57275 100687 57278
rect 102461 57338 102527 57341
rect 135029 57338 135095 57341
rect 102461 57336 104932 57338
rect 102461 57280 102466 57336
rect 102522 57280 104932 57336
rect 102461 57278 104932 57280
rect 132716 57336 135095 57338
rect 132716 57280 135034 57336
rect 135090 57280 135095 57336
rect 132716 57278 135095 57280
rect 102461 57275 102527 57278
rect 135029 57275 135095 57278
rect 136869 57338 136935 57341
rect 140046 57338 140106 57648
rect 169854 57474 169914 57716
rect 172657 57474 172723 57477
rect 169854 57472 172723 57474
rect 169854 57416 172662 57472
rect 172718 57416 172723 57472
rect 169854 57414 172723 57416
rect 172657 57411 172723 57414
rect 172657 57338 172723 57341
rect 136869 57336 140106 57338
rect 136869 57280 136874 57336
rect 136930 57280 140106 57336
rect 136869 57278 140106 57280
rect 169670 57336 172723 57338
rect 169670 57280 172662 57336
rect 172718 57280 172723 57336
rect 169670 57278 172723 57280
rect 136869 57275 136935 57278
rect 66397 57202 66463 57205
rect 100529 57202 100595 57205
rect 66397 57200 67948 57202
rect 66397 57144 66402 57200
rect 66458 57144 67948 57200
rect 66397 57142 67948 57144
rect 97756 57200 100595 57202
rect 97756 57144 100534 57200
rect 100590 57144 100595 57200
rect 97756 57142 100595 57144
rect 66397 57139 66463 57142
rect 100529 57139 100595 57142
rect 136961 57202 137027 57205
rect 136961 57200 140076 57202
rect 136961 57144 136966 57200
rect 137022 57144 140076 57200
rect 169670 57172 169730 57278
rect 172657 57275 172723 57278
rect 174589 57338 174655 57341
rect 174589 57336 177060 57338
rect 174589 57280 174594 57336
rect 174650 57280 177060 57336
rect 174589 57278 177060 57280
rect 174589 57275 174655 57278
rect 136961 57142 140076 57144
rect 136961 57139 137027 57142
rect 62809 57066 62875 57069
rect 60772 57064 62875 57066
rect 60772 57008 62814 57064
rect 62870 57008 62875 57064
rect 60772 57006 62875 57008
rect 62809 57003 62875 57006
rect 102645 56658 102711 56661
rect 135305 56658 135371 56661
rect 102645 56656 104932 56658
rect 102645 56600 102650 56656
rect 102706 56600 104932 56656
rect 102645 56598 104932 56600
rect 132716 56656 135371 56658
rect 132716 56600 135310 56656
rect 135366 56600 135371 56656
rect 132716 56598 135371 56600
rect 102645 56595 102711 56598
rect 135305 56595 135371 56598
rect 174221 56658 174287 56661
rect 174221 56656 177060 56658
rect 174221 56600 174226 56656
rect 174282 56600 177060 56656
rect 174221 56598 177060 56600
rect 174221 56595 174287 56598
rect 66397 56522 66463 56525
rect 66397 56520 67948 56522
rect 66397 56464 66402 56520
rect 66458 56464 67948 56520
rect 66397 56462 67948 56464
rect 66397 56459 66463 56462
rect 62901 56386 62967 56389
rect 60772 56384 62967 56386
rect 60772 56328 62906 56384
rect 62962 56328 62967 56384
rect 60772 56326 62967 56328
rect 62901 56323 62967 56326
rect 97726 56114 97786 56424
rect 100621 56114 100687 56117
rect 97726 56112 100687 56114
rect 97726 56056 100626 56112
rect 100682 56056 100687 56112
rect 97726 56054 100687 56056
rect 100621 56051 100687 56054
rect 102369 56114 102435 56117
rect 135029 56114 135095 56117
rect 102369 56112 104932 56114
rect 102369 56056 102374 56112
rect 102430 56056 104932 56112
rect 102369 56054 104932 56056
rect 132716 56112 135095 56114
rect 132716 56056 135034 56112
rect 135090 56056 135095 56112
rect 132716 56054 135095 56056
rect 102369 56051 102435 56054
rect 135029 56051 135095 56054
rect 136777 56114 136843 56117
rect 140046 56114 140106 56424
rect 136777 56112 140106 56114
rect 136777 56056 136782 56112
rect 136838 56056 140106 56112
rect 136777 56054 140106 56056
rect 169854 56114 169914 56492
rect 172657 56114 172723 56117
rect 169854 56112 172723 56114
rect 169854 56056 172662 56112
rect 172718 56056 172723 56112
rect 169854 56054 172723 56056
rect 136777 56051 136843 56054
rect 172657 56051 172723 56054
rect 174129 56114 174195 56117
rect 174129 56112 177060 56114
rect 174129 56056 174134 56112
rect 174190 56056 177060 56112
rect 174129 56054 177060 56056
rect 174129 56051 174195 56054
rect 66397 55978 66463 55981
rect 66397 55976 67948 55978
rect 66397 55920 66402 55976
rect 66458 55920 67948 55976
rect 66397 55918 67948 55920
rect 66397 55915 66463 55918
rect 62533 55842 62599 55845
rect 60772 55840 62599 55842
rect 60772 55784 62538 55840
rect 62594 55784 62599 55840
rect 60772 55782 62599 55784
rect 97726 55842 97786 55880
rect 100897 55842 100963 55845
rect 97726 55840 100963 55842
rect 97726 55784 100902 55840
rect 100958 55784 100963 55840
rect 97726 55782 100963 55784
rect 62533 55779 62599 55782
rect 100897 55779 100963 55782
rect 136869 55842 136935 55845
rect 140046 55842 140106 55880
rect 136869 55840 140106 55842
rect 136869 55784 136874 55840
rect 136930 55784 140106 55840
rect 136869 55782 140106 55784
rect 169854 55842 169914 55948
rect 172657 55842 172723 55845
rect 169854 55840 172723 55842
rect 169854 55784 172662 55840
rect 172718 55784 172723 55840
rect 169854 55782 172723 55784
rect 136869 55779 136935 55782
rect 172657 55779 172723 55782
rect 102461 55570 102527 55573
rect 134753 55570 134819 55573
rect 102461 55568 104932 55570
rect 102461 55512 102466 55568
rect 102522 55512 104932 55568
rect 102461 55510 104932 55512
rect 132716 55568 134819 55570
rect 132716 55512 134758 55568
rect 134814 55512 134819 55568
rect 132716 55510 134819 55512
rect 102461 55507 102527 55510
rect 134753 55507 134819 55510
rect 174313 55570 174379 55573
rect 174313 55568 177060 55570
rect 174313 55512 174318 55568
rect 174374 55512 177060 55568
rect 174313 55510 177060 55512
rect 174313 55507 174379 55510
rect 62717 55298 62783 55301
rect 60772 55296 62783 55298
rect 60772 55240 62722 55296
rect 62778 55240 62783 55296
rect 60772 55238 62783 55240
rect 62717 55235 62783 55238
rect 66305 55298 66371 55301
rect 66305 55296 67948 55298
rect 66305 55240 66310 55296
rect 66366 55240 67948 55296
rect 66305 55238 67948 55240
rect 66305 55235 66371 55238
rect 97726 54890 97786 55200
rect 102553 55026 102619 55029
rect 135397 55026 135463 55029
rect 102553 55024 104932 55026
rect 102553 54968 102558 55024
rect 102614 54968 104932 55024
rect 102553 54966 104932 54968
rect 132716 55024 135463 55026
rect 132716 54968 135402 55024
rect 135458 54968 135463 55024
rect 132716 54966 135463 54968
rect 102553 54963 102619 54966
rect 135397 54963 135463 54966
rect 100621 54890 100687 54893
rect 97726 54888 100687 54890
rect 97726 54832 100626 54888
rect 100682 54832 100687 54888
rect 97726 54830 100687 54832
rect 100621 54827 100687 54830
rect 136777 54890 136843 54893
rect 140046 54890 140106 55200
rect 136777 54888 140106 54890
rect 136777 54832 136782 54888
rect 136838 54832 140106 54888
rect 136777 54830 140106 54832
rect 169854 54890 169914 55268
rect 174405 55026 174471 55029
rect 174405 55024 177060 55026
rect 174405 54968 174410 55024
rect 174466 54968 177060 55024
rect 174405 54966 177060 54968
rect 174405 54963 174471 54966
rect 172105 54890 172171 54893
rect 169854 54888 172171 54890
rect 169854 54832 172110 54888
rect 172166 54832 172171 54888
rect 169854 54830 172171 54832
rect 136777 54827 136843 54830
rect 172105 54827 172171 54830
rect 62625 54754 62691 54757
rect 60772 54752 62691 54754
rect 60772 54696 62630 54752
rect 62686 54696 62691 54752
rect 60772 54694 62691 54696
rect 62625 54691 62691 54694
rect 66397 54754 66463 54757
rect 66397 54752 67948 54754
rect 66397 54696 66402 54752
rect 66458 54696 67948 54752
rect 66397 54694 67948 54696
rect 66397 54691 66463 54694
rect 97726 54618 97786 54656
rect 100805 54618 100871 54621
rect 97726 54616 100871 54618
rect 97726 54560 100810 54616
rect 100866 54560 100871 54616
rect 97726 54558 100871 54560
rect 100805 54555 100871 54558
rect 137145 54618 137211 54621
rect 140046 54618 140106 54656
rect 137145 54616 140106 54618
rect 137145 54560 137150 54616
rect 137206 54560 140106 54616
rect 137145 54558 140106 54560
rect 169854 54618 169914 54724
rect 172657 54618 172723 54621
rect 169854 54616 172723 54618
rect 169854 54560 172662 54616
rect 172718 54560 172723 54616
rect 169854 54558 172723 54560
rect 137145 54555 137211 54558
rect 172657 54555 172723 54558
rect 102369 54482 102435 54485
rect 135029 54482 135095 54485
rect 102369 54480 104932 54482
rect 102369 54424 102374 54480
rect 102430 54424 104932 54480
rect 102369 54422 104932 54424
rect 132716 54480 135095 54482
rect 132716 54424 135034 54480
rect 135090 54424 135095 54480
rect 132716 54422 135095 54424
rect 102369 54419 102435 54422
rect 135029 54419 135095 54422
rect 174221 54482 174287 54485
rect 174221 54480 177060 54482
rect 174221 54424 174226 54480
rect 174282 54424 177060 54480
rect 174221 54422 177060 54424
rect 174221 54419 174287 54422
rect 63637 54210 63703 54213
rect 60772 54208 63703 54210
rect 60772 54152 63642 54208
rect 63698 54152 63703 54208
rect 60772 54150 63703 54152
rect 63637 54147 63703 54150
rect 66397 54210 66463 54213
rect 66397 54208 67948 54210
rect 66397 54152 66402 54208
rect 66458 54152 67948 54208
rect 66397 54150 67948 54152
rect 66397 54147 66463 54150
rect 97726 53666 97786 54112
rect 102645 53802 102711 53805
rect 134201 53802 134267 53805
rect 102645 53800 104932 53802
rect 102645 53744 102650 53800
rect 102706 53744 104932 53800
rect 102645 53742 104932 53744
rect 132716 53800 134267 53802
rect 132716 53744 134206 53800
rect 134262 53744 134267 53800
rect 132716 53742 134267 53744
rect 102645 53739 102711 53742
rect 134201 53739 134267 53742
rect 100621 53666 100687 53669
rect 97726 53664 100687 53666
rect 97726 53608 100626 53664
rect 100682 53608 100687 53664
rect 97726 53606 100687 53608
rect 100621 53603 100687 53606
rect 136777 53666 136843 53669
rect 140046 53666 140106 54112
rect 136777 53664 140106 53666
rect 136777 53608 136782 53664
rect 136838 53608 140106 53664
rect 136777 53606 140106 53608
rect 169854 53666 169914 54180
rect 174957 53802 175023 53805
rect 174957 53800 177060 53802
rect 174957 53744 174962 53800
rect 175018 53744 177060 53800
rect 174957 53742 177060 53744
rect 174957 53739 175023 53742
rect 171645 53666 171711 53669
rect 169854 53664 171711 53666
rect 169854 53608 171650 53664
rect 171706 53608 171711 53664
rect 169854 53606 171711 53608
rect 136777 53603 136843 53606
rect 171645 53603 171711 53606
rect 30517 53530 30583 53533
rect 63269 53530 63335 53533
rect 30517 53528 32988 53530
rect 30517 53472 30522 53528
rect 30578 53472 32988 53528
rect 30517 53470 32988 53472
rect 60772 53528 63335 53530
rect 60772 53472 63274 53528
rect 63330 53472 63335 53528
rect 60772 53470 63335 53472
rect 30517 53467 30583 53470
rect 63269 53467 63335 53470
rect 65293 53530 65359 53533
rect 65293 53528 67948 53530
rect 65293 53472 65298 53528
rect 65354 53472 67948 53528
rect 65293 53470 67948 53472
rect 65293 53467 65359 53470
rect 97726 53122 97786 53432
rect 102461 53258 102527 53261
rect 135121 53258 135187 53261
rect 102461 53256 104932 53258
rect 102461 53200 102466 53256
rect 102522 53200 104932 53256
rect 102461 53198 104932 53200
rect 132716 53256 135187 53258
rect 132716 53200 135126 53256
rect 135182 53200 135187 53256
rect 132716 53198 135187 53200
rect 102461 53195 102527 53198
rect 135121 53195 135187 53198
rect 100621 53122 100687 53125
rect 97726 53120 100687 53122
rect 97726 53064 100626 53120
rect 100682 53064 100687 53120
rect 97726 53062 100687 53064
rect 100621 53059 100687 53062
rect 136869 53122 136935 53125
rect 140046 53122 140106 53432
rect 169854 53258 169914 53500
rect 172657 53258 172723 53261
rect 169854 53256 172723 53258
rect 169854 53200 172662 53256
rect 172718 53200 172723 53256
rect 169854 53198 172723 53200
rect 172657 53195 172723 53198
rect 174773 53258 174839 53261
rect 174773 53256 177060 53258
rect 174773 53200 174778 53256
rect 174834 53200 177060 53256
rect 174773 53198 177060 53200
rect 174773 53195 174839 53198
rect 136869 53120 140106 53122
rect 136869 53064 136874 53120
rect 136930 53064 140106 53120
rect 136869 53062 140106 53064
rect 136869 53059 136935 53062
rect 63545 52986 63611 52989
rect 60772 52984 63611 52986
rect 60772 52928 63550 52984
rect 63606 52928 63611 52984
rect 60772 52926 63611 52928
rect 63545 52923 63611 52926
rect 66305 52986 66371 52989
rect 66305 52984 67948 52986
rect 66305 52928 66310 52984
rect 66366 52928 67948 52984
rect 66305 52926 67948 52928
rect 66305 52923 66371 52926
rect 63361 52442 63427 52445
rect 60772 52440 63427 52442
rect 60772 52384 63366 52440
rect 63422 52384 63427 52440
rect 60772 52382 63427 52384
rect 97726 52442 97786 52888
rect 102553 52714 102619 52717
rect 134293 52714 134359 52717
rect 102553 52712 104932 52714
rect 102553 52656 102558 52712
rect 102614 52656 104932 52712
rect 102553 52654 104932 52656
rect 132716 52712 134359 52714
rect 132716 52656 134298 52712
rect 134354 52656 134359 52712
rect 132716 52654 134359 52656
rect 102553 52651 102619 52654
rect 134293 52651 134359 52654
rect 100621 52442 100687 52445
rect 97726 52440 100687 52442
rect 97726 52384 100626 52440
rect 100682 52384 100687 52440
rect 97726 52382 100687 52384
rect 63361 52379 63427 52382
rect 100621 52379 100687 52382
rect 136685 52442 136751 52445
rect 140046 52442 140106 52888
rect 136685 52440 140106 52442
rect 136685 52384 136690 52440
rect 136746 52384 140106 52440
rect 136685 52382 140106 52384
rect 169854 52442 169914 52956
rect 175325 52714 175391 52717
rect 175325 52712 177060 52714
rect 175325 52656 175330 52712
rect 175386 52656 177060 52712
rect 175325 52654 177060 52656
rect 175325 52651 175391 52654
rect 172013 52442 172079 52445
rect 169854 52440 172079 52442
rect 169854 52384 172018 52440
rect 172074 52384 172079 52440
rect 169854 52382 172079 52384
rect 136685 52379 136751 52382
rect 172013 52379 172079 52382
rect 65293 52306 65359 52309
rect 65293 52304 67948 52306
rect 65293 52248 65298 52304
rect 65354 52248 67948 52304
rect 65293 52246 67948 52248
rect 65293 52243 65359 52246
rect 63729 51898 63795 51901
rect 60772 51896 63795 51898
rect 60772 51840 63734 51896
rect 63790 51840 63795 51896
rect 60772 51838 63795 51840
rect 97726 51898 97786 52208
rect 102737 52170 102803 52173
rect 135121 52170 135187 52173
rect 102737 52168 104932 52170
rect 102737 52112 102742 52168
rect 102798 52112 104932 52168
rect 102737 52110 104932 52112
rect 132716 52168 135187 52170
rect 132716 52112 135126 52168
rect 135182 52112 135187 52168
rect 132716 52110 135187 52112
rect 102737 52107 102803 52110
rect 135121 52107 135187 52110
rect 100621 51898 100687 51901
rect 97726 51896 100687 51898
rect 97726 51840 100626 51896
rect 100682 51840 100687 51896
rect 97726 51838 100687 51840
rect 63729 51835 63795 51838
rect 100621 51835 100687 51838
rect 136777 51898 136843 51901
rect 140046 51898 140106 52208
rect 169854 52034 169914 52276
rect 174129 52170 174195 52173
rect 174129 52168 177060 52170
rect 174129 52112 174134 52168
rect 174190 52112 177060 52168
rect 174129 52110 177060 52112
rect 174129 52107 174195 52110
rect 172565 52034 172631 52037
rect 169854 52032 172631 52034
rect 169854 51976 172570 52032
rect 172626 51976 172631 52032
rect 169854 51974 172631 51976
rect 172565 51971 172631 51974
rect 172657 51898 172723 51901
rect 136777 51896 140106 51898
rect 136777 51840 136782 51896
rect 136838 51840 140106 51896
rect 136777 51838 140106 51840
rect 169670 51896 172723 51898
rect 169670 51840 172662 51896
rect 172718 51840 172723 51896
rect 169670 51838 172723 51840
rect 136777 51835 136843 51838
rect 65661 51762 65727 51765
rect 100529 51762 100595 51765
rect 65661 51760 67948 51762
rect 65661 51704 65666 51760
rect 65722 51704 67948 51760
rect 65661 51702 67948 51704
rect 97756 51760 100595 51762
rect 97756 51704 100534 51760
rect 100590 51704 100595 51760
rect 97756 51702 100595 51704
rect 65661 51699 65727 51702
rect 100529 51699 100595 51702
rect 136869 51762 136935 51765
rect 136869 51760 140076 51762
rect 136869 51704 136874 51760
rect 136930 51704 140076 51760
rect 169670 51732 169730 51838
rect 172657 51835 172723 51838
rect 136869 51702 140076 51704
rect 136869 51699 136935 51702
rect 102369 51626 102435 51629
rect 135397 51626 135463 51629
rect 102369 51624 104932 51626
rect 102369 51568 102374 51624
rect 102430 51568 104932 51624
rect 102369 51566 104932 51568
rect 132716 51624 135463 51626
rect 132716 51568 135402 51624
rect 135458 51568 135463 51624
rect 132716 51566 135463 51568
rect 102369 51563 102435 51566
rect 135397 51563 135463 51566
rect 174497 51626 174563 51629
rect 174497 51624 177060 51626
rect 174497 51568 174502 51624
rect 174558 51568 177060 51624
rect 174497 51566 177060 51568
rect 174497 51563 174563 51566
rect 62809 51354 62875 51357
rect 60772 51352 62875 51354
rect 60772 51296 62814 51352
rect 62870 51296 62875 51352
rect 60772 51294 62875 51296
rect 62809 51291 62875 51294
rect 66397 51218 66463 51221
rect 66397 51216 67948 51218
rect 66397 51160 66402 51216
rect 66458 51160 67948 51216
rect 66397 51158 67948 51160
rect 66397 51155 66463 51158
rect 63729 50674 63795 50677
rect 60772 50672 63795 50674
rect 60772 50616 63734 50672
rect 63790 50616 63795 50672
rect 60772 50614 63795 50616
rect 97726 50674 97786 51120
rect 102645 50946 102711 50949
rect 135397 50946 135463 50949
rect 102645 50944 104932 50946
rect 102645 50888 102650 50944
rect 102706 50888 104932 50944
rect 102645 50886 104932 50888
rect 132716 50944 135463 50946
rect 132716 50888 135402 50944
rect 135458 50888 135463 50944
rect 132716 50886 135463 50888
rect 102645 50883 102711 50886
rect 135397 50883 135463 50886
rect 100621 50674 100687 50677
rect 97726 50672 100687 50674
rect 97726 50616 100626 50672
rect 100682 50616 100687 50672
rect 97726 50614 100687 50616
rect 63729 50611 63795 50614
rect 100621 50611 100687 50614
rect 136777 50674 136843 50677
rect 140046 50674 140106 51120
rect 169854 50810 169914 51188
rect 174221 50946 174287 50949
rect 174221 50944 177060 50946
rect 174221 50888 174226 50944
rect 174282 50888 177060 50944
rect 174221 50886 177060 50888
rect 174221 50883 174287 50886
rect 172197 50810 172263 50813
rect 169854 50808 172263 50810
rect 169854 50752 172202 50808
rect 172258 50752 172263 50808
rect 169854 50750 172263 50752
rect 172197 50747 172263 50750
rect 136777 50672 140106 50674
rect 136777 50616 136782 50672
rect 136838 50616 140106 50672
rect 136777 50614 140106 50616
rect 136777 50611 136843 50614
rect 65661 50538 65727 50541
rect 65661 50536 67948 50538
rect 65661 50480 65666 50536
rect 65722 50480 67948 50536
rect 65661 50478 67948 50480
rect 65661 50475 65727 50478
rect 97726 50402 97786 50440
rect 100621 50402 100687 50405
rect 97726 50400 100687 50402
rect 97726 50344 100626 50400
rect 100682 50344 100687 50400
rect 97726 50342 100687 50344
rect 100621 50339 100687 50342
rect 102461 50402 102527 50405
rect 135029 50402 135095 50405
rect 102461 50400 104932 50402
rect 102461 50344 102466 50400
rect 102522 50344 104932 50400
rect 102461 50342 104932 50344
rect 132716 50400 135095 50402
rect 132716 50344 135034 50400
rect 135090 50344 135095 50400
rect 132716 50342 135095 50344
rect 102461 50339 102527 50342
rect 135029 50339 135095 50342
rect 136869 50402 136935 50405
rect 140046 50402 140106 50440
rect 136869 50400 140106 50402
rect 136869 50344 136874 50400
rect 136930 50344 140106 50400
rect 136869 50342 140106 50344
rect 169854 50402 169914 50508
rect 172657 50402 172723 50405
rect 169854 50400 172723 50402
rect 169854 50344 172662 50400
rect 172718 50344 172723 50400
rect 169854 50342 172723 50344
rect 136869 50339 136935 50342
rect 172657 50339 172723 50342
rect 174313 50402 174379 50405
rect 174313 50400 177060 50402
rect 174313 50344 174318 50400
rect 174374 50344 177060 50400
rect 174313 50342 177060 50344
rect 174313 50339 174379 50342
rect 63361 50130 63427 50133
rect 60772 50128 63427 50130
rect 60772 50072 63366 50128
rect 63422 50072 63427 50128
rect 60772 50070 63427 50072
rect 63361 50067 63427 50070
rect 65477 49994 65543 49997
rect 65477 49992 67948 49994
rect 65477 49936 65482 49992
rect 65538 49936 67948 49992
rect 65477 49934 67948 49936
rect 65477 49931 65543 49934
rect 62717 49586 62783 49589
rect 60772 49584 62783 49586
rect 60772 49528 62722 49584
rect 62778 49528 62783 49584
rect 60772 49526 62783 49528
rect 62717 49523 62783 49526
rect 97726 49450 97786 49896
rect 102553 49858 102619 49861
rect 135305 49858 135371 49861
rect 102553 49856 104932 49858
rect 102553 49800 102558 49856
rect 102614 49800 104932 49856
rect 102553 49798 104932 49800
rect 132716 49856 135371 49858
rect 132716 49800 135310 49856
rect 135366 49800 135371 49856
rect 132716 49798 135371 49800
rect 102553 49795 102619 49798
rect 135305 49795 135371 49798
rect 100621 49450 100687 49453
rect 97726 49448 100687 49450
rect 97726 49392 100626 49448
rect 100682 49392 100687 49448
rect 97726 49390 100687 49392
rect 100621 49387 100687 49390
rect 136869 49450 136935 49453
rect 140046 49450 140106 49896
rect 136869 49448 140106 49450
rect 136869 49392 136874 49448
rect 136930 49392 140106 49448
rect 136869 49390 140106 49392
rect 169854 49450 169914 49964
rect 174405 49858 174471 49861
rect 174405 49856 177060 49858
rect 174405 49800 174410 49856
rect 174466 49800 177060 49856
rect 174405 49798 177060 49800
rect 174405 49795 174471 49798
rect 172657 49450 172723 49453
rect 169854 49448 172723 49450
rect 169854 49392 172662 49448
rect 172718 49392 172723 49448
rect 169854 49390 172723 49392
rect 136869 49387 136935 49390
rect 172657 49387 172723 49390
rect 66397 49314 66463 49317
rect 102645 49314 102711 49317
rect 134845 49314 134911 49317
rect 66397 49312 67948 49314
rect 66397 49256 66402 49312
rect 66458 49256 67948 49312
rect 66397 49254 67948 49256
rect 102645 49312 104932 49314
rect 102645 49256 102650 49312
rect 102706 49256 104932 49312
rect 102645 49254 104932 49256
rect 132716 49312 134911 49314
rect 132716 49256 134850 49312
rect 134906 49256 134911 49312
rect 174129 49314 174195 49317
rect 174129 49312 177060 49314
rect 132716 49254 134911 49256
rect 66397 49251 66463 49254
rect 102645 49251 102711 49254
rect 134845 49251 134911 49254
rect 63821 49042 63887 49045
rect 60772 49040 63887 49042
rect 60772 48984 63826 49040
rect 63882 48984 63887 49040
rect 60772 48982 63887 48984
rect 97726 49042 97786 49216
rect 100621 49042 100687 49045
rect 97726 49040 100687 49042
rect 97726 48984 100626 49040
rect 100682 48984 100687 49040
rect 97726 48982 100687 48984
rect 63821 48979 63887 48982
rect 100621 48979 100687 48982
rect 136777 48906 136843 48909
rect 140046 48906 140106 49216
rect 169854 49178 169914 49284
rect 174129 49256 174134 49312
rect 174190 49256 177060 49312
rect 174129 49254 177060 49256
rect 174129 49251 174195 49254
rect 171829 49178 171895 49181
rect 169854 49176 171895 49178
rect 169854 49120 171834 49176
rect 171890 49120 171895 49176
rect 169854 49118 171895 49120
rect 171829 49115 171895 49118
rect 136777 48904 140106 48906
rect 136777 48848 136782 48904
rect 136838 48848 140106 48904
rect 136777 48846 140106 48848
rect 136777 48843 136843 48846
rect 64925 48770 64991 48773
rect 102369 48770 102435 48773
rect 135397 48770 135463 48773
rect 64925 48768 67948 48770
rect 64925 48712 64930 48768
rect 64986 48712 67948 48768
rect 64925 48710 67948 48712
rect 102369 48768 104932 48770
rect 102369 48712 102374 48768
rect 102430 48712 104932 48768
rect 102369 48710 104932 48712
rect 132716 48768 135463 48770
rect 132716 48712 135402 48768
rect 135458 48712 135463 48768
rect 174313 48770 174379 48773
rect 174313 48768 177060 48770
rect 132716 48710 135463 48712
rect 64925 48707 64991 48710
rect 102369 48707 102435 48710
rect 135397 48707 135463 48710
rect 62809 48498 62875 48501
rect 60772 48496 62875 48498
rect 60772 48440 62814 48496
rect 62870 48440 62875 48496
rect 60772 48438 62875 48440
rect 62809 48435 62875 48438
rect 97726 48362 97786 48672
rect 100621 48362 100687 48365
rect 97726 48360 100687 48362
rect 97726 48304 100626 48360
rect 100682 48304 100687 48360
rect 97726 48302 100687 48304
rect 100621 48299 100687 48302
rect 136685 48362 136751 48365
rect 140046 48362 140106 48672
rect 136685 48360 140106 48362
rect 136685 48304 136690 48360
rect 136746 48304 140106 48360
rect 136685 48302 140106 48304
rect 169854 48362 169914 48740
rect 174313 48712 174318 48768
rect 174374 48712 177060 48768
rect 174313 48710 177060 48712
rect 174313 48707 174379 48710
rect 172565 48362 172631 48365
rect 169854 48360 172631 48362
rect 169854 48304 172570 48360
rect 172626 48304 172631 48360
rect 169854 48302 172631 48304
rect 136685 48299 136751 48302
rect 172565 48299 172631 48302
rect 63729 47818 63795 47821
rect 60772 47816 63795 47818
rect 60772 47760 63734 47816
rect 63790 47760 63795 47816
rect 60772 47758 63795 47760
rect 63729 47755 63795 47758
rect 65017 47818 65083 47821
rect 67918 47818 67978 48196
rect 65017 47816 67978 47818
rect 65017 47760 65022 47816
rect 65078 47760 67978 47816
rect 65017 47758 67978 47760
rect 65017 47755 65083 47758
rect 97726 47682 97786 48128
rect 102461 48090 102527 48093
rect 135305 48090 135371 48093
rect 102461 48088 104932 48090
rect 102461 48032 102466 48088
rect 102522 48032 104932 48088
rect 102461 48030 104932 48032
rect 132716 48088 135371 48090
rect 132716 48032 135310 48088
rect 135366 48032 135371 48088
rect 132716 48030 135371 48032
rect 102461 48027 102527 48030
rect 135305 48027 135371 48030
rect 100621 47682 100687 47685
rect 97726 47680 100687 47682
rect 97726 47624 100626 47680
rect 100682 47624 100687 47680
rect 97726 47622 100687 47624
rect 100621 47619 100687 47622
rect 136777 47682 136843 47685
rect 140046 47682 140106 48128
rect 169854 47954 169914 48196
rect 174221 48090 174287 48093
rect 174221 48088 177060 48090
rect 174221 48032 174226 48088
rect 174282 48032 177060 48088
rect 174221 48030 177060 48032
rect 174221 48027 174287 48030
rect 172657 47954 172723 47957
rect 169854 47952 172723 47954
rect 169854 47896 172662 47952
rect 172718 47896 172723 47952
rect 169854 47894 172723 47896
rect 172657 47891 172723 47894
rect 172657 47682 172723 47685
rect 136777 47680 140106 47682
rect 136777 47624 136782 47680
rect 136838 47624 140106 47680
rect 136777 47622 140106 47624
rect 169670 47680 172723 47682
rect 169670 47624 172662 47680
rect 172718 47624 172723 47680
rect 169670 47622 172723 47624
rect 136777 47619 136843 47622
rect 65661 47546 65727 47549
rect 100621 47546 100687 47549
rect 65661 47544 67948 47546
rect 65661 47488 65666 47544
rect 65722 47488 67948 47544
rect 65661 47486 67948 47488
rect 97756 47544 100687 47546
rect 97756 47488 100626 47544
rect 100682 47488 100687 47544
rect 97756 47486 100687 47488
rect 65661 47483 65727 47486
rect 100621 47483 100687 47486
rect 102553 47546 102619 47549
rect 134753 47546 134819 47549
rect 102553 47544 104932 47546
rect 102553 47488 102558 47544
rect 102614 47488 104932 47544
rect 102553 47486 104932 47488
rect 132716 47544 134819 47546
rect 132716 47488 134758 47544
rect 134814 47488 134819 47544
rect 132716 47486 134819 47488
rect 102553 47483 102619 47486
rect 134753 47483 134819 47486
rect 136869 47546 136935 47549
rect 136869 47544 140076 47546
rect 136869 47488 136874 47544
rect 136930 47488 140076 47544
rect 169670 47516 169730 47622
rect 172657 47619 172723 47622
rect 174405 47546 174471 47549
rect 174405 47544 177060 47546
rect 136869 47486 140076 47488
rect 174405 47488 174410 47544
rect 174466 47488 177060 47544
rect 174405 47486 177060 47488
rect 136869 47483 136935 47486
rect 174405 47483 174471 47486
rect 63361 47274 63427 47277
rect 60772 47272 63427 47274
rect 60772 47216 63366 47272
rect 63422 47216 63427 47272
rect 60772 47214 63427 47216
rect 63361 47211 63427 47214
rect 66397 47002 66463 47005
rect 102645 47002 102711 47005
rect 135305 47002 135371 47005
rect 66397 47000 67948 47002
rect 66397 46944 66402 47000
rect 66458 46944 67948 47000
rect 66397 46942 67948 46944
rect 102645 47000 104932 47002
rect 102645 46944 102650 47000
rect 102706 46944 104932 47000
rect 102645 46942 104932 46944
rect 132716 47000 135371 47002
rect 132716 46944 135310 47000
rect 135366 46944 135371 47000
rect 174221 47002 174287 47005
rect 174221 47000 177060 47002
rect 132716 46942 135371 46944
rect 66397 46939 66463 46942
rect 102645 46939 102711 46942
rect 135305 46939 135371 46942
rect 62901 46730 62967 46733
rect 60772 46728 62967 46730
rect 60772 46672 62906 46728
rect 62962 46672 62967 46728
rect 60772 46670 62967 46672
rect 62901 46667 62967 46670
rect 97726 46458 97786 46904
rect 100621 46458 100687 46461
rect 97726 46456 100687 46458
rect 97726 46400 100626 46456
rect 100682 46400 100687 46456
rect 97726 46398 100687 46400
rect 100621 46395 100687 46398
rect 102369 46458 102435 46461
rect 134845 46458 134911 46461
rect 102369 46456 104932 46458
rect 102369 46400 102374 46456
rect 102430 46400 104932 46456
rect 102369 46398 104932 46400
rect 132716 46456 134911 46458
rect 132716 46400 134850 46456
rect 134906 46400 134911 46456
rect 132716 46398 134911 46400
rect 102369 46395 102435 46398
rect 134845 46395 134911 46398
rect 136777 46458 136843 46461
rect 140046 46458 140106 46904
rect 169854 46594 169914 46972
rect 174221 46944 174226 47000
rect 174282 46944 177060 47000
rect 174221 46942 177060 46944
rect 174221 46939 174287 46942
rect 172657 46594 172723 46597
rect 169854 46592 172723 46594
rect 169854 46536 172662 46592
rect 172718 46536 172723 46592
rect 169854 46534 172723 46536
rect 172657 46531 172723 46534
rect 136777 46456 140106 46458
rect 136777 46400 136782 46456
rect 136838 46400 140106 46456
rect 136777 46398 140106 46400
rect 174129 46458 174195 46461
rect 174129 46456 177060 46458
rect 174129 46400 174134 46456
rect 174190 46400 177060 46456
rect 174129 46398 177060 46400
rect 136777 46395 136843 46398
rect 174129 46395 174195 46398
rect 65201 46322 65267 46325
rect 65201 46320 67948 46322
rect 65201 46264 65206 46320
rect 65262 46264 67948 46320
rect 65201 46262 67948 46264
rect 65201 46259 65267 46262
rect 62717 46186 62783 46189
rect 60772 46184 62783 46186
rect 60772 46128 62722 46184
rect 62778 46128 62783 46184
rect 60772 46126 62783 46128
rect 97726 46186 97786 46224
rect 100897 46186 100963 46189
rect 97726 46184 100963 46186
rect 97726 46128 100902 46184
rect 100958 46128 100963 46184
rect 97726 46126 100963 46128
rect 62717 46123 62783 46126
rect 100897 46123 100963 46126
rect 137513 46186 137579 46189
rect 140046 46186 140106 46224
rect 137513 46184 140106 46186
rect 137513 46128 137518 46184
rect 137574 46128 140106 46184
rect 137513 46126 140106 46128
rect 169854 46186 169914 46292
rect 172657 46186 172723 46189
rect 169854 46184 172723 46186
rect 169854 46128 172662 46184
rect 172718 46128 172723 46184
rect 169854 46126 172723 46128
rect 137513 46123 137579 46126
rect 172657 46123 172723 46126
rect 102461 45914 102527 45917
rect 135397 45914 135463 45917
rect 102461 45912 104932 45914
rect 102461 45856 102466 45912
rect 102522 45856 104932 45912
rect 102461 45854 104932 45856
rect 132716 45912 135463 45914
rect 132716 45856 135402 45912
rect 135458 45856 135463 45912
rect 132716 45854 135463 45856
rect 102461 45851 102527 45854
rect 135397 45851 135463 45854
rect 174313 45914 174379 45917
rect 174313 45912 177060 45914
rect 174313 45856 174318 45912
rect 174374 45856 177060 45912
rect 174313 45854 177060 45856
rect 174313 45851 174379 45854
rect 66305 45778 66371 45781
rect 66305 45776 67948 45778
rect 66305 45720 66310 45776
rect 66366 45720 67948 45776
rect 66305 45718 67948 45720
rect 66305 45715 66371 45718
rect 62809 45642 62875 45645
rect 60772 45640 62875 45642
rect 60772 45584 62814 45640
rect 62870 45584 62875 45640
rect 60772 45582 62875 45584
rect 62809 45579 62875 45582
rect 97726 45370 97786 45680
rect 100529 45370 100595 45373
rect 97726 45368 100595 45370
rect 97726 45312 100534 45368
rect 100590 45312 100595 45368
rect 97726 45310 100595 45312
rect 100529 45307 100595 45310
rect 136685 45370 136751 45373
rect 140046 45370 140106 45680
rect 136685 45368 140106 45370
rect 136685 45312 136690 45368
rect 136746 45312 140106 45368
rect 136685 45310 140106 45312
rect 169854 45370 169914 45748
rect 171645 45370 171711 45373
rect 169854 45368 171711 45370
rect 169854 45312 171650 45368
rect 171706 45312 171711 45368
rect 169854 45310 171711 45312
rect 136685 45307 136751 45310
rect 171645 45307 171711 45310
rect 66397 45234 66463 45237
rect 102553 45234 102619 45237
rect 134661 45234 134727 45237
rect 66397 45232 67948 45234
rect 66397 45176 66402 45232
rect 66458 45176 67948 45232
rect 66397 45174 67948 45176
rect 102553 45232 104932 45234
rect 102553 45176 102558 45232
rect 102614 45176 104932 45232
rect 102553 45174 104932 45176
rect 132716 45232 134727 45234
rect 132716 45176 134666 45232
rect 134722 45176 134727 45232
rect 174221 45234 174287 45237
rect 174221 45232 177060 45234
rect 132716 45174 134727 45176
rect 66397 45171 66463 45174
rect 102553 45171 102619 45174
rect 134661 45171 134727 45174
rect 97726 45098 97786 45136
rect 99977 45098 100043 45101
rect 97726 45096 100043 45098
rect 97726 45040 99982 45096
rect 100038 45040 100043 45096
rect 97726 45038 100043 45040
rect 99977 45035 100043 45038
rect 63729 44962 63795 44965
rect 60772 44960 63795 44962
rect 60772 44904 63734 44960
rect 63790 44904 63795 44960
rect 60772 44902 63795 44904
rect 63729 44899 63795 44902
rect 136777 44962 136843 44965
rect 140046 44962 140106 45136
rect 136777 44960 140106 44962
rect 136777 44904 136782 44960
rect 136838 44904 140106 44960
rect 136777 44902 140106 44904
rect 169854 44962 169914 45204
rect 174221 45176 174226 45232
rect 174282 45176 177060 45232
rect 174221 45174 177060 45176
rect 174221 45171 174287 45174
rect 171829 44962 171895 44965
rect 169854 44960 171895 44962
rect 169854 44904 171834 44960
rect 171890 44904 171895 44960
rect 169854 44902 171895 44904
rect 136777 44899 136843 44902
rect 171829 44899 171895 44902
rect 102369 44690 102435 44693
rect 135029 44690 135095 44693
rect 102369 44688 104932 44690
rect 102369 44632 102374 44688
rect 102430 44632 104932 44688
rect 102369 44630 104932 44632
rect 132716 44688 135095 44690
rect 132716 44632 135034 44688
rect 135090 44632 135095 44688
rect 132716 44630 135095 44632
rect 102369 44627 102435 44630
rect 135029 44627 135095 44630
rect 175325 44690 175391 44693
rect 175325 44688 177060 44690
rect 175325 44632 175330 44688
rect 175386 44632 177060 44688
rect 175325 44630 177060 44632
rect 175325 44627 175391 44630
rect 66213 44554 66279 44557
rect 222521 44554 222587 44557
rect 227416 44554 227896 44584
rect 66213 44552 67948 44554
rect 66213 44496 66218 44552
rect 66274 44496 67948 44552
rect 222521 44552 227896 44554
rect 66213 44494 67948 44496
rect 66213 44491 66279 44494
rect 62809 44418 62875 44421
rect 60772 44416 62875 44418
rect 60772 44360 62814 44416
rect 62870 44360 62875 44416
rect 60772 44358 62875 44360
rect 62809 44355 62875 44358
rect 31846 44220 31852 44284
rect 31916 44282 31922 44284
rect 31916 44222 32988 44282
rect 31916 44220 31922 44222
rect 97726 44146 97786 44456
rect 99885 44146 99951 44149
rect 97726 44144 99951 44146
rect 97726 44088 99890 44144
rect 99946 44088 99951 44144
rect 97726 44086 99951 44088
rect 99885 44083 99951 44086
rect 102461 44146 102527 44149
rect 135397 44146 135463 44149
rect 102461 44144 104932 44146
rect 102461 44088 102466 44144
rect 102522 44088 104932 44144
rect 102461 44086 104932 44088
rect 132716 44144 135463 44146
rect 132716 44088 135402 44144
rect 135458 44088 135463 44144
rect 132716 44086 135463 44088
rect 102461 44083 102527 44086
rect 135397 44083 135463 44086
rect 136777 44146 136843 44149
rect 140046 44146 140106 44456
rect 136777 44144 140106 44146
rect 136777 44088 136782 44144
rect 136838 44088 140106 44144
rect 136777 44086 140106 44088
rect 169854 44146 169914 44524
rect 222521 44496 222526 44552
rect 222582 44496 227896 44552
rect 222521 44494 227896 44496
rect 222521 44491 222587 44494
rect 227416 44464 227896 44494
rect 172657 44146 172723 44149
rect 169854 44144 172723 44146
rect 169854 44088 172662 44144
rect 172718 44088 172723 44144
rect 169854 44086 172723 44088
rect 136777 44083 136843 44086
rect 172657 44083 172723 44086
rect 175417 44146 175483 44149
rect 175417 44144 177060 44146
rect 175417 44088 175422 44144
rect 175478 44088 177060 44144
rect 175417 44086 177060 44088
rect 175417 44083 175483 44086
rect 66397 44010 66463 44013
rect 66397 44008 67948 44010
rect 66397 43952 66402 44008
rect 66458 43952 67948 44008
rect 66397 43950 67948 43952
rect 66397 43947 66463 43950
rect 63729 43874 63795 43877
rect 60772 43872 63795 43874
rect 60772 43816 63734 43872
rect 63790 43816 63795 43872
rect 60772 43814 63795 43816
rect 63729 43811 63795 43814
rect 97726 43466 97786 43912
rect 102553 43602 102619 43605
rect 135029 43602 135095 43605
rect 102553 43600 104932 43602
rect 102553 43544 102558 43600
rect 102614 43544 104932 43600
rect 102553 43542 104932 43544
rect 132716 43600 135095 43602
rect 132716 43544 135034 43600
rect 135090 43544 135095 43600
rect 132716 43542 135095 43544
rect 102553 43539 102619 43542
rect 135029 43539 135095 43542
rect 100621 43466 100687 43469
rect 97726 43464 100687 43466
rect 97726 43408 100626 43464
rect 100682 43408 100687 43464
rect 97726 43406 100687 43408
rect 100621 43403 100687 43406
rect 136869 43466 136935 43469
rect 140046 43466 140106 43912
rect 169854 43602 169914 43980
rect 172565 43602 172631 43605
rect 169854 43600 172631 43602
rect 169854 43544 172570 43600
rect 172626 43544 172631 43600
rect 169854 43542 172631 43544
rect 172565 43539 172631 43542
rect 174773 43602 174839 43605
rect 174773 43600 177060 43602
rect 174773 43544 174778 43600
rect 174834 43544 177060 43600
rect 174773 43542 177060 43544
rect 174773 43539 174839 43542
rect 136869 43464 140106 43466
rect 136869 43408 136874 43464
rect 136930 43408 140106 43464
rect 136869 43406 140106 43408
rect 136869 43403 136935 43406
rect 63637 43330 63703 43333
rect 60772 43328 63703 43330
rect 60772 43272 63642 43328
rect 63698 43272 63703 43328
rect 60772 43270 63703 43272
rect 63637 43267 63703 43270
rect 66305 43330 66371 43333
rect 66305 43328 67948 43330
rect 66305 43272 66310 43328
rect 66366 43272 67948 43328
rect 66305 43270 67948 43272
rect 66305 43267 66371 43270
rect 97726 42922 97786 43232
rect 102277 43058 102343 43061
rect 135397 43058 135463 43061
rect 102277 43056 104932 43058
rect 102277 43000 102282 43056
rect 102338 43000 104932 43056
rect 102277 42998 104932 43000
rect 132716 43056 135463 43058
rect 132716 43000 135402 43056
rect 135458 43000 135463 43056
rect 132716 42998 135463 43000
rect 102277 42995 102343 42998
rect 135397 42995 135463 42998
rect 100621 42922 100687 42925
rect 97726 42920 100687 42922
rect 97726 42864 100626 42920
rect 100682 42864 100687 42920
rect 97726 42862 100687 42864
rect 100621 42859 100687 42862
rect 136685 42922 136751 42925
rect 140046 42922 140106 43232
rect 136685 42920 140106 42922
rect 136685 42864 136690 42920
rect 136746 42864 140106 42920
rect 136685 42862 140106 42864
rect 169854 42922 169914 43300
rect 174037 43058 174103 43061
rect 174037 43056 177060 43058
rect 174037 43000 174042 43056
rect 174098 43000 177060 43056
rect 174037 42998 177060 43000
rect 174037 42995 174103 42998
rect 172197 42922 172263 42925
rect 169854 42920 172263 42922
rect 169854 42864 172202 42920
rect 172258 42864 172263 42920
rect 169854 42862 172263 42864
rect 136685 42859 136751 42862
rect 172197 42859 172263 42862
rect 63729 42786 63795 42789
rect 60772 42784 63795 42786
rect 60772 42728 63734 42784
rect 63790 42728 63795 42784
rect 60772 42726 63795 42728
rect 63729 42723 63795 42726
rect 66397 42786 66463 42789
rect 66397 42784 67948 42786
rect 66397 42728 66402 42784
rect 66458 42728 67948 42784
rect 66397 42726 67948 42728
rect 66397 42723 66463 42726
rect 63821 42514 63887 42517
rect 60742 42512 63887 42514
rect 60742 42456 63826 42512
rect 63882 42456 63887 42512
rect 60742 42454 63887 42456
rect 60742 42076 60802 42454
rect 63821 42451 63887 42454
rect 97726 42378 97786 42688
rect 100621 42378 100687 42381
rect 97726 42376 100687 42378
rect 97726 42320 100626 42376
rect 100682 42320 100687 42376
rect 97726 42318 100687 42320
rect 100621 42315 100687 42318
rect 102369 42378 102435 42381
rect 134937 42378 135003 42381
rect 102369 42376 104932 42378
rect 102369 42320 102374 42376
rect 102430 42320 104932 42376
rect 102369 42318 104932 42320
rect 132716 42376 135003 42378
rect 132716 42320 134942 42376
rect 134998 42320 135003 42376
rect 132716 42318 135003 42320
rect 102369 42315 102435 42318
rect 134937 42315 135003 42318
rect 136869 42378 136935 42381
rect 140046 42378 140106 42688
rect 136869 42376 140106 42378
rect 136869 42320 136874 42376
rect 136930 42320 140106 42376
rect 136869 42318 140106 42320
rect 169854 42378 169914 42756
rect 172657 42378 172723 42381
rect 169854 42376 172723 42378
rect 169854 42320 172662 42376
rect 172718 42320 172723 42376
rect 169854 42318 172723 42320
rect 136869 42315 136935 42318
rect 172657 42315 172723 42318
rect 174129 42378 174195 42381
rect 174129 42376 177060 42378
rect 174129 42320 174134 42376
rect 174190 42320 177060 42376
rect 174129 42318 177060 42320
rect 174129 42315 174195 42318
rect 66397 42242 66463 42245
rect 66397 42240 67948 42242
rect 66397 42184 66402 42240
rect 66458 42184 67948 42240
rect 66397 42182 67948 42184
rect 66397 42179 66463 42182
rect 97726 42106 97786 42144
rect 100621 42106 100687 42109
rect 97726 42104 100687 42106
rect 97726 42048 100626 42104
rect 100682 42048 100687 42104
rect 97726 42046 100687 42048
rect 100621 42043 100687 42046
rect 136777 42106 136843 42109
rect 140046 42106 140106 42144
rect 136777 42104 140106 42106
rect 136777 42048 136782 42104
rect 136838 42048 140106 42104
rect 136777 42046 140106 42048
rect 169854 42106 169914 42212
rect 172657 42106 172723 42109
rect 169854 42104 172723 42106
rect 169854 42048 172662 42104
rect 172718 42048 172723 42104
rect 169854 42046 172723 42048
rect 136777 42043 136843 42046
rect 172657 42043 172723 42046
rect 102553 41834 102619 41837
rect 135305 41834 135371 41837
rect 102553 41832 104932 41834
rect 102553 41776 102558 41832
rect 102614 41776 104932 41832
rect 102553 41774 104932 41776
rect 132716 41832 135371 41834
rect 132716 41776 135310 41832
rect 135366 41776 135371 41832
rect 132716 41774 135371 41776
rect 102553 41771 102619 41774
rect 135305 41771 135371 41774
rect 174221 41834 174287 41837
rect 174221 41832 177060 41834
rect 174221 41776 174226 41832
rect 174282 41776 177060 41832
rect 174221 41774 177060 41776
rect 174221 41771 174287 41774
rect 63729 41562 63795 41565
rect 60772 41560 63795 41562
rect 60772 41504 63734 41560
rect 63790 41504 63795 41560
rect 60772 41502 63795 41504
rect 63729 41499 63795 41502
rect 9896 41290 10376 41320
rect 11933 41290 11999 41293
rect 9896 41288 11999 41290
rect 9896 41232 11938 41288
rect 11994 41232 11999 41288
rect 9896 41230 11999 41232
rect 9896 41200 10376 41230
rect 11933 41227 11999 41230
rect 102461 41290 102527 41293
rect 135397 41290 135463 41293
rect 102461 41288 104932 41290
rect 102461 41232 102466 41288
rect 102522 41232 104932 41288
rect 102461 41230 104932 41232
rect 132716 41288 135463 41290
rect 132716 41232 135402 41288
rect 135458 41232 135463 41288
rect 132716 41230 135463 41232
rect 102461 41227 102527 41230
rect 135397 41227 135463 41230
rect 174313 41290 174379 41293
rect 174313 41288 177060 41290
rect 174313 41232 174318 41288
rect 174374 41232 177060 41288
rect 174313 41230 177060 41232
rect 174313 41227 174379 41230
rect 63821 41018 63887 41021
rect 60772 41016 63887 41018
rect 60772 40960 63826 41016
rect 63882 40960 63887 41016
rect 60772 40958 63887 40960
rect 63821 40955 63887 40958
rect 102369 40746 102435 40749
rect 134845 40746 134911 40749
rect 102369 40744 104932 40746
rect 102369 40688 102374 40744
rect 102430 40688 104932 40744
rect 102369 40686 104932 40688
rect 132716 40744 134911 40746
rect 132716 40688 134850 40744
rect 134906 40688 134911 40744
rect 132716 40686 134911 40688
rect 102369 40683 102435 40686
rect 134845 40683 134911 40686
rect 174129 40746 174195 40749
rect 174129 40744 177060 40746
rect 174129 40688 174134 40744
rect 174190 40688 177060 40744
rect 174129 40686 177060 40688
rect 174129 40683 174195 40686
rect 63177 40474 63243 40477
rect 60772 40472 63243 40474
rect 60772 40416 63182 40472
rect 63238 40416 63243 40472
rect 60772 40414 63243 40416
rect 63177 40411 63243 40414
rect 66254 40412 66260 40476
rect 66324 40474 66330 40476
rect 66397 40474 66463 40477
rect 93854 40474 93860 40476
rect 66324 40472 93860 40474
rect 66324 40416 66402 40472
rect 66458 40416 93860 40472
rect 66324 40414 93860 40416
rect 66324 40412 66330 40414
rect 66397 40411 66463 40414
rect 93854 40412 93860 40414
rect 93924 40474 93930 40476
rect 93997 40474 94063 40477
rect 93924 40472 94063 40474
rect 93924 40416 94002 40472
rect 94058 40416 94063 40472
rect 93924 40414 94063 40416
rect 93924 40412 93930 40414
rect 93997 40411 94063 40414
rect 102369 40202 102435 40205
rect 102369 40200 104932 40202
rect 102369 40144 102374 40200
rect 102430 40144 104932 40200
rect 102369 40142 104932 40144
rect 102369 40139 102435 40142
rect 109637 40068 109703 40069
rect 109637 40066 109684 40068
rect 109592 40064 109684 40066
rect 109592 40008 109642 40064
rect 109592 40006 109684 40008
rect 109637 40004 109684 40006
rect 109748 40004 109754 40068
rect 109637 40003 109703 40004
rect 60742 39522 60802 39832
rect 132686 39658 132746 40104
rect 136910 39732 136916 39796
rect 136980 39794 136986 39796
rect 138157 39794 138223 39797
rect 166033 39794 166099 39797
rect 166166 39794 166172 39796
rect 136980 39792 166172 39794
rect 136980 39736 138162 39792
rect 138218 39736 166038 39792
rect 166094 39736 166172 39792
rect 136980 39734 166172 39736
rect 136980 39732 136986 39734
rect 138157 39731 138223 39734
rect 166033 39731 166099 39734
rect 166166 39732 166172 39734
rect 166236 39732 166242 39796
rect 134477 39658 134543 39661
rect 132686 39656 134543 39658
rect 132686 39600 134482 39656
rect 134538 39600 134543 39656
rect 132686 39598 134543 39600
rect 134477 39595 134543 39598
rect 62809 39522 62875 39525
rect 60742 39520 62875 39522
rect 60742 39464 62814 39520
rect 62870 39464 62875 39520
rect 60742 39462 62875 39464
rect 62809 39459 62875 39462
rect 174129 39522 174195 39525
rect 177030 39522 177090 40104
rect 181397 40068 181463 40069
rect 181397 40066 181444 40068
rect 181352 40064 181444 40066
rect 181352 40008 181402 40064
rect 181352 40006 181444 40008
rect 181397 40004 181444 40006
rect 181508 40004 181514 40068
rect 181397 40003 181463 40004
rect 174129 39520 177090 39522
rect 174129 39464 174134 39520
rect 174190 39464 177090 39520
rect 174129 39462 177090 39464
rect 174129 39459 174195 39462
rect 136869 33402 136935 33405
rect 136869 33400 140106 33402
rect 136869 33344 136874 33400
rect 136930 33344 140106 33400
rect 136869 33342 140106 33344
rect 136869 33339 136935 33342
rect 140046 32760 140106 33342
rect 66213 32722 66279 32725
rect 66213 32720 67948 32722
rect 66213 32664 66218 32720
rect 66274 32664 67948 32720
rect 66213 32662 67948 32664
rect 66213 32659 66279 32662
rect 138065 25106 138131 25109
rect 138065 25104 140106 25106
rect 138065 25048 138070 25104
rect 138126 25048 140106 25104
rect 138065 25046 140106 25048
rect 138065 25043 138131 25046
rect 140046 24736 140106 25046
rect 66305 24698 66371 24701
rect 66305 24696 67948 24698
rect 66305 24640 66310 24696
rect 66366 24640 67948 24696
rect 66305 24638 67948 24640
rect 66305 24635 66371 24638
rect 222705 20754 222771 20757
rect 227416 20754 227896 20784
rect 222705 20752 227896 20754
rect 222705 20696 222710 20752
rect 222766 20696 227896 20752
rect 222705 20694 227896 20696
rect 222705 20691 222771 20694
rect 227416 20664 227896 20694
rect 9896 19666 10376 19696
rect 13313 19666 13379 19669
rect 9896 19664 13379 19666
rect 9896 19608 13318 19664
rect 13374 19608 13379 19664
rect 9896 19606 13379 19608
rect 9896 19576 10376 19606
rect 13313 19603 13379 19606
rect 138157 17082 138223 17085
rect 138157 17080 140106 17082
rect 138157 17024 138162 17080
rect 138218 17024 140106 17080
rect 138157 17022 140106 17024
rect 138157 17019 138223 17022
rect 140046 16848 140106 17022
rect 66397 16810 66463 16813
rect 66397 16808 67948 16810
rect 66397 16752 66402 16808
rect 66458 16752 67948 16808
rect 66397 16750 67948 16752
rect 66397 16747 66463 16750
<< via3 >>
rect 37924 217212 37988 217276
rect 204260 215852 204324 215916
rect 204812 211636 204876 211700
rect 207572 192460 207636 192524
rect 207572 192324 207636 192388
rect 207204 182804 207268 182868
rect 207388 172876 207452 172940
rect 207572 172876 207636 172940
rect 207572 163220 207636 163284
rect 207388 153760 207452 153764
rect 207388 153704 207438 153760
rect 207438 153704 207452 153760
rect 207388 153700 207452 153704
rect 207388 152264 207452 152268
rect 207388 152208 207438 152264
rect 207438 152208 207452 152264
rect 207388 152204 207452 152208
rect 37924 151524 37988 151588
rect 207756 142684 207820 142748
rect 101036 142548 101100 142612
rect 167276 142548 167340 142612
rect 207756 142548 207820 142612
rect 71044 141868 71108 141932
rect 146300 141868 146364 141932
rect 31852 141384 31916 141388
rect 31852 141328 31866 141384
rect 31866 141328 31916 141384
rect 31852 141324 31916 141328
rect 94228 141324 94292 141388
rect 101404 131396 101468 131460
rect 21548 127588 21612 127652
rect 31852 118476 31916 118540
rect 71044 113580 71108 113644
rect 142988 113580 143052 113644
rect 167276 113580 167340 113644
rect 56876 113232 56940 113236
rect 56876 113176 56926 113232
rect 56926 113176 56940 113232
rect 56876 113172 56940 113176
rect 73068 113172 73132 113236
rect 94228 112628 94292 112692
rect 129740 77540 129804 77604
rect 101404 71208 101468 71212
rect 101404 71152 101418 71208
rect 101418 71152 101468 71208
rect 101404 71148 101468 71152
rect 101036 71012 101100 71076
rect 31852 69440 31916 69444
rect 31852 69384 31902 69440
rect 31902 69384 31916 69440
rect 31852 69380 31916 69384
rect 201500 69244 201564 69308
rect 31852 44220 31916 44284
rect 66260 40412 66324 40476
rect 93860 40412 93924 40476
rect 109684 40064 109748 40068
rect 109684 40008 109698 40064
rect 109698 40008 109748 40064
rect 109684 40004 109748 40008
rect 136916 39732 136980 39796
rect 166172 39732 166236 39796
rect 181444 40064 181508 40068
rect 181444 40008 181458 40064
rect 181458 40008 181508 40064
rect 181444 40004 181508 40008
<< metal4 >>
rect 0 255254 4000 255376
rect 0 255018 122 255254
rect 358 255018 442 255254
rect 678 255018 762 255254
rect 998 255018 1082 255254
rect 1318 255018 1402 255254
rect 1638 255018 1722 255254
rect 1958 255018 2042 255254
rect 2278 255018 2362 255254
rect 2598 255018 2682 255254
rect 2918 255018 3002 255254
rect 3238 255018 3322 255254
rect 3558 255018 3642 255254
rect 3878 255018 4000 255254
rect 0 254934 4000 255018
rect 0 254698 122 254934
rect 358 254698 442 254934
rect 678 254698 762 254934
rect 998 254698 1082 254934
rect 1318 254698 1402 254934
rect 1638 254698 1722 254934
rect 1958 254698 2042 254934
rect 2278 254698 2362 254934
rect 2598 254698 2682 254934
rect 2918 254698 3002 254934
rect 3238 254698 3322 254934
rect 3558 254698 3642 254934
rect 3878 254698 4000 254934
rect 0 254614 4000 254698
rect 0 254378 122 254614
rect 358 254378 442 254614
rect 678 254378 762 254614
rect 998 254378 1082 254614
rect 1318 254378 1402 254614
rect 1638 254378 1722 254614
rect 1958 254378 2042 254614
rect 2278 254378 2362 254614
rect 2598 254378 2682 254614
rect 2918 254378 3002 254614
rect 3238 254378 3322 254614
rect 3558 254378 3642 254614
rect 3878 254378 4000 254614
rect 0 254294 4000 254378
rect 0 254058 122 254294
rect 358 254058 442 254294
rect 678 254058 762 254294
rect 998 254058 1082 254294
rect 1318 254058 1402 254294
rect 1638 254058 1722 254294
rect 1958 254058 2042 254294
rect 2278 254058 2362 254294
rect 2598 254058 2682 254294
rect 2918 254058 3002 254294
rect 3238 254058 3322 254294
rect 3558 254058 3642 254294
rect 3878 254058 4000 254294
rect 0 253974 4000 254058
rect 0 253738 122 253974
rect 358 253738 442 253974
rect 678 253738 762 253974
rect 998 253738 1082 253974
rect 1318 253738 1402 253974
rect 1638 253738 1722 253974
rect 1958 253738 2042 253974
rect 2278 253738 2362 253974
rect 2598 253738 2682 253974
rect 2918 253738 3002 253974
rect 3238 253738 3322 253974
rect 3558 253738 3642 253974
rect 3878 253738 4000 253974
rect 0 253654 4000 253738
rect 0 253418 122 253654
rect 358 253418 442 253654
rect 678 253418 762 253654
rect 998 253418 1082 253654
rect 1318 253418 1402 253654
rect 1638 253418 1722 253654
rect 1958 253418 2042 253654
rect 2278 253418 2362 253654
rect 2598 253418 2682 253654
rect 2918 253418 3002 253654
rect 3238 253418 3322 253654
rect 3558 253418 3642 253654
rect 3878 253418 4000 253654
rect 0 253334 4000 253418
rect 0 253098 122 253334
rect 358 253098 442 253334
rect 678 253098 762 253334
rect 998 253098 1082 253334
rect 1318 253098 1402 253334
rect 1638 253098 1722 253334
rect 1958 253098 2042 253334
rect 2278 253098 2362 253334
rect 2598 253098 2682 253334
rect 2918 253098 3002 253334
rect 3238 253098 3322 253334
rect 3558 253098 3642 253334
rect 3878 253098 4000 253334
rect 0 253014 4000 253098
rect 0 252778 122 253014
rect 358 252778 442 253014
rect 678 252778 762 253014
rect 998 252778 1082 253014
rect 1318 252778 1402 253014
rect 1638 252778 1722 253014
rect 1958 252778 2042 253014
rect 2278 252778 2362 253014
rect 2598 252778 2682 253014
rect 2918 252778 3002 253014
rect 3238 252778 3322 253014
rect 3558 252778 3642 253014
rect 3878 252778 4000 253014
rect 0 252694 4000 252778
rect 0 252458 122 252694
rect 358 252458 442 252694
rect 678 252458 762 252694
rect 998 252458 1082 252694
rect 1318 252458 1402 252694
rect 1638 252458 1722 252694
rect 1958 252458 2042 252694
rect 2278 252458 2362 252694
rect 2598 252458 2682 252694
rect 2918 252458 3002 252694
rect 3238 252458 3322 252694
rect 3558 252458 3642 252694
rect 3878 252458 4000 252694
rect 0 252374 4000 252458
rect 0 252138 122 252374
rect 358 252138 442 252374
rect 678 252138 762 252374
rect 998 252138 1082 252374
rect 1318 252138 1402 252374
rect 1638 252138 1722 252374
rect 1958 252138 2042 252374
rect 2278 252138 2362 252374
rect 2598 252138 2682 252374
rect 2918 252138 3002 252374
rect 3238 252138 3322 252374
rect 3558 252138 3642 252374
rect 3878 252138 4000 252374
rect 0 252054 4000 252138
rect 0 251818 122 252054
rect 358 251818 442 252054
rect 678 251818 762 252054
rect 998 251818 1082 252054
rect 1318 251818 1402 252054
rect 1638 251818 1722 252054
rect 1958 251818 2042 252054
rect 2278 251818 2362 252054
rect 2598 251818 2682 252054
rect 2918 251818 3002 252054
rect 3238 251818 3322 252054
rect 3558 251818 3642 252054
rect 3878 251818 4000 252054
rect 0 251734 4000 251818
rect 0 251498 122 251734
rect 358 251498 442 251734
rect 678 251498 762 251734
rect 998 251498 1082 251734
rect 1318 251498 1402 251734
rect 1638 251498 1722 251734
rect 1958 251498 2042 251734
rect 2278 251498 2362 251734
rect 2598 251498 2682 251734
rect 2918 251498 3002 251734
rect 3238 251498 3322 251734
rect 3558 251498 3642 251734
rect 3878 251498 4000 251734
rect 0 228918 4000 251498
rect 233740 255254 237740 255376
rect 233740 255018 233862 255254
rect 234098 255018 234182 255254
rect 234418 255018 234502 255254
rect 234738 255018 234822 255254
rect 235058 255018 235142 255254
rect 235378 255018 235462 255254
rect 235698 255018 235782 255254
rect 236018 255018 236102 255254
rect 236338 255018 236422 255254
rect 236658 255018 236742 255254
rect 236978 255018 237062 255254
rect 237298 255018 237382 255254
rect 237618 255018 237740 255254
rect 233740 254934 237740 255018
rect 233740 254698 233862 254934
rect 234098 254698 234182 254934
rect 234418 254698 234502 254934
rect 234738 254698 234822 254934
rect 235058 254698 235142 254934
rect 235378 254698 235462 254934
rect 235698 254698 235782 254934
rect 236018 254698 236102 254934
rect 236338 254698 236422 254934
rect 236658 254698 236742 254934
rect 236978 254698 237062 254934
rect 237298 254698 237382 254934
rect 237618 254698 237740 254934
rect 233740 254614 237740 254698
rect 233740 254378 233862 254614
rect 234098 254378 234182 254614
rect 234418 254378 234502 254614
rect 234738 254378 234822 254614
rect 235058 254378 235142 254614
rect 235378 254378 235462 254614
rect 235698 254378 235782 254614
rect 236018 254378 236102 254614
rect 236338 254378 236422 254614
rect 236658 254378 236742 254614
rect 236978 254378 237062 254614
rect 237298 254378 237382 254614
rect 237618 254378 237740 254614
rect 233740 254294 237740 254378
rect 233740 254058 233862 254294
rect 234098 254058 234182 254294
rect 234418 254058 234502 254294
rect 234738 254058 234822 254294
rect 235058 254058 235142 254294
rect 235378 254058 235462 254294
rect 235698 254058 235782 254294
rect 236018 254058 236102 254294
rect 236338 254058 236422 254294
rect 236658 254058 236742 254294
rect 236978 254058 237062 254294
rect 237298 254058 237382 254294
rect 237618 254058 237740 254294
rect 233740 253974 237740 254058
rect 233740 253738 233862 253974
rect 234098 253738 234182 253974
rect 234418 253738 234502 253974
rect 234738 253738 234822 253974
rect 235058 253738 235142 253974
rect 235378 253738 235462 253974
rect 235698 253738 235782 253974
rect 236018 253738 236102 253974
rect 236338 253738 236422 253974
rect 236658 253738 236742 253974
rect 236978 253738 237062 253974
rect 237298 253738 237382 253974
rect 237618 253738 237740 253974
rect 233740 253654 237740 253738
rect 233740 253418 233862 253654
rect 234098 253418 234182 253654
rect 234418 253418 234502 253654
rect 234738 253418 234822 253654
rect 235058 253418 235142 253654
rect 235378 253418 235462 253654
rect 235698 253418 235782 253654
rect 236018 253418 236102 253654
rect 236338 253418 236422 253654
rect 236658 253418 236742 253654
rect 236978 253418 237062 253654
rect 237298 253418 237382 253654
rect 237618 253418 237740 253654
rect 233740 253334 237740 253418
rect 233740 253098 233862 253334
rect 234098 253098 234182 253334
rect 234418 253098 234502 253334
rect 234738 253098 234822 253334
rect 235058 253098 235142 253334
rect 235378 253098 235462 253334
rect 235698 253098 235782 253334
rect 236018 253098 236102 253334
rect 236338 253098 236422 253334
rect 236658 253098 236742 253334
rect 236978 253098 237062 253334
rect 237298 253098 237382 253334
rect 237618 253098 237740 253334
rect 233740 253014 237740 253098
rect 233740 252778 233862 253014
rect 234098 252778 234182 253014
rect 234418 252778 234502 253014
rect 234738 252778 234822 253014
rect 235058 252778 235142 253014
rect 235378 252778 235462 253014
rect 235698 252778 235782 253014
rect 236018 252778 236102 253014
rect 236338 252778 236422 253014
rect 236658 252778 236742 253014
rect 236978 252778 237062 253014
rect 237298 252778 237382 253014
rect 237618 252778 237740 253014
rect 233740 252694 237740 252778
rect 233740 252458 233862 252694
rect 234098 252458 234182 252694
rect 234418 252458 234502 252694
rect 234738 252458 234822 252694
rect 235058 252458 235142 252694
rect 235378 252458 235462 252694
rect 235698 252458 235782 252694
rect 236018 252458 236102 252694
rect 236338 252458 236422 252694
rect 236658 252458 236742 252694
rect 236978 252458 237062 252694
rect 237298 252458 237382 252694
rect 237618 252458 237740 252694
rect 233740 252374 237740 252458
rect 233740 252138 233862 252374
rect 234098 252138 234182 252374
rect 234418 252138 234502 252374
rect 234738 252138 234822 252374
rect 235058 252138 235142 252374
rect 235378 252138 235462 252374
rect 235698 252138 235782 252374
rect 236018 252138 236102 252374
rect 236338 252138 236422 252374
rect 236658 252138 236742 252374
rect 236978 252138 237062 252374
rect 237298 252138 237382 252374
rect 237618 252138 237740 252374
rect 233740 252054 237740 252138
rect 233740 251818 233862 252054
rect 234098 251818 234182 252054
rect 234418 251818 234502 252054
rect 234738 251818 234822 252054
rect 235058 251818 235142 252054
rect 235378 251818 235462 252054
rect 235698 251818 235782 252054
rect 236018 251818 236102 252054
rect 236338 251818 236422 252054
rect 236658 251818 236742 252054
rect 236978 251818 237062 252054
rect 237298 251818 237382 252054
rect 237618 251818 237740 252054
rect 233740 251734 237740 251818
rect 233740 251498 233862 251734
rect 234098 251498 234182 251734
rect 234418 251498 234502 251734
rect 234738 251498 234822 251734
rect 235058 251498 235142 251734
rect 235378 251498 235462 251734
rect 235698 251498 235782 251734
rect 236018 251498 236102 251734
rect 236338 251498 236422 251734
rect 236658 251498 236742 251734
rect 236978 251498 237062 251734
rect 237298 251498 237382 251734
rect 237618 251498 237740 251734
rect 0 228682 122 228918
rect 358 228682 442 228918
rect 678 228682 762 228918
rect 998 228682 1082 228918
rect 1318 228682 1402 228918
rect 1638 228682 1722 228918
rect 1958 228682 2042 228918
rect 2278 228682 2362 228918
rect 2598 228682 2682 228918
rect 2918 228682 3002 228918
rect 3238 228682 3322 228918
rect 3558 228682 3642 228918
rect 3878 228682 4000 228918
rect 0 206518 4000 228682
rect 0 206282 122 206518
rect 358 206282 442 206518
rect 678 206282 762 206518
rect 998 206282 1082 206518
rect 1318 206282 1402 206518
rect 1638 206282 1722 206518
rect 1958 206282 2042 206518
rect 2278 206282 2362 206518
rect 2598 206282 2682 206518
rect 2918 206282 3002 206518
rect 3238 206282 3322 206518
rect 3558 206282 3642 206518
rect 3878 206282 4000 206518
rect 0 184118 4000 206282
rect 0 183882 122 184118
rect 358 183882 442 184118
rect 678 183882 762 184118
rect 998 183882 1082 184118
rect 1318 183882 1402 184118
rect 1638 183882 1722 184118
rect 1958 183882 2042 184118
rect 2278 183882 2362 184118
rect 2598 183882 2682 184118
rect 2918 183882 3002 184118
rect 3238 183882 3322 184118
rect 3558 183882 3642 184118
rect 3878 183882 4000 184118
rect 0 161718 4000 183882
rect 0 161482 122 161718
rect 358 161482 442 161718
rect 678 161482 762 161718
rect 998 161482 1082 161718
rect 1318 161482 1402 161718
rect 1638 161482 1722 161718
rect 1958 161482 2042 161718
rect 2278 161482 2362 161718
rect 2598 161482 2682 161718
rect 2918 161482 3002 161718
rect 3238 161482 3322 161718
rect 3558 161482 3642 161718
rect 3878 161482 4000 161718
rect 0 139318 4000 161482
rect 0 139082 122 139318
rect 358 139082 442 139318
rect 678 139082 762 139318
rect 998 139082 1082 139318
rect 1318 139082 1402 139318
rect 1638 139082 1722 139318
rect 1958 139082 2042 139318
rect 2278 139082 2362 139318
rect 2598 139082 2682 139318
rect 2918 139082 3002 139318
rect 3238 139082 3322 139318
rect 3558 139082 3642 139318
rect 3878 139082 4000 139318
rect 0 116918 4000 139082
rect 0 116682 122 116918
rect 358 116682 442 116918
rect 678 116682 762 116918
rect 998 116682 1082 116918
rect 1318 116682 1402 116918
rect 1638 116682 1722 116918
rect 1958 116682 2042 116918
rect 2278 116682 2362 116918
rect 2598 116682 2682 116918
rect 2918 116682 3002 116918
rect 3238 116682 3322 116918
rect 3558 116682 3642 116918
rect 3878 116682 4000 116918
rect 0 94518 4000 116682
rect 0 94282 122 94518
rect 358 94282 442 94518
rect 678 94282 762 94518
rect 998 94282 1082 94518
rect 1318 94282 1402 94518
rect 1638 94282 1722 94518
rect 1958 94282 2042 94518
rect 2278 94282 2362 94518
rect 2598 94282 2682 94518
rect 2918 94282 3002 94518
rect 3238 94282 3322 94518
rect 3558 94282 3642 94518
rect 3878 94282 4000 94518
rect 0 72118 4000 94282
rect 0 71882 122 72118
rect 358 71882 442 72118
rect 678 71882 762 72118
rect 998 71882 1082 72118
rect 1318 71882 1402 72118
rect 1638 71882 1722 72118
rect 1958 71882 2042 72118
rect 2278 71882 2362 72118
rect 2598 71882 2682 72118
rect 2918 71882 3002 72118
rect 3238 71882 3322 72118
rect 3558 71882 3642 72118
rect 3878 71882 4000 72118
rect 0 49718 4000 71882
rect 0 49482 122 49718
rect 358 49482 442 49718
rect 678 49482 762 49718
rect 998 49482 1082 49718
rect 1318 49482 1402 49718
rect 1638 49482 1722 49718
rect 1958 49482 2042 49718
rect 2278 49482 2362 49718
rect 2598 49482 2682 49718
rect 2918 49482 3002 49718
rect 3238 49482 3322 49718
rect 3558 49482 3642 49718
rect 3878 49482 4000 49718
rect 0 27318 4000 49482
rect 0 27082 122 27318
rect 358 27082 442 27318
rect 678 27082 762 27318
rect 998 27082 1082 27318
rect 1318 27082 1402 27318
rect 1638 27082 1722 27318
rect 1958 27082 2042 27318
rect 2278 27082 2362 27318
rect 2598 27082 2682 27318
rect 2918 27082 3002 27318
rect 3238 27082 3322 27318
rect 3558 27082 3642 27318
rect 3878 27082 4000 27318
rect 0 3878 4000 27082
rect 5000 250254 9000 250376
rect 5000 250018 5122 250254
rect 5358 250018 5442 250254
rect 5678 250018 5762 250254
rect 5998 250018 6082 250254
rect 6318 250018 6402 250254
rect 6638 250018 6722 250254
rect 6958 250018 7042 250254
rect 7278 250018 7362 250254
rect 7598 250018 7682 250254
rect 7918 250018 8002 250254
rect 8238 250018 8322 250254
rect 8558 250018 8642 250254
rect 8878 250018 9000 250254
rect 5000 249934 9000 250018
rect 5000 249698 5122 249934
rect 5358 249698 5442 249934
rect 5678 249698 5762 249934
rect 5998 249698 6082 249934
rect 6318 249698 6402 249934
rect 6638 249698 6722 249934
rect 6958 249698 7042 249934
rect 7278 249698 7362 249934
rect 7598 249698 7682 249934
rect 7918 249698 8002 249934
rect 8238 249698 8322 249934
rect 8558 249698 8642 249934
rect 8878 249698 9000 249934
rect 5000 249614 9000 249698
rect 5000 249378 5122 249614
rect 5358 249378 5442 249614
rect 5678 249378 5762 249614
rect 5998 249378 6082 249614
rect 6318 249378 6402 249614
rect 6638 249378 6722 249614
rect 6958 249378 7042 249614
rect 7278 249378 7362 249614
rect 7598 249378 7682 249614
rect 7918 249378 8002 249614
rect 8238 249378 8322 249614
rect 8558 249378 8642 249614
rect 8878 249378 9000 249614
rect 5000 249294 9000 249378
rect 5000 249058 5122 249294
rect 5358 249058 5442 249294
rect 5678 249058 5762 249294
rect 5998 249058 6082 249294
rect 6318 249058 6402 249294
rect 6638 249058 6722 249294
rect 6958 249058 7042 249294
rect 7278 249058 7362 249294
rect 7598 249058 7682 249294
rect 7918 249058 8002 249294
rect 8238 249058 8322 249294
rect 8558 249058 8642 249294
rect 8878 249058 9000 249294
rect 5000 248974 9000 249058
rect 5000 248738 5122 248974
rect 5358 248738 5442 248974
rect 5678 248738 5762 248974
rect 5998 248738 6082 248974
rect 6318 248738 6402 248974
rect 6638 248738 6722 248974
rect 6958 248738 7042 248974
rect 7278 248738 7362 248974
rect 7598 248738 7682 248974
rect 7918 248738 8002 248974
rect 8238 248738 8322 248974
rect 8558 248738 8642 248974
rect 8878 248738 9000 248974
rect 5000 248654 9000 248738
rect 5000 248418 5122 248654
rect 5358 248418 5442 248654
rect 5678 248418 5762 248654
rect 5998 248418 6082 248654
rect 6318 248418 6402 248654
rect 6638 248418 6722 248654
rect 6958 248418 7042 248654
rect 7278 248418 7362 248654
rect 7598 248418 7682 248654
rect 7918 248418 8002 248654
rect 8238 248418 8322 248654
rect 8558 248418 8642 248654
rect 8878 248418 9000 248654
rect 5000 248334 9000 248418
rect 5000 248098 5122 248334
rect 5358 248098 5442 248334
rect 5678 248098 5762 248334
rect 5998 248098 6082 248334
rect 6318 248098 6402 248334
rect 6638 248098 6722 248334
rect 6958 248098 7042 248334
rect 7278 248098 7362 248334
rect 7598 248098 7682 248334
rect 7918 248098 8002 248334
rect 8238 248098 8322 248334
rect 8558 248098 8642 248334
rect 8878 248098 9000 248334
rect 5000 248014 9000 248098
rect 5000 247778 5122 248014
rect 5358 247778 5442 248014
rect 5678 247778 5762 248014
rect 5998 247778 6082 248014
rect 6318 247778 6402 248014
rect 6638 247778 6722 248014
rect 6958 247778 7042 248014
rect 7278 247778 7362 248014
rect 7598 247778 7682 248014
rect 7918 247778 8002 248014
rect 8238 247778 8322 248014
rect 8558 247778 8642 248014
rect 8878 247778 9000 248014
rect 5000 247694 9000 247778
rect 5000 247458 5122 247694
rect 5358 247458 5442 247694
rect 5678 247458 5762 247694
rect 5998 247458 6082 247694
rect 6318 247458 6402 247694
rect 6638 247458 6722 247694
rect 6958 247458 7042 247694
rect 7278 247458 7362 247694
rect 7598 247458 7682 247694
rect 7918 247458 8002 247694
rect 8238 247458 8322 247694
rect 8558 247458 8642 247694
rect 8878 247458 9000 247694
rect 5000 247374 9000 247458
rect 5000 247138 5122 247374
rect 5358 247138 5442 247374
rect 5678 247138 5762 247374
rect 5998 247138 6082 247374
rect 6318 247138 6402 247374
rect 6638 247138 6722 247374
rect 6958 247138 7042 247374
rect 7278 247138 7362 247374
rect 7598 247138 7682 247374
rect 7918 247138 8002 247374
rect 8238 247138 8322 247374
rect 8558 247138 8642 247374
rect 8878 247138 9000 247374
rect 5000 247054 9000 247138
rect 5000 246818 5122 247054
rect 5358 246818 5442 247054
rect 5678 246818 5762 247054
rect 5998 246818 6082 247054
rect 6318 246818 6402 247054
rect 6638 246818 6722 247054
rect 6958 246818 7042 247054
rect 7278 246818 7362 247054
rect 7598 246818 7682 247054
rect 7918 246818 8002 247054
rect 8238 246818 8322 247054
rect 8558 246818 8642 247054
rect 8878 246818 9000 247054
rect 5000 246734 9000 246818
rect 5000 246498 5122 246734
rect 5358 246498 5442 246734
rect 5678 246498 5762 246734
rect 5998 246498 6082 246734
rect 6318 246498 6402 246734
rect 6638 246498 6722 246734
rect 6958 246498 7042 246734
rect 7278 246498 7362 246734
rect 7598 246498 7682 246734
rect 7918 246498 8002 246734
rect 8238 246498 8322 246734
rect 8558 246498 8642 246734
rect 8878 246498 9000 246734
rect 5000 240118 9000 246498
rect 228740 250254 232740 250376
rect 228740 250018 228862 250254
rect 229098 250018 229182 250254
rect 229418 250018 229502 250254
rect 229738 250018 229822 250254
rect 230058 250018 230142 250254
rect 230378 250018 230462 250254
rect 230698 250018 230782 250254
rect 231018 250018 231102 250254
rect 231338 250018 231422 250254
rect 231658 250018 231742 250254
rect 231978 250018 232062 250254
rect 232298 250018 232382 250254
rect 232618 250018 232740 250254
rect 228740 249934 232740 250018
rect 228740 249698 228862 249934
rect 229098 249698 229182 249934
rect 229418 249698 229502 249934
rect 229738 249698 229822 249934
rect 230058 249698 230142 249934
rect 230378 249698 230462 249934
rect 230698 249698 230782 249934
rect 231018 249698 231102 249934
rect 231338 249698 231422 249934
rect 231658 249698 231742 249934
rect 231978 249698 232062 249934
rect 232298 249698 232382 249934
rect 232618 249698 232740 249934
rect 228740 249614 232740 249698
rect 228740 249378 228862 249614
rect 229098 249378 229182 249614
rect 229418 249378 229502 249614
rect 229738 249378 229822 249614
rect 230058 249378 230142 249614
rect 230378 249378 230462 249614
rect 230698 249378 230782 249614
rect 231018 249378 231102 249614
rect 231338 249378 231422 249614
rect 231658 249378 231742 249614
rect 231978 249378 232062 249614
rect 232298 249378 232382 249614
rect 232618 249378 232740 249614
rect 228740 249294 232740 249378
rect 228740 249058 228862 249294
rect 229098 249058 229182 249294
rect 229418 249058 229502 249294
rect 229738 249058 229822 249294
rect 230058 249058 230142 249294
rect 230378 249058 230462 249294
rect 230698 249058 230782 249294
rect 231018 249058 231102 249294
rect 231338 249058 231422 249294
rect 231658 249058 231742 249294
rect 231978 249058 232062 249294
rect 232298 249058 232382 249294
rect 232618 249058 232740 249294
rect 228740 248974 232740 249058
rect 228740 248738 228862 248974
rect 229098 248738 229182 248974
rect 229418 248738 229502 248974
rect 229738 248738 229822 248974
rect 230058 248738 230142 248974
rect 230378 248738 230462 248974
rect 230698 248738 230782 248974
rect 231018 248738 231102 248974
rect 231338 248738 231422 248974
rect 231658 248738 231742 248974
rect 231978 248738 232062 248974
rect 232298 248738 232382 248974
rect 232618 248738 232740 248974
rect 228740 248654 232740 248738
rect 228740 248418 228862 248654
rect 229098 248418 229182 248654
rect 229418 248418 229502 248654
rect 229738 248418 229822 248654
rect 230058 248418 230142 248654
rect 230378 248418 230462 248654
rect 230698 248418 230782 248654
rect 231018 248418 231102 248654
rect 231338 248418 231422 248654
rect 231658 248418 231742 248654
rect 231978 248418 232062 248654
rect 232298 248418 232382 248654
rect 232618 248418 232740 248654
rect 228740 248334 232740 248418
rect 228740 248098 228862 248334
rect 229098 248098 229182 248334
rect 229418 248098 229502 248334
rect 229738 248098 229822 248334
rect 230058 248098 230142 248334
rect 230378 248098 230462 248334
rect 230698 248098 230782 248334
rect 231018 248098 231102 248334
rect 231338 248098 231422 248334
rect 231658 248098 231742 248334
rect 231978 248098 232062 248334
rect 232298 248098 232382 248334
rect 232618 248098 232740 248334
rect 228740 248014 232740 248098
rect 228740 247778 228862 248014
rect 229098 247778 229182 248014
rect 229418 247778 229502 248014
rect 229738 247778 229822 248014
rect 230058 247778 230142 248014
rect 230378 247778 230462 248014
rect 230698 247778 230782 248014
rect 231018 247778 231102 248014
rect 231338 247778 231422 248014
rect 231658 247778 231742 248014
rect 231978 247778 232062 248014
rect 232298 247778 232382 248014
rect 232618 247778 232740 248014
rect 228740 247694 232740 247778
rect 228740 247458 228862 247694
rect 229098 247458 229182 247694
rect 229418 247458 229502 247694
rect 229738 247458 229822 247694
rect 230058 247458 230142 247694
rect 230378 247458 230462 247694
rect 230698 247458 230782 247694
rect 231018 247458 231102 247694
rect 231338 247458 231422 247694
rect 231658 247458 231742 247694
rect 231978 247458 232062 247694
rect 232298 247458 232382 247694
rect 232618 247458 232740 247694
rect 228740 247374 232740 247458
rect 228740 247138 228862 247374
rect 229098 247138 229182 247374
rect 229418 247138 229502 247374
rect 229738 247138 229822 247374
rect 230058 247138 230142 247374
rect 230378 247138 230462 247374
rect 230698 247138 230782 247374
rect 231018 247138 231102 247374
rect 231338 247138 231422 247374
rect 231658 247138 231742 247374
rect 231978 247138 232062 247374
rect 232298 247138 232382 247374
rect 232618 247138 232740 247374
rect 228740 247054 232740 247138
rect 228740 246818 228862 247054
rect 229098 246818 229182 247054
rect 229418 246818 229502 247054
rect 229738 246818 229822 247054
rect 230058 246818 230142 247054
rect 230378 246818 230462 247054
rect 230698 246818 230782 247054
rect 231018 246818 231102 247054
rect 231338 246818 231422 247054
rect 231658 246818 231742 247054
rect 231978 246818 232062 247054
rect 232298 246818 232382 247054
rect 232618 246818 232740 247054
rect 228740 246734 232740 246818
rect 228740 246498 228862 246734
rect 229098 246498 229182 246734
rect 229418 246498 229502 246734
rect 229738 246498 229822 246734
rect 230058 246498 230142 246734
rect 230378 246498 230462 246734
rect 230698 246498 230782 246734
rect 231018 246498 231102 246734
rect 231338 246498 231422 246734
rect 231658 246498 231742 246734
rect 231978 246498 232062 246734
rect 232298 246498 232382 246734
rect 232618 246498 232740 246734
rect 5000 239882 5122 240118
rect 5358 239882 5442 240118
rect 5678 239882 5762 240118
rect 5998 239882 6082 240118
rect 6318 239882 6402 240118
rect 6638 239882 6722 240118
rect 6958 239882 7042 240118
rect 7278 239882 7362 240118
rect 7598 239882 7682 240118
rect 7918 239882 8002 240118
rect 8238 239882 8322 240118
rect 8558 239882 8642 240118
rect 8878 239882 9000 240118
rect 5000 217718 9000 239882
rect 72774 240118 73094 240160
rect 72774 239882 72816 240118
rect 73052 239882 73094 240118
rect 72774 239840 73094 239882
rect 144774 240118 145094 240160
rect 144774 239882 144816 240118
rect 145052 239882 145094 240118
rect 144774 239840 145094 239882
rect 228740 240118 232740 246498
rect 228740 239882 228862 240118
rect 229098 239882 229182 240118
rect 229418 239882 229502 240118
rect 229738 239882 229822 240118
rect 230058 239882 230142 240118
rect 230378 239882 230462 240118
rect 230698 239882 230782 240118
rect 231018 239882 231102 240118
rect 231338 239882 231422 240118
rect 231658 239882 231742 240118
rect 231978 239882 232062 240118
rect 232298 239882 232382 240118
rect 232618 239882 232740 240118
rect 77774 228918 78094 228960
rect 77774 228682 77816 228918
rect 78052 228682 78094 228918
rect 77774 228640 78094 228682
rect 149774 228918 150094 228960
rect 149774 228682 149816 228918
rect 150052 228682 150094 228918
rect 149774 228640 150094 228682
rect 5000 217482 5122 217718
rect 5358 217482 5442 217718
rect 5678 217482 5762 217718
rect 5998 217482 6082 217718
rect 6318 217482 6402 217718
rect 6638 217482 6722 217718
rect 6958 217482 7042 217718
rect 7278 217482 7362 217718
rect 7598 217482 7682 217718
rect 7918 217482 8002 217718
rect 8238 217482 8322 217718
rect 8558 217482 8642 217718
rect 8878 217482 9000 217718
rect 5000 195318 9000 217482
rect 228740 217718 232740 239882
rect 228740 217482 228862 217718
rect 229098 217482 229182 217718
rect 229418 217482 229502 217718
rect 229738 217482 229822 217718
rect 230058 217482 230142 217718
rect 230378 217482 230462 217718
rect 230698 217482 230782 217718
rect 231018 217482 231102 217718
rect 231338 217482 231422 217718
rect 231658 217482 231742 217718
rect 231978 217482 232062 217718
rect 232298 217482 232382 217718
rect 232618 217482 232740 217718
rect 37923 217276 37989 217277
rect 37923 217212 37924 217276
rect 37988 217212 37989 217276
rect 37923 217211 37989 217212
rect 5000 195082 5122 195318
rect 5358 195082 5442 195318
rect 5678 195082 5762 195318
rect 5998 195082 6082 195318
rect 6318 195082 6402 195318
rect 6638 195082 6722 195318
rect 6958 195082 7042 195318
rect 7278 195082 7362 195318
rect 7598 195082 7682 195318
rect 7918 195082 8002 195318
rect 8238 195082 8322 195318
rect 8558 195082 8642 195318
rect 8878 195082 9000 195318
rect 5000 172918 9000 195082
rect 5000 172682 5122 172918
rect 5358 172682 5442 172918
rect 5678 172682 5762 172918
rect 5998 172682 6082 172918
rect 6318 172682 6402 172918
rect 6638 172682 6722 172918
rect 6958 172682 7042 172918
rect 7278 172682 7362 172918
rect 7598 172682 7682 172918
rect 7918 172682 8002 172918
rect 8238 172682 8322 172918
rect 8558 172682 8642 172918
rect 8878 172682 9000 172918
rect 5000 150518 9000 172682
rect 17507 172918 17827 172960
rect 17507 172682 17549 172918
rect 17785 172682 17827 172918
rect 17507 172640 17827 172682
rect 20173 161718 20493 161760
rect 20173 161482 20215 161718
rect 20451 161482 20493 161718
rect 20173 161440 20493 161482
rect 37926 151589 37986 217211
rect 204259 215916 204325 215917
rect 204259 215852 204260 215916
rect 204324 215852 204325 215916
rect 204259 215851 204325 215852
rect 204262 211834 204322 215851
rect 204262 211774 204874 211834
rect 204814 211701 204874 211774
rect 204811 211700 204877 211701
rect 204811 211636 204812 211700
rect 204876 211636 204877 211700
rect 204811 211635 204877 211636
rect 42885 206518 43205 206560
rect 42885 206282 42927 206518
rect 43163 206282 43205 206518
rect 42885 206240 43205 206282
rect 78840 206518 79160 206560
rect 78840 206282 78882 206518
rect 79118 206282 79160 206518
rect 78840 206240 79160 206282
rect 115173 206518 115493 206560
rect 115173 206282 115215 206518
rect 115451 206282 115493 206518
rect 115173 206240 115493 206282
rect 150840 206518 151160 206560
rect 150840 206282 150882 206518
rect 151118 206282 151160 206518
rect 150840 206240 151160 206282
rect 187173 206518 187493 206560
rect 187173 206282 187215 206518
rect 187451 206282 187493 206518
rect 187173 206240 187493 206282
rect 38219 195318 38539 195360
rect 38219 195082 38261 195318
rect 38497 195082 38539 195318
rect 38219 195040 38539 195082
rect 73840 195318 74160 195360
rect 73840 195082 73882 195318
rect 74118 195082 74160 195318
rect 73840 195040 74160 195082
rect 110507 195318 110827 195360
rect 110507 195082 110549 195318
rect 110785 195082 110827 195318
rect 110507 195040 110827 195082
rect 145840 195318 146160 195360
rect 145840 195082 145882 195318
rect 146118 195082 146160 195318
rect 145840 195040 146160 195082
rect 182507 195318 182827 195360
rect 182507 195082 182549 195318
rect 182785 195082 182827 195318
rect 182507 195040 182827 195082
rect 228740 195318 232740 217482
rect 228740 195082 228862 195318
rect 229098 195082 229182 195318
rect 229418 195082 229502 195318
rect 229738 195082 229822 195318
rect 230058 195082 230142 195318
rect 230378 195082 230462 195318
rect 230698 195082 230782 195318
rect 231018 195082 231102 195318
rect 231338 195082 231422 195318
rect 231658 195082 231742 195318
rect 231978 195082 232062 195318
rect 232298 195082 232382 195318
rect 232618 195082 232740 195318
rect 207571 192524 207637 192525
rect 207571 192460 207572 192524
rect 207636 192460 207637 192524
rect 207571 192459 207637 192460
rect 207574 192389 207634 192459
rect 207571 192388 207637 192389
rect 207571 192324 207572 192388
rect 207636 192324 207637 192388
rect 207571 192323 207637 192324
rect 207203 182868 207269 182869
rect 207203 182804 207204 182868
rect 207268 182804 207269 182868
rect 207203 182803 207269 182804
rect 207206 175794 207266 182803
rect 207206 175734 207450 175794
rect 42507 172918 42827 172960
rect 42507 172682 42549 172918
rect 42785 172682 42827 172918
rect 42507 172640 42827 172682
rect 67104 172918 67424 172960
rect 67104 172682 67146 172918
rect 67382 172682 67424 172918
rect 67104 172640 67424 172682
rect 114507 172918 114827 172960
rect 114507 172682 114549 172918
rect 114785 172682 114827 172918
rect 114507 172640 114827 172682
rect 139104 172918 139424 172960
rect 139104 172682 139146 172918
rect 139382 172682 139424 172918
rect 139104 172640 139424 172682
rect 186507 172918 186827 172960
rect 207390 172941 207450 175734
rect 186507 172682 186549 172918
rect 186785 172682 186827 172918
rect 207387 172940 207453 172941
rect 207387 172876 207388 172940
rect 207452 172876 207453 172940
rect 207387 172875 207453 172876
rect 207571 172940 207637 172941
rect 207571 172876 207572 172940
rect 207636 172876 207637 172940
rect 207571 172875 207637 172876
rect 211507 172918 211827 172960
rect 186507 172640 186827 172682
rect 207574 163285 207634 172875
rect 211507 172682 211549 172918
rect 211785 172682 211827 172918
rect 211507 172640 211827 172682
rect 228740 172918 232740 195082
rect 228740 172682 228862 172918
rect 229098 172682 229182 172918
rect 229418 172682 229502 172918
rect 229738 172682 229822 172918
rect 230058 172682 230142 172918
rect 230378 172682 230462 172918
rect 230698 172682 230782 172918
rect 231018 172682 231102 172918
rect 231338 172682 231422 172918
rect 231658 172682 231742 172918
rect 231978 172682 232062 172918
rect 232298 172682 232382 172918
rect 232618 172682 232740 172918
rect 207571 163284 207637 163285
rect 207571 163220 207572 163284
rect 207636 163220 207637 163284
rect 207571 163219 207637 163220
rect 45173 161718 45493 161760
rect 45173 161482 45215 161718
rect 45451 161482 45493 161718
rect 45173 161440 45493 161482
rect 82464 161718 82784 161760
rect 82464 161482 82506 161718
rect 82742 161482 82784 161718
rect 82464 161440 82784 161482
rect 117173 161718 117493 161760
rect 117173 161482 117215 161718
rect 117451 161482 117493 161718
rect 117173 161440 117493 161482
rect 154464 161718 154784 161760
rect 154464 161482 154506 161718
rect 154742 161482 154784 161718
rect 154464 161440 154784 161482
rect 189173 161718 189493 161760
rect 189173 161482 189215 161718
rect 189451 161482 189493 161718
rect 189173 161440 189493 161482
rect 214173 161718 214493 161760
rect 214173 161482 214215 161718
rect 214451 161482 214493 161718
rect 214173 161440 214493 161482
rect 207387 153764 207453 153765
rect 207387 153700 207388 153764
rect 207452 153700 207453 153764
rect 207387 153699 207453 153700
rect 207390 152269 207450 153699
rect 207387 152268 207453 152269
rect 207387 152204 207388 152268
rect 207452 152204 207453 152268
rect 207387 152203 207453 152204
rect 37923 151588 37989 151589
rect 37923 151524 37924 151588
rect 37988 151524 37989 151588
rect 37923 151523 37989 151524
rect 5000 150282 5122 150518
rect 5358 150282 5442 150518
rect 5678 150282 5762 150518
rect 5998 150282 6082 150518
rect 6318 150282 6402 150518
rect 6638 150282 6722 150518
rect 6958 150282 7042 150518
rect 7278 150282 7362 150518
rect 7598 150282 7682 150518
rect 7918 150282 8002 150518
rect 8238 150282 8322 150518
rect 8558 150282 8642 150518
rect 8878 150282 9000 150518
rect 5000 128118 9000 150282
rect 17507 150518 17827 150560
rect 17507 150282 17549 150518
rect 17785 150282 17827 150518
rect 17507 150240 17827 150282
rect 42507 150518 42827 150560
rect 42507 150282 42549 150518
rect 42785 150282 42827 150518
rect 42507 150240 42827 150282
rect 67104 150518 67424 150560
rect 67104 150282 67146 150518
rect 67382 150282 67424 150518
rect 67104 150240 67424 150282
rect 114507 150518 114827 150560
rect 114507 150282 114549 150518
rect 114785 150282 114827 150518
rect 114507 150240 114827 150282
rect 139104 150518 139424 150560
rect 139104 150282 139146 150518
rect 139382 150282 139424 150518
rect 139104 150240 139424 150282
rect 186507 150518 186827 150560
rect 186507 150282 186549 150518
rect 186785 150282 186827 150518
rect 186507 150240 186827 150282
rect 211507 150518 211827 150560
rect 211507 150282 211549 150518
rect 211785 150282 211827 150518
rect 211507 150240 211827 150282
rect 228740 150518 232740 172682
rect 228740 150282 228862 150518
rect 229098 150282 229182 150518
rect 229418 150282 229502 150518
rect 229738 150282 229822 150518
rect 230058 150282 230142 150518
rect 230378 150282 230462 150518
rect 230698 150282 230782 150518
rect 231018 150282 231102 150518
rect 231338 150282 231422 150518
rect 231658 150282 231742 150518
rect 231978 150282 232062 150518
rect 232298 150282 232382 150518
rect 232618 150282 232740 150518
rect 207755 142748 207821 142749
rect 207755 142684 207756 142748
rect 207820 142684 207821 142748
rect 207755 142683 207821 142684
rect 207758 142613 207818 142683
rect 101035 142612 101101 142613
rect 101035 142548 101036 142612
rect 101100 142548 101101 142612
rect 101035 142547 101101 142548
rect 167275 142612 167341 142613
rect 167275 142548 167276 142612
rect 167340 142548 167341 142612
rect 167275 142547 167341 142548
rect 207755 142612 207821 142613
rect 207755 142548 207756 142612
rect 207820 142548 207821 142612
rect 207755 142547 207821 142548
rect 71043 141932 71109 141933
rect 71043 141868 71044 141932
rect 71108 141868 71109 141932
rect 71043 141867 71109 141868
rect 31851 141388 31917 141389
rect 31851 141324 31852 141388
rect 31916 141324 31917 141388
rect 31851 141323 31917 141324
rect 5000 127882 5122 128118
rect 5358 127882 5442 128118
rect 5678 127882 5762 128118
rect 5998 127882 6082 128118
rect 6318 127882 6402 128118
rect 6638 127882 6722 128118
rect 6958 127882 7042 128118
rect 7278 127882 7362 128118
rect 7598 127882 7682 128118
rect 7918 127882 8002 128118
rect 8238 127882 8322 128118
rect 8558 127882 8642 128118
rect 8878 127882 9000 128118
rect 5000 105718 9000 127882
rect 21550 127653 21610 128726
rect 21547 127652 21613 127653
rect 21547 127588 21548 127652
rect 21612 127588 21613 127652
rect 21547 127587 21613 127588
rect 31854 118541 31914 141323
rect 43173 139318 43493 139360
rect 43173 139082 43215 139318
rect 43451 139082 43493 139318
rect 43173 139040 43493 139082
rect 71046 137034 71106 141867
rect 94227 141388 94293 141389
rect 94227 141324 94228 141388
rect 94292 141324 94293 141388
rect 94227 141323 94293 141324
rect 70862 136974 71106 137034
rect 70862 134994 70922 136974
rect 70862 134934 71106 134994
rect 67734 128962 67794 131446
rect 71046 129554 71106 134934
rect 70678 129494 71106 129554
rect 38507 128118 38827 128160
rect 38507 127882 38549 128118
rect 38785 127882 38827 128118
rect 38507 127840 38827 127882
rect 31851 118540 31917 118541
rect 31851 118476 31852 118540
rect 31916 118476 31917 118540
rect 31851 118475 31917 118476
rect 31854 114002 31914 118475
rect 70678 117994 70738 129494
rect 73840 128118 74160 128160
rect 73840 127882 73882 128118
rect 74118 127882 74160 128118
rect 73840 127840 74160 127882
rect 70678 117934 71106 117994
rect 43173 116918 43493 116960
rect 43173 116682 43215 116918
rect 43451 116682 43493 116918
rect 43173 116640 43493 116682
rect 56878 113237 56938 113766
rect 71046 113645 71106 117934
rect 71043 113644 71109 113645
rect 71043 113580 71044 113644
rect 71108 113580 71109 113644
rect 71043 113579 71109 113580
rect 56875 113236 56941 113237
rect 56875 113172 56876 113236
rect 56940 113172 56941 113236
rect 56875 113171 56941 113172
rect 94230 112693 94290 141323
rect 94227 112692 94293 112693
rect 94227 112628 94228 112692
rect 94292 112628 94293 112692
rect 94227 112627 94293 112628
rect 5000 105482 5122 105718
rect 5358 105482 5442 105718
rect 5678 105482 5762 105718
rect 5998 105482 6082 105718
rect 6318 105482 6402 105718
rect 6638 105482 6722 105718
rect 6958 105482 7042 105718
rect 7278 105482 7362 105718
rect 7598 105482 7682 105718
rect 7918 105482 8002 105718
rect 8238 105482 8322 105718
rect 8558 105482 8642 105718
rect 8878 105482 9000 105718
rect 5000 83318 9000 105482
rect 17507 105718 17827 105760
rect 17507 105482 17549 105718
rect 17785 105482 17827 105718
rect 17507 105440 17827 105482
rect 42507 105718 42827 105760
rect 42507 105482 42549 105718
rect 42785 105482 42827 105718
rect 42507 105440 42827 105482
rect 67104 105718 67424 105760
rect 67104 105482 67146 105718
rect 67382 105482 67424 105718
rect 67104 105440 67424 105482
rect 20173 94518 20493 94560
rect 20173 94282 20215 94518
rect 20451 94282 20493 94518
rect 20173 94240 20493 94282
rect 45173 94518 45493 94560
rect 45173 94282 45215 94518
rect 45451 94282 45493 94518
rect 45173 94240 45493 94282
rect 82464 94518 82784 94560
rect 82464 94282 82506 94518
rect 82742 94282 82784 94518
rect 82464 94240 82784 94282
rect 5000 83082 5122 83318
rect 5358 83082 5442 83318
rect 5678 83082 5762 83318
rect 5998 83082 6082 83318
rect 6318 83082 6402 83318
rect 6638 83082 6722 83318
rect 6958 83082 7042 83318
rect 7278 83082 7362 83318
rect 7598 83082 7682 83318
rect 7918 83082 8002 83318
rect 8238 83082 8322 83318
rect 8558 83082 8642 83318
rect 8878 83082 9000 83318
rect 5000 60918 9000 83082
rect 17507 83318 17827 83360
rect 17507 83082 17549 83318
rect 17785 83082 17827 83318
rect 17507 83040 17827 83082
rect 42507 83318 42827 83360
rect 42507 83082 42549 83318
rect 42785 83082 42827 83318
rect 42507 83040 42827 83082
rect 67104 83318 67424 83360
rect 67104 83082 67146 83318
rect 67382 83082 67424 83318
rect 67104 83040 67424 83082
rect 101038 71077 101098 142547
rect 146299 141932 146365 141933
rect 146299 141868 146300 141932
rect 146364 141868 146365 141932
rect 146299 141867 146365 141868
rect 115173 139318 115493 139360
rect 115173 139082 115215 139318
rect 115451 139082 115493 139318
rect 115173 139040 115493 139082
rect 146302 138482 146362 141867
rect 101403 131396 101404 131446
rect 101468 131396 101469 131446
rect 101403 131395 101469 131396
rect 101406 71213 101466 131395
rect 110507 128118 110827 128160
rect 110507 127882 110549 128118
rect 110785 127882 110827 128118
rect 110507 127840 110827 127882
rect 142622 117994 142682 136886
rect 145840 128118 146160 128160
rect 145840 127882 145882 128118
rect 146118 127882 146160 128118
rect 145840 127840 146160 127882
rect 142622 117934 143050 117994
rect 115173 116918 115493 116960
rect 115173 116682 115215 116918
rect 115451 116682 115493 116918
rect 115173 116640 115493 116682
rect 142990 113645 143050 117934
rect 167278 113645 167338 142547
rect 187173 139318 187493 139360
rect 187173 139082 187215 139318
rect 187451 139082 187493 139318
rect 187173 139040 187493 139082
rect 182507 128118 182827 128160
rect 182507 127882 182549 128118
rect 182785 127882 182827 128118
rect 182507 127840 182827 127882
rect 228740 128118 232740 150282
rect 228740 127882 228862 128118
rect 229098 127882 229182 128118
rect 229418 127882 229502 128118
rect 229738 127882 229822 128118
rect 230058 127882 230142 128118
rect 230378 127882 230462 128118
rect 230698 127882 230782 128118
rect 231018 127882 231102 128118
rect 231338 127882 231422 128118
rect 231658 127882 231742 128118
rect 231978 127882 232062 128118
rect 232298 127882 232382 128118
rect 232618 127882 232740 128118
rect 187173 116918 187493 116960
rect 187173 116682 187215 116918
rect 187451 116682 187493 116918
rect 187173 116640 187493 116682
rect 142987 113644 143053 113645
rect 142987 113580 142988 113644
rect 143052 113580 143053 113644
rect 142987 113579 143053 113580
rect 167275 113644 167341 113645
rect 167275 113580 167276 113644
rect 167340 113580 167341 113644
rect 167275 113579 167341 113580
rect 114507 105718 114827 105760
rect 114507 105482 114549 105718
rect 114785 105482 114827 105718
rect 114507 105440 114827 105482
rect 139104 105718 139424 105760
rect 139104 105482 139146 105718
rect 139382 105482 139424 105718
rect 139104 105440 139424 105482
rect 186507 105718 186827 105760
rect 186507 105482 186549 105718
rect 186785 105482 186827 105718
rect 186507 105440 186827 105482
rect 211507 105718 211827 105760
rect 211507 105482 211549 105718
rect 211785 105482 211827 105718
rect 211507 105440 211827 105482
rect 228740 105718 232740 127882
rect 228740 105482 228862 105718
rect 229098 105482 229182 105718
rect 229418 105482 229502 105718
rect 229738 105482 229822 105718
rect 230058 105482 230142 105718
rect 230378 105482 230462 105718
rect 230698 105482 230782 105718
rect 231018 105482 231102 105718
rect 231338 105482 231422 105718
rect 231658 105482 231742 105718
rect 231978 105482 232062 105718
rect 232298 105482 232382 105718
rect 232618 105482 232740 105718
rect 117173 94518 117493 94560
rect 117173 94282 117215 94518
rect 117451 94282 117493 94518
rect 117173 94240 117493 94282
rect 154464 94518 154784 94560
rect 154464 94282 154506 94518
rect 154742 94282 154784 94518
rect 154464 94240 154784 94282
rect 189173 94518 189493 94560
rect 189173 94282 189215 94518
rect 189451 94282 189493 94518
rect 189173 94240 189493 94282
rect 214173 94518 214493 94560
rect 214173 94282 214215 94518
rect 214451 94282 214493 94518
rect 214173 94240 214493 94282
rect 114507 83318 114827 83360
rect 114507 83082 114549 83318
rect 114785 83082 114827 83318
rect 114507 83040 114827 83082
rect 139104 83318 139424 83360
rect 139104 83082 139146 83318
rect 139382 83082 139424 83318
rect 139104 83040 139424 83082
rect 186507 83318 186827 83360
rect 186507 83082 186549 83318
rect 186785 83082 186827 83318
rect 186507 83040 186827 83082
rect 211507 83318 211827 83360
rect 211507 83082 211549 83318
rect 211785 83082 211827 83318
rect 211507 83040 211827 83082
rect 228740 83318 232740 105482
rect 228740 83082 228862 83318
rect 229098 83082 229182 83318
rect 229418 83082 229502 83318
rect 229738 83082 229822 83318
rect 230058 83082 230142 83318
rect 230378 83082 230462 83318
rect 230698 83082 230782 83318
rect 231018 83082 231102 83318
rect 231338 83082 231422 83318
rect 231658 83082 231742 83318
rect 231978 83082 232062 83318
rect 232298 83082 232382 83318
rect 232618 83082 232740 83318
rect 129739 77604 129805 77605
rect 129739 77540 129740 77604
rect 129804 77540 129805 77604
rect 129739 77539 129805 77540
rect 101403 71212 101469 71213
rect 101403 71148 101404 71212
rect 101468 71148 101469 71212
rect 101403 71147 101469 71148
rect 101035 71076 101101 71077
rect 101035 71012 101036 71076
rect 101100 71012 101101 71076
rect 101035 71011 101101 71012
rect 31851 69444 31917 69445
rect 31851 69380 31852 69444
rect 31916 69380 31917 69444
rect 31851 69379 31917 69380
rect 5000 60682 5122 60918
rect 5358 60682 5442 60918
rect 5678 60682 5762 60918
rect 5998 60682 6082 60918
rect 6318 60682 6402 60918
rect 6638 60682 6722 60918
rect 6958 60682 7042 60918
rect 7278 60682 7362 60918
rect 7598 60682 7682 60918
rect 7918 60682 8002 60918
rect 8238 60682 8322 60918
rect 8558 60682 8642 60918
rect 8878 60682 9000 60918
rect 5000 38518 9000 60682
rect 31854 44285 31914 69379
rect 38507 60918 38827 60960
rect 38507 60682 38549 60918
rect 38785 60682 38827 60918
rect 38507 60640 38827 60682
rect 73840 60918 74160 60960
rect 73840 60682 73882 60918
rect 74118 60682 74160 60918
rect 73840 60640 74160 60682
rect 110507 60918 110827 60960
rect 110507 60682 110549 60918
rect 110785 60682 110827 60918
rect 110507 60640 110827 60682
rect 43173 49718 43493 49760
rect 43173 49482 43215 49718
rect 43451 49482 43493 49718
rect 43173 49440 43493 49482
rect 78840 49718 79160 49760
rect 78840 49482 78882 49718
rect 79118 49482 79160 49718
rect 78840 49440 79160 49482
rect 115173 49718 115493 49760
rect 115173 49482 115215 49718
rect 115451 49482 115493 49718
rect 115173 49440 115493 49482
rect 31851 44284 31917 44285
rect 31851 44220 31852 44284
rect 31916 44220 31917 44284
rect 31851 44219 31917 44220
rect 31854 41242 31914 44219
rect 66262 40477 66322 41006
rect 129742 40562 129802 77539
rect 201499 69308 201565 69309
rect 201499 69244 201500 69308
rect 201564 69244 201565 69308
rect 201499 69243 201565 69244
rect 201502 65634 201562 69243
rect 201502 65574 201746 65634
rect 145840 60918 146160 60960
rect 145840 60682 145882 60918
rect 146118 60682 146160 60918
rect 145840 60640 146160 60682
rect 182507 60918 182827 60960
rect 182507 60682 182549 60918
rect 182785 60682 182827 60918
rect 182507 60640 182827 60682
rect 150840 49718 151160 49760
rect 150840 49482 150882 49718
rect 151118 49482 151160 49718
rect 150840 49440 151160 49482
rect 187173 49718 187493 49760
rect 187173 49482 187215 49718
rect 187451 49482 187493 49718
rect 187173 49440 187493 49482
rect 201686 41834 201746 65574
rect 201502 41774 201746 41834
rect 228740 60918 232740 83082
rect 228740 60682 228862 60918
rect 229098 60682 229182 60918
rect 229418 60682 229502 60918
rect 229738 60682 229822 60918
rect 230058 60682 230142 60918
rect 230378 60682 230462 60918
rect 230698 60682 230782 60918
rect 231018 60682 231102 60918
rect 231338 60682 231422 60918
rect 231658 60682 231742 60918
rect 231978 60682 232062 60918
rect 232298 60682 232382 60918
rect 232618 60682 232740 60918
rect 66259 40476 66325 40477
rect 66259 40412 66260 40476
rect 66324 40412 66325 40476
rect 66259 40411 66325 40412
rect 108914 40414 109598 40474
rect 109686 40069 109746 40326
rect 109683 40068 109749 40069
rect 109683 40004 109684 40068
rect 109748 40004 109749 40068
rect 109683 40003 109749 40004
rect 136918 39797 136978 40326
rect 181446 40069 181506 40326
rect 181443 40068 181509 40069
rect 181443 40004 181444 40068
rect 181508 40004 181509 40068
rect 181443 40003 181509 40004
rect 136915 39796 136981 39797
rect 136915 39732 136916 39796
rect 136980 39732 136981 39796
rect 136915 39731 136981 39732
rect 201502 39202 201562 41774
rect 5000 38282 5122 38518
rect 5358 38282 5442 38518
rect 5678 38282 5762 38518
rect 5998 38282 6082 38518
rect 6318 38282 6402 38518
rect 6638 38282 6722 38518
rect 6958 38282 7042 38518
rect 7278 38282 7362 38518
rect 7598 38282 7682 38518
rect 7918 38282 8002 38518
rect 8238 38282 8322 38518
rect 8558 38282 8642 38518
rect 8878 38282 9000 38518
rect 5000 16118 9000 38282
rect 228740 38518 232740 60682
rect 228740 38282 228862 38518
rect 229098 38282 229182 38518
rect 229418 38282 229502 38518
rect 229738 38282 229822 38518
rect 230058 38282 230142 38518
rect 230378 38282 230462 38518
rect 230698 38282 230782 38518
rect 231018 38282 231102 38518
rect 231338 38282 231422 38518
rect 231658 38282 231742 38518
rect 231978 38282 232062 38518
rect 232298 38282 232382 38518
rect 232618 38282 232740 38518
rect 78840 27318 79160 27360
rect 78840 27082 78882 27318
rect 79118 27082 79160 27318
rect 78840 27040 79160 27082
rect 150840 27318 151160 27360
rect 150840 27082 150882 27318
rect 151118 27082 151160 27318
rect 150840 27040 151160 27082
rect 5000 15882 5122 16118
rect 5358 15882 5442 16118
rect 5678 15882 5762 16118
rect 5998 15882 6082 16118
rect 6318 15882 6402 16118
rect 6638 15882 6722 16118
rect 6958 15882 7042 16118
rect 7278 15882 7362 16118
rect 7598 15882 7682 16118
rect 7918 15882 8002 16118
rect 8238 15882 8322 16118
rect 8558 15882 8642 16118
rect 8878 15882 9000 16118
rect 5000 8878 9000 15882
rect 73840 16118 74160 16160
rect 73840 15882 73882 16118
rect 74118 15882 74160 16118
rect 73840 15840 74160 15882
rect 145840 16118 146160 16160
rect 145840 15882 145882 16118
rect 146118 15882 146160 16118
rect 145840 15840 146160 15882
rect 228740 16118 232740 38282
rect 228740 15882 228862 16118
rect 229098 15882 229182 16118
rect 229418 15882 229502 16118
rect 229738 15882 229822 16118
rect 230058 15882 230142 16118
rect 230378 15882 230462 16118
rect 230698 15882 230782 16118
rect 231018 15882 231102 16118
rect 231338 15882 231422 16118
rect 231658 15882 231742 16118
rect 231978 15882 232062 16118
rect 232298 15882 232382 16118
rect 232618 15882 232740 16118
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 9000 8878
rect 5000 8558 9000 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 9000 8558
rect 5000 8238 9000 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 9000 8238
rect 5000 7918 9000 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 9000 7918
rect 5000 7598 9000 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 9000 7598
rect 5000 7278 9000 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 9000 7278
rect 5000 6958 9000 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 9000 6958
rect 5000 6638 9000 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 9000 6638
rect 5000 6318 9000 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 9000 6318
rect 5000 5998 9000 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 9000 5998
rect 5000 5678 9000 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 9000 5678
rect 5000 5358 9000 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 9000 5358
rect 5000 5000 9000 5122
rect 228740 8878 232740 15882
rect 228740 8642 228862 8878
rect 229098 8642 229182 8878
rect 229418 8642 229502 8878
rect 229738 8642 229822 8878
rect 230058 8642 230142 8878
rect 230378 8642 230462 8878
rect 230698 8642 230782 8878
rect 231018 8642 231102 8878
rect 231338 8642 231422 8878
rect 231658 8642 231742 8878
rect 231978 8642 232062 8878
rect 232298 8642 232382 8878
rect 232618 8642 232740 8878
rect 228740 8558 232740 8642
rect 228740 8322 228862 8558
rect 229098 8322 229182 8558
rect 229418 8322 229502 8558
rect 229738 8322 229822 8558
rect 230058 8322 230142 8558
rect 230378 8322 230462 8558
rect 230698 8322 230782 8558
rect 231018 8322 231102 8558
rect 231338 8322 231422 8558
rect 231658 8322 231742 8558
rect 231978 8322 232062 8558
rect 232298 8322 232382 8558
rect 232618 8322 232740 8558
rect 228740 8238 232740 8322
rect 228740 8002 228862 8238
rect 229098 8002 229182 8238
rect 229418 8002 229502 8238
rect 229738 8002 229822 8238
rect 230058 8002 230142 8238
rect 230378 8002 230462 8238
rect 230698 8002 230782 8238
rect 231018 8002 231102 8238
rect 231338 8002 231422 8238
rect 231658 8002 231742 8238
rect 231978 8002 232062 8238
rect 232298 8002 232382 8238
rect 232618 8002 232740 8238
rect 228740 7918 232740 8002
rect 228740 7682 228862 7918
rect 229098 7682 229182 7918
rect 229418 7682 229502 7918
rect 229738 7682 229822 7918
rect 230058 7682 230142 7918
rect 230378 7682 230462 7918
rect 230698 7682 230782 7918
rect 231018 7682 231102 7918
rect 231338 7682 231422 7918
rect 231658 7682 231742 7918
rect 231978 7682 232062 7918
rect 232298 7682 232382 7918
rect 232618 7682 232740 7918
rect 228740 7598 232740 7682
rect 228740 7362 228862 7598
rect 229098 7362 229182 7598
rect 229418 7362 229502 7598
rect 229738 7362 229822 7598
rect 230058 7362 230142 7598
rect 230378 7362 230462 7598
rect 230698 7362 230782 7598
rect 231018 7362 231102 7598
rect 231338 7362 231422 7598
rect 231658 7362 231742 7598
rect 231978 7362 232062 7598
rect 232298 7362 232382 7598
rect 232618 7362 232740 7598
rect 228740 7278 232740 7362
rect 228740 7042 228862 7278
rect 229098 7042 229182 7278
rect 229418 7042 229502 7278
rect 229738 7042 229822 7278
rect 230058 7042 230142 7278
rect 230378 7042 230462 7278
rect 230698 7042 230782 7278
rect 231018 7042 231102 7278
rect 231338 7042 231422 7278
rect 231658 7042 231742 7278
rect 231978 7042 232062 7278
rect 232298 7042 232382 7278
rect 232618 7042 232740 7278
rect 228740 6958 232740 7042
rect 228740 6722 228862 6958
rect 229098 6722 229182 6958
rect 229418 6722 229502 6958
rect 229738 6722 229822 6958
rect 230058 6722 230142 6958
rect 230378 6722 230462 6958
rect 230698 6722 230782 6958
rect 231018 6722 231102 6958
rect 231338 6722 231422 6958
rect 231658 6722 231742 6958
rect 231978 6722 232062 6958
rect 232298 6722 232382 6958
rect 232618 6722 232740 6958
rect 228740 6638 232740 6722
rect 228740 6402 228862 6638
rect 229098 6402 229182 6638
rect 229418 6402 229502 6638
rect 229738 6402 229822 6638
rect 230058 6402 230142 6638
rect 230378 6402 230462 6638
rect 230698 6402 230782 6638
rect 231018 6402 231102 6638
rect 231338 6402 231422 6638
rect 231658 6402 231742 6638
rect 231978 6402 232062 6638
rect 232298 6402 232382 6638
rect 232618 6402 232740 6638
rect 228740 6318 232740 6402
rect 228740 6082 228862 6318
rect 229098 6082 229182 6318
rect 229418 6082 229502 6318
rect 229738 6082 229822 6318
rect 230058 6082 230142 6318
rect 230378 6082 230462 6318
rect 230698 6082 230782 6318
rect 231018 6082 231102 6318
rect 231338 6082 231422 6318
rect 231658 6082 231742 6318
rect 231978 6082 232062 6318
rect 232298 6082 232382 6318
rect 232618 6082 232740 6318
rect 228740 5998 232740 6082
rect 228740 5762 228862 5998
rect 229098 5762 229182 5998
rect 229418 5762 229502 5998
rect 229738 5762 229822 5998
rect 230058 5762 230142 5998
rect 230378 5762 230462 5998
rect 230698 5762 230782 5998
rect 231018 5762 231102 5998
rect 231338 5762 231422 5998
rect 231658 5762 231742 5998
rect 231978 5762 232062 5998
rect 232298 5762 232382 5998
rect 232618 5762 232740 5998
rect 228740 5678 232740 5762
rect 228740 5442 228862 5678
rect 229098 5442 229182 5678
rect 229418 5442 229502 5678
rect 229738 5442 229822 5678
rect 230058 5442 230142 5678
rect 230378 5442 230462 5678
rect 230698 5442 230782 5678
rect 231018 5442 231102 5678
rect 231338 5442 231422 5678
rect 231658 5442 231742 5678
rect 231978 5442 232062 5678
rect 232298 5442 232382 5678
rect 232618 5442 232740 5678
rect 228740 5358 232740 5442
rect 228740 5122 228862 5358
rect 229098 5122 229182 5358
rect 229418 5122 229502 5358
rect 229738 5122 229822 5358
rect 230058 5122 230142 5358
rect 230378 5122 230462 5358
rect 230698 5122 230782 5358
rect 231018 5122 231102 5358
rect 231338 5122 231422 5358
rect 231658 5122 231742 5358
rect 231978 5122 232062 5358
rect 232298 5122 232382 5358
rect 232618 5122 232740 5358
rect 228740 5000 232740 5122
rect 233740 228918 237740 251498
rect 233740 228682 233862 228918
rect 234098 228682 234182 228918
rect 234418 228682 234502 228918
rect 234738 228682 234822 228918
rect 235058 228682 235142 228918
rect 235378 228682 235462 228918
rect 235698 228682 235782 228918
rect 236018 228682 236102 228918
rect 236338 228682 236422 228918
rect 236658 228682 236742 228918
rect 236978 228682 237062 228918
rect 237298 228682 237382 228918
rect 237618 228682 237740 228918
rect 233740 206518 237740 228682
rect 233740 206282 233862 206518
rect 234098 206282 234182 206518
rect 234418 206282 234502 206518
rect 234738 206282 234822 206518
rect 235058 206282 235142 206518
rect 235378 206282 235462 206518
rect 235698 206282 235782 206518
rect 236018 206282 236102 206518
rect 236338 206282 236422 206518
rect 236658 206282 236742 206518
rect 236978 206282 237062 206518
rect 237298 206282 237382 206518
rect 237618 206282 237740 206518
rect 233740 184118 237740 206282
rect 233740 183882 233862 184118
rect 234098 183882 234182 184118
rect 234418 183882 234502 184118
rect 234738 183882 234822 184118
rect 235058 183882 235142 184118
rect 235378 183882 235462 184118
rect 235698 183882 235782 184118
rect 236018 183882 236102 184118
rect 236338 183882 236422 184118
rect 236658 183882 236742 184118
rect 236978 183882 237062 184118
rect 237298 183882 237382 184118
rect 237618 183882 237740 184118
rect 233740 161718 237740 183882
rect 233740 161482 233862 161718
rect 234098 161482 234182 161718
rect 234418 161482 234502 161718
rect 234738 161482 234822 161718
rect 235058 161482 235142 161718
rect 235378 161482 235462 161718
rect 235698 161482 235782 161718
rect 236018 161482 236102 161718
rect 236338 161482 236422 161718
rect 236658 161482 236742 161718
rect 236978 161482 237062 161718
rect 237298 161482 237382 161718
rect 237618 161482 237740 161718
rect 233740 139318 237740 161482
rect 233740 139082 233862 139318
rect 234098 139082 234182 139318
rect 234418 139082 234502 139318
rect 234738 139082 234822 139318
rect 235058 139082 235142 139318
rect 235378 139082 235462 139318
rect 235698 139082 235782 139318
rect 236018 139082 236102 139318
rect 236338 139082 236422 139318
rect 236658 139082 236742 139318
rect 236978 139082 237062 139318
rect 237298 139082 237382 139318
rect 237618 139082 237740 139318
rect 233740 116918 237740 139082
rect 233740 116682 233862 116918
rect 234098 116682 234182 116918
rect 234418 116682 234502 116918
rect 234738 116682 234822 116918
rect 235058 116682 235142 116918
rect 235378 116682 235462 116918
rect 235698 116682 235782 116918
rect 236018 116682 236102 116918
rect 236338 116682 236422 116918
rect 236658 116682 236742 116918
rect 236978 116682 237062 116918
rect 237298 116682 237382 116918
rect 237618 116682 237740 116918
rect 233740 94518 237740 116682
rect 233740 94282 233862 94518
rect 234098 94282 234182 94518
rect 234418 94282 234502 94518
rect 234738 94282 234822 94518
rect 235058 94282 235142 94518
rect 235378 94282 235462 94518
rect 235698 94282 235782 94518
rect 236018 94282 236102 94518
rect 236338 94282 236422 94518
rect 236658 94282 236742 94518
rect 236978 94282 237062 94518
rect 237298 94282 237382 94518
rect 237618 94282 237740 94518
rect 233740 72118 237740 94282
rect 233740 71882 233862 72118
rect 234098 71882 234182 72118
rect 234418 71882 234502 72118
rect 234738 71882 234822 72118
rect 235058 71882 235142 72118
rect 235378 71882 235462 72118
rect 235698 71882 235782 72118
rect 236018 71882 236102 72118
rect 236338 71882 236422 72118
rect 236658 71882 236742 72118
rect 236978 71882 237062 72118
rect 237298 71882 237382 72118
rect 237618 71882 237740 72118
rect 233740 49718 237740 71882
rect 233740 49482 233862 49718
rect 234098 49482 234182 49718
rect 234418 49482 234502 49718
rect 234738 49482 234822 49718
rect 235058 49482 235142 49718
rect 235378 49482 235462 49718
rect 235698 49482 235782 49718
rect 236018 49482 236102 49718
rect 236338 49482 236422 49718
rect 236658 49482 236742 49718
rect 236978 49482 237062 49718
rect 237298 49482 237382 49718
rect 237618 49482 237740 49718
rect 233740 27318 237740 49482
rect 233740 27082 233862 27318
rect 234098 27082 234182 27318
rect 234418 27082 234502 27318
rect 234738 27082 234822 27318
rect 235058 27082 235142 27318
rect 235378 27082 235462 27318
rect 235698 27082 235782 27318
rect 236018 27082 236102 27318
rect 236338 27082 236422 27318
rect 236658 27082 236742 27318
rect 236978 27082 237062 27318
rect 237298 27082 237382 27318
rect 237618 27082 237740 27318
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 4000 3878
rect 0 3558 4000 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 4000 3558
rect 0 3238 4000 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 4000 3238
rect 0 2918 4000 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 4000 2918
rect 0 2598 4000 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 4000 2598
rect 0 2278 4000 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 4000 2278
rect 0 1958 4000 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 4000 1958
rect 0 1638 4000 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 4000 1638
rect 0 1318 4000 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 4000 1318
rect 0 998 4000 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 4000 998
rect 0 678 4000 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 4000 678
rect 0 358 4000 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 4000 358
rect 0 0 4000 122
rect 233740 3878 237740 27082
rect 233740 3642 233862 3878
rect 234098 3642 234182 3878
rect 234418 3642 234502 3878
rect 234738 3642 234822 3878
rect 235058 3642 235142 3878
rect 235378 3642 235462 3878
rect 235698 3642 235782 3878
rect 236018 3642 236102 3878
rect 236338 3642 236422 3878
rect 236658 3642 236742 3878
rect 236978 3642 237062 3878
rect 237298 3642 237382 3878
rect 237618 3642 237740 3878
rect 233740 3558 237740 3642
rect 233740 3322 233862 3558
rect 234098 3322 234182 3558
rect 234418 3322 234502 3558
rect 234738 3322 234822 3558
rect 235058 3322 235142 3558
rect 235378 3322 235462 3558
rect 235698 3322 235782 3558
rect 236018 3322 236102 3558
rect 236338 3322 236422 3558
rect 236658 3322 236742 3558
rect 236978 3322 237062 3558
rect 237298 3322 237382 3558
rect 237618 3322 237740 3558
rect 233740 3238 237740 3322
rect 233740 3002 233862 3238
rect 234098 3002 234182 3238
rect 234418 3002 234502 3238
rect 234738 3002 234822 3238
rect 235058 3002 235142 3238
rect 235378 3002 235462 3238
rect 235698 3002 235782 3238
rect 236018 3002 236102 3238
rect 236338 3002 236422 3238
rect 236658 3002 236742 3238
rect 236978 3002 237062 3238
rect 237298 3002 237382 3238
rect 237618 3002 237740 3238
rect 233740 2918 237740 3002
rect 233740 2682 233862 2918
rect 234098 2682 234182 2918
rect 234418 2682 234502 2918
rect 234738 2682 234822 2918
rect 235058 2682 235142 2918
rect 235378 2682 235462 2918
rect 235698 2682 235782 2918
rect 236018 2682 236102 2918
rect 236338 2682 236422 2918
rect 236658 2682 236742 2918
rect 236978 2682 237062 2918
rect 237298 2682 237382 2918
rect 237618 2682 237740 2918
rect 233740 2598 237740 2682
rect 233740 2362 233862 2598
rect 234098 2362 234182 2598
rect 234418 2362 234502 2598
rect 234738 2362 234822 2598
rect 235058 2362 235142 2598
rect 235378 2362 235462 2598
rect 235698 2362 235782 2598
rect 236018 2362 236102 2598
rect 236338 2362 236422 2598
rect 236658 2362 236742 2598
rect 236978 2362 237062 2598
rect 237298 2362 237382 2598
rect 237618 2362 237740 2598
rect 233740 2278 237740 2362
rect 233740 2042 233862 2278
rect 234098 2042 234182 2278
rect 234418 2042 234502 2278
rect 234738 2042 234822 2278
rect 235058 2042 235142 2278
rect 235378 2042 235462 2278
rect 235698 2042 235782 2278
rect 236018 2042 236102 2278
rect 236338 2042 236422 2278
rect 236658 2042 236742 2278
rect 236978 2042 237062 2278
rect 237298 2042 237382 2278
rect 237618 2042 237740 2278
rect 233740 1958 237740 2042
rect 233740 1722 233862 1958
rect 234098 1722 234182 1958
rect 234418 1722 234502 1958
rect 234738 1722 234822 1958
rect 235058 1722 235142 1958
rect 235378 1722 235462 1958
rect 235698 1722 235782 1958
rect 236018 1722 236102 1958
rect 236338 1722 236422 1958
rect 236658 1722 236742 1958
rect 236978 1722 237062 1958
rect 237298 1722 237382 1958
rect 237618 1722 237740 1958
rect 233740 1638 237740 1722
rect 233740 1402 233862 1638
rect 234098 1402 234182 1638
rect 234418 1402 234502 1638
rect 234738 1402 234822 1638
rect 235058 1402 235142 1638
rect 235378 1402 235462 1638
rect 235698 1402 235782 1638
rect 236018 1402 236102 1638
rect 236338 1402 236422 1638
rect 236658 1402 236742 1638
rect 236978 1402 237062 1638
rect 237298 1402 237382 1638
rect 237618 1402 237740 1638
rect 233740 1318 237740 1402
rect 233740 1082 233862 1318
rect 234098 1082 234182 1318
rect 234418 1082 234502 1318
rect 234738 1082 234822 1318
rect 235058 1082 235142 1318
rect 235378 1082 235462 1318
rect 235698 1082 235782 1318
rect 236018 1082 236102 1318
rect 236338 1082 236422 1318
rect 236658 1082 236742 1318
rect 236978 1082 237062 1318
rect 237298 1082 237382 1318
rect 237618 1082 237740 1318
rect 233740 998 237740 1082
rect 233740 762 233862 998
rect 234098 762 234182 998
rect 234418 762 234502 998
rect 234738 762 234822 998
rect 235058 762 235142 998
rect 235378 762 235462 998
rect 235698 762 235782 998
rect 236018 762 236102 998
rect 236338 762 236422 998
rect 236658 762 236742 998
rect 236978 762 237062 998
rect 237298 762 237382 998
rect 237618 762 237740 998
rect 233740 678 237740 762
rect 233740 442 233862 678
rect 234098 442 234182 678
rect 234418 442 234502 678
rect 234738 442 234822 678
rect 235058 442 235142 678
rect 235378 442 235462 678
rect 235698 442 235782 678
rect 236018 442 236102 678
rect 236338 442 236422 678
rect 236658 442 236742 678
rect 236978 442 237062 678
rect 237298 442 237382 678
rect 237618 442 237740 678
rect 233740 358 237740 442
rect 233740 122 233862 358
rect 234098 122 234182 358
rect 234418 122 234502 358
rect 234738 122 234822 358
rect 235058 122 235142 358
rect 235378 122 235462 358
rect 235698 122 235782 358
rect 236018 122 236102 358
rect 236338 122 236422 358
rect 236658 122 236742 358
rect 236978 122 237062 358
rect 237298 122 237382 358
rect 237618 122 237740 358
rect 233740 0 237740 122
<< via4 >>
rect 122 255018 358 255254
rect 442 255018 678 255254
rect 762 255018 998 255254
rect 1082 255018 1318 255254
rect 1402 255018 1638 255254
rect 1722 255018 1958 255254
rect 2042 255018 2278 255254
rect 2362 255018 2598 255254
rect 2682 255018 2918 255254
rect 3002 255018 3238 255254
rect 3322 255018 3558 255254
rect 3642 255018 3878 255254
rect 122 254698 358 254934
rect 442 254698 678 254934
rect 762 254698 998 254934
rect 1082 254698 1318 254934
rect 1402 254698 1638 254934
rect 1722 254698 1958 254934
rect 2042 254698 2278 254934
rect 2362 254698 2598 254934
rect 2682 254698 2918 254934
rect 3002 254698 3238 254934
rect 3322 254698 3558 254934
rect 3642 254698 3878 254934
rect 122 254378 358 254614
rect 442 254378 678 254614
rect 762 254378 998 254614
rect 1082 254378 1318 254614
rect 1402 254378 1638 254614
rect 1722 254378 1958 254614
rect 2042 254378 2278 254614
rect 2362 254378 2598 254614
rect 2682 254378 2918 254614
rect 3002 254378 3238 254614
rect 3322 254378 3558 254614
rect 3642 254378 3878 254614
rect 122 254058 358 254294
rect 442 254058 678 254294
rect 762 254058 998 254294
rect 1082 254058 1318 254294
rect 1402 254058 1638 254294
rect 1722 254058 1958 254294
rect 2042 254058 2278 254294
rect 2362 254058 2598 254294
rect 2682 254058 2918 254294
rect 3002 254058 3238 254294
rect 3322 254058 3558 254294
rect 3642 254058 3878 254294
rect 122 253738 358 253974
rect 442 253738 678 253974
rect 762 253738 998 253974
rect 1082 253738 1318 253974
rect 1402 253738 1638 253974
rect 1722 253738 1958 253974
rect 2042 253738 2278 253974
rect 2362 253738 2598 253974
rect 2682 253738 2918 253974
rect 3002 253738 3238 253974
rect 3322 253738 3558 253974
rect 3642 253738 3878 253974
rect 122 253418 358 253654
rect 442 253418 678 253654
rect 762 253418 998 253654
rect 1082 253418 1318 253654
rect 1402 253418 1638 253654
rect 1722 253418 1958 253654
rect 2042 253418 2278 253654
rect 2362 253418 2598 253654
rect 2682 253418 2918 253654
rect 3002 253418 3238 253654
rect 3322 253418 3558 253654
rect 3642 253418 3878 253654
rect 122 253098 358 253334
rect 442 253098 678 253334
rect 762 253098 998 253334
rect 1082 253098 1318 253334
rect 1402 253098 1638 253334
rect 1722 253098 1958 253334
rect 2042 253098 2278 253334
rect 2362 253098 2598 253334
rect 2682 253098 2918 253334
rect 3002 253098 3238 253334
rect 3322 253098 3558 253334
rect 3642 253098 3878 253334
rect 122 252778 358 253014
rect 442 252778 678 253014
rect 762 252778 998 253014
rect 1082 252778 1318 253014
rect 1402 252778 1638 253014
rect 1722 252778 1958 253014
rect 2042 252778 2278 253014
rect 2362 252778 2598 253014
rect 2682 252778 2918 253014
rect 3002 252778 3238 253014
rect 3322 252778 3558 253014
rect 3642 252778 3878 253014
rect 122 252458 358 252694
rect 442 252458 678 252694
rect 762 252458 998 252694
rect 1082 252458 1318 252694
rect 1402 252458 1638 252694
rect 1722 252458 1958 252694
rect 2042 252458 2278 252694
rect 2362 252458 2598 252694
rect 2682 252458 2918 252694
rect 3002 252458 3238 252694
rect 3322 252458 3558 252694
rect 3642 252458 3878 252694
rect 122 252138 358 252374
rect 442 252138 678 252374
rect 762 252138 998 252374
rect 1082 252138 1318 252374
rect 1402 252138 1638 252374
rect 1722 252138 1958 252374
rect 2042 252138 2278 252374
rect 2362 252138 2598 252374
rect 2682 252138 2918 252374
rect 3002 252138 3238 252374
rect 3322 252138 3558 252374
rect 3642 252138 3878 252374
rect 122 251818 358 252054
rect 442 251818 678 252054
rect 762 251818 998 252054
rect 1082 251818 1318 252054
rect 1402 251818 1638 252054
rect 1722 251818 1958 252054
rect 2042 251818 2278 252054
rect 2362 251818 2598 252054
rect 2682 251818 2918 252054
rect 3002 251818 3238 252054
rect 3322 251818 3558 252054
rect 3642 251818 3878 252054
rect 122 251498 358 251734
rect 442 251498 678 251734
rect 762 251498 998 251734
rect 1082 251498 1318 251734
rect 1402 251498 1638 251734
rect 1722 251498 1958 251734
rect 2042 251498 2278 251734
rect 2362 251498 2598 251734
rect 2682 251498 2918 251734
rect 3002 251498 3238 251734
rect 3322 251498 3558 251734
rect 3642 251498 3878 251734
rect 233862 255018 234098 255254
rect 234182 255018 234418 255254
rect 234502 255018 234738 255254
rect 234822 255018 235058 255254
rect 235142 255018 235378 255254
rect 235462 255018 235698 255254
rect 235782 255018 236018 255254
rect 236102 255018 236338 255254
rect 236422 255018 236658 255254
rect 236742 255018 236978 255254
rect 237062 255018 237298 255254
rect 237382 255018 237618 255254
rect 233862 254698 234098 254934
rect 234182 254698 234418 254934
rect 234502 254698 234738 254934
rect 234822 254698 235058 254934
rect 235142 254698 235378 254934
rect 235462 254698 235698 254934
rect 235782 254698 236018 254934
rect 236102 254698 236338 254934
rect 236422 254698 236658 254934
rect 236742 254698 236978 254934
rect 237062 254698 237298 254934
rect 237382 254698 237618 254934
rect 233862 254378 234098 254614
rect 234182 254378 234418 254614
rect 234502 254378 234738 254614
rect 234822 254378 235058 254614
rect 235142 254378 235378 254614
rect 235462 254378 235698 254614
rect 235782 254378 236018 254614
rect 236102 254378 236338 254614
rect 236422 254378 236658 254614
rect 236742 254378 236978 254614
rect 237062 254378 237298 254614
rect 237382 254378 237618 254614
rect 233862 254058 234098 254294
rect 234182 254058 234418 254294
rect 234502 254058 234738 254294
rect 234822 254058 235058 254294
rect 235142 254058 235378 254294
rect 235462 254058 235698 254294
rect 235782 254058 236018 254294
rect 236102 254058 236338 254294
rect 236422 254058 236658 254294
rect 236742 254058 236978 254294
rect 237062 254058 237298 254294
rect 237382 254058 237618 254294
rect 233862 253738 234098 253974
rect 234182 253738 234418 253974
rect 234502 253738 234738 253974
rect 234822 253738 235058 253974
rect 235142 253738 235378 253974
rect 235462 253738 235698 253974
rect 235782 253738 236018 253974
rect 236102 253738 236338 253974
rect 236422 253738 236658 253974
rect 236742 253738 236978 253974
rect 237062 253738 237298 253974
rect 237382 253738 237618 253974
rect 233862 253418 234098 253654
rect 234182 253418 234418 253654
rect 234502 253418 234738 253654
rect 234822 253418 235058 253654
rect 235142 253418 235378 253654
rect 235462 253418 235698 253654
rect 235782 253418 236018 253654
rect 236102 253418 236338 253654
rect 236422 253418 236658 253654
rect 236742 253418 236978 253654
rect 237062 253418 237298 253654
rect 237382 253418 237618 253654
rect 233862 253098 234098 253334
rect 234182 253098 234418 253334
rect 234502 253098 234738 253334
rect 234822 253098 235058 253334
rect 235142 253098 235378 253334
rect 235462 253098 235698 253334
rect 235782 253098 236018 253334
rect 236102 253098 236338 253334
rect 236422 253098 236658 253334
rect 236742 253098 236978 253334
rect 237062 253098 237298 253334
rect 237382 253098 237618 253334
rect 233862 252778 234098 253014
rect 234182 252778 234418 253014
rect 234502 252778 234738 253014
rect 234822 252778 235058 253014
rect 235142 252778 235378 253014
rect 235462 252778 235698 253014
rect 235782 252778 236018 253014
rect 236102 252778 236338 253014
rect 236422 252778 236658 253014
rect 236742 252778 236978 253014
rect 237062 252778 237298 253014
rect 237382 252778 237618 253014
rect 233862 252458 234098 252694
rect 234182 252458 234418 252694
rect 234502 252458 234738 252694
rect 234822 252458 235058 252694
rect 235142 252458 235378 252694
rect 235462 252458 235698 252694
rect 235782 252458 236018 252694
rect 236102 252458 236338 252694
rect 236422 252458 236658 252694
rect 236742 252458 236978 252694
rect 237062 252458 237298 252694
rect 237382 252458 237618 252694
rect 233862 252138 234098 252374
rect 234182 252138 234418 252374
rect 234502 252138 234738 252374
rect 234822 252138 235058 252374
rect 235142 252138 235378 252374
rect 235462 252138 235698 252374
rect 235782 252138 236018 252374
rect 236102 252138 236338 252374
rect 236422 252138 236658 252374
rect 236742 252138 236978 252374
rect 237062 252138 237298 252374
rect 237382 252138 237618 252374
rect 233862 251818 234098 252054
rect 234182 251818 234418 252054
rect 234502 251818 234738 252054
rect 234822 251818 235058 252054
rect 235142 251818 235378 252054
rect 235462 251818 235698 252054
rect 235782 251818 236018 252054
rect 236102 251818 236338 252054
rect 236422 251818 236658 252054
rect 236742 251818 236978 252054
rect 237062 251818 237298 252054
rect 237382 251818 237618 252054
rect 233862 251498 234098 251734
rect 234182 251498 234418 251734
rect 234502 251498 234738 251734
rect 234822 251498 235058 251734
rect 235142 251498 235378 251734
rect 235462 251498 235698 251734
rect 235782 251498 236018 251734
rect 236102 251498 236338 251734
rect 236422 251498 236658 251734
rect 236742 251498 236978 251734
rect 237062 251498 237298 251734
rect 237382 251498 237618 251734
rect 122 228682 358 228918
rect 442 228682 678 228918
rect 762 228682 998 228918
rect 1082 228682 1318 228918
rect 1402 228682 1638 228918
rect 1722 228682 1958 228918
rect 2042 228682 2278 228918
rect 2362 228682 2598 228918
rect 2682 228682 2918 228918
rect 3002 228682 3238 228918
rect 3322 228682 3558 228918
rect 3642 228682 3878 228918
rect 122 206282 358 206518
rect 442 206282 678 206518
rect 762 206282 998 206518
rect 1082 206282 1318 206518
rect 1402 206282 1638 206518
rect 1722 206282 1958 206518
rect 2042 206282 2278 206518
rect 2362 206282 2598 206518
rect 2682 206282 2918 206518
rect 3002 206282 3238 206518
rect 3322 206282 3558 206518
rect 3642 206282 3878 206518
rect 122 183882 358 184118
rect 442 183882 678 184118
rect 762 183882 998 184118
rect 1082 183882 1318 184118
rect 1402 183882 1638 184118
rect 1722 183882 1958 184118
rect 2042 183882 2278 184118
rect 2362 183882 2598 184118
rect 2682 183882 2918 184118
rect 3002 183882 3238 184118
rect 3322 183882 3558 184118
rect 3642 183882 3878 184118
rect 122 161482 358 161718
rect 442 161482 678 161718
rect 762 161482 998 161718
rect 1082 161482 1318 161718
rect 1402 161482 1638 161718
rect 1722 161482 1958 161718
rect 2042 161482 2278 161718
rect 2362 161482 2598 161718
rect 2682 161482 2918 161718
rect 3002 161482 3238 161718
rect 3322 161482 3558 161718
rect 3642 161482 3878 161718
rect 122 139082 358 139318
rect 442 139082 678 139318
rect 762 139082 998 139318
rect 1082 139082 1318 139318
rect 1402 139082 1638 139318
rect 1722 139082 1958 139318
rect 2042 139082 2278 139318
rect 2362 139082 2598 139318
rect 2682 139082 2918 139318
rect 3002 139082 3238 139318
rect 3322 139082 3558 139318
rect 3642 139082 3878 139318
rect 122 116682 358 116918
rect 442 116682 678 116918
rect 762 116682 998 116918
rect 1082 116682 1318 116918
rect 1402 116682 1638 116918
rect 1722 116682 1958 116918
rect 2042 116682 2278 116918
rect 2362 116682 2598 116918
rect 2682 116682 2918 116918
rect 3002 116682 3238 116918
rect 3322 116682 3558 116918
rect 3642 116682 3878 116918
rect 122 94282 358 94518
rect 442 94282 678 94518
rect 762 94282 998 94518
rect 1082 94282 1318 94518
rect 1402 94282 1638 94518
rect 1722 94282 1958 94518
rect 2042 94282 2278 94518
rect 2362 94282 2598 94518
rect 2682 94282 2918 94518
rect 3002 94282 3238 94518
rect 3322 94282 3558 94518
rect 3642 94282 3878 94518
rect 122 71882 358 72118
rect 442 71882 678 72118
rect 762 71882 998 72118
rect 1082 71882 1318 72118
rect 1402 71882 1638 72118
rect 1722 71882 1958 72118
rect 2042 71882 2278 72118
rect 2362 71882 2598 72118
rect 2682 71882 2918 72118
rect 3002 71882 3238 72118
rect 3322 71882 3558 72118
rect 3642 71882 3878 72118
rect 122 49482 358 49718
rect 442 49482 678 49718
rect 762 49482 998 49718
rect 1082 49482 1318 49718
rect 1402 49482 1638 49718
rect 1722 49482 1958 49718
rect 2042 49482 2278 49718
rect 2362 49482 2598 49718
rect 2682 49482 2918 49718
rect 3002 49482 3238 49718
rect 3322 49482 3558 49718
rect 3642 49482 3878 49718
rect 122 27082 358 27318
rect 442 27082 678 27318
rect 762 27082 998 27318
rect 1082 27082 1318 27318
rect 1402 27082 1638 27318
rect 1722 27082 1958 27318
rect 2042 27082 2278 27318
rect 2362 27082 2598 27318
rect 2682 27082 2918 27318
rect 3002 27082 3238 27318
rect 3322 27082 3558 27318
rect 3642 27082 3878 27318
rect 5122 250018 5358 250254
rect 5442 250018 5678 250254
rect 5762 250018 5998 250254
rect 6082 250018 6318 250254
rect 6402 250018 6638 250254
rect 6722 250018 6958 250254
rect 7042 250018 7278 250254
rect 7362 250018 7598 250254
rect 7682 250018 7918 250254
rect 8002 250018 8238 250254
rect 8322 250018 8558 250254
rect 8642 250018 8878 250254
rect 5122 249698 5358 249934
rect 5442 249698 5678 249934
rect 5762 249698 5998 249934
rect 6082 249698 6318 249934
rect 6402 249698 6638 249934
rect 6722 249698 6958 249934
rect 7042 249698 7278 249934
rect 7362 249698 7598 249934
rect 7682 249698 7918 249934
rect 8002 249698 8238 249934
rect 8322 249698 8558 249934
rect 8642 249698 8878 249934
rect 5122 249378 5358 249614
rect 5442 249378 5678 249614
rect 5762 249378 5998 249614
rect 6082 249378 6318 249614
rect 6402 249378 6638 249614
rect 6722 249378 6958 249614
rect 7042 249378 7278 249614
rect 7362 249378 7598 249614
rect 7682 249378 7918 249614
rect 8002 249378 8238 249614
rect 8322 249378 8558 249614
rect 8642 249378 8878 249614
rect 5122 249058 5358 249294
rect 5442 249058 5678 249294
rect 5762 249058 5998 249294
rect 6082 249058 6318 249294
rect 6402 249058 6638 249294
rect 6722 249058 6958 249294
rect 7042 249058 7278 249294
rect 7362 249058 7598 249294
rect 7682 249058 7918 249294
rect 8002 249058 8238 249294
rect 8322 249058 8558 249294
rect 8642 249058 8878 249294
rect 5122 248738 5358 248974
rect 5442 248738 5678 248974
rect 5762 248738 5998 248974
rect 6082 248738 6318 248974
rect 6402 248738 6638 248974
rect 6722 248738 6958 248974
rect 7042 248738 7278 248974
rect 7362 248738 7598 248974
rect 7682 248738 7918 248974
rect 8002 248738 8238 248974
rect 8322 248738 8558 248974
rect 8642 248738 8878 248974
rect 5122 248418 5358 248654
rect 5442 248418 5678 248654
rect 5762 248418 5998 248654
rect 6082 248418 6318 248654
rect 6402 248418 6638 248654
rect 6722 248418 6958 248654
rect 7042 248418 7278 248654
rect 7362 248418 7598 248654
rect 7682 248418 7918 248654
rect 8002 248418 8238 248654
rect 8322 248418 8558 248654
rect 8642 248418 8878 248654
rect 5122 248098 5358 248334
rect 5442 248098 5678 248334
rect 5762 248098 5998 248334
rect 6082 248098 6318 248334
rect 6402 248098 6638 248334
rect 6722 248098 6958 248334
rect 7042 248098 7278 248334
rect 7362 248098 7598 248334
rect 7682 248098 7918 248334
rect 8002 248098 8238 248334
rect 8322 248098 8558 248334
rect 8642 248098 8878 248334
rect 5122 247778 5358 248014
rect 5442 247778 5678 248014
rect 5762 247778 5998 248014
rect 6082 247778 6318 248014
rect 6402 247778 6638 248014
rect 6722 247778 6958 248014
rect 7042 247778 7278 248014
rect 7362 247778 7598 248014
rect 7682 247778 7918 248014
rect 8002 247778 8238 248014
rect 8322 247778 8558 248014
rect 8642 247778 8878 248014
rect 5122 247458 5358 247694
rect 5442 247458 5678 247694
rect 5762 247458 5998 247694
rect 6082 247458 6318 247694
rect 6402 247458 6638 247694
rect 6722 247458 6958 247694
rect 7042 247458 7278 247694
rect 7362 247458 7598 247694
rect 7682 247458 7918 247694
rect 8002 247458 8238 247694
rect 8322 247458 8558 247694
rect 8642 247458 8878 247694
rect 5122 247138 5358 247374
rect 5442 247138 5678 247374
rect 5762 247138 5998 247374
rect 6082 247138 6318 247374
rect 6402 247138 6638 247374
rect 6722 247138 6958 247374
rect 7042 247138 7278 247374
rect 7362 247138 7598 247374
rect 7682 247138 7918 247374
rect 8002 247138 8238 247374
rect 8322 247138 8558 247374
rect 8642 247138 8878 247374
rect 5122 246818 5358 247054
rect 5442 246818 5678 247054
rect 5762 246818 5998 247054
rect 6082 246818 6318 247054
rect 6402 246818 6638 247054
rect 6722 246818 6958 247054
rect 7042 246818 7278 247054
rect 7362 246818 7598 247054
rect 7682 246818 7918 247054
rect 8002 246818 8238 247054
rect 8322 246818 8558 247054
rect 8642 246818 8878 247054
rect 5122 246498 5358 246734
rect 5442 246498 5678 246734
rect 5762 246498 5998 246734
rect 6082 246498 6318 246734
rect 6402 246498 6638 246734
rect 6722 246498 6958 246734
rect 7042 246498 7278 246734
rect 7362 246498 7598 246734
rect 7682 246498 7918 246734
rect 8002 246498 8238 246734
rect 8322 246498 8558 246734
rect 8642 246498 8878 246734
rect 228862 250018 229098 250254
rect 229182 250018 229418 250254
rect 229502 250018 229738 250254
rect 229822 250018 230058 250254
rect 230142 250018 230378 250254
rect 230462 250018 230698 250254
rect 230782 250018 231018 250254
rect 231102 250018 231338 250254
rect 231422 250018 231658 250254
rect 231742 250018 231978 250254
rect 232062 250018 232298 250254
rect 232382 250018 232618 250254
rect 228862 249698 229098 249934
rect 229182 249698 229418 249934
rect 229502 249698 229738 249934
rect 229822 249698 230058 249934
rect 230142 249698 230378 249934
rect 230462 249698 230698 249934
rect 230782 249698 231018 249934
rect 231102 249698 231338 249934
rect 231422 249698 231658 249934
rect 231742 249698 231978 249934
rect 232062 249698 232298 249934
rect 232382 249698 232618 249934
rect 228862 249378 229098 249614
rect 229182 249378 229418 249614
rect 229502 249378 229738 249614
rect 229822 249378 230058 249614
rect 230142 249378 230378 249614
rect 230462 249378 230698 249614
rect 230782 249378 231018 249614
rect 231102 249378 231338 249614
rect 231422 249378 231658 249614
rect 231742 249378 231978 249614
rect 232062 249378 232298 249614
rect 232382 249378 232618 249614
rect 228862 249058 229098 249294
rect 229182 249058 229418 249294
rect 229502 249058 229738 249294
rect 229822 249058 230058 249294
rect 230142 249058 230378 249294
rect 230462 249058 230698 249294
rect 230782 249058 231018 249294
rect 231102 249058 231338 249294
rect 231422 249058 231658 249294
rect 231742 249058 231978 249294
rect 232062 249058 232298 249294
rect 232382 249058 232618 249294
rect 228862 248738 229098 248974
rect 229182 248738 229418 248974
rect 229502 248738 229738 248974
rect 229822 248738 230058 248974
rect 230142 248738 230378 248974
rect 230462 248738 230698 248974
rect 230782 248738 231018 248974
rect 231102 248738 231338 248974
rect 231422 248738 231658 248974
rect 231742 248738 231978 248974
rect 232062 248738 232298 248974
rect 232382 248738 232618 248974
rect 228862 248418 229098 248654
rect 229182 248418 229418 248654
rect 229502 248418 229738 248654
rect 229822 248418 230058 248654
rect 230142 248418 230378 248654
rect 230462 248418 230698 248654
rect 230782 248418 231018 248654
rect 231102 248418 231338 248654
rect 231422 248418 231658 248654
rect 231742 248418 231978 248654
rect 232062 248418 232298 248654
rect 232382 248418 232618 248654
rect 228862 248098 229098 248334
rect 229182 248098 229418 248334
rect 229502 248098 229738 248334
rect 229822 248098 230058 248334
rect 230142 248098 230378 248334
rect 230462 248098 230698 248334
rect 230782 248098 231018 248334
rect 231102 248098 231338 248334
rect 231422 248098 231658 248334
rect 231742 248098 231978 248334
rect 232062 248098 232298 248334
rect 232382 248098 232618 248334
rect 228862 247778 229098 248014
rect 229182 247778 229418 248014
rect 229502 247778 229738 248014
rect 229822 247778 230058 248014
rect 230142 247778 230378 248014
rect 230462 247778 230698 248014
rect 230782 247778 231018 248014
rect 231102 247778 231338 248014
rect 231422 247778 231658 248014
rect 231742 247778 231978 248014
rect 232062 247778 232298 248014
rect 232382 247778 232618 248014
rect 228862 247458 229098 247694
rect 229182 247458 229418 247694
rect 229502 247458 229738 247694
rect 229822 247458 230058 247694
rect 230142 247458 230378 247694
rect 230462 247458 230698 247694
rect 230782 247458 231018 247694
rect 231102 247458 231338 247694
rect 231422 247458 231658 247694
rect 231742 247458 231978 247694
rect 232062 247458 232298 247694
rect 232382 247458 232618 247694
rect 228862 247138 229098 247374
rect 229182 247138 229418 247374
rect 229502 247138 229738 247374
rect 229822 247138 230058 247374
rect 230142 247138 230378 247374
rect 230462 247138 230698 247374
rect 230782 247138 231018 247374
rect 231102 247138 231338 247374
rect 231422 247138 231658 247374
rect 231742 247138 231978 247374
rect 232062 247138 232298 247374
rect 232382 247138 232618 247374
rect 228862 246818 229098 247054
rect 229182 246818 229418 247054
rect 229502 246818 229738 247054
rect 229822 246818 230058 247054
rect 230142 246818 230378 247054
rect 230462 246818 230698 247054
rect 230782 246818 231018 247054
rect 231102 246818 231338 247054
rect 231422 246818 231658 247054
rect 231742 246818 231978 247054
rect 232062 246818 232298 247054
rect 232382 246818 232618 247054
rect 228862 246498 229098 246734
rect 229182 246498 229418 246734
rect 229502 246498 229738 246734
rect 229822 246498 230058 246734
rect 230142 246498 230378 246734
rect 230462 246498 230698 246734
rect 230782 246498 231018 246734
rect 231102 246498 231338 246734
rect 231422 246498 231658 246734
rect 231742 246498 231978 246734
rect 232062 246498 232298 246734
rect 232382 246498 232618 246734
rect 5122 239882 5358 240118
rect 5442 239882 5678 240118
rect 5762 239882 5998 240118
rect 6082 239882 6318 240118
rect 6402 239882 6638 240118
rect 6722 239882 6958 240118
rect 7042 239882 7278 240118
rect 7362 239882 7598 240118
rect 7682 239882 7918 240118
rect 8002 239882 8238 240118
rect 8322 239882 8558 240118
rect 8642 239882 8878 240118
rect 72816 239882 73052 240118
rect 144816 239882 145052 240118
rect 228862 239882 229098 240118
rect 229182 239882 229418 240118
rect 229502 239882 229738 240118
rect 229822 239882 230058 240118
rect 230142 239882 230378 240118
rect 230462 239882 230698 240118
rect 230782 239882 231018 240118
rect 231102 239882 231338 240118
rect 231422 239882 231658 240118
rect 231742 239882 231978 240118
rect 232062 239882 232298 240118
rect 232382 239882 232618 240118
rect 77816 228682 78052 228918
rect 149816 228682 150052 228918
rect 5122 217482 5358 217718
rect 5442 217482 5678 217718
rect 5762 217482 5998 217718
rect 6082 217482 6318 217718
rect 6402 217482 6638 217718
rect 6722 217482 6958 217718
rect 7042 217482 7278 217718
rect 7362 217482 7598 217718
rect 7682 217482 7918 217718
rect 8002 217482 8238 217718
rect 8322 217482 8558 217718
rect 8642 217482 8878 217718
rect 228862 217482 229098 217718
rect 229182 217482 229418 217718
rect 229502 217482 229738 217718
rect 229822 217482 230058 217718
rect 230142 217482 230378 217718
rect 230462 217482 230698 217718
rect 230782 217482 231018 217718
rect 231102 217482 231338 217718
rect 231422 217482 231658 217718
rect 231742 217482 231978 217718
rect 232062 217482 232298 217718
rect 232382 217482 232618 217718
rect 5122 195082 5358 195318
rect 5442 195082 5678 195318
rect 5762 195082 5998 195318
rect 6082 195082 6318 195318
rect 6402 195082 6638 195318
rect 6722 195082 6958 195318
rect 7042 195082 7278 195318
rect 7362 195082 7598 195318
rect 7682 195082 7918 195318
rect 8002 195082 8238 195318
rect 8322 195082 8558 195318
rect 8642 195082 8878 195318
rect 5122 172682 5358 172918
rect 5442 172682 5678 172918
rect 5762 172682 5998 172918
rect 6082 172682 6318 172918
rect 6402 172682 6638 172918
rect 6722 172682 6958 172918
rect 7042 172682 7278 172918
rect 7362 172682 7598 172918
rect 7682 172682 7918 172918
rect 8002 172682 8238 172918
rect 8322 172682 8558 172918
rect 8642 172682 8878 172918
rect 17549 172682 17785 172918
rect 20215 161482 20451 161718
rect 42927 206282 43163 206518
rect 78882 206282 79118 206518
rect 115215 206282 115451 206518
rect 150882 206282 151118 206518
rect 187215 206282 187451 206518
rect 38261 195082 38497 195318
rect 73882 195082 74118 195318
rect 110549 195082 110785 195318
rect 145882 195082 146118 195318
rect 182549 195082 182785 195318
rect 228862 195082 229098 195318
rect 229182 195082 229418 195318
rect 229502 195082 229738 195318
rect 229822 195082 230058 195318
rect 230142 195082 230378 195318
rect 230462 195082 230698 195318
rect 230782 195082 231018 195318
rect 231102 195082 231338 195318
rect 231422 195082 231658 195318
rect 231742 195082 231978 195318
rect 232062 195082 232298 195318
rect 232382 195082 232618 195318
rect 42549 172682 42785 172918
rect 67146 172682 67382 172918
rect 114549 172682 114785 172918
rect 139146 172682 139382 172918
rect 186549 172682 186785 172918
rect 211549 172682 211785 172918
rect 228862 172682 229098 172918
rect 229182 172682 229418 172918
rect 229502 172682 229738 172918
rect 229822 172682 230058 172918
rect 230142 172682 230378 172918
rect 230462 172682 230698 172918
rect 230782 172682 231018 172918
rect 231102 172682 231338 172918
rect 231422 172682 231658 172918
rect 231742 172682 231978 172918
rect 232062 172682 232298 172918
rect 232382 172682 232618 172918
rect 45215 161482 45451 161718
rect 82506 161482 82742 161718
rect 117215 161482 117451 161718
rect 154506 161482 154742 161718
rect 189215 161482 189451 161718
rect 214215 161482 214451 161718
rect 5122 150282 5358 150518
rect 5442 150282 5678 150518
rect 5762 150282 5998 150518
rect 6082 150282 6318 150518
rect 6402 150282 6638 150518
rect 6722 150282 6958 150518
rect 7042 150282 7278 150518
rect 7362 150282 7598 150518
rect 7682 150282 7918 150518
rect 8002 150282 8238 150518
rect 8322 150282 8558 150518
rect 8642 150282 8878 150518
rect 17549 150282 17785 150518
rect 42549 150282 42785 150518
rect 67146 150282 67382 150518
rect 114549 150282 114785 150518
rect 139146 150282 139382 150518
rect 186549 150282 186785 150518
rect 211549 150282 211785 150518
rect 228862 150282 229098 150518
rect 229182 150282 229418 150518
rect 229502 150282 229738 150518
rect 229822 150282 230058 150518
rect 230142 150282 230378 150518
rect 230462 150282 230698 150518
rect 230782 150282 231018 150518
rect 231102 150282 231338 150518
rect 231422 150282 231658 150518
rect 231742 150282 231978 150518
rect 232062 150282 232298 150518
rect 232382 150282 232618 150518
rect 21462 128726 21698 128962
rect 5122 127882 5358 128118
rect 5442 127882 5678 128118
rect 5762 127882 5998 128118
rect 6082 127882 6318 128118
rect 6402 127882 6638 128118
rect 6722 127882 6958 128118
rect 7042 127882 7278 128118
rect 7362 127882 7598 128118
rect 7682 127882 7918 128118
rect 8002 127882 8238 128118
rect 8322 127882 8558 128118
rect 8642 127882 8878 128118
rect 43215 139082 43451 139318
rect 67646 131446 67882 131682
rect 67646 128726 67882 128962
rect 38549 127882 38785 128118
rect 73882 127882 74118 128118
rect 43215 116682 43451 116918
rect 31766 113766 32002 114002
rect 56790 113766 57026 114002
rect 72982 113236 73218 113322
rect 72982 113172 73068 113236
rect 73068 113172 73132 113236
rect 73132 113172 73218 113236
rect 72982 113086 73218 113172
rect 5122 105482 5358 105718
rect 5442 105482 5678 105718
rect 5762 105482 5998 105718
rect 6082 105482 6318 105718
rect 6402 105482 6638 105718
rect 6722 105482 6958 105718
rect 7042 105482 7278 105718
rect 7362 105482 7598 105718
rect 7682 105482 7918 105718
rect 8002 105482 8238 105718
rect 8322 105482 8558 105718
rect 8642 105482 8878 105718
rect 17549 105482 17785 105718
rect 42549 105482 42785 105718
rect 67146 105482 67382 105718
rect 20215 94282 20451 94518
rect 45215 94282 45451 94518
rect 82506 94282 82742 94518
rect 5122 83082 5358 83318
rect 5442 83082 5678 83318
rect 5762 83082 5998 83318
rect 6082 83082 6318 83318
rect 6402 83082 6638 83318
rect 6722 83082 6958 83318
rect 7042 83082 7278 83318
rect 7362 83082 7598 83318
rect 7682 83082 7918 83318
rect 8002 83082 8238 83318
rect 8322 83082 8558 83318
rect 8642 83082 8878 83318
rect 17549 83082 17785 83318
rect 42549 83082 42785 83318
rect 67146 83082 67382 83318
rect 115215 139082 115451 139318
rect 146214 138246 146450 138482
rect 142534 136886 142770 137122
rect 101318 131460 101554 131682
rect 101318 131446 101404 131460
rect 101404 131446 101468 131460
rect 101468 131446 101554 131460
rect 110549 127882 110785 128118
rect 145882 127882 146118 128118
rect 115215 116682 115451 116918
rect 187215 139082 187451 139318
rect 182549 127882 182785 128118
rect 228862 127882 229098 128118
rect 229182 127882 229418 128118
rect 229502 127882 229738 128118
rect 229822 127882 230058 128118
rect 230142 127882 230378 128118
rect 230462 127882 230698 128118
rect 230782 127882 231018 128118
rect 231102 127882 231338 128118
rect 231422 127882 231658 128118
rect 231742 127882 231978 128118
rect 232062 127882 232298 128118
rect 232382 127882 232618 128118
rect 187215 116682 187451 116918
rect 114549 105482 114785 105718
rect 139146 105482 139382 105718
rect 186549 105482 186785 105718
rect 211549 105482 211785 105718
rect 228862 105482 229098 105718
rect 229182 105482 229418 105718
rect 229502 105482 229738 105718
rect 229822 105482 230058 105718
rect 230142 105482 230378 105718
rect 230462 105482 230698 105718
rect 230782 105482 231018 105718
rect 231102 105482 231338 105718
rect 231422 105482 231658 105718
rect 231742 105482 231978 105718
rect 232062 105482 232298 105718
rect 232382 105482 232618 105718
rect 117215 94282 117451 94518
rect 154506 94282 154742 94518
rect 189215 94282 189451 94518
rect 214215 94282 214451 94518
rect 114549 83082 114785 83318
rect 139146 83082 139382 83318
rect 186549 83082 186785 83318
rect 211549 83082 211785 83318
rect 228862 83082 229098 83318
rect 229182 83082 229418 83318
rect 229502 83082 229738 83318
rect 229822 83082 230058 83318
rect 230142 83082 230378 83318
rect 230462 83082 230698 83318
rect 230782 83082 231018 83318
rect 231102 83082 231338 83318
rect 231422 83082 231658 83318
rect 231742 83082 231978 83318
rect 232062 83082 232298 83318
rect 232382 83082 232618 83318
rect 5122 60682 5358 60918
rect 5442 60682 5678 60918
rect 5762 60682 5998 60918
rect 6082 60682 6318 60918
rect 6402 60682 6638 60918
rect 6722 60682 6958 60918
rect 7042 60682 7278 60918
rect 7362 60682 7598 60918
rect 7682 60682 7918 60918
rect 8002 60682 8238 60918
rect 8322 60682 8558 60918
rect 8642 60682 8878 60918
rect 38549 60682 38785 60918
rect 73882 60682 74118 60918
rect 110549 60682 110785 60918
rect 43215 49482 43451 49718
rect 78882 49482 79118 49718
rect 115215 49482 115451 49718
rect 31766 41006 32002 41242
rect 66174 41006 66410 41242
rect 145882 60682 146118 60918
rect 182549 60682 182785 60918
rect 150882 49482 151118 49718
rect 187215 49482 187451 49718
rect 228862 60682 229098 60918
rect 229182 60682 229418 60918
rect 229502 60682 229738 60918
rect 229822 60682 230058 60918
rect 230142 60682 230378 60918
rect 230462 60682 230698 60918
rect 230782 60682 231018 60918
rect 231102 60682 231338 60918
rect 231422 60682 231658 60918
rect 231742 60682 231978 60918
rect 232062 60682 232298 60918
rect 232382 60682 232618 60918
rect 93774 40476 94010 40562
rect 93774 40412 93860 40476
rect 93860 40412 93924 40476
rect 93924 40412 94010 40476
rect 93774 40326 94010 40412
rect 108678 40326 108914 40562
rect 109598 40326 109834 40562
rect 129654 40326 129890 40562
rect 136830 40326 137066 40562
rect 181358 40326 181594 40562
rect 166086 39796 166322 39882
rect 166086 39732 166172 39796
rect 166172 39732 166236 39796
rect 166236 39732 166322 39796
rect 166086 39646 166322 39732
rect 201414 38966 201650 39202
rect 5122 38282 5358 38518
rect 5442 38282 5678 38518
rect 5762 38282 5998 38518
rect 6082 38282 6318 38518
rect 6402 38282 6638 38518
rect 6722 38282 6958 38518
rect 7042 38282 7278 38518
rect 7362 38282 7598 38518
rect 7682 38282 7918 38518
rect 8002 38282 8238 38518
rect 8322 38282 8558 38518
rect 8642 38282 8878 38518
rect 228862 38282 229098 38518
rect 229182 38282 229418 38518
rect 229502 38282 229738 38518
rect 229822 38282 230058 38518
rect 230142 38282 230378 38518
rect 230462 38282 230698 38518
rect 230782 38282 231018 38518
rect 231102 38282 231338 38518
rect 231422 38282 231658 38518
rect 231742 38282 231978 38518
rect 232062 38282 232298 38518
rect 232382 38282 232618 38518
rect 78882 27082 79118 27318
rect 150882 27082 151118 27318
rect 5122 15882 5358 16118
rect 5442 15882 5678 16118
rect 5762 15882 5998 16118
rect 6082 15882 6318 16118
rect 6402 15882 6638 16118
rect 6722 15882 6958 16118
rect 7042 15882 7278 16118
rect 7362 15882 7598 16118
rect 7682 15882 7918 16118
rect 8002 15882 8238 16118
rect 8322 15882 8558 16118
rect 8642 15882 8878 16118
rect 73882 15882 74118 16118
rect 145882 15882 146118 16118
rect 228862 15882 229098 16118
rect 229182 15882 229418 16118
rect 229502 15882 229738 16118
rect 229822 15882 230058 16118
rect 230142 15882 230378 16118
rect 230462 15882 230698 16118
rect 230782 15882 231018 16118
rect 231102 15882 231338 16118
rect 231422 15882 231658 16118
rect 231742 15882 231978 16118
rect 232062 15882 232298 16118
rect 232382 15882 232618 16118
rect 5122 8642 5358 8878
rect 5442 8642 5678 8878
rect 5762 8642 5998 8878
rect 6082 8642 6318 8878
rect 6402 8642 6638 8878
rect 6722 8642 6958 8878
rect 7042 8642 7278 8878
rect 7362 8642 7598 8878
rect 7682 8642 7918 8878
rect 8002 8642 8238 8878
rect 8322 8642 8558 8878
rect 8642 8642 8878 8878
rect 5122 8322 5358 8558
rect 5442 8322 5678 8558
rect 5762 8322 5998 8558
rect 6082 8322 6318 8558
rect 6402 8322 6638 8558
rect 6722 8322 6958 8558
rect 7042 8322 7278 8558
rect 7362 8322 7598 8558
rect 7682 8322 7918 8558
rect 8002 8322 8238 8558
rect 8322 8322 8558 8558
rect 8642 8322 8878 8558
rect 5122 8002 5358 8238
rect 5442 8002 5678 8238
rect 5762 8002 5998 8238
rect 6082 8002 6318 8238
rect 6402 8002 6638 8238
rect 6722 8002 6958 8238
rect 7042 8002 7278 8238
rect 7362 8002 7598 8238
rect 7682 8002 7918 8238
rect 8002 8002 8238 8238
rect 8322 8002 8558 8238
rect 8642 8002 8878 8238
rect 5122 7682 5358 7918
rect 5442 7682 5678 7918
rect 5762 7682 5998 7918
rect 6082 7682 6318 7918
rect 6402 7682 6638 7918
rect 6722 7682 6958 7918
rect 7042 7682 7278 7918
rect 7362 7682 7598 7918
rect 7682 7682 7918 7918
rect 8002 7682 8238 7918
rect 8322 7682 8558 7918
rect 8642 7682 8878 7918
rect 5122 7362 5358 7598
rect 5442 7362 5678 7598
rect 5762 7362 5998 7598
rect 6082 7362 6318 7598
rect 6402 7362 6638 7598
rect 6722 7362 6958 7598
rect 7042 7362 7278 7598
rect 7362 7362 7598 7598
rect 7682 7362 7918 7598
rect 8002 7362 8238 7598
rect 8322 7362 8558 7598
rect 8642 7362 8878 7598
rect 5122 7042 5358 7278
rect 5442 7042 5678 7278
rect 5762 7042 5998 7278
rect 6082 7042 6318 7278
rect 6402 7042 6638 7278
rect 6722 7042 6958 7278
rect 7042 7042 7278 7278
rect 7362 7042 7598 7278
rect 7682 7042 7918 7278
rect 8002 7042 8238 7278
rect 8322 7042 8558 7278
rect 8642 7042 8878 7278
rect 5122 6722 5358 6958
rect 5442 6722 5678 6958
rect 5762 6722 5998 6958
rect 6082 6722 6318 6958
rect 6402 6722 6638 6958
rect 6722 6722 6958 6958
rect 7042 6722 7278 6958
rect 7362 6722 7598 6958
rect 7682 6722 7918 6958
rect 8002 6722 8238 6958
rect 8322 6722 8558 6958
rect 8642 6722 8878 6958
rect 5122 6402 5358 6638
rect 5442 6402 5678 6638
rect 5762 6402 5998 6638
rect 6082 6402 6318 6638
rect 6402 6402 6638 6638
rect 6722 6402 6958 6638
rect 7042 6402 7278 6638
rect 7362 6402 7598 6638
rect 7682 6402 7918 6638
rect 8002 6402 8238 6638
rect 8322 6402 8558 6638
rect 8642 6402 8878 6638
rect 5122 6082 5358 6318
rect 5442 6082 5678 6318
rect 5762 6082 5998 6318
rect 6082 6082 6318 6318
rect 6402 6082 6638 6318
rect 6722 6082 6958 6318
rect 7042 6082 7278 6318
rect 7362 6082 7598 6318
rect 7682 6082 7918 6318
rect 8002 6082 8238 6318
rect 8322 6082 8558 6318
rect 8642 6082 8878 6318
rect 5122 5762 5358 5998
rect 5442 5762 5678 5998
rect 5762 5762 5998 5998
rect 6082 5762 6318 5998
rect 6402 5762 6638 5998
rect 6722 5762 6958 5998
rect 7042 5762 7278 5998
rect 7362 5762 7598 5998
rect 7682 5762 7918 5998
rect 8002 5762 8238 5998
rect 8322 5762 8558 5998
rect 8642 5762 8878 5998
rect 5122 5442 5358 5678
rect 5442 5442 5678 5678
rect 5762 5442 5998 5678
rect 6082 5442 6318 5678
rect 6402 5442 6638 5678
rect 6722 5442 6958 5678
rect 7042 5442 7278 5678
rect 7362 5442 7598 5678
rect 7682 5442 7918 5678
rect 8002 5442 8238 5678
rect 8322 5442 8558 5678
rect 8642 5442 8878 5678
rect 5122 5122 5358 5358
rect 5442 5122 5678 5358
rect 5762 5122 5998 5358
rect 6082 5122 6318 5358
rect 6402 5122 6638 5358
rect 6722 5122 6958 5358
rect 7042 5122 7278 5358
rect 7362 5122 7598 5358
rect 7682 5122 7918 5358
rect 8002 5122 8238 5358
rect 8322 5122 8558 5358
rect 8642 5122 8878 5358
rect 228862 8642 229098 8878
rect 229182 8642 229418 8878
rect 229502 8642 229738 8878
rect 229822 8642 230058 8878
rect 230142 8642 230378 8878
rect 230462 8642 230698 8878
rect 230782 8642 231018 8878
rect 231102 8642 231338 8878
rect 231422 8642 231658 8878
rect 231742 8642 231978 8878
rect 232062 8642 232298 8878
rect 232382 8642 232618 8878
rect 228862 8322 229098 8558
rect 229182 8322 229418 8558
rect 229502 8322 229738 8558
rect 229822 8322 230058 8558
rect 230142 8322 230378 8558
rect 230462 8322 230698 8558
rect 230782 8322 231018 8558
rect 231102 8322 231338 8558
rect 231422 8322 231658 8558
rect 231742 8322 231978 8558
rect 232062 8322 232298 8558
rect 232382 8322 232618 8558
rect 228862 8002 229098 8238
rect 229182 8002 229418 8238
rect 229502 8002 229738 8238
rect 229822 8002 230058 8238
rect 230142 8002 230378 8238
rect 230462 8002 230698 8238
rect 230782 8002 231018 8238
rect 231102 8002 231338 8238
rect 231422 8002 231658 8238
rect 231742 8002 231978 8238
rect 232062 8002 232298 8238
rect 232382 8002 232618 8238
rect 228862 7682 229098 7918
rect 229182 7682 229418 7918
rect 229502 7682 229738 7918
rect 229822 7682 230058 7918
rect 230142 7682 230378 7918
rect 230462 7682 230698 7918
rect 230782 7682 231018 7918
rect 231102 7682 231338 7918
rect 231422 7682 231658 7918
rect 231742 7682 231978 7918
rect 232062 7682 232298 7918
rect 232382 7682 232618 7918
rect 228862 7362 229098 7598
rect 229182 7362 229418 7598
rect 229502 7362 229738 7598
rect 229822 7362 230058 7598
rect 230142 7362 230378 7598
rect 230462 7362 230698 7598
rect 230782 7362 231018 7598
rect 231102 7362 231338 7598
rect 231422 7362 231658 7598
rect 231742 7362 231978 7598
rect 232062 7362 232298 7598
rect 232382 7362 232618 7598
rect 228862 7042 229098 7278
rect 229182 7042 229418 7278
rect 229502 7042 229738 7278
rect 229822 7042 230058 7278
rect 230142 7042 230378 7278
rect 230462 7042 230698 7278
rect 230782 7042 231018 7278
rect 231102 7042 231338 7278
rect 231422 7042 231658 7278
rect 231742 7042 231978 7278
rect 232062 7042 232298 7278
rect 232382 7042 232618 7278
rect 228862 6722 229098 6958
rect 229182 6722 229418 6958
rect 229502 6722 229738 6958
rect 229822 6722 230058 6958
rect 230142 6722 230378 6958
rect 230462 6722 230698 6958
rect 230782 6722 231018 6958
rect 231102 6722 231338 6958
rect 231422 6722 231658 6958
rect 231742 6722 231978 6958
rect 232062 6722 232298 6958
rect 232382 6722 232618 6958
rect 228862 6402 229098 6638
rect 229182 6402 229418 6638
rect 229502 6402 229738 6638
rect 229822 6402 230058 6638
rect 230142 6402 230378 6638
rect 230462 6402 230698 6638
rect 230782 6402 231018 6638
rect 231102 6402 231338 6638
rect 231422 6402 231658 6638
rect 231742 6402 231978 6638
rect 232062 6402 232298 6638
rect 232382 6402 232618 6638
rect 228862 6082 229098 6318
rect 229182 6082 229418 6318
rect 229502 6082 229738 6318
rect 229822 6082 230058 6318
rect 230142 6082 230378 6318
rect 230462 6082 230698 6318
rect 230782 6082 231018 6318
rect 231102 6082 231338 6318
rect 231422 6082 231658 6318
rect 231742 6082 231978 6318
rect 232062 6082 232298 6318
rect 232382 6082 232618 6318
rect 228862 5762 229098 5998
rect 229182 5762 229418 5998
rect 229502 5762 229738 5998
rect 229822 5762 230058 5998
rect 230142 5762 230378 5998
rect 230462 5762 230698 5998
rect 230782 5762 231018 5998
rect 231102 5762 231338 5998
rect 231422 5762 231658 5998
rect 231742 5762 231978 5998
rect 232062 5762 232298 5998
rect 232382 5762 232618 5998
rect 228862 5442 229098 5678
rect 229182 5442 229418 5678
rect 229502 5442 229738 5678
rect 229822 5442 230058 5678
rect 230142 5442 230378 5678
rect 230462 5442 230698 5678
rect 230782 5442 231018 5678
rect 231102 5442 231338 5678
rect 231422 5442 231658 5678
rect 231742 5442 231978 5678
rect 232062 5442 232298 5678
rect 232382 5442 232618 5678
rect 228862 5122 229098 5358
rect 229182 5122 229418 5358
rect 229502 5122 229738 5358
rect 229822 5122 230058 5358
rect 230142 5122 230378 5358
rect 230462 5122 230698 5358
rect 230782 5122 231018 5358
rect 231102 5122 231338 5358
rect 231422 5122 231658 5358
rect 231742 5122 231978 5358
rect 232062 5122 232298 5358
rect 232382 5122 232618 5358
rect 233862 228682 234098 228918
rect 234182 228682 234418 228918
rect 234502 228682 234738 228918
rect 234822 228682 235058 228918
rect 235142 228682 235378 228918
rect 235462 228682 235698 228918
rect 235782 228682 236018 228918
rect 236102 228682 236338 228918
rect 236422 228682 236658 228918
rect 236742 228682 236978 228918
rect 237062 228682 237298 228918
rect 237382 228682 237618 228918
rect 233862 206282 234098 206518
rect 234182 206282 234418 206518
rect 234502 206282 234738 206518
rect 234822 206282 235058 206518
rect 235142 206282 235378 206518
rect 235462 206282 235698 206518
rect 235782 206282 236018 206518
rect 236102 206282 236338 206518
rect 236422 206282 236658 206518
rect 236742 206282 236978 206518
rect 237062 206282 237298 206518
rect 237382 206282 237618 206518
rect 233862 183882 234098 184118
rect 234182 183882 234418 184118
rect 234502 183882 234738 184118
rect 234822 183882 235058 184118
rect 235142 183882 235378 184118
rect 235462 183882 235698 184118
rect 235782 183882 236018 184118
rect 236102 183882 236338 184118
rect 236422 183882 236658 184118
rect 236742 183882 236978 184118
rect 237062 183882 237298 184118
rect 237382 183882 237618 184118
rect 233862 161482 234098 161718
rect 234182 161482 234418 161718
rect 234502 161482 234738 161718
rect 234822 161482 235058 161718
rect 235142 161482 235378 161718
rect 235462 161482 235698 161718
rect 235782 161482 236018 161718
rect 236102 161482 236338 161718
rect 236422 161482 236658 161718
rect 236742 161482 236978 161718
rect 237062 161482 237298 161718
rect 237382 161482 237618 161718
rect 233862 139082 234098 139318
rect 234182 139082 234418 139318
rect 234502 139082 234738 139318
rect 234822 139082 235058 139318
rect 235142 139082 235378 139318
rect 235462 139082 235698 139318
rect 235782 139082 236018 139318
rect 236102 139082 236338 139318
rect 236422 139082 236658 139318
rect 236742 139082 236978 139318
rect 237062 139082 237298 139318
rect 237382 139082 237618 139318
rect 233862 116682 234098 116918
rect 234182 116682 234418 116918
rect 234502 116682 234738 116918
rect 234822 116682 235058 116918
rect 235142 116682 235378 116918
rect 235462 116682 235698 116918
rect 235782 116682 236018 116918
rect 236102 116682 236338 116918
rect 236422 116682 236658 116918
rect 236742 116682 236978 116918
rect 237062 116682 237298 116918
rect 237382 116682 237618 116918
rect 233862 94282 234098 94518
rect 234182 94282 234418 94518
rect 234502 94282 234738 94518
rect 234822 94282 235058 94518
rect 235142 94282 235378 94518
rect 235462 94282 235698 94518
rect 235782 94282 236018 94518
rect 236102 94282 236338 94518
rect 236422 94282 236658 94518
rect 236742 94282 236978 94518
rect 237062 94282 237298 94518
rect 237382 94282 237618 94518
rect 233862 71882 234098 72118
rect 234182 71882 234418 72118
rect 234502 71882 234738 72118
rect 234822 71882 235058 72118
rect 235142 71882 235378 72118
rect 235462 71882 235698 72118
rect 235782 71882 236018 72118
rect 236102 71882 236338 72118
rect 236422 71882 236658 72118
rect 236742 71882 236978 72118
rect 237062 71882 237298 72118
rect 237382 71882 237618 72118
rect 233862 49482 234098 49718
rect 234182 49482 234418 49718
rect 234502 49482 234738 49718
rect 234822 49482 235058 49718
rect 235142 49482 235378 49718
rect 235462 49482 235698 49718
rect 235782 49482 236018 49718
rect 236102 49482 236338 49718
rect 236422 49482 236658 49718
rect 236742 49482 236978 49718
rect 237062 49482 237298 49718
rect 237382 49482 237618 49718
rect 233862 27082 234098 27318
rect 234182 27082 234418 27318
rect 234502 27082 234738 27318
rect 234822 27082 235058 27318
rect 235142 27082 235378 27318
rect 235462 27082 235698 27318
rect 235782 27082 236018 27318
rect 236102 27082 236338 27318
rect 236422 27082 236658 27318
rect 236742 27082 236978 27318
rect 237062 27082 237298 27318
rect 237382 27082 237618 27318
rect 122 3642 358 3878
rect 442 3642 678 3878
rect 762 3642 998 3878
rect 1082 3642 1318 3878
rect 1402 3642 1638 3878
rect 1722 3642 1958 3878
rect 2042 3642 2278 3878
rect 2362 3642 2598 3878
rect 2682 3642 2918 3878
rect 3002 3642 3238 3878
rect 3322 3642 3558 3878
rect 3642 3642 3878 3878
rect 122 3322 358 3558
rect 442 3322 678 3558
rect 762 3322 998 3558
rect 1082 3322 1318 3558
rect 1402 3322 1638 3558
rect 1722 3322 1958 3558
rect 2042 3322 2278 3558
rect 2362 3322 2598 3558
rect 2682 3322 2918 3558
rect 3002 3322 3238 3558
rect 3322 3322 3558 3558
rect 3642 3322 3878 3558
rect 122 3002 358 3238
rect 442 3002 678 3238
rect 762 3002 998 3238
rect 1082 3002 1318 3238
rect 1402 3002 1638 3238
rect 1722 3002 1958 3238
rect 2042 3002 2278 3238
rect 2362 3002 2598 3238
rect 2682 3002 2918 3238
rect 3002 3002 3238 3238
rect 3322 3002 3558 3238
rect 3642 3002 3878 3238
rect 122 2682 358 2918
rect 442 2682 678 2918
rect 762 2682 998 2918
rect 1082 2682 1318 2918
rect 1402 2682 1638 2918
rect 1722 2682 1958 2918
rect 2042 2682 2278 2918
rect 2362 2682 2598 2918
rect 2682 2682 2918 2918
rect 3002 2682 3238 2918
rect 3322 2682 3558 2918
rect 3642 2682 3878 2918
rect 122 2362 358 2598
rect 442 2362 678 2598
rect 762 2362 998 2598
rect 1082 2362 1318 2598
rect 1402 2362 1638 2598
rect 1722 2362 1958 2598
rect 2042 2362 2278 2598
rect 2362 2362 2598 2598
rect 2682 2362 2918 2598
rect 3002 2362 3238 2598
rect 3322 2362 3558 2598
rect 3642 2362 3878 2598
rect 122 2042 358 2278
rect 442 2042 678 2278
rect 762 2042 998 2278
rect 1082 2042 1318 2278
rect 1402 2042 1638 2278
rect 1722 2042 1958 2278
rect 2042 2042 2278 2278
rect 2362 2042 2598 2278
rect 2682 2042 2918 2278
rect 3002 2042 3238 2278
rect 3322 2042 3558 2278
rect 3642 2042 3878 2278
rect 122 1722 358 1958
rect 442 1722 678 1958
rect 762 1722 998 1958
rect 1082 1722 1318 1958
rect 1402 1722 1638 1958
rect 1722 1722 1958 1958
rect 2042 1722 2278 1958
rect 2362 1722 2598 1958
rect 2682 1722 2918 1958
rect 3002 1722 3238 1958
rect 3322 1722 3558 1958
rect 3642 1722 3878 1958
rect 122 1402 358 1638
rect 442 1402 678 1638
rect 762 1402 998 1638
rect 1082 1402 1318 1638
rect 1402 1402 1638 1638
rect 1722 1402 1958 1638
rect 2042 1402 2278 1638
rect 2362 1402 2598 1638
rect 2682 1402 2918 1638
rect 3002 1402 3238 1638
rect 3322 1402 3558 1638
rect 3642 1402 3878 1638
rect 122 1082 358 1318
rect 442 1082 678 1318
rect 762 1082 998 1318
rect 1082 1082 1318 1318
rect 1402 1082 1638 1318
rect 1722 1082 1958 1318
rect 2042 1082 2278 1318
rect 2362 1082 2598 1318
rect 2682 1082 2918 1318
rect 3002 1082 3238 1318
rect 3322 1082 3558 1318
rect 3642 1082 3878 1318
rect 122 762 358 998
rect 442 762 678 998
rect 762 762 998 998
rect 1082 762 1318 998
rect 1402 762 1638 998
rect 1722 762 1958 998
rect 2042 762 2278 998
rect 2362 762 2598 998
rect 2682 762 2918 998
rect 3002 762 3238 998
rect 3322 762 3558 998
rect 3642 762 3878 998
rect 122 442 358 678
rect 442 442 678 678
rect 762 442 998 678
rect 1082 442 1318 678
rect 1402 442 1638 678
rect 1722 442 1958 678
rect 2042 442 2278 678
rect 2362 442 2598 678
rect 2682 442 2918 678
rect 3002 442 3238 678
rect 3322 442 3558 678
rect 3642 442 3878 678
rect 122 122 358 358
rect 442 122 678 358
rect 762 122 998 358
rect 1082 122 1318 358
rect 1402 122 1638 358
rect 1722 122 1958 358
rect 2042 122 2278 358
rect 2362 122 2598 358
rect 2682 122 2918 358
rect 3002 122 3238 358
rect 3322 122 3558 358
rect 3642 122 3878 358
rect 233862 3642 234098 3878
rect 234182 3642 234418 3878
rect 234502 3642 234738 3878
rect 234822 3642 235058 3878
rect 235142 3642 235378 3878
rect 235462 3642 235698 3878
rect 235782 3642 236018 3878
rect 236102 3642 236338 3878
rect 236422 3642 236658 3878
rect 236742 3642 236978 3878
rect 237062 3642 237298 3878
rect 237382 3642 237618 3878
rect 233862 3322 234098 3558
rect 234182 3322 234418 3558
rect 234502 3322 234738 3558
rect 234822 3322 235058 3558
rect 235142 3322 235378 3558
rect 235462 3322 235698 3558
rect 235782 3322 236018 3558
rect 236102 3322 236338 3558
rect 236422 3322 236658 3558
rect 236742 3322 236978 3558
rect 237062 3322 237298 3558
rect 237382 3322 237618 3558
rect 233862 3002 234098 3238
rect 234182 3002 234418 3238
rect 234502 3002 234738 3238
rect 234822 3002 235058 3238
rect 235142 3002 235378 3238
rect 235462 3002 235698 3238
rect 235782 3002 236018 3238
rect 236102 3002 236338 3238
rect 236422 3002 236658 3238
rect 236742 3002 236978 3238
rect 237062 3002 237298 3238
rect 237382 3002 237618 3238
rect 233862 2682 234098 2918
rect 234182 2682 234418 2918
rect 234502 2682 234738 2918
rect 234822 2682 235058 2918
rect 235142 2682 235378 2918
rect 235462 2682 235698 2918
rect 235782 2682 236018 2918
rect 236102 2682 236338 2918
rect 236422 2682 236658 2918
rect 236742 2682 236978 2918
rect 237062 2682 237298 2918
rect 237382 2682 237618 2918
rect 233862 2362 234098 2598
rect 234182 2362 234418 2598
rect 234502 2362 234738 2598
rect 234822 2362 235058 2598
rect 235142 2362 235378 2598
rect 235462 2362 235698 2598
rect 235782 2362 236018 2598
rect 236102 2362 236338 2598
rect 236422 2362 236658 2598
rect 236742 2362 236978 2598
rect 237062 2362 237298 2598
rect 237382 2362 237618 2598
rect 233862 2042 234098 2278
rect 234182 2042 234418 2278
rect 234502 2042 234738 2278
rect 234822 2042 235058 2278
rect 235142 2042 235378 2278
rect 235462 2042 235698 2278
rect 235782 2042 236018 2278
rect 236102 2042 236338 2278
rect 236422 2042 236658 2278
rect 236742 2042 236978 2278
rect 237062 2042 237298 2278
rect 237382 2042 237618 2278
rect 233862 1722 234098 1958
rect 234182 1722 234418 1958
rect 234502 1722 234738 1958
rect 234822 1722 235058 1958
rect 235142 1722 235378 1958
rect 235462 1722 235698 1958
rect 235782 1722 236018 1958
rect 236102 1722 236338 1958
rect 236422 1722 236658 1958
rect 236742 1722 236978 1958
rect 237062 1722 237298 1958
rect 237382 1722 237618 1958
rect 233862 1402 234098 1638
rect 234182 1402 234418 1638
rect 234502 1402 234738 1638
rect 234822 1402 235058 1638
rect 235142 1402 235378 1638
rect 235462 1402 235698 1638
rect 235782 1402 236018 1638
rect 236102 1402 236338 1638
rect 236422 1402 236658 1638
rect 236742 1402 236978 1638
rect 237062 1402 237298 1638
rect 237382 1402 237618 1638
rect 233862 1082 234098 1318
rect 234182 1082 234418 1318
rect 234502 1082 234738 1318
rect 234822 1082 235058 1318
rect 235142 1082 235378 1318
rect 235462 1082 235698 1318
rect 235782 1082 236018 1318
rect 236102 1082 236338 1318
rect 236422 1082 236658 1318
rect 236742 1082 236978 1318
rect 237062 1082 237298 1318
rect 237382 1082 237618 1318
rect 233862 762 234098 998
rect 234182 762 234418 998
rect 234502 762 234738 998
rect 234822 762 235058 998
rect 235142 762 235378 998
rect 235462 762 235698 998
rect 235782 762 236018 998
rect 236102 762 236338 998
rect 236422 762 236658 998
rect 236742 762 236978 998
rect 237062 762 237298 998
rect 237382 762 237618 998
rect 233862 442 234098 678
rect 234182 442 234418 678
rect 234502 442 234738 678
rect 234822 442 235058 678
rect 235142 442 235378 678
rect 235462 442 235698 678
rect 235782 442 236018 678
rect 236102 442 236338 678
rect 236422 442 236658 678
rect 236742 442 236978 678
rect 237062 442 237298 678
rect 237382 442 237618 678
rect 233862 122 234098 358
rect 234182 122 234418 358
rect 234502 122 234738 358
rect 234822 122 235058 358
rect 235142 122 235378 358
rect 235462 122 235698 358
rect 235782 122 236018 358
rect 236102 122 236338 358
rect 236422 122 236658 358
rect 236742 122 236978 358
rect 237062 122 237298 358
rect 237382 122 237618 358
<< metal5 >>
rect 0 255254 237740 255376
rect 0 255018 122 255254
rect 358 255018 442 255254
rect 678 255018 762 255254
rect 998 255018 1082 255254
rect 1318 255018 1402 255254
rect 1638 255018 1722 255254
rect 1958 255018 2042 255254
rect 2278 255018 2362 255254
rect 2598 255018 2682 255254
rect 2918 255018 3002 255254
rect 3238 255018 3322 255254
rect 3558 255018 3642 255254
rect 3878 255018 233862 255254
rect 234098 255018 234182 255254
rect 234418 255018 234502 255254
rect 234738 255018 234822 255254
rect 235058 255018 235142 255254
rect 235378 255018 235462 255254
rect 235698 255018 235782 255254
rect 236018 255018 236102 255254
rect 236338 255018 236422 255254
rect 236658 255018 236742 255254
rect 236978 255018 237062 255254
rect 237298 255018 237382 255254
rect 237618 255018 237740 255254
rect 0 254934 237740 255018
rect 0 254698 122 254934
rect 358 254698 442 254934
rect 678 254698 762 254934
rect 998 254698 1082 254934
rect 1318 254698 1402 254934
rect 1638 254698 1722 254934
rect 1958 254698 2042 254934
rect 2278 254698 2362 254934
rect 2598 254698 2682 254934
rect 2918 254698 3002 254934
rect 3238 254698 3322 254934
rect 3558 254698 3642 254934
rect 3878 254698 233862 254934
rect 234098 254698 234182 254934
rect 234418 254698 234502 254934
rect 234738 254698 234822 254934
rect 235058 254698 235142 254934
rect 235378 254698 235462 254934
rect 235698 254698 235782 254934
rect 236018 254698 236102 254934
rect 236338 254698 236422 254934
rect 236658 254698 236742 254934
rect 236978 254698 237062 254934
rect 237298 254698 237382 254934
rect 237618 254698 237740 254934
rect 0 254614 237740 254698
rect 0 254378 122 254614
rect 358 254378 442 254614
rect 678 254378 762 254614
rect 998 254378 1082 254614
rect 1318 254378 1402 254614
rect 1638 254378 1722 254614
rect 1958 254378 2042 254614
rect 2278 254378 2362 254614
rect 2598 254378 2682 254614
rect 2918 254378 3002 254614
rect 3238 254378 3322 254614
rect 3558 254378 3642 254614
rect 3878 254378 233862 254614
rect 234098 254378 234182 254614
rect 234418 254378 234502 254614
rect 234738 254378 234822 254614
rect 235058 254378 235142 254614
rect 235378 254378 235462 254614
rect 235698 254378 235782 254614
rect 236018 254378 236102 254614
rect 236338 254378 236422 254614
rect 236658 254378 236742 254614
rect 236978 254378 237062 254614
rect 237298 254378 237382 254614
rect 237618 254378 237740 254614
rect 0 254294 237740 254378
rect 0 254058 122 254294
rect 358 254058 442 254294
rect 678 254058 762 254294
rect 998 254058 1082 254294
rect 1318 254058 1402 254294
rect 1638 254058 1722 254294
rect 1958 254058 2042 254294
rect 2278 254058 2362 254294
rect 2598 254058 2682 254294
rect 2918 254058 3002 254294
rect 3238 254058 3322 254294
rect 3558 254058 3642 254294
rect 3878 254058 233862 254294
rect 234098 254058 234182 254294
rect 234418 254058 234502 254294
rect 234738 254058 234822 254294
rect 235058 254058 235142 254294
rect 235378 254058 235462 254294
rect 235698 254058 235782 254294
rect 236018 254058 236102 254294
rect 236338 254058 236422 254294
rect 236658 254058 236742 254294
rect 236978 254058 237062 254294
rect 237298 254058 237382 254294
rect 237618 254058 237740 254294
rect 0 253974 237740 254058
rect 0 253738 122 253974
rect 358 253738 442 253974
rect 678 253738 762 253974
rect 998 253738 1082 253974
rect 1318 253738 1402 253974
rect 1638 253738 1722 253974
rect 1958 253738 2042 253974
rect 2278 253738 2362 253974
rect 2598 253738 2682 253974
rect 2918 253738 3002 253974
rect 3238 253738 3322 253974
rect 3558 253738 3642 253974
rect 3878 253738 233862 253974
rect 234098 253738 234182 253974
rect 234418 253738 234502 253974
rect 234738 253738 234822 253974
rect 235058 253738 235142 253974
rect 235378 253738 235462 253974
rect 235698 253738 235782 253974
rect 236018 253738 236102 253974
rect 236338 253738 236422 253974
rect 236658 253738 236742 253974
rect 236978 253738 237062 253974
rect 237298 253738 237382 253974
rect 237618 253738 237740 253974
rect 0 253654 237740 253738
rect 0 253418 122 253654
rect 358 253418 442 253654
rect 678 253418 762 253654
rect 998 253418 1082 253654
rect 1318 253418 1402 253654
rect 1638 253418 1722 253654
rect 1958 253418 2042 253654
rect 2278 253418 2362 253654
rect 2598 253418 2682 253654
rect 2918 253418 3002 253654
rect 3238 253418 3322 253654
rect 3558 253418 3642 253654
rect 3878 253418 233862 253654
rect 234098 253418 234182 253654
rect 234418 253418 234502 253654
rect 234738 253418 234822 253654
rect 235058 253418 235142 253654
rect 235378 253418 235462 253654
rect 235698 253418 235782 253654
rect 236018 253418 236102 253654
rect 236338 253418 236422 253654
rect 236658 253418 236742 253654
rect 236978 253418 237062 253654
rect 237298 253418 237382 253654
rect 237618 253418 237740 253654
rect 0 253334 237740 253418
rect 0 253098 122 253334
rect 358 253098 442 253334
rect 678 253098 762 253334
rect 998 253098 1082 253334
rect 1318 253098 1402 253334
rect 1638 253098 1722 253334
rect 1958 253098 2042 253334
rect 2278 253098 2362 253334
rect 2598 253098 2682 253334
rect 2918 253098 3002 253334
rect 3238 253098 3322 253334
rect 3558 253098 3642 253334
rect 3878 253098 233862 253334
rect 234098 253098 234182 253334
rect 234418 253098 234502 253334
rect 234738 253098 234822 253334
rect 235058 253098 235142 253334
rect 235378 253098 235462 253334
rect 235698 253098 235782 253334
rect 236018 253098 236102 253334
rect 236338 253098 236422 253334
rect 236658 253098 236742 253334
rect 236978 253098 237062 253334
rect 237298 253098 237382 253334
rect 237618 253098 237740 253334
rect 0 253014 237740 253098
rect 0 252778 122 253014
rect 358 252778 442 253014
rect 678 252778 762 253014
rect 998 252778 1082 253014
rect 1318 252778 1402 253014
rect 1638 252778 1722 253014
rect 1958 252778 2042 253014
rect 2278 252778 2362 253014
rect 2598 252778 2682 253014
rect 2918 252778 3002 253014
rect 3238 252778 3322 253014
rect 3558 252778 3642 253014
rect 3878 252778 233862 253014
rect 234098 252778 234182 253014
rect 234418 252778 234502 253014
rect 234738 252778 234822 253014
rect 235058 252778 235142 253014
rect 235378 252778 235462 253014
rect 235698 252778 235782 253014
rect 236018 252778 236102 253014
rect 236338 252778 236422 253014
rect 236658 252778 236742 253014
rect 236978 252778 237062 253014
rect 237298 252778 237382 253014
rect 237618 252778 237740 253014
rect 0 252694 237740 252778
rect 0 252458 122 252694
rect 358 252458 442 252694
rect 678 252458 762 252694
rect 998 252458 1082 252694
rect 1318 252458 1402 252694
rect 1638 252458 1722 252694
rect 1958 252458 2042 252694
rect 2278 252458 2362 252694
rect 2598 252458 2682 252694
rect 2918 252458 3002 252694
rect 3238 252458 3322 252694
rect 3558 252458 3642 252694
rect 3878 252458 233862 252694
rect 234098 252458 234182 252694
rect 234418 252458 234502 252694
rect 234738 252458 234822 252694
rect 235058 252458 235142 252694
rect 235378 252458 235462 252694
rect 235698 252458 235782 252694
rect 236018 252458 236102 252694
rect 236338 252458 236422 252694
rect 236658 252458 236742 252694
rect 236978 252458 237062 252694
rect 237298 252458 237382 252694
rect 237618 252458 237740 252694
rect 0 252374 237740 252458
rect 0 252138 122 252374
rect 358 252138 442 252374
rect 678 252138 762 252374
rect 998 252138 1082 252374
rect 1318 252138 1402 252374
rect 1638 252138 1722 252374
rect 1958 252138 2042 252374
rect 2278 252138 2362 252374
rect 2598 252138 2682 252374
rect 2918 252138 3002 252374
rect 3238 252138 3322 252374
rect 3558 252138 3642 252374
rect 3878 252138 233862 252374
rect 234098 252138 234182 252374
rect 234418 252138 234502 252374
rect 234738 252138 234822 252374
rect 235058 252138 235142 252374
rect 235378 252138 235462 252374
rect 235698 252138 235782 252374
rect 236018 252138 236102 252374
rect 236338 252138 236422 252374
rect 236658 252138 236742 252374
rect 236978 252138 237062 252374
rect 237298 252138 237382 252374
rect 237618 252138 237740 252374
rect 0 252054 237740 252138
rect 0 251818 122 252054
rect 358 251818 442 252054
rect 678 251818 762 252054
rect 998 251818 1082 252054
rect 1318 251818 1402 252054
rect 1638 251818 1722 252054
rect 1958 251818 2042 252054
rect 2278 251818 2362 252054
rect 2598 251818 2682 252054
rect 2918 251818 3002 252054
rect 3238 251818 3322 252054
rect 3558 251818 3642 252054
rect 3878 251818 233862 252054
rect 234098 251818 234182 252054
rect 234418 251818 234502 252054
rect 234738 251818 234822 252054
rect 235058 251818 235142 252054
rect 235378 251818 235462 252054
rect 235698 251818 235782 252054
rect 236018 251818 236102 252054
rect 236338 251818 236422 252054
rect 236658 251818 236742 252054
rect 236978 251818 237062 252054
rect 237298 251818 237382 252054
rect 237618 251818 237740 252054
rect 0 251734 237740 251818
rect 0 251498 122 251734
rect 358 251498 442 251734
rect 678 251498 762 251734
rect 998 251498 1082 251734
rect 1318 251498 1402 251734
rect 1638 251498 1722 251734
rect 1958 251498 2042 251734
rect 2278 251498 2362 251734
rect 2598 251498 2682 251734
rect 2918 251498 3002 251734
rect 3238 251498 3322 251734
rect 3558 251498 3642 251734
rect 3878 251498 233862 251734
rect 234098 251498 234182 251734
rect 234418 251498 234502 251734
rect 234738 251498 234822 251734
rect 235058 251498 235142 251734
rect 235378 251498 235462 251734
rect 235698 251498 235782 251734
rect 236018 251498 236102 251734
rect 236338 251498 236422 251734
rect 236658 251498 236742 251734
rect 236978 251498 237062 251734
rect 237298 251498 237382 251734
rect 237618 251498 237740 251734
rect 0 251376 237740 251498
rect 5000 250254 232740 250376
rect 5000 250018 5122 250254
rect 5358 250018 5442 250254
rect 5678 250018 5762 250254
rect 5998 250018 6082 250254
rect 6318 250018 6402 250254
rect 6638 250018 6722 250254
rect 6958 250018 7042 250254
rect 7278 250018 7362 250254
rect 7598 250018 7682 250254
rect 7918 250018 8002 250254
rect 8238 250018 8322 250254
rect 8558 250018 8642 250254
rect 8878 250018 228862 250254
rect 229098 250018 229182 250254
rect 229418 250018 229502 250254
rect 229738 250018 229822 250254
rect 230058 250018 230142 250254
rect 230378 250018 230462 250254
rect 230698 250018 230782 250254
rect 231018 250018 231102 250254
rect 231338 250018 231422 250254
rect 231658 250018 231742 250254
rect 231978 250018 232062 250254
rect 232298 250018 232382 250254
rect 232618 250018 232740 250254
rect 5000 249934 232740 250018
rect 5000 249698 5122 249934
rect 5358 249698 5442 249934
rect 5678 249698 5762 249934
rect 5998 249698 6082 249934
rect 6318 249698 6402 249934
rect 6638 249698 6722 249934
rect 6958 249698 7042 249934
rect 7278 249698 7362 249934
rect 7598 249698 7682 249934
rect 7918 249698 8002 249934
rect 8238 249698 8322 249934
rect 8558 249698 8642 249934
rect 8878 249698 228862 249934
rect 229098 249698 229182 249934
rect 229418 249698 229502 249934
rect 229738 249698 229822 249934
rect 230058 249698 230142 249934
rect 230378 249698 230462 249934
rect 230698 249698 230782 249934
rect 231018 249698 231102 249934
rect 231338 249698 231422 249934
rect 231658 249698 231742 249934
rect 231978 249698 232062 249934
rect 232298 249698 232382 249934
rect 232618 249698 232740 249934
rect 5000 249614 232740 249698
rect 5000 249378 5122 249614
rect 5358 249378 5442 249614
rect 5678 249378 5762 249614
rect 5998 249378 6082 249614
rect 6318 249378 6402 249614
rect 6638 249378 6722 249614
rect 6958 249378 7042 249614
rect 7278 249378 7362 249614
rect 7598 249378 7682 249614
rect 7918 249378 8002 249614
rect 8238 249378 8322 249614
rect 8558 249378 8642 249614
rect 8878 249378 228862 249614
rect 229098 249378 229182 249614
rect 229418 249378 229502 249614
rect 229738 249378 229822 249614
rect 230058 249378 230142 249614
rect 230378 249378 230462 249614
rect 230698 249378 230782 249614
rect 231018 249378 231102 249614
rect 231338 249378 231422 249614
rect 231658 249378 231742 249614
rect 231978 249378 232062 249614
rect 232298 249378 232382 249614
rect 232618 249378 232740 249614
rect 5000 249294 232740 249378
rect 5000 249058 5122 249294
rect 5358 249058 5442 249294
rect 5678 249058 5762 249294
rect 5998 249058 6082 249294
rect 6318 249058 6402 249294
rect 6638 249058 6722 249294
rect 6958 249058 7042 249294
rect 7278 249058 7362 249294
rect 7598 249058 7682 249294
rect 7918 249058 8002 249294
rect 8238 249058 8322 249294
rect 8558 249058 8642 249294
rect 8878 249058 228862 249294
rect 229098 249058 229182 249294
rect 229418 249058 229502 249294
rect 229738 249058 229822 249294
rect 230058 249058 230142 249294
rect 230378 249058 230462 249294
rect 230698 249058 230782 249294
rect 231018 249058 231102 249294
rect 231338 249058 231422 249294
rect 231658 249058 231742 249294
rect 231978 249058 232062 249294
rect 232298 249058 232382 249294
rect 232618 249058 232740 249294
rect 5000 248974 232740 249058
rect 5000 248738 5122 248974
rect 5358 248738 5442 248974
rect 5678 248738 5762 248974
rect 5998 248738 6082 248974
rect 6318 248738 6402 248974
rect 6638 248738 6722 248974
rect 6958 248738 7042 248974
rect 7278 248738 7362 248974
rect 7598 248738 7682 248974
rect 7918 248738 8002 248974
rect 8238 248738 8322 248974
rect 8558 248738 8642 248974
rect 8878 248738 228862 248974
rect 229098 248738 229182 248974
rect 229418 248738 229502 248974
rect 229738 248738 229822 248974
rect 230058 248738 230142 248974
rect 230378 248738 230462 248974
rect 230698 248738 230782 248974
rect 231018 248738 231102 248974
rect 231338 248738 231422 248974
rect 231658 248738 231742 248974
rect 231978 248738 232062 248974
rect 232298 248738 232382 248974
rect 232618 248738 232740 248974
rect 5000 248654 232740 248738
rect 5000 248418 5122 248654
rect 5358 248418 5442 248654
rect 5678 248418 5762 248654
rect 5998 248418 6082 248654
rect 6318 248418 6402 248654
rect 6638 248418 6722 248654
rect 6958 248418 7042 248654
rect 7278 248418 7362 248654
rect 7598 248418 7682 248654
rect 7918 248418 8002 248654
rect 8238 248418 8322 248654
rect 8558 248418 8642 248654
rect 8878 248418 228862 248654
rect 229098 248418 229182 248654
rect 229418 248418 229502 248654
rect 229738 248418 229822 248654
rect 230058 248418 230142 248654
rect 230378 248418 230462 248654
rect 230698 248418 230782 248654
rect 231018 248418 231102 248654
rect 231338 248418 231422 248654
rect 231658 248418 231742 248654
rect 231978 248418 232062 248654
rect 232298 248418 232382 248654
rect 232618 248418 232740 248654
rect 5000 248334 232740 248418
rect 5000 248098 5122 248334
rect 5358 248098 5442 248334
rect 5678 248098 5762 248334
rect 5998 248098 6082 248334
rect 6318 248098 6402 248334
rect 6638 248098 6722 248334
rect 6958 248098 7042 248334
rect 7278 248098 7362 248334
rect 7598 248098 7682 248334
rect 7918 248098 8002 248334
rect 8238 248098 8322 248334
rect 8558 248098 8642 248334
rect 8878 248098 228862 248334
rect 229098 248098 229182 248334
rect 229418 248098 229502 248334
rect 229738 248098 229822 248334
rect 230058 248098 230142 248334
rect 230378 248098 230462 248334
rect 230698 248098 230782 248334
rect 231018 248098 231102 248334
rect 231338 248098 231422 248334
rect 231658 248098 231742 248334
rect 231978 248098 232062 248334
rect 232298 248098 232382 248334
rect 232618 248098 232740 248334
rect 5000 248014 232740 248098
rect 5000 247778 5122 248014
rect 5358 247778 5442 248014
rect 5678 247778 5762 248014
rect 5998 247778 6082 248014
rect 6318 247778 6402 248014
rect 6638 247778 6722 248014
rect 6958 247778 7042 248014
rect 7278 247778 7362 248014
rect 7598 247778 7682 248014
rect 7918 247778 8002 248014
rect 8238 247778 8322 248014
rect 8558 247778 8642 248014
rect 8878 247778 228862 248014
rect 229098 247778 229182 248014
rect 229418 247778 229502 248014
rect 229738 247778 229822 248014
rect 230058 247778 230142 248014
rect 230378 247778 230462 248014
rect 230698 247778 230782 248014
rect 231018 247778 231102 248014
rect 231338 247778 231422 248014
rect 231658 247778 231742 248014
rect 231978 247778 232062 248014
rect 232298 247778 232382 248014
rect 232618 247778 232740 248014
rect 5000 247694 232740 247778
rect 5000 247458 5122 247694
rect 5358 247458 5442 247694
rect 5678 247458 5762 247694
rect 5998 247458 6082 247694
rect 6318 247458 6402 247694
rect 6638 247458 6722 247694
rect 6958 247458 7042 247694
rect 7278 247458 7362 247694
rect 7598 247458 7682 247694
rect 7918 247458 8002 247694
rect 8238 247458 8322 247694
rect 8558 247458 8642 247694
rect 8878 247458 228862 247694
rect 229098 247458 229182 247694
rect 229418 247458 229502 247694
rect 229738 247458 229822 247694
rect 230058 247458 230142 247694
rect 230378 247458 230462 247694
rect 230698 247458 230782 247694
rect 231018 247458 231102 247694
rect 231338 247458 231422 247694
rect 231658 247458 231742 247694
rect 231978 247458 232062 247694
rect 232298 247458 232382 247694
rect 232618 247458 232740 247694
rect 5000 247374 232740 247458
rect 5000 247138 5122 247374
rect 5358 247138 5442 247374
rect 5678 247138 5762 247374
rect 5998 247138 6082 247374
rect 6318 247138 6402 247374
rect 6638 247138 6722 247374
rect 6958 247138 7042 247374
rect 7278 247138 7362 247374
rect 7598 247138 7682 247374
rect 7918 247138 8002 247374
rect 8238 247138 8322 247374
rect 8558 247138 8642 247374
rect 8878 247138 228862 247374
rect 229098 247138 229182 247374
rect 229418 247138 229502 247374
rect 229738 247138 229822 247374
rect 230058 247138 230142 247374
rect 230378 247138 230462 247374
rect 230698 247138 230782 247374
rect 231018 247138 231102 247374
rect 231338 247138 231422 247374
rect 231658 247138 231742 247374
rect 231978 247138 232062 247374
rect 232298 247138 232382 247374
rect 232618 247138 232740 247374
rect 5000 247054 232740 247138
rect 5000 246818 5122 247054
rect 5358 246818 5442 247054
rect 5678 246818 5762 247054
rect 5998 246818 6082 247054
rect 6318 246818 6402 247054
rect 6638 246818 6722 247054
rect 6958 246818 7042 247054
rect 7278 246818 7362 247054
rect 7598 246818 7682 247054
rect 7918 246818 8002 247054
rect 8238 246818 8322 247054
rect 8558 246818 8642 247054
rect 8878 246818 228862 247054
rect 229098 246818 229182 247054
rect 229418 246818 229502 247054
rect 229738 246818 229822 247054
rect 230058 246818 230142 247054
rect 230378 246818 230462 247054
rect 230698 246818 230782 247054
rect 231018 246818 231102 247054
rect 231338 246818 231422 247054
rect 231658 246818 231742 247054
rect 231978 246818 232062 247054
rect 232298 246818 232382 247054
rect 232618 246818 232740 247054
rect 5000 246734 232740 246818
rect 5000 246498 5122 246734
rect 5358 246498 5442 246734
rect 5678 246498 5762 246734
rect 5998 246498 6082 246734
rect 6318 246498 6402 246734
rect 6638 246498 6722 246734
rect 6958 246498 7042 246734
rect 7278 246498 7362 246734
rect 7598 246498 7682 246734
rect 7918 246498 8002 246734
rect 8238 246498 8322 246734
rect 8558 246498 8642 246734
rect 8878 246498 228862 246734
rect 229098 246498 229182 246734
rect 229418 246498 229502 246734
rect 229738 246498 229822 246734
rect 230058 246498 230142 246734
rect 230378 246498 230462 246734
rect 230698 246498 230782 246734
rect 231018 246498 231102 246734
rect 231338 246498 231422 246734
rect 231658 246498 231742 246734
rect 231978 246498 232062 246734
rect 232298 246498 232382 246734
rect 232618 246498 232740 246734
rect 5000 246376 232740 246498
rect 0 240118 237740 240160
rect 0 239882 5122 240118
rect 5358 239882 5442 240118
rect 5678 239882 5762 240118
rect 5998 239882 6082 240118
rect 6318 239882 6402 240118
rect 6638 239882 6722 240118
rect 6958 239882 7042 240118
rect 7278 239882 7362 240118
rect 7598 239882 7682 240118
rect 7918 239882 8002 240118
rect 8238 239882 8322 240118
rect 8558 239882 8642 240118
rect 8878 239882 72816 240118
rect 73052 239882 144816 240118
rect 145052 239882 228862 240118
rect 229098 239882 229182 240118
rect 229418 239882 229502 240118
rect 229738 239882 229822 240118
rect 230058 239882 230142 240118
rect 230378 239882 230462 240118
rect 230698 239882 230782 240118
rect 231018 239882 231102 240118
rect 231338 239882 231422 240118
rect 231658 239882 231742 240118
rect 231978 239882 232062 240118
rect 232298 239882 232382 240118
rect 232618 239882 237740 240118
rect 0 239840 237740 239882
rect 0 228918 237740 228960
rect 0 228682 122 228918
rect 358 228682 442 228918
rect 678 228682 762 228918
rect 998 228682 1082 228918
rect 1318 228682 1402 228918
rect 1638 228682 1722 228918
rect 1958 228682 2042 228918
rect 2278 228682 2362 228918
rect 2598 228682 2682 228918
rect 2918 228682 3002 228918
rect 3238 228682 3322 228918
rect 3558 228682 3642 228918
rect 3878 228682 77816 228918
rect 78052 228682 149816 228918
rect 150052 228682 233862 228918
rect 234098 228682 234182 228918
rect 234418 228682 234502 228918
rect 234738 228682 234822 228918
rect 235058 228682 235142 228918
rect 235378 228682 235462 228918
rect 235698 228682 235782 228918
rect 236018 228682 236102 228918
rect 236338 228682 236422 228918
rect 236658 228682 236742 228918
rect 236978 228682 237062 228918
rect 237298 228682 237382 228918
rect 237618 228682 237740 228918
rect 0 228640 237740 228682
rect 0 217718 237740 217760
rect 0 217482 5122 217718
rect 5358 217482 5442 217718
rect 5678 217482 5762 217718
rect 5998 217482 6082 217718
rect 6318 217482 6402 217718
rect 6638 217482 6722 217718
rect 6958 217482 7042 217718
rect 7278 217482 7362 217718
rect 7598 217482 7682 217718
rect 7918 217482 8002 217718
rect 8238 217482 8322 217718
rect 8558 217482 8642 217718
rect 8878 217482 228862 217718
rect 229098 217482 229182 217718
rect 229418 217482 229502 217718
rect 229738 217482 229822 217718
rect 230058 217482 230142 217718
rect 230378 217482 230462 217718
rect 230698 217482 230782 217718
rect 231018 217482 231102 217718
rect 231338 217482 231422 217718
rect 231658 217482 231742 217718
rect 231978 217482 232062 217718
rect 232298 217482 232382 217718
rect 232618 217482 237740 217718
rect 0 217440 237740 217482
rect 0 206518 237740 206560
rect 0 206282 122 206518
rect 358 206282 442 206518
rect 678 206282 762 206518
rect 998 206282 1082 206518
rect 1318 206282 1402 206518
rect 1638 206282 1722 206518
rect 1958 206282 2042 206518
rect 2278 206282 2362 206518
rect 2598 206282 2682 206518
rect 2918 206282 3002 206518
rect 3238 206282 3322 206518
rect 3558 206282 3642 206518
rect 3878 206282 42927 206518
rect 43163 206282 78882 206518
rect 79118 206282 115215 206518
rect 115451 206282 150882 206518
rect 151118 206282 187215 206518
rect 187451 206282 233862 206518
rect 234098 206282 234182 206518
rect 234418 206282 234502 206518
rect 234738 206282 234822 206518
rect 235058 206282 235142 206518
rect 235378 206282 235462 206518
rect 235698 206282 235782 206518
rect 236018 206282 236102 206518
rect 236338 206282 236422 206518
rect 236658 206282 236742 206518
rect 236978 206282 237062 206518
rect 237298 206282 237382 206518
rect 237618 206282 237740 206518
rect 0 206240 237740 206282
rect 0 195318 237740 195360
rect 0 195082 5122 195318
rect 5358 195082 5442 195318
rect 5678 195082 5762 195318
rect 5998 195082 6082 195318
rect 6318 195082 6402 195318
rect 6638 195082 6722 195318
rect 6958 195082 7042 195318
rect 7278 195082 7362 195318
rect 7598 195082 7682 195318
rect 7918 195082 8002 195318
rect 8238 195082 8322 195318
rect 8558 195082 8642 195318
rect 8878 195082 38261 195318
rect 38497 195082 73882 195318
rect 74118 195082 110549 195318
rect 110785 195082 145882 195318
rect 146118 195082 182549 195318
rect 182785 195082 228862 195318
rect 229098 195082 229182 195318
rect 229418 195082 229502 195318
rect 229738 195082 229822 195318
rect 230058 195082 230142 195318
rect 230378 195082 230462 195318
rect 230698 195082 230782 195318
rect 231018 195082 231102 195318
rect 231338 195082 231422 195318
rect 231658 195082 231742 195318
rect 231978 195082 232062 195318
rect 232298 195082 232382 195318
rect 232618 195082 237740 195318
rect 0 195040 237740 195082
rect 0 184118 237740 184160
rect 0 183882 122 184118
rect 358 183882 442 184118
rect 678 183882 762 184118
rect 998 183882 1082 184118
rect 1318 183882 1402 184118
rect 1638 183882 1722 184118
rect 1958 183882 2042 184118
rect 2278 183882 2362 184118
rect 2598 183882 2682 184118
rect 2918 183882 3002 184118
rect 3238 183882 3322 184118
rect 3558 183882 3642 184118
rect 3878 183882 233862 184118
rect 234098 183882 234182 184118
rect 234418 183882 234502 184118
rect 234738 183882 234822 184118
rect 235058 183882 235142 184118
rect 235378 183882 235462 184118
rect 235698 183882 235782 184118
rect 236018 183882 236102 184118
rect 236338 183882 236422 184118
rect 236658 183882 236742 184118
rect 236978 183882 237062 184118
rect 237298 183882 237382 184118
rect 237618 183882 237740 184118
rect 0 183840 237740 183882
rect 0 172918 237740 172960
rect 0 172682 5122 172918
rect 5358 172682 5442 172918
rect 5678 172682 5762 172918
rect 5998 172682 6082 172918
rect 6318 172682 6402 172918
rect 6638 172682 6722 172918
rect 6958 172682 7042 172918
rect 7278 172682 7362 172918
rect 7598 172682 7682 172918
rect 7918 172682 8002 172918
rect 8238 172682 8322 172918
rect 8558 172682 8642 172918
rect 8878 172682 17549 172918
rect 17785 172682 42549 172918
rect 42785 172682 67146 172918
rect 67382 172682 114549 172918
rect 114785 172682 139146 172918
rect 139382 172682 186549 172918
rect 186785 172682 211549 172918
rect 211785 172682 228862 172918
rect 229098 172682 229182 172918
rect 229418 172682 229502 172918
rect 229738 172682 229822 172918
rect 230058 172682 230142 172918
rect 230378 172682 230462 172918
rect 230698 172682 230782 172918
rect 231018 172682 231102 172918
rect 231338 172682 231422 172918
rect 231658 172682 231742 172918
rect 231978 172682 232062 172918
rect 232298 172682 232382 172918
rect 232618 172682 237740 172918
rect 0 172640 237740 172682
rect 0 161718 237740 161760
rect 0 161482 122 161718
rect 358 161482 442 161718
rect 678 161482 762 161718
rect 998 161482 1082 161718
rect 1318 161482 1402 161718
rect 1638 161482 1722 161718
rect 1958 161482 2042 161718
rect 2278 161482 2362 161718
rect 2598 161482 2682 161718
rect 2918 161482 3002 161718
rect 3238 161482 3322 161718
rect 3558 161482 3642 161718
rect 3878 161482 20215 161718
rect 20451 161482 45215 161718
rect 45451 161482 82506 161718
rect 82742 161482 117215 161718
rect 117451 161482 154506 161718
rect 154742 161482 189215 161718
rect 189451 161482 214215 161718
rect 214451 161482 233862 161718
rect 234098 161482 234182 161718
rect 234418 161482 234502 161718
rect 234738 161482 234822 161718
rect 235058 161482 235142 161718
rect 235378 161482 235462 161718
rect 235698 161482 235782 161718
rect 236018 161482 236102 161718
rect 236338 161482 236422 161718
rect 236658 161482 236742 161718
rect 236978 161482 237062 161718
rect 237298 161482 237382 161718
rect 237618 161482 237740 161718
rect 0 161440 237740 161482
rect 0 150518 237740 150560
rect 0 150282 5122 150518
rect 5358 150282 5442 150518
rect 5678 150282 5762 150518
rect 5998 150282 6082 150518
rect 6318 150282 6402 150518
rect 6638 150282 6722 150518
rect 6958 150282 7042 150518
rect 7278 150282 7362 150518
rect 7598 150282 7682 150518
rect 7918 150282 8002 150518
rect 8238 150282 8322 150518
rect 8558 150282 8642 150518
rect 8878 150282 17549 150518
rect 17785 150282 42549 150518
rect 42785 150282 67146 150518
rect 67382 150282 114549 150518
rect 114785 150282 139146 150518
rect 139382 150282 186549 150518
rect 186785 150282 211549 150518
rect 211785 150282 228862 150518
rect 229098 150282 229182 150518
rect 229418 150282 229502 150518
rect 229738 150282 229822 150518
rect 230058 150282 230142 150518
rect 230378 150282 230462 150518
rect 230698 150282 230782 150518
rect 231018 150282 231102 150518
rect 231338 150282 231422 150518
rect 231658 150282 231742 150518
rect 231978 150282 232062 150518
rect 232298 150282 232382 150518
rect 232618 150282 237740 150518
rect 0 150240 237740 150282
rect 0 139318 237740 139360
rect 0 139082 122 139318
rect 358 139082 442 139318
rect 678 139082 762 139318
rect 998 139082 1082 139318
rect 1318 139082 1402 139318
rect 1638 139082 1722 139318
rect 1958 139082 2042 139318
rect 2278 139082 2362 139318
rect 2598 139082 2682 139318
rect 2918 139082 3002 139318
rect 3238 139082 3322 139318
rect 3558 139082 3642 139318
rect 3878 139082 43215 139318
rect 43451 139082 115215 139318
rect 115451 139082 187215 139318
rect 187451 139082 233862 139318
rect 234098 139082 234182 139318
rect 234418 139082 234502 139318
rect 234738 139082 234822 139318
rect 235058 139082 235142 139318
rect 235378 139082 235462 139318
rect 235698 139082 235782 139318
rect 236018 139082 236102 139318
rect 236338 139082 236422 139318
rect 236658 139082 236742 139318
rect 236978 139082 237062 139318
rect 237298 139082 237382 139318
rect 237618 139082 237740 139318
rect 0 139040 237740 139082
rect 145988 138482 146492 138524
rect 145988 138246 146214 138482
rect 146450 138246 146492 138482
rect 145988 138204 146492 138246
rect 145988 137164 146308 138204
rect 142492 137122 146308 137164
rect 142492 136886 142534 137122
rect 142770 136886 146308 137122
rect 142492 136844 146308 136886
rect 67604 131682 101596 131724
rect 67604 131446 67646 131682
rect 67882 131446 101318 131682
rect 101554 131446 101596 131682
rect 67604 131404 101596 131446
rect 21420 128962 67924 129004
rect 21420 128726 21462 128962
rect 21698 128726 67646 128962
rect 67882 128726 67924 128962
rect 21420 128684 67924 128726
rect 0 128118 237740 128160
rect 0 127882 5122 128118
rect 5358 127882 5442 128118
rect 5678 127882 5762 128118
rect 5998 127882 6082 128118
rect 6318 127882 6402 128118
rect 6638 127882 6722 128118
rect 6958 127882 7042 128118
rect 7278 127882 7362 128118
rect 7598 127882 7682 128118
rect 7918 127882 8002 128118
rect 8238 127882 8322 128118
rect 8558 127882 8642 128118
rect 8878 127882 38549 128118
rect 38785 127882 73882 128118
rect 74118 127882 110549 128118
rect 110785 127882 145882 128118
rect 146118 127882 182549 128118
rect 182785 127882 228862 128118
rect 229098 127882 229182 128118
rect 229418 127882 229502 128118
rect 229738 127882 229822 128118
rect 230058 127882 230142 128118
rect 230378 127882 230462 128118
rect 230698 127882 230782 128118
rect 231018 127882 231102 128118
rect 231338 127882 231422 128118
rect 231658 127882 231742 128118
rect 231978 127882 232062 128118
rect 232298 127882 232382 128118
rect 232618 127882 237740 128118
rect 0 127840 237740 127882
rect 0 116918 237740 116960
rect 0 116682 122 116918
rect 358 116682 442 116918
rect 678 116682 762 116918
rect 998 116682 1082 116918
rect 1318 116682 1402 116918
rect 1638 116682 1722 116918
rect 1958 116682 2042 116918
rect 2278 116682 2362 116918
rect 2598 116682 2682 116918
rect 2918 116682 3002 116918
rect 3238 116682 3322 116918
rect 3558 116682 3642 116918
rect 3878 116682 43215 116918
rect 43451 116682 115215 116918
rect 115451 116682 187215 116918
rect 187451 116682 233862 116918
rect 234098 116682 234182 116918
rect 234418 116682 234502 116918
rect 234738 116682 234822 116918
rect 235058 116682 235142 116918
rect 235378 116682 235462 116918
rect 235698 116682 235782 116918
rect 236018 116682 236102 116918
rect 236338 116682 236422 116918
rect 236658 116682 236742 116918
rect 236978 116682 237062 116918
rect 237298 116682 237382 116918
rect 237618 116682 237740 116918
rect 0 116640 237740 116682
rect 31724 114002 58172 114044
rect 31724 113766 31766 114002
rect 32002 113766 56790 114002
rect 57026 113766 58172 114002
rect 31724 113724 58172 113766
rect 57852 113364 58172 113724
rect 57852 113322 73260 113364
rect 57852 113086 72982 113322
rect 73218 113086 73260 113322
rect 57852 113044 73260 113086
rect 0 105718 237740 105760
rect 0 105482 5122 105718
rect 5358 105482 5442 105718
rect 5678 105482 5762 105718
rect 5998 105482 6082 105718
rect 6318 105482 6402 105718
rect 6638 105482 6722 105718
rect 6958 105482 7042 105718
rect 7278 105482 7362 105718
rect 7598 105482 7682 105718
rect 7918 105482 8002 105718
rect 8238 105482 8322 105718
rect 8558 105482 8642 105718
rect 8878 105482 17549 105718
rect 17785 105482 42549 105718
rect 42785 105482 67146 105718
rect 67382 105482 114549 105718
rect 114785 105482 139146 105718
rect 139382 105482 186549 105718
rect 186785 105482 211549 105718
rect 211785 105482 228862 105718
rect 229098 105482 229182 105718
rect 229418 105482 229502 105718
rect 229738 105482 229822 105718
rect 230058 105482 230142 105718
rect 230378 105482 230462 105718
rect 230698 105482 230782 105718
rect 231018 105482 231102 105718
rect 231338 105482 231422 105718
rect 231658 105482 231742 105718
rect 231978 105482 232062 105718
rect 232298 105482 232382 105718
rect 232618 105482 237740 105718
rect 0 105440 237740 105482
rect 0 94518 237740 94560
rect 0 94282 122 94518
rect 358 94282 442 94518
rect 678 94282 762 94518
rect 998 94282 1082 94518
rect 1318 94282 1402 94518
rect 1638 94282 1722 94518
rect 1958 94282 2042 94518
rect 2278 94282 2362 94518
rect 2598 94282 2682 94518
rect 2918 94282 3002 94518
rect 3238 94282 3322 94518
rect 3558 94282 3642 94518
rect 3878 94282 20215 94518
rect 20451 94282 45215 94518
rect 45451 94282 82506 94518
rect 82742 94282 117215 94518
rect 117451 94282 154506 94518
rect 154742 94282 189215 94518
rect 189451 94282 214215 94518
rect 214451 94282 233862 94518
rect 234098 94282 234182 94518
rect 234418 94282 234502 94518
rect 234738 94282 234822 94518
rect 235058 94282 235142 94518
rect 235378 94282 235462 94518
rect 235698 94282 235782 94518
rect 236018 94282 236102 94518
rect 236338 94282 236422 94518
rect 236658 94282 236742 94518
rect 236978 94282 237062 94518
rect 237298 94282 237382 94518
rect 237618 94282 237740 94518
rect 0 94240 237740 94282
rect 0 83318 237740 83360
rect 0 83082 5122 83318
rect 5358 83082 5442 83318
rect 5678 83082 5762 83318
rect 5998 83082 6082 83318
rect 6318 83082 6402 83318
rect 6638 83082 6722 83318
rect 6958 83082 7042 83318
rect 7278 83082 7362 83318
rect 7598 83082 7682 83318
rect 7918 83082 8002 83318
rect 8238 83082 8322 83318
rect 8558 83082 8642 83318
rect 8878 83082 17549 83318
rect 17785 83082 42549 83318
rect 42785 83082 67146 83318
rect 67382 83082 114549 83318
rect 114785 83082 139146 83318
rect 139382 83082 186549 83318
rect 186785 83082 211549 83318
rect 211785 83082 228862 83318
rect 229098 83082 229182 83318
rect 229418 83082 229502 83318
rect 229738 83082 229822 83318
rect 230058 83082 230142 83318
rect 230378 83082 230462 83318
rect 230698 83082 230782 83318
rect 231018 83082 231102 83318
rect 231338 83082 231422 83318
rect 231658 83082 231742 83318
rect 231978 83082 232062 83318
rect 232298 83082 232382 83318
rect 232618 83082 237740 83318
rect 0 83040 237740 83082
rect 0 72118 237740 72160
rect 0 71882 122 72118
rect 358 71882 442 72118
rect 678 71882 762 72118
rect 998 71882 1082 72118
rect 1318 71882 1402 72118
rect 1638 71882 1722 72118
rect 1958 71882 2042 72118
rect 2278 71882 2362 72118
rect 2598 71882 2682 72118
rect 2918 71882 3002 72118
rect 3238 71882 3322 72118
rect 3558 71882 3642 72118
rect 3878 71882 233862 72118
rect 234098 71882 234182 72118
rect 234418 71882 234502 72118
rect 234738 71882 234822 72118
rect 235058 71882 235142 72118
rect 235378 71882 235462 72118
rect 235698 71882 235782 72118
rect 236018 71882 236102 72118
rect 236338 71882 236422 72118
rect 236658 71882 236742 72118
rect 236978 71882 237062 72118
rect 237298 71882 237382 72118
rect 237618 71882 237740 72118
rect 0 71840 237740 71882
rect 0 60918 237740 60960
rect 0 60682 5122 60918
rect 5358 60682 5442 60918
rect 5678 60682 5762 60918
rect 5998 60682 6082 60918
rect 6318 60682 6402 60918
rect 6638 60682 6722 60918
rect 6958 60682 7042 60918
rect 7278 60682 7362 60918
rect 7598 60682 7682 60918
rect 7918 60682 8002 60918
rect 8238 60682 8322 60918
rect 8558 60682 8642 60918
rect 8878 60682 38549 60918
rect 38785 60682 73882 60918
rect 74118 60682 110549 60918
rect 110785 60682 145882 60918
rect 146118 60682 182549 60918
rect 182785 60682 228862 60918
rect 229098 60682 229182 60918
rect 229418 60682 229502 60918
rect 229738 60682 229822 60918
rect 230058 60682 230142 60918
rect 230378 60682 230462 60918
rect 230698 60682 230782 60918
rect 231018 60682 231102 60918
rect 231338 60682 231422 60918
rect 231658 60682 231742 60918
rect 231978 60682 232062 60918
rect 232298 60682 232382 60918
rect 232618 60682 237740 60918
rect 0 60640 237740 60682
rect 0 49718 237740 49760
rect 0 49482 122 49718
rect 358 49482 442 49718
rect 678 49482 762 49718
rect 998 49482 1082 49718
rect 1318 49482 1402 49718
rect 1638 49482 1722 49718
rect 1958 49482 2042 49718
rect 2278 49482 2362 49718
rect 2598 49482 2682 49718
rect 2918 49482 3002 49718
rect 3238 49482 3322 49718
rect 3558 49482 3642 49718
rect 3878 49482 43215 49718
rect 43451 49482 78882 49718
rect 79118 49482 115215 49718
rect 115451 49482 150882 49718
rect 151118 49482 187215 49718
rect 187451 49482 233862 49718
rect 234098 49482 234182 49718
rect 234418 49482 234502 49718
rect 234738 49482 234822 49718
rect 235058 49482 235142 49718
rect 235378 49482 235462 49718
rect 235698 49482 235782 49718
rect 236018 49482 236102 49718
rect 236338 49482 236422 49718
rect 236658 49482 236742 49718
rect 236978 49482 237062 49718
rect 237298 49482 237382 49718
rect 237618 49482 237740 49718
rect 0 49440 237740 49482
rect 31724 41242 66452 41284
rect 31724 41006 31766 41242
rect 32002 41006 66174 41242
rect 66410 41006 66452 41242
rect 31724 40964 66452 41006
rect 93732 40562 108956 40604
rect 93732 40326 93774 40562
rect 94010 40326 108678 40562
rect 108914 40326 108956 40562
rect 93732 40284 108956 40326
rect 109556 40562 118708 40604
rect 109556 40326 109598 40562
rect 109834 40326 118708 40562
rect 109556 40284 118708 40326
rect 99252 38924 99756 40284
rect 118388 39244 118708 40284
rect 128508 40562 137108 40604
rect 128508 40326 129654 40562
rect 129890 40326 136830 40562
rect 137066 40326 137108 40562
rect 128508 40284 137108 40326
rect 171380 40562 190652 40604
rect 171380 40326 181358 40562
rect 181594 40326 190652 40562
rect 171380 40284 190652 40326
rect 128508 39244 128828 40284
rect 171380 39924 171700 40284
rect 166044 39882 171700 39924
rect 166044 39646 166086 39882
rect 166322 39646 171700 39882
rect 166044 39604 171700 39646
rect 118388 38924 128828 39244
rect 190332 39244 190652 40284
rect 190332 39202 201692 39244
rect 190332 38966 201414 39202
rect 201650 38966 201692 39202
rect 190332 38924 201692 38966
rect 0 38518 237740 38560
rect 0 38282 5122 38518
rect 5358 38282 5442 38518
rect 5678 38282 5762 38518
rect 5998 38282 6082 38518
rect 6318 38282 6402 38518
rect 6638 38282 6722 38518
rect 6958 38282 7042 38518
rect 7278 38282 7362 38518
rect 7598 38282 7682 38518
rect 7918 38282 8002 38518
rect 8238 38282 8322 38518
rect 8558 38282 8642 38518
rect 8878 38282 228862 38518
rect 229098 38282 229182 38518
rect 229418 38282 229502 38518
rect 229738 38282 229822 38518
rect 230058 38282 230142 38518
rect 230378 38282 230462 38518
rect 230698 38282 230782 38518
rect 231018 38282 231102 38518
rect 231338 38282 231422 38518
rect 231658 38282 231742 38518
rect 231978 38282 232062 38518
rect 232298 38282 232382 38518
rect 232618 38282 237740 38518
rect 0 38240 237740 38282
rect 0 27318 237740 27360
rect 0 27082 122 27318
rect 358 27082 442 27318
rect 678 27082 762 27318
rect 998 27082 1082 27318
rect 1318 27082 1402 27318
rect 1638 27082 1722 27318
rect 1958 27082 2042 27318
rect 2278 27082 2362 27318
rect 2598 27082 2682 27318
rect 2918 27082 3002 27318
rect 3238 27082 3322 27318
rect 3558 27082 3642 27318
rect 3878 27082 78882 27318
rect 79118 27082 150882 27318
rect 151118 27082 233862 27318
rect 234098 27082 234182 27318
rect 234418 27082 234502 27318
rect 234738 27082 234822 27318
rect 235058 27082 235142 27318
rect 235378 27082 235462 27318
rect 235698 27082 235782 27318
rect 236018 27082 236102 27318
rect 236338 27082 236422 27318
rect 236658 27082 236742 27318
rect 236978 27082 237062 27318
rect 237298 27082 237382 27318
rect 237618 27082 237740 27318
rect 0 27040 237740 27082
rect 0 16118 237740 16160
rect 0 15882 5122 16118
rect 5358 15882 5442 16118
rect 5678 15882 5762 16118
rect 5998 15882 6082 16118
rect 6318 15882 6402 16118
rect 6638 15882 6722 16118
rect 6958 15882 7042 16118
rect 7278 15882 7362 16118
rect 7598 15882 7682 16118
rect 7918 15882 8002 16118
rect 8238 15882 8322 16118
rect 8558 15882 8642 16118
rect 8878 15882 73882 16118
rect 74118 15882 145882 16118
rect 146118 15882 228862 16118
rect 229098 15882 229182 16118
rect 229418 15882 229502 16118
rect 229738 15882 229822 16118
rect 230058 15882 230142 16118
rect 230378 15882 230462 16118
rect 230698 15882 230782 16118
rect 231018 15882 231102 16118
rect 231338 15882 231422 16118
rect 231658 15882 231742 16118
rect 231978 15882 232062 16118
rect 232298 15882 232382 16118
rect 232618 15882 237740 16118
rect 0 15840 237740 15882
rect 5000 8878 232740 9000
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 228862 8878
rect 229098 8642 229182 8878
rect 229418 8642 229502 8878
rect 229738 8642 229822 8878
rect 230058 8642 230142 8878
rect 230378 8642 230462 8878
rect 230698 8642 230782 8878
rect 231018 8642 231102 8878
rect 231338 8642 231422 8878
rect 231658 8642 231742 8878
rect 231978 8642 232062 8878
rect 232298 8642 232382 8878
rect 232618 8642 232740 8878
rect 5000 8558 232740 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 228862 8558
rect 229098 8322 229182 8558
rect 229418 8322 229502 8558
rect 229738 8322 229822 8558
rect 230058 8322 230142 8558
rect 230378 8322 230462 8558
rect 230698 8322 230782 8558
rect 231018 8322 231102 8558
rect 231338 8322 231422 8558
rect 231658 8322 231742 8558
rect 231978 8322 232062 8558
rect 232298 8322 232382 8558
rect 232618 8322 232740 8558
rect 5000 8238 232740 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 228862 8238
rect 229098 8002 229182 8238
rect 229418 8002 229502 8238
rect 229738 8002 229822 8238
rect 230058 8002 230142 8238
rect 230378 8002 230462 8238
rect 230698 8002 230782 8238
rect 231018 8002 231102 8238
rect 231338 8002 231422 8238
rect 231658 8002 231742 8238
rect 231978 8002 232062 8238
rect 232298 8002 232382 8238
rect 232618 8002 232740 8238
rect 5000 7918 232740 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 228862 7918
rect 229098 7682 229182 7918
rect 229418 7682 229502 7918
rect 229738 7682 229822 7918
rect 230058 7682 230142 7918
rect 230378 7682 230462 7918
rect 230698 7682 230782 7918
rect 231018 7682 231102 7918
rect 231338 7682 231422 7918
rect 231658 7682 231742 7918
rect 231978 7682 232062 7918
rect 232298 7682 232382 7918
rect 232618 7682 232740 7918
rect 5000 7598 232740 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 228862 7598
rect 229098 7362 229182 7598
rect 229418 7362 229502 7598
rect 229738 7362 229822 7598
rect 230058 7362 230142 7598
rect 230378 7362 230462 7598
rect 230698 7362 230782 7598
rect 231018 7362 231102 7598
rect 231338 7362 231422 7598
rect 231658 7362 231742 7598
rect 231978 7362 232062 7598
rect 232298 7362 232382 7598
rect 232618 7362 232740 7598
rect 5000 7278 232740 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 228862 7278
rect 229098 7042 229182 7278
rect 229418 7042 229502 7278
rect 229738 7042 229822 7278
rect 230058 7042 230142 7278
rect 230378 7042 230462 7278
rect 230698 7042 230782 7278
rect 231018 7042 231102 7278
rect 231338 7042 231422 7278
rect 231658 7042 231742 7278
rect 231978 7042 232062 7278
rect 232298 7042 232382 7278
rect 232618 7042 232740 7278
rect 5000 6958 232740 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 228862 6958
rect 229098 6722 229182 6958
rect 229418 6722 229502 6958
rect 229738 6722 229822 6958
rect 230058 6722 230142 6958
rect 230378 6722 230462 6958
rect 230698 6722 230782 6958
rect 231018 6722 231102 6958
rect 231338 6722 231422 6958
rect 231658 6722 231742 6958
rect 231978 6722 232062 6958
rect 232298 6722 232382 6958
rect 232618 6722 232740 6958
rect 5000 6638 232740 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 228862 6638
rect 229098 6402 229182 6638
rect 229418 6402 229502 6638
rect 229738 6402 229822 6638
rect 230058 6402 230142 6638
rect 230378 6402 230462 6638
rect 230698 6402 230782 6638
rect 231018 6402 231102 6638
rect 231338 6402 231422 6638
rect 231658 6402 231742 6638
rect 231978 6402 232062 6638
rect 232298 6402 232382 6638
rect 232618 6402 232740 6638
rect 5000 6318 232740 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 228862 6318
rect 229098 6082 229182 6318
rect 229418 6082 229502 6318
rect 229738 6082 229822 6318
rect 230058 6082 230142 6318
rect 230378 6082 230462 6318
rect 230698 6082 230782 6318
rect 231018 6082 231102 6318
rect 231338 6082 231422 6318
rect 231658 6082 231742 6318
rect 231978 6082 232062 6318
rect 232298 6082 232382 6318
rect 232618 6082 232740 6318
rect 5000 5998 232740 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 228862 5998
rect 229098 5762 229182 5998
rect 229418 5762 229502 5998
rect 229738 5762 229822 5998
rect 230058 5762 230142 5998
rect 230378 5762 230462 5998
rect 230698 5762 230782 5998
rect 231018 5762 231102 5998
rect 231338 5762 231422 5998
rect 231658 5762 231742 5998
rect 231978 5762 232062 5998
rect 232298 5762 232382 5998
rect 232618 5762 232740 5998
rect 5000 5678 232740 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 228862 5678
rect 229098 5442 229182 5678
rect 229418 5442 229502 5678
rect 229738 5442 229822 5678
rect 230058 5442 230142 5678
rect 230378 5442 230462 5678
rect 230698 5442 230782 5678
rect 231018 5442 231102 5678
rect 231338 5442 231422 5678
rect 231658 5442 231742 5678
rect 231978 5442 232062 5678
rect 232298 5442 232382 5678
rect 232618 5442 232740 5678
rect 5000 5358 232740 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 228862 5358
rect 229098 5122 229182 5358
rect 229418 5122 229502 5358
rect 229738 5122 229822 5358
rect 230058 5122 230142 5358
rect 230378 5122 230462 5358
rect 230698 5122 230782 5358
rect 231018 5122 231102 5358
rect 231338 5122 231422 5358
rect 231658 5122 231742 5358
rect 231978 5122 232062 5358
rect 232298 5122 232382 5358
rect 232618 5122 232740 5358
rect 5000 5000 232740 5122
rect 0 3878 237740 4000
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 233862 3878
rect 234098 3642 234182 3878
rect 234418 3642 234502 3878
rect 234738 3642 234822 3878
rect 235058 3642 235142 3878
rect 235378 3642 235462 3878
rect 235698 3642 235782 3878
rect 236018 3642 236102 3878
rect 236338 3642 236422 3878
rect 236658 3642 236742 3878
rect 236978 3642 237062 3878
rect 237298 3642 237382 3878
rect 237618 3642 237740 3878
rect 0 3558 237740 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 233862 3558
rect 234098 3322 234182 3558
rect 234418 3322 234502 3558
rect 234738 3322 234822 3558
rect 235058 3322 235142 3558
rect 235378 3322 235462 3558
rect 235698 3322 235782 3558
rect 236018 3322 236102 3558
rect 236338 3322 236422 3558
rect 236658 3322 236742 3558
rect 236978 3322 237062 3558
rect 237298 3322 237382 3558
rect 237618 3322 237740 3558
rect 0 3238 237740 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 233862 3238
rect 234098 3002 234182 3238
rect 234418 3002 234502 3238
rect 234738 3002 234822 3238
rect 235058 3002 235142 3238
rect 235378 3002 235462 3238
rect 235698 3002 235782 3238
rect 236018 3002 236102 3238
rect 236338 3002 236422 3238
rect 236658 3002 236742 3238
rect 236978 3002 237062 3238
rect 237298 3002 237382 3238
rect 237618 3002 237740 3238
rect 0 2918 237740 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 233862 2918
rect 234098 2682 234182 2918
rect 234418 2682 234502 2918
rect 234738 2682 234822 2918
rect 235058 2682 235142 2918
rect 235378 2682 235462 2918
rect 235698 2682 235782 2918
rect 236018 2682 236102 2918
rect 236338 2682 236422 2918
rect 236658 2682 236742 2918
rect 236978 2682 237062 2918
rect 237298 2682 237382 2918
rect 237618 2682 237740 2918
rect 0 2598 237740 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 233862 2598
rect 234098 2362 234182 2598
rect 234418 2362 234502 2598
rect 234738 2362 234822 2598
rect 235058 2362 235142 2598
rect 235378 2362 235462 2598
rect 235698 2362 235782 2598
rect 236018 2362 236102 2598
rect 236338 2362 236422 2598
rect 236658 2362 236742 2598
rect 236978 2362 237062 2598
rect 237298 2362 237382 2598
rect 237618 2362 237740 2598
rect 0 2278 237740 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 233862 2278
rect 234098 2042 234182 2278
rect 234418 2042 234502 2278
rect 234738 2042 234822 2278
rect 235058 2042 235142 2278
rect 235378 2042 235462 2278
rect 235698 2042 235782 2278
rect 236018 2042 236102 2278
rect 236338 2042 236422 2278
rect 236658 2042 236742 2278
rect 236978 2042 237062 2278
rect 237298 2042 237382 2278
rect 237618 2042 237740 2278
rect 0 1958 237740 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 233862 1958
rect 234098 1722 234182 1958
rect 234418 1722 234502 1958
rect 234738 1722 234822 1958
rect 235058 1722 235142 1958
rect 235378 1722 235462 1958
rect 235698 1722 235782 1958
rect 236018 1722 236102 1958
rect 236338 1722 236422 1958
rect 236658 1722 236742 1958
rect 236978 1722 237062 1958
rect 237298 1722 237382 1958
rect 237618 1722 237740 1958
rect 0 1638 237740 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 233862 1638
rect 234098 1402 234182 1638
rect 234418 1402 234502 1638
rect 234738 1402 234822 1638
rect 235058 1402 235142 1638
rect 235378 1402 235462 1638
rect 235698 1402 235782 1638
rect 236018 1402 236102 1638
rect 236338 1402 236422 1638
rect 236658 1402 236742 1638
rect 236978 1402 237062 1638
rect 237298 1402 237382 1638
rect 237618 1402 237740 1638
rect 0 1318 237740 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 233862 1318
rect 234098 1082 234182 1318
rect 234418 1082 234502 1318
rect 234738 1082 234822 1318
rect 235058 1082 235142 1318
rect 235378 1082 235462 1318
rect 235698 1082 235782 1318
rect 236018 1082 236102 1318
rect 236338 1082 236422 1318
rect 236658 1082 236742 1318
rect 236978 1082 237062 1318
rect 237298 1082 237382 1318
rect 237618 1082 237740 1318
rect 0 998 237740 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 233862 998
rect 234098 762 234182 998
rect 234418 762 234502 998
rect 234738 762 234822 998
rect 235058 762 235142 998
rect 235378 762 235462 998
rect 235698 762 235782 998
rect 236018 762 236102 998
rect 236338 762 236422 998
rect 236658 762 236742 998
rect 236978 762 237062 998
rect 237298 762 237382 998
rect 237618 762 237740 998
rect 0 678 237740 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 233862 678
rect 234098 442 234182 678
rect 234418 442 234502 678
rect 234738 442 234822 678
rect 235058 442 235142 678
rect 235378 442 235462 678
rect 235698 442 235782 678
rect 236018 442 236102 678
rect 236338 442 236422 678
rect 236658 442 236742 678
rect 236978 442 237062 678
rect 237298 442 237382 678
rect 237618 442 237740 678
rect 0 358 237740 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 233862 358
rect 234098 122 234182 358
rect 234418 122 234502 358
rect 234738 122 234822 358
rect 235058 122 235142 358
rect 235378 122 235462 358
rect 235698 122 235782 358
rect 236018 122 236102 358
rect 236338 122 236422 358
rect 236658 122 236742 358
rect 236978 122 237062 358
rect 237298 122 237382 358
rect 237618 122 237740 358
rect 0 0 237740 122
use sb_0__0_  sb_0__0_
timestamp 1604675407
transform 1 0 32896 0 1 39824
box 0 0 28000 27720
use grid_io_bottom  grid_io_bottom_1__0_
timestamp 1604675407
transform 1 0 67896 0 1 12824
box 0 0 28926 24000
use cbx_1__0_  cbx_1__0_
timestamp 1604675407
transform 1 0 67896 0 1 41824
box 0 0 30000 24000
use sb_1__0_  sb_1__0_
timestamp 1604675407
transform 1 0 104896 0 1 39824
box 0 0 28000 28000
use grid_io_bottom  grid_io_bottom_2__0_
timestamp 1604675407
transform 1 0 139896 0 1 12824
box 0 0 28926 24000
use cbx_1__0_  cbx_2__0_
timestamp 1604675407
transform 1 0 139896 0 1 41824
box 0 0 30000 24000
use sb_2__0_  sb_2__0_
timestamp 1604675407
transform 1 0 176896 0 1 39824
box 0 0 27679 28000
use grid_io_left  grid_io_left_0__1_
timestamp 1604675407
transform 1 0 13896 0 1 70824
box 0 0 16000 37584
use cby_0__1_  cby_0__1_
timestamp 1604675407
transform 1 0 38896 0 1 70824
box 0 0 16000 40000
use grid_clb  grid_clb_1__1_
timestamp 1604675407
transform 1 0 62896 0 1 70824
box 0 0 40000 40000
use cby_1__1_  cby_1__1_
timestamp 1604675407
transform 1 0 110896 0 1 70824
box 0 0 16000 40000
use grid_clb  grid_clb_2__1_
timestamp 1604675407
transform 1 0 134896 0 1 70824
box 0 0 40000 40000
use grid_io_right  grid_io_right_3__1_
timestamp 1604675407
transform 1 0 207896 0 1 70824
box 0 0 16000 37584
use cby_1__1_  cby_2__1_
timestamp 1604675407
transform 1 0 182896 0 1 70824
box 0 0 16000 40000
use grid_io_left  grid_io_left_0__2_
timestamp 1604675407
transform 1 0 13896 0 1 144824
box 0 0 16000 37584
use sb_0__1_  sb_0__1_
timestamp 1604675407
transform 1 0 32896 0 1 113824
box 0 0 28000 28000
use cby_0__1_  cby_0__2_
timestamp 1604675407
transform 1 0 38896 0 1 144824
box 0 0 16000 40000
use grid_clb  grid_clb_1__2_
timestamp 1604675407
transform 1 0 62896 0 1 144824
box 0 0 40000 40000
use cbx_1__1_  cbx_1__1_
timestamp 1604675407
transform 1 0 67896 0 1 115824
box 0 0 30000 24000
use sb_1__1_  sb_1__1_
timestamp 1604675407
transform 1 0 104896 0 1 113824
box 0 0 28000 28000
use cby_1__1_  cby_1__2_
timestamp 1604675407
transform 1 0 110896 0 1 144824
box 0 0 16000 40000
use grid_clb  grid_clb_2__2_
timestamp 1604675407
transform 1 0 134896 0 1 144824
box 0 0 40000 40000
use cbx_1__1_  cbx_2__1_
timestamp 1604675407
transform 1 0 139896 0 1 115824
box 0 0 30000 24000
use grid_io_right  grid_io_right_3__2_
timestamp 1604675407
transform 1 0 207896 0 1 144824
box 0 0 16000 37584
use sb_2__1_  sb_2__1_
timestamp 1604675407
transform 1 0 176896 0 1 113824
box 0 0 28000 28000
use cby_1__1_  cby_2__2_
timestamp 1604675407
transform 1 0 182896 0 1 144824
box 0 0 16000 40000
use sb_0__2_  sb_0__2_
timestamp 1604675407
transform 1 0 32895 0 1 187824
box 1 0 27712 28000
use cbx_1__2_  cbx_1__2_
timestamp 1604675407
transform 1 0 67896 0 1 189824
box 0 0 30000 23826
use sb_1__2_  sb_1__2_
timestamp 1604675407
transform 1 0 104896 0 1 187824
box 0 0 28000 28000
use cbx_1__2_  cbx_2__2_
timestamp 1604675407
transform 1 0 139896 0 1 189824
box 0 0 30000 23826
use sb_2__2_  sb_2__2_
timestamp 1604675407
transform 1 0 176896 0 1 187824
box 0 0 28000 27600
use grid_io_top  grid_io_top_1__3_
timestamp 1604675407
transform 1 0 67896 0 1 218824
box 0 0 28934 24000
use grid_io_top  grid_io_top_2__3_
timestamp 1604675407
transform 1 0 139896 0 1 218824
box 0 0 28934 24000
<< labels >>
rlabel metal3 s 9896 127696 10376 127816 6 Test_en
port 0 nsew default input
rlabel metal3 s 227416 211064 227896 211184 6 ccff_head
port 1 nsew default input
rlabel metal3 s 9896 19576 10376 19696 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 9896 149320 10376 149440 6 clk
port 3 nsew default input
rlabel metal2 s 23530 246344 23586 246824 6 gfpga_pad_GPIO_A[0]
port 4 nsew default tristate
rlabel metal2 s 50762 246344 50818 246824 6 gfpga_pad_GPIO_A[1]
port 5 nsew default tristate
rlabel metal3 s 227416 20664 227896 20784 6 gfpga_pad_GPIO_A[2]
port 6 nsew default tristate
rlabel metal3 s 227416 44464 227896 44584 6 gfpga_pad_GPIO_A[3]
port 7 nsew default tristate
rlabel metal2 s 23530 8824 23586 9304 6 gfpga_pad_GPIO_A[4]
port 8 nsew default tristate
rlabel metal2 s 50762 8824 50818 9304 6 gfpga_pad_GPIO_A[5]
port 9 nsew default tristate
rlabel metal3 s 9896 41200 10376 41320 6 gfpga_pad_GPIO_A[6]
port 10 nsew default tristate
rlabel metal3 s 9896 62824 10376 62944 6 gfpga_pad_GPIO_A[7]
port 11 nsew default tristate
rlabel metal2 s 77994 246344 78050 246824 6 gfpga_pad_GPIO_IE[0]
port 12 nsew default tristate
rlabel metal2 s 105226 246344 105282 246824 6 gfpga_pad_GPIO_IE[1]
port 13 nsew default tristate
rlabel metal3 s 227416 68264 227896 68384 6 gfpga_pad_GPIO_IE[2]
port 14 nsew default tristate
rlabel metal3 s 227416 92064 227896 92184 6 gfpga_pad_GPIO_IE[3]
port 15 nsew default tristate
rlabel metal2 s 77994 8824 78050 9304 6 gfpga_pad_GPIO_IE[4]
port 16 nsew default tristate
rlabel metal2 s 105226 8824 105282 9304 6 gfpga_pad_GPIO_IE[5]
port 17 nsew default tristate
rlabel metal3 s 9896 84448 10376 84568 6 gfpga_pad_GPIO_IE[6]
port 18 nsew default tristate
rlabel metal3 s 9896 106072 10376 106192 6 gfpga_pad_GPIO_IE[7]
port 19 nsew default tristate
rlabel metal2 s 132550 246344 132606 246824 6 gfpga_pad_GPIO_OE[0]
port 20 nsew default tristate
rlabel metal2 s 159782 246344 159838 246824 6 gfpga_pad_GPIO_OE[1]
port 21 nsew default tristate
rlabel metal3 s 227416 115864 227896 115984 6 gfpga_pad_GPIO_OE[2]
port 22 nsew default tristate
rlabel metal3 s 227416 139664 227896 139784 6 gfpga_pad_GPIO_OE[3]
port 23 nsew default tristate
rlabel metal2 s 132550 8824 132606 9304 6 gfpga_pad_GPIO_OE[4]
port 24 nsew default tristate
rlabel metal2 s 159782 8824 159838 9304 6 gfpga_pad_GPIO_OE[5]
port 25 nsew default tristate
rlabel metal3 s 9896 170944 10376 171064 6 gfpga_pad_GPIO_OE[6]
port 26 nsew default tristate
rlabel metal3 s 9896 192568 10376 192688 6 gfpga_pad_GPIO_OE[7]
port 27 nsew default tristate
rlabel metal2 s 187014 246344 187070 246824 6 gfpga_pad_GPIO_Y[0]
port 28 nsew default bidirectional
rlabel metal2 s 214246 246344 214302 246824 6 gfpga_pad_GPIO_Y[1]
port 29 nsew default bidirectional
rlabel metal3 s 227416 163464 227896 163584 6 gfpga_pad_GPIO_Y[2]
port 30 nsew default bidirectional
rlabel metal3 s 227416 187264 227896 187384 6 gfpga_pad_GPIO_Y[3]
port 31 nsew default bidirectional
rlabel metal2 s 187014 8824 187070 9304 6 gfpga_pad_GPIO_Y[4]
port 32 nsew default bidirectional
rlabel metal2 s 214246 8824 214302 9304 6 gfpga_pad_GPIO_Y[5]
port 33 nsew default bidirectional
rlabel metal3 s 9896 214192 10376 214312 6 gfpga_pad_GPIO_Y[6]
port 34 nsew default bidirectional
rlabel metal3 s 9896 235816 10376 235936 6 gfpga_pad_GPIO_Y[7]
port 35 nsew default bidirectional
rlabel metal3 s 227416 234864 227896 234984 6 prog_clk
port 36 nsew default input
rlabel metal5 s 5000 5000 232740 9000 8 VPWR
port 37 nsew default input
rlabel metal5 s 0 0 237740 4000 8 VGND
port 38 nsew default input
<< properties >>
string FIXED_BBOX 0 0 237740 255376
<< end >>
