* NGSPICE file created from cbx_1__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

.subckt cbx_1__0_ SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP bottom_grid_pin_0_ bottom_grid_pin_10_
+ bottom_grid_pin_2_ bottom_grid_pin_4_ bottom_grid_pin_6_ bottom_grid_pin_8_ ccff_head
+ ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] gfpga_pad_EMBEDDED_IO_SOC_DIR[0] gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
+ gfpga_pad_EMBEDDED_IO_SOC_DIR[2] gfpga_pad_EMBEDDED_IO_SOC_DIR[3] gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
+ gfpga_pad_EMBEDDED_IO_SOC_DIR[5] gfpga_pad_EMBEDDED_IO_SOC_IN[0] gfpga_pad_EMBEDDED_IO_SOC_IN[1]
+ gfpga_pad_EMBEDDED_IO_SOC_IN[2] gfpga_pad_EMBEDDED_IO_SOC_IN[3] gfpga_pad_EMBEDDED_IO_SOC_IN[4]
+ gfpga_pad_EMBEDDED_IO_SOC_IN[5] gfpga_pad_EMBEDDED_IO_SOC_OUT[0] gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
+ gfpga_pad_EMBEDDED_IO_SOC_OUT[2] gfpga_pad_EMBEDDED_IO_SOC_OUT[3] gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
+ gfpga_pad_EMBEDDED_IO_SOC_OUT[5] prog_clk top_width_0_height_0__pin_0_ top_width_0_height_0__pin_10_
+ top_width_0_height_0__pin_11_lower top_width_0_height_0__pin_11_upper top_width_0_height_0__pin_1_lower
+ top_width_0_height_0__pin_1_upper top_width_0_height_0__pin_2_ top_width_0_height_0__pin_3_lower
+ top_width_0_height_0__pin_3_upper top_width_0_height_0__pin_4_ top_width_0_height_0__pin_5_lower
+ top_width_0_height_0__pin_5_upper top_width_0_height_0__pin_6_ top_width_0_height_0__pin_7_lower
+ top_width_0_height_0__pin_7_upper top_width_0_height_0__pin_8_ top_width_0_height_0__pin_9_lower
+ top_width_0_height_0__pin_9_upper VPWR VGND
Xmux_top_ipin_1.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_1.mux_l1_in_2_/S
+ mux_top_ipin_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_66_ gfpga_pad_EMBEDDED_IO_SOC_IN[3] top_width_0_height_0__pin_7_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_49_ _49_/A gfpga_pad_EMBEDDED_IO_SOC_DIR[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_1.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_1.mux_l1_in_2_/S
+ mux_top_ipin_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_65_ gfpga_pad_EMBEDDED_IO_SOC_IN[3] top_width_0_height_0__pin_7_lower VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
X_48_ _48_/A gfpga_pad_EMBEDDED_IO_SOC_DIR[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_64_ gfpga_pad_EMBEDDED_IO_SOC_IN[2] top_width_0_height_0__pin_5_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_4.mux_l4_in_0_/X bottom_grid_pin_8_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_47_ _47_/A gfpga_pad_EMBEDDED_IO_SOC_DIR[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_1_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_2_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_13_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_63_ gfpga_pad_EMBEDDED_IO_SOC_IN[2] top_width_0_height_0__pin_5_lower VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_46_ _46_/A gfpga_pad_EMBEDDED_IO_SOC_DIR[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29_ chanx_left_in[15] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_2.mux_l2_in_3_ _08_/HI chanx_right_in[18] mux_top_ipin_2.mux_l2_in_1_/S
+ mux_top_ipin_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_62_ gfpga_pad_EMBEDDED_IO_SOC_IN[1] top_width_0_height_0__pin_3_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_2.mux_l4_in_0_ mux_top_ipin_2.mux_l3_in_1_/X mux_top_ipin_2.mux_l3_in_0_/X
+ mux_top_ipin_2.mux_l4_in_0_/S mux_top_ipin_2.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_45_ ccff_tail gfpga_pad_EMBEDDED_IO_SOC_DIR[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_io_mode_io__3.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ _48_/A _47_/A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28_ chanx_left_in[16] chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_2.mux_l3_in_1_ mux_top_ipin_2.mux_l2_in_3_/X mux_top_ipin_2.mux_l2_in_2_/X
+ mux_top_ipin_2.mux_l3_in_0_/S mux_top_ipin_2.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_2.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_2.mux_l2_in_1_/S
+ mux_top_ipin_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_61_ gfpga_pad_EMBEDDED_IO_SOC_IN[1] top_width_0_height_0__pin_3_lower VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_44_ chanx_left_in[0] chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27_ chanx_left_in[17] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_2.mux_l3_in_0_ mux_top_ipin_2.mux_l2_in_1_/X mux_top_ipin_2.mux_l2_in_0_/X
+ mux_top_ipin_2.mux_l3_in_0_/S mux_top_ipin_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_2.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_2.mux_l1_in_2_/X mux_top_ipin_2.mux_l2_in_1_/S
+ mux_top_ipin_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_60_ gfpga_pad_EMBEDDED_IO_SOC_IN[0] top_width_0_height_0__pin_1_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xclkbuf_2_0_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_2.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_2.mux_l1_in_2_/S
+ mux_top_ipin_2.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_43_ chanx_left_in[1] chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26_ chanx_left_in[18] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09_ _09_/HI _09_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_2.mux_l2_in_0_ mux_top_ipin_2.mux_l1_in_1_/X mux_top_ipin_2.mux_l1_in_0_/X
+ mux_top_ipin_2.mux_l2_in_1_/S mux_top_ipin_2.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_2.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_2.mux_l1_in_2_/S
+ mux_top_ipin_2.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_1.mux_l3_in_0_/S mux_top_ipin_1.mux_l4_in_0_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_42_ chanx_left_in[2] chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25_ chanx_left_in[19] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08_ _08_/HI _08_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_4.mux_l3_in_0_/S mux_top_ipin_4.mux_l4_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_1.mux_l2_in_1_/S mux_top_ipin_1.mux_l3_in_0_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_2.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_2.mux_l1_in_2_/S
+ mux_top_ipin_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_41_ chanx_left_in[3] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_24_ chanx_right_in[0] chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_0.mux_l4_in_0_/X bottom_grid_pin_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_07_ _07_/HI _07_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_4.mux_l2_in_0_/S mux_top_ipin_4.mux_l3_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_1.mux_l1_in_2_/S mux_top_ipin_1.mux_l2_in_1_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_40_ chanx_left_in[4] chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mux_top_ipin_5.mux_l4_in_0_/S _50_/A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23_ chanx_right_in[1] chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06_ _06_/HI _06_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_4.mux_l1_in_1_/S mux_top_ipin_4.mux_l2_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_0.mux_l4_in_0_/S mux_top_ipin_1.mux_l1_in_2_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22_ chanx_right_in[2] chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_3.mux_l4_in_0_/S mux_top_ipin_4.mux_l1_in_1_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_3.mux_l2_in_3_ _09_/HI chanx_right_in[19] mux_top_ipin_3.mux_l2_in_2_/S
+ mux_top_ipin_3.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_21_ chanx_right_in[3] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_3.mux_l4_in_0_ mux_top_ipin_3.mux_l3_in_1_/X mux_top_ipin_3.mux_l3_in_0_/X
+ mux_top_ipin_3.mux_l4_in_0_/S mux_top_ipin_3.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_3.mux_l3_in_1_ mux_top_ipin_3.mux_l2_in_3_/X mux_top_ipin_3.mux_l2_in_2_/X
+ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_3.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[13] mux_top_ipin_3.mux_l2_in_2_/S
+ mux_top_ipin_3.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20_ chanx_right_in[4] chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_3.mux_l4_in_0_/X bottom_grid_pin_6_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_ipin_3.mux_l3_in_0_ mux_top_ipin_3.mux_l2_in_1_/X mux_top_ipin_3.mux_l2_in_0_/X
+ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_3.mux_l1_in_2_/X mux_top_ipin_3.mux_l2_in_2_/S
+ mux_top_ipin_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_3.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_3.mux_l1_in_0_/S
+ mux_top_ipin_3.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_3.mux_l2_in_0_ mux_top_ipin_3.mux_l1_in_1_/X mux_top_ipin_3.mux_l1_in_0_/X
+ mux_top_ipin_3.mux_l2_in_2_/S mux_top_ipin_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_78_ chanx_right_in[11] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_3.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_3.mux_l1_in_0_/S
+ mux_top_ipin_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_io_mode_io__4.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ _47_/A _46_/A ltile_io_mode_io__4.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_77_ chanx_right_in[12] chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_3.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_3.mux_l1_in_0_/S
+ mux_top_ipin_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_76_ chanx_right_in[13] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_59_ gfpga_pad_EMBEDDED_IO_SOC_IN[0] top_width_0_height_0__pin_1_lower VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_75_ chanx_right_in[14] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_58_ gfpga_pad_EMBEDDED_IO_SOC_IN[5] top_width_0_height_0__pin_11_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_74_ chanx_right_in[15] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_3_ _10_/HI chanx_right_in[14] mux_top_ipin_4.mux_l2_in_0_/S
+ mux_top_ipin_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_57_ gfpga_pad_EMBEDDED_IO_SOC_IN[5] top_width_0_height_0__pin_11_lower VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_4.mux_l4_in_0_ mux_top_ipin_4.mux_l3_in_1_/X mux_top_ipin_4.mux_l3_in_0_/X
+ mux_top_ipin_4.mux_l4_in_0_/S mux_top_ipin_4.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l4_in_0_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_4.mux_l3_in_1_ mux_top_ipin_4.mux_l2_in_3_/X mux_top_ipin_4.mux_l2_in_2_/X
+ mux_top_ipin_4.mux_l3_in_0_/S mux_top_ipin_4.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_73_ chanx_right_in[16] chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[8] mux_top_ipin_4.mux_l2_in_0_/S
+ mux_top_ipin_4.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_io_mode_io__1.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ _50_/A _49_/A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l4_in_0_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_56_ top_width_0_height_0__pin_0_ gfpga_pad_EMBEDDED_IO_SOC_OUT[0] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
XFILLER_16_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_39_ chanx_left_in[5] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_0.mux_l2_in_2_/S mux_top_ipin_0.mux_l3_in_1_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_4.mux_l3_in_0_ mux_top_ipin_4.mux_l2_in_1_/X mux_top_ipin_4.mux_l2_in_0_/X
+ mux_top_ipin_4.mux_l3_in_0_/S mux_top_ipin_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_72_ chanx_right_in[17] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_4.mux_l2_in_1_ chanx_left_in[8] mux_top_ipin_4.mux_l1_in_2_/X mux_top_ipin_4.mux_l2_in_0_/S
+ mux_top_ipin_4.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_55_ top_width_0_height_0__pin_2_ gfpga_pad_EMBEDDED_IO_SOC_OUT[1] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_3.mux_l2_in_2_/S mux_top_ipin_3.mux_l3_in_1_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_4.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_4.mux_l1_in_1_/S
+ mux_top_ipin_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_38_ chanx_left_in[6] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_0.mux_l1_in_0_/S mux_top_ipin_0.mux_l2_in_2_/S
+ clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_71_ chanx_right_in[18] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_0_ mux_top_ipin_4.mux_l1_in_1_/X mux_top_ipin_4.mux_l1_in_0_/X
+ mux_top_ipin_4.mux_l2_in_0_/S mux_top_ipin_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_54_ top_width_0_height_0__pin_4_ gfpga_pad_EMBEDDED_IO_SOC_OUT[2] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_3.mux_l1_in_0_/S mux_top_ipin_3.mux_l2_in_2_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_4.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_4.mux_l1_in_1_/S
+ mux_top_ipin_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_37_ chanx_left_in[7] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_top_ipin_0.mux_l1_in_0_/S
+ mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_70_ chanx_right_in[19] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_2.mux_l4_in_0_/S mux_top_ipin_3.mux_l1_in_0_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_53_ top_width_0_height_0__pin_6_ gfpga_pad_EMBEDDED_IO_SOC_OUT[3] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
XPHY_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_4.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_4.mux_l1_in_1_/S
+ mux_top_ipin_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36_ chanx_left_in[8] chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_19_ chanx_right_in[5] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_2.mux_l4_in_0_/X bottom_grid_pin_4_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_52_ top_width_0_height_0__pin_8_ gfpga_pad_EMBEDDED_IO_SOC_OUT[4] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
XPHY_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35_ chanx_left_in[9] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_18_ chanx_right_in[6] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_51_ top_width_0_height_0__pin_10_ gfpga_pad_EMBEDDED_IO_SOC_OUT[5] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34_ chanx_left_in[10] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17_ chanx_right_in[7] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_io_mode_io__5.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ _46_/A ccff_tail clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_0.mux_l2_in_3_ _06_/HI chanx_right_in[16] mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_0.mux_l4_in_0_ mux_top_ipin_0.mux_l3_in_1_/X mux_top_ipin_0.mux_l3_in_0_/X
+ mux_top_ipin_0.mux_l4_in_0_/S mux_top_ipin_0.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_50_ _50_/A gfpga_pad_EMBEDDED_IO_SOC_DIR[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_33_ chanx_left_in[11] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_3_ _11_/HI chanx_right_in[15] mux_top_ipin_5.mux_l2_in_3_/S
+ mux_top_ipin_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_0.mux_l3_in_1_ mux_top_ipin_0.mux_l2_in_3_/X mux_top_ipin_0.mux_l2_in_2_/X
+ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16_ chanx_right_in[8] chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_5.mux_l4_in_0_ mux_top_ipin_5.mux_l3_in_1_/X mux_top_ipin_5.mux_l3_in_0_/X
+ mux_top_ipin_5.mux_l4_in_0_/S mux_top_ipin_5.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_5.mux_l3_in_1_ mux_top_ipin_5.mux_l2_in_3_/X mux_top_ipin_5.mux_l2_in_2_/X
+ mux_top_ipin_5.mux_l3_in_1_/S mux_top_ipin_5.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32_ chanx_left_in[12] chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[9] mux_top_ipin_5.mux_l2_in_3_/S
+ mux_top_ipin_5.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.mux_l3_in_0_ mux_top_ipin_0.mux_l2_in_1_/X mux_top_ipin_0.mux_l2_in_0_/X
+ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15_ chanx_right_in[9] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_0.mux_l1_in_2_/X mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_0.mux_l1_in_0_/S
+ mux_top_ipin_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.mux_l3_in_0_ mux_top_ipin_5.mux_l2_in_1_/X mux_top_ipin_5.mux_l2_in_0_/X
+ mux_top_ipin_5.mux_l3_in_1_/S mux_top_ipin_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_5.mux_l4_in_0_/X bottom_grid_pin_10_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31_ chanx_left_in[13] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_1_ chanx_left_in[9] mux_top_ipin_5.mux_l1_in_2_/X mux_top_ipin_5.mux_l2_in_3_/S
+ mux_top_ipin_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14_ chanx_right_in[10] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_5.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_5.mux_l1_in_2_/S
+ mux_top_ipin_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.mux_l2_in_0_ mux_top_ipin_0.mux_l1_in_1_/X mux_top_ipin_0.mux_l1_in_0_/X
+ mux_top_ipin_0.mux_l2_in_2_/S mux_top_ipin_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_0.mux_l1_in_0_/S
+ mux_top_ipin_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_5.mux_l2_in_0_ mux_top_ipin_5.mux_l1_in_1_/X mux_top_ipin_5.mux_l1_in_0_/X
+ mux_top_ipin_5.mux_l2_in_3_/S mux_top_ipin_5.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_30_ chanx_left_in[14] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13_ _13_/HI SC_OUT_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_3_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_5.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_5.mux_l1_in_2_/S
+ mux_top_ipin_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_0.mux_l1_in_0_/S
+ mux_top_ipin_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12_ _12_/HI SC_OUT_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_io_mode_io__2.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ _49_/A _48_/A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_5.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_5.mux_l1_in_2_/S
+ mux_top_ipin_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11_ _11_/HI _11_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_1_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_2.mux_l3_in_0_/S mux_top_ipin_2.mux_l4_in_0_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10_ _10_/HI _10_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_5.mux_l3_in_1_/S mux_top_ipin_5.mux_l4_in_0_/S
+ clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_prog_clk clkbuf_1_1_0_prog_clk/X clkbuf_2_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_2.mux_l2_in_1_/S mux_top_ipin_2.mux_l3_in_0_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_1.mux_l2_in_3_ _07_/HI chanx_right_in[17] mux_top_ipin_1.mux_l2_in_1_/S
+ mux_top_ipin_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_1.mux_l4_in_0_ mux_top_ipin_1.mux_l3_in_1_/X mux_top_ipin_1.mux_l3_in_0_/X
+ mux_top_ipin_1.mux_l4_in_0_/S mux_top_ipin_1.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_69_ SC_IN_BOT SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_5.mux_l2_in_3_/S mux_top_ipin_5.mux_l3_in_1_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_1.mux_l3_in_1_ mux_top_ipin_1.mux_l2_in_3_/X mux_top_ipin_1.mux_l2_in_2_/X
+ mux_top_ipin_1.mux_l3_in_0_/S mux_top_ipin_1.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_2.mux_l1_in_2_/S mux_top_ipin_2.mux_l2_in_1_/S
+ clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_1.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_1.mux_l2_in_1_/S
+ mux_top_ipin_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_1.mux_l4_in_0_/X bottom_grid_pin_2_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_68_ gfpga_pad_EMBEDDED_IO_SOC_IN[4] top_width_0_height_0__pin_9_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_5.mux_l1_in_2_/S mux_top_ipin_5.mux_l2_in_3_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_1.mux_l3_in_0_ mux_top_ipin_1.mux_l2_in_1_/X mux_top_ipin_1.mux_l2_in_0_/X
+ mux_top_ipin_1.mux_l3_in_0_/S mux_top_ipin_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_1.mux_l4_in_0_/S mux_top_ipin_2.mux_l1_in_2_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_1.mux_l1_in_2_/X mux_top_ipin_1.mux_l2_in_1_/S
+ mux_top_ipin_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_1.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_1.mux_l1_in_2_/S
+ mux_top_ipin_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_67_ gfpga_pad_EMBEDDED_IO_SOC_IN[4] top_width_0_height_0__pin_9_lower VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_4.mux_l4_in_0_/S mux_top_ipin_5.mux_l1_in_2_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_2_0_prog_clk clkbuf_1_1_0_prog_clk/X clkbuf_2_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_1.mux_l2_in_0_ mux_top_ipin_1.mux_l1_in_1_/X mux_top_ipin_1.mux_l1_in_0_/X
+ mux_top_ipin_1.mux_l2_in_1_/S mux_top_ipin_1.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

