magic
tech sky130A
magscale 1 2
timestamp 1605004653
<< locali >>
rect 2789 13855 2823 13957
rect 14933 6647 14967 6885
rect 2421 6103 2455 6205
rect 2973 3927 3007 4097
<< viali >>
rect 1593 25449 1627 25483
rect 1593 24905 1627 24939
rect 1409 24701 1443 24735
rect 2053 24565 2087 24599
rect 1593 24361 1627 24395
rect 2697 24361 2731 24395
rect 1409 24225 1443 24259
rect 2513 24225 2547 24259
rect 2053 24089 2087 24123
rect 2513 23817 2547 23851
rect 3249 23817 3283 23851
rect 24777 23817 24811 23851
rect 2053 23681 2087 23715
rect 3709 23681 3743 23715
rect 1777 23613 1811 23647
rect 3065 23613 3099 23647
rect 1685 23477 1719 23511
rect 2053 23205 2087 23239
rect 12725 23205 12759 23239
rect 1777 23137 1811 23171
rect 12449 23137 12483 23171
rect 3249 22729 3283 22763
rect 1961 22593 1995 22627
rect 1685 22525 1719 22559
rect 1777 22525 1811 22559
rect 3065 22525 3099 22559
rect 2605 22389 2639 22423
rect 3709 22389 3743 22423
rect 12725 22389 12759 22423
rect 1409 22049 1443 22083
rect 2513 22049 2547 22083
rect 2697 21913 2731 21947
rect 1593 21845 1627 21879
rect 1593 21641 1627 21675
rect 8585 21641 8619 21675
rect 2697 21573 2731 21607
rect 7297 21505 7331 21539
rect 1409 21437 1443 21471
rect 2513 21437 2547 21471
rect 3065 21437 3099 21471
rect 7113 21437 7147 21471
rect 8401 21437 8435 21471
rect 8953 21437 8987 21471
rect 2421 21369 2455 21403
rect 2053 21301 2087 21335
rect 7849 21301 7883 21335
rect 1777 20961 1811 20995
rect 7941 20961 7975 20995
rect 1685 20893 1719 20927
rect 2053 20893 2087 20927
rect 8125 20893 8159 20927
rect 2605 20553 2639 20587
rect 4353 20553 4387 20587
rect 2053 20417 2087 20451
rect 8769 20417 8803 20451
rect 1777 20349 1811 20383
rect 3065 20349 3099 20383
rect 3617 20349 3651 20383
rect 4169 20349 4203 20383
rect 4721 20349 4755 20383
rect 8585 20349 8619 20383
rect 1685 20213 1719 20247
rect 3249 20213 3283 20247
rect 7941 20213 7975 20247
rect 9413 20213 9447 20247
rect 4261 20009 4295 20043
rect 1869 19941 1903 19975
rect 7941 19941 7975 19975
rect 1593 19873 1627 19907
rect 2881 19873 2915 19907
rect 4077 19873 4111 19907
rect 7665 19873 7699 19907
rect 5181 19805 5215 19839
rect 3065 19669 3099 19703
rect 6929 19669 6963 19703
rect 4077 19465 4111 19499
rect 3341 19329 3375 19363
rect 7389 19329 7423 19363
rect 1869 19261 1903 19295
rect 2145 19261 2179 19295
rect 3157 19261 3191 19295
rect 4445 19261 4479 19295
rect 4997 19261 5031 19295
rect 7297 19261 7331 19295
rect 5733 19193 5767 19227
rect 6561 19193 6595 19227
rect 7205 19193 7239 19227
rect 1685 19125 1719 19159
rect 2697 19125 2731 19159
rect 3065 19125 3099 19159
rect 4629 19125 4663 19159
rect 6285 19125 6319 19159
rect 6837 19125 6871 19159
rect 7849 19125 7883 19159
rect 10977 19125 11011 19159
rect 2789 18921 2823 18955
rect 5610 18853 5644 18887
rect 10670 18853 10704 18887
rect 1593 18785 1627 18819
rect 2881 18785 2915 18819
rect 4077 18785 4111 18819
rect 1869 18717 1903 18751
rect 5365 18717 5399 18751
rect 8585 18717 8619 18751
rect 10425 18717 10459 18751
rect 3433 18649 3467 18683
rect 4261 18649 4295 18683
rect 2329 18581 2363 18615
rect 3065 18581 3099 18615
rect 3893 18581 3927 18615
rect 4629 18581 4663 18615
rect 6745 18581 6779 18615
rect 7757 18581 7791 18615
rect 9321 18581 9355 18615
rect 11805 18581 11839 18615
rect 12541 18581 12575 18615
rect 3709 18377 3743 18411
rect 7665 18377 7699 18411
rect 12173 18377 12207 18411
rect 10609 18309 10643 18343
rect 11161 18309 11195 18343
rect 1777 18241 1811 18275
rect 2329 18241 2363 18275
rect 3065 18241 3099 18275
rect 8217 18241 8251 18275
rect 13001 18241 13035 18275
rect 1501 18173 1535 18207
rect 2789 18173 2823 18207
rect 4261 18173 4295 18207
rect 7573 18173 7607 18207
rect 8033 18173 8067 18207
rect 9229 18173 9263 18207
rect 12817 18173 12851 18207
rect 4169 18105 4203 18139
rect 4506 18105 4540 18139
rect 9137 18105 9171 18139
rect 9474 18105 9508 18139
rect 12909 18105 12943 18139
rect 2697 18037 2731 18071
rect 5641 18037 5675 18071
rect 6193 18037 6227 18071
rect 7205 18037 7239 18071
rect 8125 18037 8159 18071
rect 11805 18037 11839 18071
rect 12449 18037 12483 18071
rect 2145 17833 2179 17867
rect 7665 17833 7699 17867
rect 9689 17833 9723 17867
rect 12725 17833 12759 17867
rect 6552 17765 6586 17799
rect 11612 17765 11646 17799
rect 2237 17697 2271 17731
rect 3249 17697 3283 17731
rect 4813 17697 4847 17731
rect 4905 17697 4939 17731
rect 10057 17697 10091 17731
rect 1685 17629 1719 17663
rect 2329 17629 2363 17663
rect 4997 17629 5031 17663
rect 6285 17629 6319 17663
rect 10149 17629 10183 17663
rect 10241 17629 10275 17663
rect 10793 17629 10827 17663
rect 11345 17629 11379 17663
rect 5457 17561 5491 17595
rect 6101 17561 6135 17595
rect 9413 17561 9447 17595
rect 1777 17493 1811 17527
rect 2881 17493 2915 17527
rect 3617 17493 3651 17527
rect 4261 17493 4295 17527
rect 4445 17493 4479 17527
rect 4721 17289 4755 17323
rect 5641 17289 5675 17323
rect 6285 17289 6319 17323
rect 9229 17289 9263 17323
rect 10701 17289 10735 17323
rect 11437 17289 11471 17323
rect 12265 17289 12299 17323
rect 2789 17221 2823 17255
rect 2237 17153 2271 17187
rect 6837 17153 6871 17187
rect 9321 17153 9355 17187
rect 2053 17085 2087 17119
rect 3341 17085 3375 17119
rect 11805 17085 11839 17119
rect 12449 17085 12483 17119
rect 3586 17017 3620 17051
rect 6653 17017 6687 17051
rect 7104 17017 7138 17051
rect 9588 17017 9622 17051
rect 12694 17017 12728 17051
rect 1685 16949 1719 16983
rect 2145 16949 2179 16983
rect 3157 16949 3191 16983
rect 5365 16949 5399 16983
rect 8217 16949 8251 16983
rect 8769 16949 8803 16983
rect 13829 16949 13863 16983
rect 1869 16745 1903 16779
rect 2421 16745 2455 16779
rect 4077 16745 4111 16779
rect 4537 16745 4571 16779
rect 5181 16745 5215 16779
rect 5917 16745 5951 16779
rect 6469 16745 6503 16779
rect 7849 16745 7883 16779
rect 8033 16745 8067 16779
rect 10241 16745 10275 16779
rect 11161 16745 11195 16779
rect 1409 16677 1443 16711
rect 2329 16677 2363 16711
rect 3801 16677 3835 16711
rect 6377 16677 6411 16711
rect 8401 16677 8435 16711
rect 9689 16677 9723 16711
rect 10609 16677 10643 16711
rect 2789 16609 2823 16643
rect 2881 16609 2915 16643
rect 3433 16609 3467 16643
rect 4445 16609 4479 16643
rect 5549 16609 5583 16643
rect 6837 16609 6871 16643
rect 8493 16609 8527 16643
rect 11529 16609 11563 16643
rect 2973 16541 3007 16575
rect 4721 16541 4755 16575
rect 6929 16541 6963 16575
rect 7021 16541 7055 16575
rect 8677 16541 8711 16575
rect 11621 16541 11655 16575
rect 11805 16541 11839 16575
rect 7481 16405 7515 16439
rect 9413 16405 9447 16439
rect 12541 16405 12575 16439
rect 2421 16201 2455 16235
rect 4629 16201 4663 16235
rect 5089 16201 5123 16235
rect 6837 16201 6871 16235
rect 8309 16201 8343 16235
rect 8677 16201 8711 16235
rect 10609 16201 10643 16235
rect 11529 16201 11563 16235
rect 11897 16201 11931 16235
rect 7297 16065 7331 16099
rect 7481 16065 7515 16099
rect 9229 16065 9263 16099
rect 1409 15997 1443 16031
rect 2697 15997 2731 16031
rect 5181 15997 5215 16031
rect 1685 15929 1719 15963
rect 2964 15929 2998 15963
rect 5457 15929 5491 15963
rect 7205 15929 7239 15963
rect 7849 15929 7883 15963
rect 9137 15929 9171 15963
rect 9474 15929 9508 15963
rect 4077 15861 4111 15895
rect 6101 15861 6135 15895
rect 6561 15861 6595 15895
rect 11253 15861 11287 15895
rect 12449 15861 12483 15895
rect 1409 15657 1443 15691
rect 2329 15657 2363 15691
rect 2421 15657 2455 15691
rect 3893 15657 3927 15691
rect 6561 15657 6595 15691
rect 7113 15657 7147 15691
rect 8217 15657 8251 15691
rect 9689 15657 9723 15691
rect 11621 15657 11655 15691
rect 11989 15657 12023 15691
rect 12725 15657 12759 15691
rect 4322 15589 4356 15623
rect 2789 15521 2823 15555
rect 6193 15521 6227 15555
rect 7021 15521 7055 15555
rect 7481 15521 7515 15555
rect 10057 15521 10091 15555
rect 11437 15521 11471 15555
rect 2881 15453 2915 15487
rect 3065 15453 3099 15487
rect 4077 15453 4111 15487
rect 7573 15453 7607 15487
rect 7757 15453 7791 15487
rect 10149 15453 10183 15487
rect 10241 15453 10275 15487
rect 12081 15453 12115 15487
rect 12265 15453 12299 15487
rect 1961 15317 1995 15351
rect 3525 15317 3559 15351
rect 5457 15317 5491 15351
rect 6837 15317 6871 15351
rect 8493 15317 8527 15351
rect 9045 15317 9079 15351
rect 9413 15317 9447 15351
rect 11253 15317 11287 15351
rect 13001 15317 13035 15351
rect 2697 15113 2731 15147
rect 3801 15113 3835 15147
rect 4169 15113 4203 15147
rect 5641 15113 5675 15147
rect 6285 15113 6319 15147
rect 8217 15113 8251 15147
rect 10701 15113 10735 15147
rect 11253 15113 11287 15147
rect 11713 15113 11747 15147
rect 1685 14977 1719 15011
rect 3341 14977 3375 15011
rect 4261 14977 4295 15011
rect 9229 14977 9263 15011
rect 1409 14909 1443 14943
rect 6837 14909 6871 14943
rect 9321 14909 9355 14943
rect 12449 14909 12483 14943
rect 12716 14909 12750 14943
rect 3157 14841 3191 14875
rect 4528 14841 4562 14875
rect 7104 14841 7138 14875
rect 9566 14841 9600 14875
rect 2513 14773 2547 14807
rect 3065 14773 3099 14807
rect 6653 14773 6687 14807
rect 8861 14773 8895 14807
rect 12081 14773 12115 14807
rect 13829 14773 13863 14807
rect 1501 14569 1535 14603
rect 4629 14569 4663 14603
rect 4905 14569 4939 14603
rect 6285 14569 6319 14603
rect 6653 14569 6687 14603
rect 8677 14569 8711 14603
rect 11161 14569 11195 14603
rect 11805 14569 11839 14603
rect 1961 14501 1995 14535
rect 2513 14501 2547 14535
rect 3249 14501 3283 14535
rect 7012 14501 7046 14535
rect 12716 14501 12750 14535
rect 1869 14433 1903 14467
rect 3617 14433 3651 14467
rect 5273 14433 5307 14467
rect 6745 14433 6779 14467
rect 9413 14433 9447 14467
rect 10048 14433 10082 14467
rect 12081 14433 12115 14467
rect 12449 14433 12483 14467
rect 2145 14365 2179 14399
rect 5365 14365 5399 14399
rect 5549 14365 5583 14399
rect 9137 14365 9171 14399
rect 9781 14365 9815 14399
rect 4353 14297 4387 14331
rect 9229 14297 9263 14331
rect 2881 14229 2915 14263
rect 8125 14229 8159 14263
rect 13829 14229 13863 14263
rect 1869 14025 1903 14059
rect 3249 14025 3283 14059
rect 4261 14025 4295 14059
rect 6561 14025 6595 14059
rect 7021 14025 7055 14059
rect 7481 14025 7515 14059
rect 7941 14025 7975 14059
rect 10885 14025 10919 14059
rect 12449 14025 12483 14059
rect 13461 14025 13495 14059
rect 2789 13957 2823 13991
rect 2973 13957 3007 13991
rect 11897 13957 11931 13991
rect 24225 13957 24259 13991
rect 1777 13889 1811 13923
rect 2329 13889 2363 13923
rect 2513 13889 2547 13923
rect 3617 13889 3651 13923
rect 4169 13889 4203 13923
rect 4905 13889 4939 13923
rect 5733 13889 5767 13923
rect 8493 13889 8527 13923
rect 8953 13889 8987 13923
rect 9413 13889 9447 13923
rect 9965 13889 9999 13923
rect 10149 13889 10183 13923
rect 13001 13889 13035 13923
rect 2789 13821 2823 13855
rect 5365 13821 5399 13855
rect 6837 13821 6871 13855
rect 7849 13821 7883 13855
rect 12265 13821 12299 13855
rect 12909 13821 12943 13855
rect 24041 13821 24075 13855
rect 24593 13821 24627 13855
rect 2237 13753 2271 13787
rect 8401 13753 8435 13787
rect 9873 13753 9907 13787
rect 12817 13753 12851 13787
rect 4629 13685 4663 13719
rect 4721 13685 4755 13719
rect 6101 13685 6135 13719
rect 8309 13685 8343 13719
rect 9505 13685 9539 13719
rect 10609 13685 10643 13719
rect 11069 13685 11103 13719
rect 14013 13685 14047 13719
rect 2881 13481 2915 13515
rect 4353 13481 4387 13515
rect 6193 13481 6227 13515
rect 7297 13481 7331 13515
rect 8401 13481 8435 13515
rect 8769 13481 8803 13515
rect 9965 13481 9999 13515
rect 11437 13481 11471 13515
rect 12449 13481 12483 13515
rect 12817 13481 12851 13515
rect 13369 13481 13403 13515
rect 1768 13413 1802 13447
rect 3801 13413 3835 13447
rect 3525 13345 3559 13379
rect 5080 13345 5114 13379
rect 7665 13345 7699 13379
rect 10324 13345 10358 13379
rect 13737 13345 13771 13379
rect 15568 13345 15602 13379
rect 23397 13345 23431 13379
rect 1501 13277 1535 13311
rect 4813 13277 4847 13311
rect 7757 13277 7791 13311
rect 7941 13277 7975 13311
rect 10057 13277 10091 13311
rect 13829 13277 13863 13311
rect 14013 13277 14047 13311
rect 15301 13277 15335 13311
rect 16681 13209 16715 13243
rect 4629 13141 4663 13175
rect 6929 13141 6963 13175
rect 9045 13141 9079 13175
rect 9505 13141 9539 13175
rect 13185 13141 13219 13175
rect 23581 13141 23615 13175
rect 1869 12937 1903 12971
rect 3249 12937 3283 12971
rect 6837 12937 6871 12971
rect 8217 12937 8251 12971
rect 9413 12937 9447 12971
rect 11897 12937 11931 12971
rect 12909 12937 12943 12971
rect 13277 12937 13311 12971
rect 15669 12937 15703 12971
rect 23397 12937 23431 12971
rect 4813 12869 4847 12903
rect 23857 12869 23891 12903
rect 2513 12801 2547 12835
rect 6561 12801 6595 12835
rect 7389 12801 7423 12835
rect 9321 12801 9355 12835
rect 10057 12801 10091 12835
rect 3433 12733 3467 12767
rect 3689 12733 3723 12767
rect 9781 12733 9815 12767
rect 13369 12733 13403 12767
rect 23673 12733 23707 12767
rect 24225 12733 24259 12767
rect 2237 12665 2271 12699
rect 2973 12665 3007 12699
rect 5733 12665 5767 12699
rect 6285 12665 6319 12699
rect 7205 12665 7239 12699
rect 10517 12665 10551 12699
rect 13636 12665 13670 12699
rect 15393 12665 15427 12699
rect 1777 12597 1811 12631
rect 2329 12597 2363 12631
rect 5457 12597 5491 12631
rect 7297 12597 7331 12631
rect 7849 12597 7883 12631
rect 8401 12597 8435 12631
rect 8861 12597 8895 12631
rect 9873 12597 9907 12631
rect 10793 12597 10827 12631
rect 11161 12597 11195 12631
rect 11345 12597 11379 12631
rect 14749 12597 14783 12631
rect 2881 12393 2915 12427
rect 3433 12393 3467 12427
rect 6009 12393 6043 12427
rect 7113 12393 7147 12427
rect 11713 12393 11747 12427
rect 12817 12393 12851 12427
rect 4896 12325 4930 12359
rect 12265 12325 12299 12359
rect 1768 12257 1802 12291
rect 4629 12257 4663 12291
rect 7481 12257 7515 12291
rect 8861 12257 8895 12291
rect 10600 12257 10634 12291
rect 13185 12257 13219 12291
rect 13921 12257 13955 12291
rect 15669 12257 15703 12291
rect 22293 12257 22327 12291
rect 1501 12189 1535 12223
rect 7573 12189 7607 12223
rect 7665 12189 7699 12223
rect 10333 12189 10367 12223
rect 12725 12189 12759 12223
rect 13277 12189 13311 12223
rect 13369 12189 13403 12223
rect 15761 12189 15795 12223
rect 15853 12189 15887 12223
rect 6929 12121 6963 12155
rect 8217 12121 8251 12155
rect 8585 12121 8619 12155
rect 9873 12121 9907 12155
rect 14289 12121 14323 12155
rect 15301 12121 15335 12155
rect 3893 12053 3927 12087
rect 4353 12053 4387 12087
rect 8677 12053 8711 12087
rect 9505 12053 9539 12087
rect 22477 12053 22511 12087
rect 2605 11849 2639 11883
rect 2973 11849 3007 11883
rect 4905 11849 4939 11883
rect 5549 11849 5583 11883
rect 6377 11849 6411 11883
rect 12173 11849 12207 11883
rect 14105 11849 14139 11883
rect 15209 11849 15243 11883
rect 22293 11849 22327 11883
rect 6469 11781 6503 11815
rect 2145 11713 2179 11747
rect 4353 11713 4387 11747
rect 5273 11713 5307 11747
rect 9689 11713 9723 11747
rect 11897 11713 11931 11747
rect 15761 11713 15795 11747
rect 16221 11713 16255 11747
rect 1961 11645 1995 11679
rect 4169 11645 4203 11679
rect 5365 11645 5399 11679
rect 5917 11645 5951 11679
rect 6653 11645 6687 11679
rect 6837 11645 6871 11679
rect 9597 11645 9631 11679
rect 12725 11645 12759 11679
rect 12992 11645 13026 11679
rect 15577 11645 15611 11679
rect 3709 11577 3743 11611
rect 7104 11577 7138 11611
rect 8769 11577 8803 11611
rect 9321 11577 9355 11611
rect 9956 11577 9990 11611
rect 15025 11577 15059 11611
rect 1593 11509 1627 11543
rect 2053 11509 2087 11543
rect 3801 11509 3835 11543
rect 4261 11509 4295 11543
rect 8217 11509 8251 11543
rect 9413 11509 9447 11543
rect 11069 11509 11103 11543
rect 14657 11509 14691 11543
rect 15669 11509 15703 11543
rect 16589 11509 16623 11543
rect 1409 11305 1443 11339
rect 1961 11305 1995 11339
rect 2421 11305 2455 11339
rect 3433 11305 3467 11339
rect 4537 11305 4571 11339
rect 5825 11305 5859 11339
rect 9689 11305 9723 11339
rect 11069 11305 11103 11339
rect 11253 11305 11287 11339
rect 12817 11305 12851 11339
rect 14013 11305 14047 11339
rect 14473 11305 14507 11339
rect 15577 11305 15611 11339
rect 15853 11305 15887 11339
rect 3893 11237 3927 11271
rect 6929 11237 6963 11271
rect 7380 11237 7414 11271
rect 12725 11237 12759 11271
rect 2789 11169 2823 11203
rect 4445 11169 4479 11203
rect 5641 11169 5675 11203
rect 10057 11169 10091 11203
rect 11621 11169 11655 11203
rect 13185 11169 13219 11203
rect 2881 11101 2915 11135
rect 2973 11101 3007 11135
rect 4629 11101 4663 11135
rect 7113 11101 7147 11135
rect 10149 11101 10183 11135
rect 10333 11101 10367 11135
rect 11713 11101 11747 11135
rect 11805 11101 11839 11135
rect 13277 11101 13311 11135
rect 13461 11101 13495 11135
rect 4077 11033 4111 11067
rect 6561 11033 6595 11067
rect 9045 11033 9079 11067
rect 9505 11033 9539 11067
rect 10793 11033 10827 11067
rect 12357 11033 12391 11067
rect 13921 11033 13955 11067
rect 2237 10965 2271 10999
rect 5089 10965 5123 10999
rect 5457 10965 5491 10999
rect 8493 10965 8527 10999
rect 1685 10761 1719 10795
rect 3157 10761 3191 10795
rect 3709 10761 3743 10795
rect 5641 10761 5675 10795
rect 6929 10761 6963 10795
rect 9873 10761 9907 10795
rect 10425 10761 10459 10795
rect 10793 10761 10827 10795
rect 11805 10761 11839 10795
rect 4261 10693 4295 10727
rect 4905 10625 4939 10659
rect 6653 10625 6687 10659
rect 7481 10625 7515 10659
rect 10977 10625 11011 10659
rect 1777 10557 1811 10591
rect 4721 10557 4755 10591
rect 8493 10557 8527 10591
rect 13185 10557 13219 10591
rect 2044 10489 2078 10523
rect 7389 10489 7423 10523
rect 8033 10489 8067 10523
rect 8401 10489 8435 10523
rect 8760 10489 8794 10523
rect 12173 10489 12207 10523
rect 4169 10421 4203 10455
rect 4629 10421 4663 10455
rect 5365 10421 5399 10455
rect 6285 10421 6319 10455
rect 7297 10421 7331 10455
rect 11437 10421 11471 10455
rect 12909 10421 12943 10455
rect 14473 10421 14507 10455
rect 2789 10217 2823 10251
rect 4077 10217 4111 10251
rect 6009 10217 6043 10251
rect 7941 10217 7975 10251
rect 8401 10217 8435 10251
rect 9689 10217 9723 10251
rect 10057 10217 10091 10251
rect 11161 10217 11195 10251
rect 11253 10217 11287 10251
rect 12449 10217 12483 10251
rect 13277 10217 13311 10251
rect 8309 10149 8343 10183
rect 11713 10149 11747 10183
rect 13737 10149 13771 10183
rect 1676 10081 1710 10115
rect 3893 10081 3927 10115
rect 4445 10081 4479 10115
rect 11621 10081 11655 10115
rect 12817 10081 12851 10115
rect 12909 10081 12943 10115
rect 13645 10081 13679 10115
rect 1409 10013 1443 10047
rect 4537 10013 4571 10047
rect 4629 10013 4663 10047
rect 5181 10013 5215 10047
rect 5549 10013 5583 10047
rect 6101 10013 6135 10047
rect 6193 10013 6227 10047
rect 8585 10013 8619 10047
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 11897 10013 11931 10047
rect 13001 10013 13035 10047
rect 13829 10013 13863 10047
rect 15301 10013 15335 10047
rect 3433 9945 3467 9979
rect 5641 9945 5675 9979
rect 7389 9945 7423 9979
rect 7665 9945 7699 9979
rect 9137 9945 9171 9979
rect 9505 9945 9539 9979
rect 6929 9877 6963 9911
rect 10701 9877 10735 9911
rect 12357 9877 12391 9911
rect 14289 9877 14323 9911
rect 14657 9877 14691 9911
rect 1685 9673 1719 9707
rect 2053 9673 2087 9707
rect 5181 9673 5215 9707
rect 5825 9673 5859 9707
rect 8769 9673 8803 9707
rect 11161 9673 11195 9707
rect 3341 9605 3375 9639
rect 9505 9605 9539 9639
rect 10517 9605 10551 9639
rect 13829 9605 13863 9639
rect 14749 9605 14783 9639
rect 15393 9605 15427 9639
rect 2881 9537 2915 9571
rect 6653 9537 6687 9571
rect 10149 9537 10183 9571
rect 2605 9469 2639 9503
rect 3801 9469 3835 9503
rect 6837 9469 6871 9503
rect 7104 9469 7138 9503
rect 9873 9469 9907 9503
rect 12449 9469 12483 9503
rect 4068 9401 4102 9435
rect 9413 9401 9447 9435
rect 9965 9401 9999 9435
rect 12694 9401 12728 9435
rect 2237 9333 2271 9367
rect 2697 9333 2731 9367
rect 3709 9333 3743 9367
rect 6101 9333 6135 9367
rect 8217 9333 8251 9367
rect 11345 9333 11379 9367
rect 11805 9333 11839 9367
rect 12173 9333 12207 9367
rect 14381 9333 14415 9367
rect 14933 9333 14967 9367
rect 1869 9129 1903 9163
rect 3893 9129 3927 9163
rect 4077 9129 4111 9163
rect 4537 9129 4571 9163
rect 5641 9129 5675 9163
rect 8309 9129 8343 9163
rect 8861 9129 8895 9163
rect 9505 9129 9539 9163
rect 9965 9129 9999 9163
rect 11713 9129 11747 9163
rect 13185 9129 13219 9163
rect 14105 9129 14139 9163
rect 2329 9061 2363 9095
rect 5089 9061 5123 9095
rect 8033 9061 8067 9095
rect 11345 9061 11379 9095
rect 13829 9061 13863 9095
rect 2237 8993 2271 9027
rect 3341 8993 3375 9027
rect 4445 8993 4479 9027
rect 5825 8993 5859 9027
rect 6092 8993 6126 9027
rect 10609 8993 10643 9027
rect 12072 8993 12106 9027
rect 15393 8993 15427 9027
rect 15660 8993 15694 9027
rect 1777 8925 1811 8959
rect 2421 8925 2455 8959
rect 4721 8925 4755 8959
rect 10701 8925 10735 8959
rect 10885 8925 10919 8959
rect 11805 8925 11839 8959
rect 2881 8857 2915 8891
rect 14473 8857 14507 8891
rect 7205 8789 7239 8823
rect 10241 8789 10275 8823
rect 14841 8789 14875 8823
rect 16773 8789 16807 8823
rect 2605 8585 2639 8619
rect 4169 8585 4203 8619
rect 4721 8585 4755 8619
rect 5181 8585 5215 8619
rect 5641 8585 5675 8619
rect 7941 8585 7975 8619
rect 10057 8585 10091 8619
rect 10701 8585 10735 8619
rect 12173 8585 12207 8619
rect 17141 8585 17175 8619
rect 6837 8517 6871 8551
rect 8401 8517 8435 8551
rect 10977 8517 11011 8551
rect 12449 8517 12483 8551
rect 13553 8517 13587 8551
rect 15853 8517 15887 8551
rect 1685 8449 1719 8483
rect 6653 8449 6687 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 11897 8449 11931 8483
rect 13001 8449 13035 8483
rect 14013 8449 14047 8483
rect 15117 8449 15151 8483
rect 16313 8449 16347 8483
rect 1409 8381 1443 8415
rect 2789 8381 2823 8415
rect 8585 8381 8619 8415
rect 8677 8381 8711 8415
rect 12909 8381 12943 8415
rect 14841 8381 14875 8415
rect 16037 8381 16071 8415
rect 16773 8381 16807 8415
rect 20913 8381 20947 8415
rect 21649 8381 21683 8415
rect 3034 8313 3068 8347
rect 5733 8313 5767 8347
rect 6285 8313 6319 8347
rect 7205 8313 7239 8347
rect 8309 8313 8343 8347
rect 8922 8313 8956 8347
rect 12817 8313 12851 8347
rect 14289 8313 14323 8347
rect 14933 8313 14967 8347
rect 15577 8313 15611 8347
rect 21189 8313 21223 8347
rect 2145 8245 2179 8279
rect 11345 8245 11379 8279
rect 14473 8245 14507 8279
rect 1409 8041 1443 8075
rect 2421 8041 2455 8075
rect 2789 8041 2823 8075
rect 3893 8041 3927 8075
rect 5089 8041 5123 8075
rect 6653 8041 6687 8075
rect 7849 8041 7883 8075
rect 8217 8041 8251 8075
rect 8861 8041 8895 8075
rect 9505 8041 9539 8075
rect 10333 8041 10367 8075
rect 4353 7973 4387 8007
rect 5733 7973 5767 8007
rect 10241 7973 10275 8007
rect 5181 7905 5215 7939
rect 8309 7905 8343 7939
rect 10977 7905 11011 7939
rect 11704 7905 11738 7939
rect 15568 7905 15602 7939
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 5273 7837 5307 7871
rect 6745 7837 6779 7871
rect 6929 7837 6963 7871
rect 8401 7837 8435 7871
rect 10517 7837 10551 7871
rect 11437 7837 11471 7871
rect 14197 7837 14231 7871
rect 15301 7837 15335 7871
rect 2237 7769 2271 7803
rect 6193 7769 6227 7803
rect 7757 7769 7791 7803
rect 9873 7769 9907 7803
rect 11253 7769 11287 7803
rect 12817 7769 12851 7803
rect 1869 7701 1903 7735
rect 3433 7701 3467 7735
rect 4721 7701 4755 7735
rect 6285 7701 6319 7735
rect 7389 7701 7423 7735
rect 13461 7701 13495 7735
rect 13829 7701 13863 7735
rect 14657 7701 14691 7735
rect 15025 7701 15059 7735
rect 16681 7701 16715 7735
rect 1409 7497 1443 7531
rect 4997 7497 5031 7531
rect 6377 7497 6411 7531
rect 7021 7497 7055 7531
rect 7481 7497 7515 7531
rect 9965 7497 9999 7531
rect 10241 7497 10275 7531
rect 12173 7497 12207 7531
rect 12725 7497 12759 7531
rect 14473 7497 14507 7531
rect 17233 7497 17267 7531
rect 17601 7497 17635 7531
rect 2881 7429 2915 7463
rect 4353 7429 4387 7463
rect 5457 7429 5491 7463
rect 10517 7429 10551 7463
rect 2053 7361 2087 7395
rect 11253 7361 11287 7395
rect 11437 7361 11471 7395
rect 13921 7361 13955 7395
rect 2973 7293 3007 7327
rect 5641 7293 5675 7327
rect 7665 7293 7699 7327
rect 7921 7293 7955 7327
rect 10701 7293 10735 7327
rect 11161 7293 11195 7327
rect 13737 7293 13771 7327
rect 14933 7293 14967 7327
rect 18061 7293 18095 7327
rect 18797 7293 18831 7327
rect 1777 7225 1811 7259
rect 3218 7225 3252 7259
rect 5365 7225 5399 7259
rect 13829 7225 13863 7259
rect 14841 7225 14875 7259
rect 15200 7225 15234 7259
rect 18337 7225 18371 7259
rect 1869 7157 1903 7191
rect 2513 7157 2547 7191
rect 5733 7157 5767 7191
rect 9045 7157 9079 7191
rect 10793 7157 10827 7191
rect 11897 7157 11931 7191
rect 13185 7157 13219 7191
rect 13369 7157 13403 7191
rect 16313 7157 16347 7191
rect 16865 7157 16899 7191
rect 3433 6953 3467 6987
rect 6377 6953 6411 6987
rect 13369 6953 13403 6987
rect 15761 6953 15795 6987
rect 17233 6953 17267 6987
rect 19165 6953 19199 6987
rect 5273 6885 5307 6919
rect 10057 6885 10091 6919
rect 14933 6885 14967 6919
rect 15025 6885 15059 6919
rect 1768 6817 1802 6851
rect 6469 6817 6503 6851
rect 6736 6817 6770 6851
rect 8401 6817 8435 6851
rect 9505 6817 9539 6851
rect 10885 6817 10919 6851
rect 11520 6817 11554 6851
rect 13921 6817 13955 6851
rect 1501 6749 1535 6783
rect 5365 6749 5399 6783
rect 5457 6749 5491 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 11253 6749 11287 6783
rect 14197 6749 14231 6783
rect 2881 6681 2915 6715
rect 12633 6681 12667 6715
rect 15853 6817 15887 6851
rect 18052 6817 18086 6851
rect 20913 6817 20947 6851
rect 16037 6749 16071 6783
rect 17785 6749 17819 6783
rect 21189 6749 21223 6783
rect 15393 6681 15427 6715
rect 3801 6613 3835 6647
rect 4261 6613 4295 6647
rect 4721 6613 4755 6647
rect 4905 6613 4939 6647
rect 6009 6613 6043 6647
rect 7849 6613 7883 6647
rect 8861 6613 8895 6647
rect 9689 6613 9723 6647
rect 13829 6613 13863 6647
rect 14657 6613 14691 6647
rect 14933 6613 14967 6647
rect 16405 6613 16439 6647
rect 16773 6613 16807 6647
rect 17601 6613 17635 6647
rect 2697 6409 2731 6443
rect 5733 6409 5767 6443
rect 7941 6409 7975 6443
rect 10517 6409 10551 6443
rect 11805 6409 11839 6443
rect 14197 6409 14231 6443
rect 16681 6409 16715 6443
rect 19073 6409 19107 6443
rect 20913 6409 20947 6443
rect 4721 6341 4755 6375
rect 10885 6341 10919 6375
rect 12449 6341 12483 6375
rect 16313 6341 16347 6375
rect 17049 6341 17083 6375
rect 2145 6273 2179 6307
rect 3065 6273 3099 6307
rect 3709 6273 3743 6307
rect 5365 6273 5399 6307
rect 6101 6273 6135 6307
rect 7297 6273 7331 6307
rect 7481 6273 7515 6307
rect 8493 6273 8527 6307
rect 13001 6273 13035 6307
rect 13461 6273 13495 6307
rect 14381 6273 14415 6307
rect 18705 6273 18739 6307
rect 19441 6273 19475 6307
rect 1961 6205 1995 6239
rect 2421 6205 2455 6239
rect 3525 6205 3559 6239
rect 5089 6205 5123 6239
rect 7205 6205 7239 6239
rect 8585 6205 8619 6239
rect 8852 6205 8886 6239
rect 14637 6205 14671 6239
rect 16865 6205 16899 6239
rect 17785 6205 17819 6239
rect 18521 6205 18555 6239
rect 3617 6137 3651 6171
rect 4261 6137 4295 6171
rect 6653 6137 6687 6171
rect 12909 6137 12943 6171
rect 13829 6137 13863 6171
rect 17509 6137 17543 6171
rect 18429 6137 18463 6171
rect 19625 6137 19659 6171
rect 1593 6069 1627 6103
rect 2053 6069 2087 6103
rect 2421 6069 2455 6103
rect 3157 6069 3191 6103
rect 4537 6069 4571 6103
rect 5181 6069 5215 6103
rect 6837 6069 6871 6103
rect 9965 6069 9999 6103
rect 11345 6069 11379 6103
rect 12173 6069 12207 6103
rect 12817 6069 12851 6103
rect 15761 6069 15795 6103
rect 18061 6069 18095 6103
rect 2145 5865 2179 5899
rect 3157 5865 3191 5899
rect 4537 5865 4571 5899
rect 6009 5865 6043 5899
rect 6561 5865 6595 5899
rect 7021 5865 7055 5899
rect 9965 5865 9999 5899
rect 10333 5865 10367 5899
rect 11805 5865 11839 5899
rect 14381 5865 14415 5899
rect 15669 5865 15703 5899
rect 15761 5865 15795 5899
rect 16313 5865 16347 5899
rect 18889 5865 18923 5899
rect 2513 5797 2547 5831
rect 3525 5797 3559 5831
rect 7380 5797 7414 5831
rect 15025 5797 15059 5831
rect 17776 5797 17810 5831
rect 4629 5729 4663 5763
rect 4896 5729 4930 5763
rect 10701 5729 10735 5763
rect 12153 5729 12187 5763
rect 20913 5729 20947 5763
rect 2605 5661 2639 5695
rect 2697 5661 2731 5695
rect 7113 5661 7147 5695
rect 10793 5661 10827 5695
rect 10885 5661 10919 5695
rect 11897 5661 11931 5695
rect 13921 5661 13955 5695
rect 15853 5661 15887 5695
rect 17509 5661 17543 5695
rect 2053 5593 2087 5627
rect 8493 5593 8527 5627
rect 15301 5593 15335 5627
rect 16865 5593 16899 5627
rect 1593 5525 1627 5559
rect 9137 5525 9171 5559
rect 9413 5525 9447 5559
rect 11345 5525 11379 5559
rect 13277 5525 13311 5559
rect 17233 5525 17267 5559
rect 21097 5525 21131 5559
rect 4261 5321 4295 5355
rect 7481 5321 7515 5355
rect 10885 5321 10919 5355
rect 11437 5321 11471 5355
rect 11805 5321 11839 5355
rect 12633 5321 12667 5355
rect 14749 5321 14783 5355
rect 15301 5321 15335 5355
rect 16865 5321 16899 5355
rect 17509 5321 17543 5355
rect 17877 5321 17911 5355
rect 20913 5321 20947 5355
rect 9045 5253 9079 5287
rect 18061 5253 18095 5287
rect 1409 5185 1443 5219
rect 5733 5185 5767 5219
rect 8401 5185 8435 5219
rect 8493 5185 8527 5219
rect 15669 5185 15703 5219
rect 16405 5185 16439 5219
rect 18705 5185 18739 5219
rect 20085 5185 20119 5219
rect 2881 5117 2915 5151
rect 3148 5117 3182 5151
rect 4905 5117 4939 5151
rect 7849 5117 7883 5151
rect 9505 5117 9539 5151
rect 12173 5117 12207 5151
rect 13369 5117 13403 5151
rect 16221 5117 16255 5151
rect 16313 5117 16347 5151
rect 19809 5117 19843 5151
rect 20545 5117 20579 5151
rect 21097 5117 21131 5151
rect 5181 5049 5215 5083
rect 5549 5049 5583 5083
rect 6285 5049 6319 5083
rect 6561 5049 6595 5083
rect 8309 5049 8343 5083
rect 9772 5049 9806 5083
rect 13277 5049 13311 5083
rect 13636 5049 13670 5083
rect 18429 5049 18463 5083
rect 19441 5049 19475 5083
rect 2237 4981 2271 5015
rect 2605 4981 2639 5015
rect 6929 4981 6963 5015
rect 7941 4981 7975 5015
rect 9321 4981 9355 5015
rect 11989 4981 12023 5015
rect 15853 4981 15887 5015
rect 18521 4981 18555 5015
rect 19073 4981 19107 5015
rect 21281 4981 21315 5015
rect 21649 4981 21683 5015
rect 2881 4777 2915 4811
rect 3433 4777 3467 4811
rect 3801 4777 3835 4811
rect 5825 4777 5859 4811
rect 7573 4777 7607 4811
rect 8309 4777 8343 4811
rect 12633 4777 12667 4811
rect 13093 4777 13127 4811
rect 15025 4777 15059 4811
rect 15761 4777 15795 4811
rect 16405 4777 16439 4811
rect 18429 4777 18463 4811
rect 10854 4709 10888 4743
rect 13001 4709 13035 4743
rect 24216 4709 24250 4743
rect 1768 4641 1802 4675
rect 4629 4641 4663 4675
rect 4721 4641 4755 4675
rect 6193 4641 6227 4675
rect 7205 4641 7239 4675
rect 7849 4641 7883 4675
rect 8953 4641 8987 4675
rect 9321 4641 9355 4675
rect 10609 4641 10643 4675
rect 13461 4641 13495 4675
rect 14105 4641 14139 4675
rect 15669 4641 15703 4675
rect 17305 4641 17339 4675
rect 19533 4641 19567 4675
rect 20913 4641 20947 4675
rect 22017 4641 22051 4675
rect 1501 4573 1535 4607
rect 4813 4573 4847 4607
rect 6285 4573 6319 4607
rect 6377 4573 6411 4607
rect 8401 4573 8435 4607
rect 8585 4573 8619 4607
rect 13553 4573 13587 4607
rect 13645 4573 13679 4607
rect 15853 4573 15887 4607
rect 17049 4573 17083 4607
rect 19809 4573 19843 4607
rect 23949 4573 23983 4607
rect 7665 4505 7699 4539
rect 7941 4505 7975 4539
rect 9965 4505 9999 4539
rect 25329 4505 25363 4539
rect 4261 4437 4295 4471
rect 5273 4437 5307 4471
rect 5641 4437 5675 4471
rect 10425 4437 10459 4471
rect 11989 4437 12023 4471
rect 14565 4437 14599 4471
rect 15301 4437 15335 4471
rect 16773 4437 16807 4471
rect 19073 4437 19107 4471
rect 21097 4437 21131 4471
rect 22201 4437 22235 4471
rect 1685 4233 1719 4267
rect 4261 4233 4295 4267
rect 6561 4233 6595 4267
rect 10241 4233 10275 4267
rect 16405 4233 16439 4267
rect 18061 4233 18095 4267
rect 19073 4233 19107 4267
rect 20821 4233 20855 4267
rect 21833 4233 21867 4267
rect 24041 4233 24075 4267
rect 4629 4165 4663 4199
rect 7941 4165 7975 4199
rect 24317 4165 24351 4199
rect 2237 4097 2271 4131
rect 2973 4097 3007 4131
rect 3065 4097 3099 4131
rect 3249 4097 3283 4131
rect 5181 4097 5215 4131
rect 5273 4097 5307 4131
rect 7021 4097 7055 4131
rect 8217 4097 8251 4131
rect 11161 4097 11195 4131
rect 11253 4097 11287 4131
rect 11897 4097 11931 4131
rect 13001 4097 13035 4131
rect 13829 4097 13863 4131
rect 18705 4097 18739 4131
rect 19901 4097 19935 4131
rect 2053 4029 2087 4063
rect 2145 3961 2179 3995
rect 2697 3961 2731 3995
rect 5825 4029 5859 4063
rect 11069 4029 11103 4063
rect 12817 4029 12851 4063
rect 14197 4029 14231 4063
rect 14473 4029 14507 4063
rect 19625 4029 19659 4063
rect 20361 4029 20395 4063
rect 20913 4029 20947 4063
rect 21465 4029 21499 4063
rect 22017 4029 22051 4063
rect 22569 4029 22603 4063
rect 3709 3961 3743 3995
rect 6193 3961 6227 3995
rect 8484 3961 8518 3995
rect 10517 3961 10551 3995
rect 12909 3961 12943 3995
rect 14718 3961 14752 3995
rect 18521 3961 18555 3995
rect 2973 3893 3007 3927
rect 4721 3893 4755 3927
rect 5089 3893 5123 3927
rect 7205 3893 7239 3927
rect 9597 3893 9631 3927
rect 10701 3893 10735 3927
rect 12173 3893 12207 3927
rect 12449 3893 12483 3927
rect 13461 3893 13495 3927
rect 14013 3893 14047 3927
rect 15853 3893 15887 3927
rect 16865 3893 16899 3927
rect 16957 3893 16991 3927
rect 17417 3893 17451 3927
rect 17785 3893 17819 3927
rect 18429 3893 18463 3927
rect 19441 3893 19475 3927
rect 21097 3893 21131 3927
rect 22201 3893 22235 3927
rect 2881 3689 2915 3723
rect 3525 3689 3559 3723
rect 5181 3689 5215 3723
rect 6745 3689 6779 3723
rect 7757 3689 7791 3723
rect 10701 3689 10735 3723
rect 11069 3689 11103 3723
rect 13277 3689 13311 3723
rect 14749 3689 14783 3723
rect 15577 3689 15611 3723
rect 18613 3689 18647 3723
rect 19349 3689 19383 3723
rect 1768 3621 1802 3655
rect 5610 3621 5644 3655
rect 8309 3621 8343 3655
rect 10149 3621 10183 3655
rect 11520 3621 11554 3655
rect 14197 3621 14231 3655
rect 16028 3621 16062 3655
rect 17693 3621 17727 3655
rect 18061 3621 18095 3655
rect 18705 3621 18739 3655
rect 5365 3553 5399 3587
rect 8217 3553 8251 3587
rect 10057 3553 10091 3587
rect 13921 3553 13955 3587
rect 15117 3553 15151 3587
rect 15761 3553 15795 3587
rect 20913 3553 20947 3587
rect 22201 3553 22235 3587
rect 23305 3553 23339 3587
rect 1501 3485 1535 3519
rect 4353 3485 4387 3519
rect 7389 3485 7423 3519
rect 8401 3485 8435 3519
rect 8953 3485 8987 3519
rect 9505 3485 9539 3519
rect 10333 3485 10367 3519
rect 11253 3485 11287 3519
rect 18797 3485 18831 3519
rect 21189 3485 21223 3519
rect 3893 3417 3927 3451
rect 7849 3417 7883 3451
rect 9689 3417 9723 3451
rect 18245 3417 18279 3451
rect 4905 3349 4939 3383
rect 12633 3349 12667 3383
rect 13645 3349 13679 3383
rect 17141 3349 17175 3383
rect 22385 3349 22419 3383
rect 23489 3349 23523 3383
rect 2053 3145 2087 3179
rect 2697 3145 2731 3179
rect 4169 3145 4203 3179
rect 5641 3145 5675 3179
rect 6193 3145 6227 3179
rect 6561 3145 6595 3179
rect 7849 3145 7883 3179
rect 10609 3145 10643 3179
rect 14381 3145 14415 3179
rect 16865 3145 16899 3179
rect 17509 3145 17543 3179
rect 19073 3145 19107 3179
rect 20729 3145 20763 3179
rect 22109 3145 22143 3179
rect 22385 3145 22419 3179
rect 23305 3145 23339 3179
rect 3709 3077 3743 3111
rect 10149 3077 10183 3111
rect 10425 3077 10459 3111
rect 13829 3077 13863 3111
rect 14749 3077 14783 3111
rect 18061 3077 18095 3111
rect 24961 3077 24995 3111
rect 3157 3009 3191 3043
rect 3341 3009 3375 3043
rect 8125 3009 8159 3043
rect 11161 3009 11195 3043
rect 12449 3009 12483 3043
rect 18613 3009 18647 3043
rect 20361 3009 20395 3043
rect 21189 3009 21223 3043
rect 2605 2941 2639 2975
rect 3065 2941 3099 2975
rect 4261 2941 4295 2975
rect 4517 2941 4551 2975
rect 11069 2941 11103 2975
rect 14933 2941 14967 2975
rect 15189 2941 15223 2975
rect 18521 2941 18555 2975
rect 19441 2941 19475 2975
rect 19625 2941 19659 2975
rect 20913 2941 20947 2975
rect 21649 2941 21683 2975
rect 22201 2941 22235 2975
rect 22753 2941 22787 2975
rect 23673 2941 23707 2975
rect 24225 2941 24259 2975
rect 24777 2941 24811 2975
rect 25329 2941 25363 2975
rect 1685 2873 1719 2907
rect 7113 2873 7147 2907
rect 8392 2873 8426 2907
rect 12265 2873 12299 2907
rect 12694 2873 12728 2907
rect 17785 2873 17819 2907
rect 18429 2873 18463 2907
rect 19901 2873 19935 2907
rect 9505 2805 9539 2839
rect 10977 2805 11011 2839
rect 11713 2805 11747 2839
rect 16313 2805 16347 2839
rect 23857 2805 23891 2839
rect 2881 2601 2915 2635
rect 6929 2601 6963 2635
rect 7941 2601 7975 2635
rect 8401 2601 8435 2635
rect 10793 2601 10827 2635
rect 11621 2601 11655 2635
rect 12909 2601 12943 2635
rect 14289 2601 14323 2635
rect 15485 2601 15519 2635
rect 16957 2601 16991 2635
rect 17693 2601 17727 2635
rect 18061 2601 18095 2635
rect 19073 2601 19107 2635
rect 22661 2601 22695 2635
rect 24777 2601 24811 2635
rect 1746 2533 1780 2567
rect 3893 2533 3927 2567
rect 4344 2533 4378 2567
rect 9505 2533 9539 2567
rect 10149 2533 10183 2567
rect 13369 2533 13403 2567
rect 15945 2533 15979 2567
rect 21465 2533 21499 2567
rect 1501 2465 1535 2499
rect 4077 2465 4111 2499
rect 6653 2465 6687 2499
rect 7297 2465 7331 2499
rect 9137 2465 9171 2499
rect 11437 2465 11471 2499
rect 12449 2465 12483 2499
rect 12725 2465 12759 2499
rect 14197 2465 14231 2499
rect 15853 2465 15887 2499
rect 17049 2465 17083 2499
rect 18337 2465 18371 2499
rect 19441 2465 19475 2499
rect 19625 2465 19659 2499
rect 20361 2465 20395 2499
rect 21189 2465 21223 2499
rect 21925 2465 21959 2499
rect 22477 2465 22511 2499
rect 23029 2465 23063 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 6377 2397 6411 2431
rect 7389 2397 7423 2431
rect 7481 2397 7515 2431
rect 8677 2397 8711 2431
rect 10241 2397 10275 2431
rect 10425 2397 10459 2431
rect 11989 2397 12023 2431
rect 14473 2397 14507 2431
rect 16037 2397 16071 2431
rect 16497 2397 16531 2431
rect 18521 2397 18555 2431
rect 19809 2397 19843 2431
rect 9781 2329 9815 2363
rect 11161 2329 11195 2363
rect 13645 2329 13679 2363
rect 13829 2329 13863 2363
rect 3525 2261 3559 2295
rect 5457 2261 5491 2295
rect 14841 2261 14875 2295
rect 15301 2261 15335 2295
rect 17233 2261 17267 2295
<< metal1 >>
rect 3326 26664 3332 26716
rect 3384 26704 3390 26716
rect 5442 26704 5448 26716
rect 3384 26676 5448 26704
rect 3384 26664 3390 26676
rect 5442 26664 5448 26676
rect 5500 26664 5506 26716
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1581 25483 1639 25489
rect 1581 25449 1593 25483
rect 1627 25480 1639 25483
rect 2774 25480 2780 25492
rect 1627 25452 2780 25480
rect 1627 25449 1639 25452
rect 1581 25443 1639 25449
rect 2774 25440 2780 25452
rect 2832 25440 2838 25492
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1578 24936 1584 24948
rect 1539 24908 1584 24936
rect 1578 24896 1584 24908
rect 1636 24896 1642 24948
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 1443 24704 2084 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 2056 24605 2084 24704
rect 2041 24599 2099 24605
rect 2041 24565 2053 24599
rect 2087 24596 2099 24599
rect 2130 24596 2136 24608
rect 2087 24568 2136 24596
rect 2087 24565 2099 24568
rect 2041 24559 2099 24565
rect 2130 24556 2136 24568
rect 2188 24556 2194 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1486 24352 1492 24404
rect 1544 24392 1550 24404
rect 1581 24395 1639 24401
rect 1581 24392 1593 24395
rect 1544 24364 1593 24392
rect 1544 24352 1550 24364
rect 1581 24361 1593 24364
rect 1627 24361 1639 24395
rect 2682 24392 2688 24404
rect 2643 24364 2688 24392
rect 1581 24355 1639 24361
rect 2682 24352 2688 24364
rect 2740 24352 2746 24404
rect 1394 24256 1400 24268
rect 1355 24228 1400 24256
rect 1394 24216 1400 24228
rect 1452 24216 1458 24268
rect 2498 24256 2504 24268
rect 2459 24228 2504 24256
rect 2498 24216 2504 24228
rect 2556 24216 2562 24268
rect 2038 24120 2044 24132
rect 1999 24092 2044 24120
rect 2038 24080 2044 24092
rect 2096 24080 2102 24132
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2498 23848 2504 23860
rect 2459 23820 2504 23848
rect 2498 23808 2504 23820
rect 2556 23808 2562 23860
rect 3234 23848 3240 23860
rect 3195 23820 3240 23848
rect 3234 23808 3240 23820
rect 3292 23808 3298 23860
rect 24762 23848 24768 23860
rect 24723 23820 24768 23848
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 2041 23715 2099 23721
rect 2041 23681 2053 23715
rect 2087 23712 2099 23715
rect 2516 23712 2544 23808
rect 3694 23712 3700 23724
rect 2087 23684 2544 23712
rect 3068 23684 3700 23712
rect 2087 23681 2099 23684
rect 2041 23675 2099 23681
rect 1765 23647 1823 23653
rect 1765 23613 1777 23647
rect 1811 23644 1823 23647
rect 1946 23644 1952 23656
rect 1811 23616 1952 23644
rect 1811 23613 1823 23616
rect 1765 23607 1823 23613
rect 1946 23604 1952 23616
rect 2004 23604 2010 23656
rect 3068 23653 3096 23684
rect 3694 23672 3700 23684
rect 3752 23672 3758 23724
rect 3053 23647 3111 23653
rect 3053 23613 3065 23647
rect 3099 23613 3111 23647
rect 3053 23607 3111 23613
rect 1394 23468 1400 23520
rect 1452 23508 1458 23520
rect 1673 23511 1731 23517
rect 1673 23508 1685 23511
rect 1452 23480 1685 23508
rect 1452 23468 1458 23480
rect 1673 23477 1685 23480
rect 1719 23508 1731 23511
rect 1946 23508 1952 23520
rect 1719 23480 1952 23508
rect 1719 23477 1731 23480
rect 1673 23471 1731 23477
rect 1946 23468 1952 23480
rect 2004 23468 2010 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2041 23239 2099 23245
rect 2041 23205 2053 23239
rect 2087 23236 2099 23239
rect 2130 23236 2136 23248
rect 2087 23208 2136 23236
rect 2087 23205 2099 23208
rect 2041 23199 2099 23205
rect 2130 23196 2136 23208
rect 2188 23196 2194 23248
rect 12710 23236 12716 23248
rect 12671 23208 12716 23236
rect 12710 23196 12716 23208
rect 12768 23196 12774 23248
rect 1670 23128 1676 23180
rect 1728 23168 1734 23180
rect 1765 23171 1823 23177
rect 1765 23168 1777 23171
rect 1728 23140 1777 23168
rect 1728 23128 1734 23140
rect 1765 23137 1777 23140
rect 1811 23137 1823 23171
rect 12434 23168 12440 23180
rect 12395 23140 12440 23168
rect 1765 23131 1823 23137
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2958 22720 2964 22772
rect 3016 22760 3022 22772
rect 3237 22763 3295 22769
rect 3237 22760 3249 22763
rect 3016 22732 3249 22760
rect 3016 22720 3022 22732
rect 3237 22729 3249 22732
rect 3283 22729 3295 22763
rect 3237 22723 3295 22729
rect 1946 22624 1952 22636
rect 1907 22596 1952 22624
rect 1946 22584 1952 22596
rect 2004 22584 2010 22636
rect 1670 22556 1676 22568
rect 1631 22528 1676 22556
rect 1670 22516 1676 22528
rect 1728 22516 1734 22568
rect 1765 22559 1823 22565
rect 1765 22525 1777 22559
rect 1811 22556 1823 22559
rect 3053 22559 3111 22565
rect 1811 22528 2636 22556
rect 1811 22525 1823 22528
rect 1765 22519 1823 22525
rect 2608 22432 2636 22528
rect 3053 22525 3065 22559
rect 3099 22556 3111 22559
rect 3099 22528 3740 22556
rect 3099 22525 3111 22528
rect 3053 22519 3111 22525
rect 3712 22432 3740 22528
rect 2590 22420 2596 22432
rect 2551 22392 2596 22420
rect 2590 22380 2596 22392
rect 2648 22380 2654 22432
rect 3694 22420 3700 22432
rect 3655 22392 3700 22420
rect 3694 22380 3700 22392
rect 3752 22380 3758 22432
rect 12434 22380 12440 22432
rect 12492 22420 12498 22432
rect 12713 22423 12771 22429
rect 12713 22420 12725 22423
rect 12492 22392 12725 22420
rect 12492 22380 12498 22392
rect 12713 22389 12725 22392
rect 12759 22420 12771 22423
rect 13354 22420 13360 22432
rect 12759 22392 13360 22420
rect 12759 22389 12771 22392
rect 12713 22383 12771 22389
rect 13354 22380 13360 22392
rect 13412 22380 13418 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1394 22080 1400 22092
rect 1355 22052 1400 22080
rect 1394 22040 1400 22052
rect 1452 22040 1458 22092
rect 2406 22040 2412 22092
rect 2464 22080 2470 22092
rect 2501 22083 2559 22089
rect 2501 22080 2513 22083
rect 2464 22052 2513 22080
rect 2464 22040 2470 22052
rect 2501 22049 2513 22052
rect 2547 22049 2559 22083
rect 2501 22043 2559 22049
rect 2682 21944 2688 21956
rect 2643 21916 2688 21944
rect 2682 21904 2688 21916
rect 2740 21904 2746 21956
rect 1578 21876 1584 21888
rect 1539 21848 1584 21876
rect 1578 21836 1584 21848
rect 1636 21836 1642 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1486 21632 1492 21684
rect 1544 21672 1550 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 1544 21644 1593 21672
rect 1544 21632 1550 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 8570 21672 8576 21684
rect 8531 21644 8576 21672
rect 1581 21635 1639 21641
rect 8570 21632 8576 21644
rect 8628 21632 8634 21684
rect 2682 21604 2688 21616
rect 2643 21576 2688 21604
rect 2682 21564 2688 21576
rect 2740 21564 2746 21616
rect 7282 21536 7288 21548
rect 7243 21508 7288 21536
rect 7282 21496 7288 21508
rect 7340 21496 7346 21548
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 1670 21468 1676 21480
rect 1443 21440 1676 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 1670 21428 1676 21440
rect 1728 21428 1734 21480
rect 2038 21428 2044 21480
rect 2096 21468 2102 21480
rect 2501 21471 2559 21477
rect 2501 21468 2513 21471
rect 2096 21440 2513 21468
rect 2096 21428 2102 21440
rect 2501 21437 2513 21440
rect 2547 21468 2559 21471
rect 3053 21471 3111 21477
rect 3053 21468 3065 21471
rect 2547 21440 3065 21468
rect 2547 21437 2559 21440
rect 2501 21431 2559 21437
rect 3053 21437 3065 21440
rect 3099 21437 3111 21471
rect 3053 21431 3111 21437
rect 7101 21471 7159 21477
rect 7101 21437 7113 21471
rect 7147 21468 7159 21471
rect 8389 21471 8447 21477
rect 7147 21440 7880 21468
rect 7147 21437 7159 21440
rect 7101 21431 7159 21437
rect 2406 21400 2412 21412
rect 2367 21372 2412 21400
rect 2406 21360 2412 21372
rect 2464 21360 2470 21412
rect 7852 21344 7880 21440
rect 8389 21437 8401 21471
rect 8435 21468 8447 21471
rect 8754 21468 8760 21480
rect 8435 21440 8760 21468
rect 8435 21437 8447 21440
rect 8389 21431 8447 21437
rect 8754 21428 8760 21440
rect 8812 21468 8818 21480
rect 8941 21471 8999 21477
rect 8941 21468 8953 21471
rect 8812 21440 8953 21468
rect 8812 21428 8818 21440
rect 8941 21437 8953 21440
rect 8987 21437 8999 21471
rect 8941 21431 8999 21437
rect 1394 21292 1400 21344
rect 1452 21332 1458 21344
rect 2041 21335 2099 21341
rect 2041 21332 2053 21335
rect 1452 21304 2053 21332
rect 1452 21292 1458 21304
rect 2041 21301 2053 21304
rect 2087 21332 2099 21335
rect 2498 21332 2504 21344
rect 2087 21304 2504 21332
rect 2087 21301 2099 21304
rect 2041 21295 2099 21301
rect 2498 21292 2504 21304
rect 2556 21292 2562 21344
rect 7834 21332 7840 21344
rect 7795 21304 7840 21332
rect 7834 21292 7840 21304
rect 7892 21292 7898 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1762 20992 1768 21004
rect 1723 20964 1768 20992
rect 1762 20952 1768 20964
rect 1820 20952 1826 21004
rect 7926 20992 7932 21004
rect 7887 20964 7932 20992
rect 7926 20952 7932 20964
rect 7984 20952 7990 21004
rect 1670 20924 1676 20936
rect 1631 20896 1676 20924
rect 1670 20884 1676 20896
rect 1728 20884 1734 20936
rect 2041 20927 2099 20933
rect 2041 20893 2053 20927
rect 2087 20924 2099 20927
rect 2682 20924 2688 20936
rect 2087 20896 2688 20924
rect 2087 20893 2099 20896
rect 2041 20887 2099 20893
rect 2682 20884 2688 20896
rect 2740 20884 2746 20936
rect 8110 20924 8116 20936
rect 8071 20896 8116 20924
rect 8110 20884 8116 20896
rect 8168 20884 8174 20936
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2590 20584 2596 20596
rect 2551 20556 2596 20584
rect 2590 20544 2596 20556
rect 2648 20544 2654 20596
rect 4154 20544 4160 20596
rect 4212 20584 4218 20596
rect 4341 20587 4399 20593
rect 4341 20584 4353 20587
rect 4212 20556 4353 20584
rect 4212 20544 4218 20556
rect 4341 20553 4353 20556
rect 4387 20553 4399 20587
rect 4341 20547 4399 20553
rect 2038 20448 2044 20460
rect 1999 20420 2044 20448
rect 2038 20408 2044 20420
rect 2096 20408 2102 20460
rect 8754 20448 8760 20460
rect 8715 20420 8760 20448
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20380 1823 20383
rect 2590 20380 2596 20392
rect 1811 20352 2596 20380
rect 1811 20349 1823 20352
rect 1765 20343 1823 20349
rect 2590 20340 2596 20352
rect 2648 20340 2654 20392
rect 2774 20340 2780 20392
rect 2832 20380 2838 20392
rect 3053 20383 3111 20389
rect 3053 20380 3065 20383
rect 2832 20352 3065 20380
rect 2832 20340 2838 20352
rect 3053 20349 3065 20352
rect 3099 20380 3111 20383
rect 3605 20383 3663 20389
rect 3605 20380 3617 20383
rect 3099 20352 3617 20380
rect 3099 20349 3111 20352
rect 3053 20343 3111 20349
rect 3605 20349 3617 20352
rect 3651 20349 3663 20383
rect 4154 20380 4160 20392
rect 4115 20352 4160 20380
rect 3605 20343 3663 20349
rect 4154 20340 4160 20352
rect 4212 20380 4218 20392
rect 4709 20383 4767 20389
rect 4709 20380 4721 20383
rect 4212 20352 4721 20380
rect 4212 20340 4218 20352
rect 4709 20349 4721 20352
rect 4755 20349 4767 20383
rect 4709 20343 4767 20349
rect 8573 20383 8631 20389
rect 8573 20349 8585 20383
rect 8619 20380 8631 20383
rect 8619 20352 9444 20380
rect 8619 20349 8631 20352
rect 8573 20343 8631 20349
rect 9416 20256 9444 20352
rect 1673 20247 1731 20253
rect 1673 20213 1685 20247
rect 1719 20244 1731 20247
rect 1762 20244 1768 20256
rect 1719 20216 1768 20244
rect 1719 20213 1731 20216
rect 1673 20207 1731 20213
rect 1762 20204 1768 20216
rect 1820 20204 1826 20256
rect 3234 20244 3240 20256
rect 3195 20216 3240 20244
rect 3234 20204 3240 20216
rect 3292 20204 3298 20256
rect 7926 20244 7932 20256
rect 7887 20216 7932 20244
rect 7926 20204 7932 20216
rect 7984 20204 7990 20256
rect 9398 20244 9404 20256
rect 9359 20216 9404 20244
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 4246 20040 4252 20052
rect 4207 20012 4252 20040
rect 4246 20000 4252 20012
rect 4304 20000 4310 20052
rect 1857 19975 1915 19981
rect 1857 19941 1869 19975
rect 1903 19972 1915 19975
rect 1903 19944 4108 19972
rect 1903 19941 1915 19944
rect 1857 19935 1915 19941
rect 4080 19916 4108 19944
rect 7374 19932 7380 19984
rect 7432 19972 7438 19984
rect 7929 19975 7987 19981
rect 7929 19972 7941 19975
rect 7432 19944 7941 19972
rect 7432 19932 7438 19944
rect 7929 19941 7941 19944
rect 7975 19941 7987 19975
rect 7929 19935 7987 19941
rect 1581 19907 1639 19913
rect 1581 19873 1593 19907
rect 1627 19904 1639 19907
rect 1670 19904 1676 19916
rect 1627 19876 1676 19904
rect 1627 19873 1639 19876
rect 1581 19867 1639 19873
rect 1670 19864 1676 19876
rect 1728 19864 1734 19916
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19904 2927 19907
rect 2958 19904 2964 19916
rect 2915 19876 2964 19904
rect 2915 19873 2927 19876
rect 2869 19867 2927 19873
rect 2958 19864 2964 19876
rect 3016 19864 3022 19916
rect 4062 19904 4068 19916
rect 3975 19876 4068 19904
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 7650 19904 7656 19916
rect 7611 19876 7656 19904
rect 7650 19864 7656 19876
rect 7708 19864 7714 19916
rect 4798 19796 4804 19848
rect 4856 19836 4862 19848
rect 5169 19839 5227 19845
rect 5169 19836 5181 19839
rect 4856 19808 5181 19836
rect 4856 19796 4862 19808
rect 5169 19805 5181 19808
rect 5215 19805 5227 19839
rect 5169 19799 5227 19805
rect 2866 19660 2872 19712
rect 2924 19700 2930 19712
rect 3053 19703 3111 19709
rect 3053 19700 3065 19703
rect 2924 19672 3065 19700
rect 2924 19660 2930 19672
rect 3053 19669 3065 19672
rect 3099 19669 3111 19703
rect 3053 19663 3111 19669
rect 6914 19660 6920 19712
rect 6972 19700 6978 19712
rect 6972 19672 7017 19700
rect 6972 19660 6978 19672
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 4062 19496 4068 19508
rect 4023 19468 4068 19496
rect 4062 19456 4068 19468
rect 4120 19456 4126 19508
rect 2498 19320 2504 19372
rect 2556 19360 2562 19372
rect 3329 19363 3387 19369
rect 3329 19360 3341 19363
rect 2556 19332 3341 19360
rect 2556 19320 2562 19332
rect 3329 19329 3341 19332
rect 3375 19329 3387 19363
rect 3329 19323 3387 19329
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 7374 19360 7380 19372
rect 6972 19332 7380 19360
rect 6972 19320 6978 19332
rect 7374 19320 7380 19332
rect 7432 19320 7438 19372
rect 1857 19295 1915 19301
rect 1857 19261 1869 19295
rect 1903 19261 1915 19295
rect 1857 19255 1915 19261
rect 2133 19295 2191 19301
rect 2133 19261 2145 19295
rect 2179 19292 2191 19295
rect 2682 19292 2688 19304
rect 2179 19264 2688 19292
rect 2179 19261 2191 19264
rect 2133 19255 2191 19261
rect 1872 19224 1900 19255
rect 2682 19252 2688 19264
rect 2740 19252 2746 19304
rect 3145 19295 3203 19301
rect 3145 19261 3157 19295
rect 3191 19261 3203 19295
rect 3145 19255 3203 19261
rect 1872 19196 2728 19224
rect 2700 19168 2728 19196
rect 1670 19156 1676 19168
rect 1631 19128 1676 19156
rect 1670 19116 1676 19128
rect 1728 19116 1734 19168
rect 2682 19156 2688 19168
rect 2643 19128 2688 19156
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 3053 19159 3111 19165
rect 3053 19125 3065 19159
rect 3099 19156 3111 19159
rect 3160 19156 3188 19255
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 4433 19295 4491 19301
rect 4433 19292 4445 19295
rect 4212 19264 4445 19292
rect 4212 19252 4218 19264
rect 4433 19261 4445 19264
rect 4479 19292 4491 19295
rect 4985 19295 5043 19301
rect 4985 19292 4997 19295
rect 4479 19264 4997 19292
rect 4479 19261 4491 19264
rect 4433 19255 4491 19261
rect 4985 19261 4997 19264
rect 5031 19261 5043 19295
rect 4985 19255 5043 19261
rect 6454 19252 6460 19304
rect 6512 19292 6518 19304
rect 7285 19295 7343 19301
rect 7285 19292 7297 19295
rect 6512 19264 7297 19292
rect 6512 19252 6518 19264
rect 7285 19261 7297 19264
rect 7331 19261 7343 19295
rect 7285 19255 7343 19261
rect 11974 19252 11980 19304
rect 12032 19292 12038 19304
rect 12986 19292 12992 19304
rect 12032 19264 12992 19292
rect 12032 19252 12038 19264
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 5721 19227 5779 19233
rect 5721 19193 5733 19227
rect 5767 19224 5779 19227
rect 6549 19227 6607 19233
rect 6549 19224 6561 19227
rect 5767 19196 6561 19224
rect 5767 19193 5779 19196
rect 5721 19187 5779 19193
rect 6549 19193 6561 19196
rect 6595 19224 6607 19227
rect 7193 19227 7251 19233
rect 7193 19224 7205 19227
rect 6595 19196 7205 19224
rect 6595 19193 6607 19196
rect 6549 19187 6607 19193
rect 7193 19193 7205 19196
rect 7239 19193 7251 19227
rect 7193 19187 7251 19193
rect 3234 19156 3240 19168
rect 3099 19128 3240 19156
rect 3099 19125 3111 19128
rect 3053 19119 3111 19125
rect 3234 19116 3240 19128
rect 3292 19116 3298 19168
rect 4614 19156 4620 19168
rect 4575 19128 4620 19156
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 6273 19159 6331 19165
rect 6273 19125 6285 19159
rect 6319 19156 6331 19159
rect 6454 19156 6460 19168
rect 6319 19128 6460 19156
rect 6319 19125 6331 19128
rect 6273 19119 6331 19125
rect 6454 19116 6460 19128
rect 6512 19116 6518 19168
rect 6822 19156 6828 19168
rect 6783 19128 6828 19156
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7650 19116 7656 19168
rect 7708 19156 7714 19168
rect 7837 19159 7895 19165
rect 7837 19156 7849 19159
rect 7708 19128 7849 19156
rect 7708 19116 7714 19128
rect 7837 19125 7849 19128
rect 7883 19125 7895 19159
rect 7837 19119 7895 19125
rect 10965 19159 11023 19165
rect 10965 19125 10977 19159
rect 11011 19156 11023 19159
rect 12158 19156 12164 19168
rect 11011 19128 12164 19156
rect 11011 19125 11023 19128
rect 10965 19119 11023 19125
rect 12158 19116 12164 19128
rect 12216 19116 12222 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1486 18912 1492 18964
rect 1544 18952 1550 18964
rect 2777 18955 2835 18961
rect 2777 18952 2789 18955
rect 1544 18924 2789 18952
rect 1544 18912 1550 18924
rect 2777 18921 2789 18924
rect 2823 18952 2835 18955
rect 4338 18952 4344 18964
rect 2823 18924 4344 18952
rect 2823 18921 2835 18924
rect 2777 18915 2835 18921
rect 4338 18912 4344 18924
rect 4396 18912 4402 18964
rect 5534 18844 5540 18896
rect 5592 18893 5598 18896
rect 5592 18887 5656 18893
rect 5592 18853 5610 18887
rect 5644 18853 5656 18887
rect 5592 18847 5656 18853
rect 5592 18844 5598 18847
rect 10594 18844 10600 18896
rect 10652 18893 10658 18896
rect 10652 18887 10716 18893
rect 10652 18853 10670 18887
rect 10704 18853 10716 18887
rect 10652 18847 10716 18853
rect 10652 18844 10658 18847
rect 1581 18819 1639 18825
rect 1581 18785 1593 18819
rect 1627 18816 1639 18819
rect 2590 18816 2596 18828
rect 1627 18788 2596 18816
rect 1627 18785 1639 18788
rect 1581 18779 1639 18785
rect 2590 18776 2596 18788
rect 2648 18776 2654 18828
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18816 2927 18819
rect 3142 18816 3148 18828
rect 2915 18788 3148 18816
rect 2915 18785 2927 18788
rect 2869 18779 2927 18785
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 3712 18788 4077 18816
rect 3712 18760 3740 18788
rect 4065 18785 4077 18788
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 1857 18751 1915 18757
rect 1857 18717 1869 18751
rect 1903 18748 1915 18751
rect 3694 18748 3700 18760
rect 1903 18720 3700 18748
rect 1903 18717 1915 18720
rect 1857 18711 1915 18717
rect 3694 18708 3700 18720
rect 3752 18708 3758 18760
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 4632 18720 5365 18748
rect 1762 18640 1768 18692
rect 1820 18680 1826 18692
rect 2958 18680 2964 18692
rect 1820 18652 2964 18680
rect 1820 18640 1826 18652
rect 2958 18640 2964 18652
rect 3016 18680 3022 18692
rect 3421 18683 3479 18689
rect 3421 18680 3433 18683
rect 3016 18652 3433 18680
rect 3016 18640 3022 18652
rect 3421 18649 3433 18652
rect 3467 18649 3479 18683
rect 4246 18680 4252 18692
rect 4207 18652 4252 18680
rect 3421 18643 3479 18649
rect 4246 18640 4252 18652
rect 4304 18640 4310 18692
rect 2314 18612 2320 18624
rect 2275 18584 2320 18612
rect 2314 18572 2320 18584
rect 2372 18572 2378 18624
rect 3050 18612 3056 18624
rect 3011 18584 3056 18612
rect 3050 18572 3056 18584
rect 3108 18572 3114 18624
rect 3878 18612 3884 18624
rect 3839 18584 3884 18612
rect 3878 18572 3884 18584
rect 3936 18612 3942 18624
rect 4632 18621 4660 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 8018 18708 8024 18760
rect 8076 18748 8082 18760
rect 8573 18751 8631 18757
rect 8573 18748 8585 18751
rect 8076 18720 8585 18748
rect 8076 18708 8082 18720
rect 8573 18717 8585 18720
rect 8619 18717 8631 18751
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 8573 18711 8631 18717
rect 9324 18720 10425 18748
rect 9324 18624 9352 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 4617 18615 4675 18621
rect 4617 18612 4629 18615
rect 3936 18584 4629 18612
rect 3936 18572 3942 18584
rect 4617 18581 4629 18584
rect 4663 18581 4675 18615
rect 6730 18612 6736 18624
rect 6691 18584 6736 18612
rect 4617 18575 4675 18581
rect 6730 18572 6736 18584
rect 6788 18572 6794 18624
rect 7745 18615 7803 18621
rect 7745 18581 7757 18615
rect 7791 18612 7803 18615
rect 8202 18612 8208 18624
rect 7791 18584 8208 18612
rect 7791 18581 7803 18584
rect 7745 18575 7803 18581
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 9306 18612 9312 18624
rect 9267 18584 9312 18612
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 11790 18612 11796 18624
rect 11751 18584 11796 18612
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 12526 18612 12532 18624
rect 12487 18584 12532 18612
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 3694 18408 3700 18420
rect 3655 18380 3700 18408
rect 3694 18368 3700 18380
rect 3752 18368 3758 18420
rect 7650 18408 7656 18420
rect 7611 18380 7656 18408
rect 7650 18368 7656 18380
rect 7708 18368 7714 18420
rect 12158 18408 12164 18420
rect 12119 18380 12164 18408
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 10594 18340 10600 18352
rect 10555 18312 10600 18340
rect 10594 18300 10600 18312
rect 10652 18340 10658 18352
rect 11149 18343 11207 18349
rect 11149 18340 11161 18343
rect 10652 18312 11161 18340
rect 10652 18300 10658 18312
rect 11149 18309 11161 18312
rect 11195 18309 11207 18343
rect 11149 18303 11207 18309
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 2590 18272 2596 18284
rect 2363 18244 2596 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 2590 18232 2596 18244
rect 2648 18232 2654 18284
rect 3053 18275 3111 18281
rect 3053 18241 3065 18275
rect 3099 18272 3111 18275
rect 4154 18272 4160 18284
rect 3099 18244 4160 18272
rect 3099 18241 3111 18244
rect 3053 18235 3111 18241
rect 4154 18232 4160 18244
rect 4212 18232 4218 18284
rect 8202 18272 8208 18284
rect 8163 18244 8208 18272
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 12989 18275 13047 18281
rect 12989 18272 13001 18275
rect 12584 18244 13001 18272
rect 12584 18232 12590 18244
rect 12989 18241 13001 18244
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 1486 18204 1492 18216
rect 1447 18176 1492 18204
rect 1486 18164 1492 18176
rect 1544 18164 1550 18216
rect 2777 18207 2835 18213
rect 2777 18204 2789 18207
rect 2700 18176 2789 18204
rect 2700 18080 2728 18176
rect 2777 18173 2789 18176
rect 2823 18173 2835 18207
rect 2777 18167 2835 18173
rect 3878 18164 3884 18216
rect 3936 18204 3942 18216
rect 4246 18204 4252 18216
rect 3936 18176 4252 18204
rect 3936 18164 3942 18176
rect 4246 18164 4252 18176
rect 4304 18164 4310 18216
rect 7561 18207 7619 18213
rect 7561 18173 7573 18207
rect 7607 18204 7619 18207
rect 8018 18204 8024 18216
rect 7607 18176 8024 18204
rect 7607 18173 7619 18176
rect 7561 18167 7619 18173
rect 8018 18164 8024 18176
rect 8076 18164 8082 18216
rect 9217 18207 9275 18213
rect 9217 18173 9229 18207
rect 9263 18204 9275 18207
rect 9306 18204 9312 18216
rect 9263 18176 9312 18204
rect 9263 18173 9275 18176
rect 9217 18167 9275 18173
rect 9306 18164 9312 18176
rect 9364 18164 9370 18216
rect 12158 18164 12164 18216
rect 12216 18204 12222 18216
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 12216 18176 12817 18204
rect 12216 18164 12222 18176
rect 12805 18173 12817 18176
rect 12851 18173 12863 18207
rect 12805 18167 12863 18173
rect 4157 18139 4215 18145
rect 4157 18105 4169 18139
rect 4203 18136 4215 18139
rect 4494 18139 4552 18145
rect 4494 18136 4506 18139
rect 4203 18108 4506 18136
rect 4203 18105 4215 18108
rect 4157 18099 4215 18105
rect 4494 18105 4506 18108
rect 4540 18136 4552 18139
rect 4982 18136 4988 18148
rect 4540 18108 4988 18136
rect 4540 18105 4552 18108
rect 4494 18099 4552 18105
rect 4982 18096 4988 18108
rect 5040 18096 5046 18148
rect 9125 18139 9183 18145
rect 9125 18105 9137 18139
rect 9171 18136 9183 18139
rect 9462 18139 9520 18145
rect 9462 18136 9474 18139
rect 9171 18108 9474 18136
rect 9171 18105 9183 18108
rect 9125 18099 9183 18105
rect 9462 18105 9474 18108
rect 9508 18136 9520 18139
rect 9766 18136 9772 18148
rect 9508 18108 9772 18136
rect 9508 18105 9520 18108
rect 9462 18099 9520 18105
rect 9766 18096 9772 18108
rect 9824 18096 9830 18148
rect 12897 18139 12955 18145
rect 12897 18136 12909 18139
rect 11808 18108 12909 18136
rect 2682 18068 2688 18080
rect 2643 18040 2688 18068
rect 2682 18028 2688 18040
rect 2740 18028 2746 18080
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 5629 18071 5687 18077
rect 5629 18068 5641 18071
rect 5592 18040 5641 18068
rect 5592 18028 5598 18040
rect 5629 18037 5641 18040
rect 5675 18068 5687 18071
rect 6181 18071 6239 18077
rect 6181 18068 6193 18071
rect 5675 18040 6193 18068
rect 5675 18037 5687 18040
rect 5629 18031 5687 18037
rect 6181 18037 6193 18040
rect 6227 18037 6239 18071
rect 6181 18031 6239 18037
rect 7193 18071 7251 18077
rect 7193 18037 7205 18071
rect 7239 18068 7251 18071
rect 8110 18068 8116 18080
rect 7239 18040 8116 18068
rect 7239 18037 7251 18040
rect 7193 18031 7251 18037
rect 8110 18028 8116 18040
rect 8168 18028 8174 18080
rect 11146 18028 11152 18080
rect 11204 18068 11210 18080
rect 11808 18077 11836 18108
rect 12897 18105 12909 18108
rect 12943 18105 12955 18139
rect 12897 18099 12955 18105
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 11204 18040 11805 18068
rect 11204 18028 11210 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 11793 18031 11851 18037
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 12492 18040 12537 18068
rect 12492 18028 12498 18040
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1854 17824 1860 17876
rect 1912 17864 1918 17876
rect 2133 17867 2191 17873
rect 2133 17864 2145 17867
rect 1912 17836 2145 17864
rect 1912 17824 1918 17836
rect 2133 17833 2145 17836
rect 2179 17864 2191 17867
rect 2314 17864 2320 17876
rect 2179 17836 2320 17864
rect 2179 17833 2191 17836
rect 2133 17827 2191 17833
rect 2314 17824 2320 17836
rect 2372 17824 2378 17876
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 7432 17836 7665 17864
rect 7432 17824 7438 17836
rect 7653 17833 7665 17836
rect 7699 17833 7711 17867
rect 7653 17827 7711 17833
rect 7834 17824 7840 17876
rect 7892 17864 7898 17876
rect 8018 17864 8024 17876
rect 7892 17836 8024 17864
rect 7892 17824 7898 17836
rect 8018 17824 8024 17836
rect 8076 17824 8082 17876
rect 9674 17864 9680 17876
rect 9635 17836 9680 17864
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 12526 17824 12532 17876
rect 12584 17864 12590 17876
rect 12713 17867 12771 17873
rect 12713 17864 12725 17867
rect 12584 17836 12725 17864
rect 12584 17824 12590 17836
rect 12713 17833 12725 17836
rect 12759 17833 12771 17867
rect 12713 17827 12771 17833
rect 6540 17799 6598 17805
rect 6540 17765 6552 17799
rect 6586 17796 6598 17799
rect 6730 17796 6736 17808
rect 6586 17768 6736 17796
rect 6586 17765 6598 17768
rect 6540 17759 6598 17765
rect 6730 17756 6736 17768
rect 6788 17756 6794 17808
rect 9766 17756 9772 17808
rect 9824 17796 9830 17808
rect 11600 17799 11658 17805
rect 9824 17768 10272 17796
rect 9824 17756 9830 17768
rect 2225 17731 2283 17737
rect 2225 17697 2237 17731
rect 2271 17728 2283 17731
rect 2498 17728 2504 17740
rect 2271 17700 2504 17728
rect 2271 17697 2283 17700
rect 2225 17691 2283 17697
rect 2498 17688 2504 17700
rect 2556 17728 2562 17740
rect 3237 17731 3295 17737
rect 3237 17728 3249 17731
rect 2556 17700 3249 17728
rect 2556 17688 2562 17700
rect 3237 17697 3249 17700
rect 3283 17697 3295 17731
rect 3237 17691 3295 17697
rect 4614 17688 4620 17740
rect 4672 17728 4678 17740
rect 4801 17731 4859 17737
rect 4801 17728 4813 17731
rect 4672 17700 4813 17728
rect 4672 17688 4678 17700
rect 4801 17697 4813 17700
rect 4847 17697 4859 17731
rect 4801 17691 4859 17697
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17728 4951 17731
rect 5350 17728 5356 17740
rect 4939 17700 5356 17728
rect 4939 17697 4951 17700
rect 4893 17691 4951 17697
rect 5350 17688 5356 17700
rect 5408 17688 5414 17740
rect 8754 17688 8760 17740
rect 8812 17728 8818 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 8812 17700 10057 17728
rect 8812 17688 8818 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 2130 17660 2136 17672
rect 1719 17632 2136 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 2130 17620 2136 17632
rect 2188 17660 2194 17672
rect 2317 17663 2375 17669
rect 2317 17660 2329 17663
rect 2188 17632 2329 17660
rect 2188 17620 2194 17632
rect 2317 17629 2329 17632
rect 2363 17629 2375 17663
rect 4982 17660 4988 17672
rect 4943 17632 4988 17660
rect 2317 17623 2375 17629
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 6273 17663 6331 17669
rect 6273 17629 6285 17663
rect 6319 17629 6331 17663
rect 10134 17660 10140 17672
rect 10095 17632 10140 17660
rect 6273 17623 6331 17629
rect 5445 17595 5503 17601
rect 5445 17592 5457 17595
rect 4264 17564 5457 17592
rect 4264 17536 4292 17564
rect 5445 17561 5457 17564
rect 5491 17592 5503 17595
rect 5994 17592 6000 17604
rect 5491 17564 6000 17592
rect 5491 17561 5503 17564
rect 5445 17555 5503 17561
rect 5994 17552 6000 17564
rect 6052 17592 6058 17604
rect 6089 17595 6147 17601
rect 6089 17592 6101 17595
rect 6052 17564 6101 17592
rect 6052 17552 6058 17564
rect 6089 17561 6101 17564
rect 6135 17592 6147 17595
rect 6288 17592 6316 17623
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10244 17669 10272 17768
rect 11600 17765 11612 17799
rect 11646 17796 11658 17799
rect 11790 17796 11796 17808
rect 11646 17768 11796 17796
rect 11646 17765 11658 17768
rect 11600 17759 11658 17765
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17660 10287 17663
rect 10686 17660 10692 17672
rect 10275 17632 10692 17660
rect 10275 17629 10287 17632
rect 10229 17623 10287 17629
rect 10686 17620 10692 17632
rect 10744 17620 10750 17672
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17660 10839 17663
rect 11330 17660 11336 17672
rect 10827 17632 11336 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 6135 17564 6316 17592
rect 6135 17561 6147 17564
rect 6089 17555 6147 17561
rect 9306 17552 9312 17604
rect 9364 17592 9370 17604
rect 9401 17595 9459 17601
rect 9401 17592 9413 17595
rect 9364 17564 9413 17592
rect 9364 17552 9370 17564
rect 9401 17561 9413 17564
rect 9447 17592 9459 17595
rect 10796 17592 10824 17623
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 9447 17564 10824 17592
rect 9447 17561 9459 17564
rect 9401 17555 9459 17561
rect 1765 17527 1823 17533
rect 1765 17493 1777 17527
rect 1811 17524 1823 17527
rect 1946 17524 1952 17536
rect 1811 17496 1952 17524
rect 1811 17493 1823 17496
rect 1765 17487 1823 17493
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 2682 17484 2688 17536
rect 2740 17524 2746 17536
rect 2869 17527 2927 17533
rect 2869 17524 2881 17527
rect 2740 17496 2881 17524
rect 2740 17484 2746 17496
rect 2869 17493 2881 17496
rect 2915 17524 2927 17527
rect 3142 17524 3148 17536
rect 2915 17496 3148 17524
rect 2915 17493 2927 17496
rect 2869 17487 2927 17493
rect 3142 17484 3148 17496
rect 3200 17484 3206 17536
rect 3418 17484 3424 17536
rect 3476 17524 3482 17536
rect 3605 17527 3663 17533
rect 3605 17524 3617 17527
rect 3476 17496 3617 17524
rect 3476 17484 3482 17496
rect 3605 17493 3617 17496
rect 3651 17524 3663 17527
rect 4246 17524 4252 17536
rect 3651 17496 4252 17524
rect 3651 17493 3663 17496
rect 3605 17487 3663 17493
rect 4246 17484 4252 17496
rect 4304 17484 4310 17536
rect 4430 17524 4436 17536
rect 4391 17496 4436 17524
rect 4430 17484 4436 17496
rect 4488 17484 4494 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 4709 17323 4767 17329
rect 4709 17289 4721 17323
rect 4755 17320 4767 17323
rect 4982 17320 4988 17332
rect 4755 17292 4988 17320
rect 4755 17289 4767 17292
rect 4709 17283 4767 17289
rect 4982 17280 4988 17292
rect 5040 17320 5046 17332
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 5040 17292 5641 17320
rect 5040 17280 5046 17292
rect 5629 17289 5641 17292
rect 5675 17289 5687 17323
rect 5629 17283 5687 17289
rect 6273 17323 6331 17329
rect 6273 17289 6285 17323
rect 6319 17320 6331 17323
rect 6730 17320 6736 17332
rect 6319 17292 6736 17320
rect 6319 17289 6331 17292
rect 6273 17283 6331 17289
rect 6730 17280 6736 17292
rect 6788 17280 6794 17332
rect 9217 17323 9275 17329
rect 9217 17289 9229 17323
rect 9263 17320 9275 17323
rect 10042 17320 10048 17332
rect 9263 17292 10048 17320
rect 9263 17289 9275 17292
rect 9217 17283 9275 17289
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 10686 17320 10692 17332
rect 10647 17292 10692 17320
rect 10686 17280 10692 17292
rect 10744 17280 10750 17332
rect 11425 17323 11483 17329
rect 11425 17289 11437 17323
rect 11471 17320 11483 17323
rect 11790 17320 11796 17332
rect 11471 17292 11796 17320
rect 11471 17289 11483 17292
rect 11425 17283 11483 17289
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 12253 17323 12311 17329
rect 12253 17289 12265 17323
rect 12299 17320 12311 17323
rect 12434 17320 12440 17332
rect 12299 17292 12440 17320
rect 12299 17289 12311 17292
rect 12253 17283 12311 17289
rect 12434 17280 12440 17292
rect 12492 17280 12498 17332
rect 2777 17255 2835 17261
rect 2777 17252 2789 17255
rect 2056 17224 2789 17252
rect 2056 17125 2084 17224
rect 2777 17221 2789 17224
rect 2823 17252 2835 17255
rect 3326 17252 3332 17264
rect 2823 17224 3332 17252
rect 2823 17221 2835 17224
rect 2777 17215 2835 17221
rect 3326 17212 3332 17224
rect 3384 17212 3390 17264
rect 2130 17144 2136 17196
rect 2188 17184 2194 17196
rect 2225 17187 2283 17193
rect 2225 17184 2237 17187
rect 2188 17156 2237 17184
rect 2188 17144 2194 17156
rect 2225 17153 2237 17156
rect 2271 17153 2283 17187
rect 2225 17147 2283 17153
rect 5994 17144 6000 17196
rect 6052 17184 6058 17196
rect 6822 17184 6828 17196
rect 6052 17156 6828 17184
rect 6052 17144 6058 17156
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 9306 17184 9312 17196
rect 9267 17156 9312 17184
rect 9306 17144 9312 17156
rect 9364 17144 9370 17196
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 3329 17119 3387 17125
rect 3329 17085 3341 17119
rect 3375 17116 3387 17119
rect 3418 17116 3424 17128
rect 3375 17088 3424 17116
rect 3375 17085 3387 17088
rect 3329 17079 3387 17085
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 11330 17076 11336 17128
rect 11388 17116 11394 17128
rect 11793 17119 11851 17125
rect 11793 17116 11805 17119
rect 11388 17088 11805 17116
rect 11388 17076 11394 17088
rect 11793 17085 11805 17088
rect 11839 17116 11851 17119
rect 12434 17116 12440 17128
rect 11839 17088 12440 17116
rect 11839 17085 11851 17088
rect 11793 17079 11851 17085
rect 12434 17076 12440 17088
rect 12492 17116 12498 17128
rect 12492 17088 12585 17116
rect 12492 17076 12498 17088
rect 3574 17051 3632 17057
rect 3574 17048 3586 17051
rect 3160 17020 3586 17048
rect 3160 16992 3188 17020
rect 3574 17017 3586 17020
rect 3620 17017 3632 17051
rect 3574 17011 3632 17017
rect 6641 17051 6699 17057
rect 6641 17017 6653 17051
rect 6687 17048 6699 17051
rect 7092 17051 7150 17057
rect 7092 17048 7104 17051
rect 6687 17020 7104 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 7092 17017 7104 17020
rect 7138 17048 7150 17051
rect 7374 17048 7380 17060
rect 7138 17020 7380 17048
rect 7138 17017 7150 17020
rect 7092 17011 7150 17017
rect 7374 17008 7380 17020
rect 7432 17008 7438 17060
rect 9582 17057 9588 17060
rect 9576 17011 9588 17057
rect 9640 17048 9646 17060
rect 9640 17020 9676 17048
rect 9582 17008 9588 17011
rect 9640 17008 9646 17020
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 12682 17051 12740 17057
rect 12682 17048 12694 17051
rect 12584 17020 12694 17048
rect 12584 17008 12590 17020
rect 12682 17017 12694 17020
rect 12728 17017 12740 17051
rect 12682 17011 12740 17017
rect 1670 16980 1676 16992
rect 1631 16952 1676 16980
rect 1670 16940 1676 16952
rect 1728 16940 1734 16992
rect 1762 16940 1768 16992
rect 1820 16980 1826 16992
rect 2130 16980 2136 16992
rect 1820 16952 2136 16980
rect 1820 16940 1826 16952
rect 2130 16940 2136 16952
rect 2188 16940 2194 16992
rect 2314 16940 2320 16992
rect 2372 16980 2378 16992
rect 2498 16980 2504 16992
rect 2372 16952 2504 16980
rect 2372 16940 2378 16952
rect 2498 16940 2504 16952
rect 2556 16940 2562 16992
rect 3142 16980 3148 16992
rect 3103 16952 3148 16980
rect 3142 16940 3148 16952
rect 3200 16940 3206 16992
rect 5350 16980 5356 16992
rect 5311 16952 5356 16980
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 7742 16940 7748 16992
rect 7800 16980 7806 16992
rect 8205 16983 8263 16989
rect 8205 16980 8217 16983
rect 7800 16952 8217 16980
rect 7800 16940 7806 16952
rect 8205 16949 8217 16952
rect 8251 16949 8263 16983
rect 8754 16980 8760 16992
rect 8715 16952 8760 16980
rect 8205 16943 8263 16949
rect 8754 16940 8760 16952
rect 8812 16940 8818 16992
rect 13814 16980 13820 16992
rect 13775 16952 13820 16980
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1762 16736 1768 16788
rect 1820 16776 1826 16788
rect 1857 16779 1915 16785
rect 1857 16776 1869 16779
rect 1820 16748 1869 16776
rect 1820 16736 1826 16748
rect 1857 16745 1869 16748
rect 1903 16745 1915 16779
rect 1857 16739 1915 16745
rect 2038 16736 2044 16788
rect 2096 16776 2102 16788
rect 2409 16779 2467 16785
rect 2096 16748 2360 16776
rect 2096 16736 2102 16748
rect 2332 16717 2360 16748
rect 2409 16745 2421 16779
rect 2455 16776 2467 16779
rect 2774 16776 2780 16788
rect 2455 16748 2780 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 2774 16736 2780 16748
rect 2832 16736 2838 16788
rect 4062 16776 4068 16788
rect 4023 16748 4068 16776
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 4430 16736 4436 16788
rect 4488 16776 4494 16788
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 4488 16748 4537 16776
rect 4488 16736 4494 16748
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 4525 16739 4583 16745
rect 4614 16736 4620 16788
rect 4672 16776 4678 16788
rect 5169 16779 5227 16785
rect 5169 16776 5181 16779
rect 4672 16748 5181 16776
rect 4672 16736 4678 16748
rect 5169 16745 5181 16748
rect 5215 16776 5227 16779
rect 5258 16776 5264 16788
rect 5215 16748 5264 16776
rect 5215 16745 5227 16748
rect 5169 16739 5227 16745
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 5905 16779 5963 16785
rect 5905 16745 5917 16779
rect 5951 16776 5963 16779
rect 5994 16776 6000 16788
rect 5951 16748 6000 16776
rect 5951 16745 5963 16748
rect 5905 16739 5963 16745
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 6454 16776 6460 16788
rect 6415 16748 6460 16776
rect 6454 16736 6460 16748
rect 6512 16736 6518 16788
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 7837 16779 7895 16785
rect 7837 16776 7849 16779
rect 6880 16748 7849 16776
rect 6880 16736 6886 16748
rect 7837 16745 7849 16748
rect 7883 16745 7895 16779
rect 8018 16776 8024 16788
rect 7979 16748 8024 16776
rect 7837 16739 7895 16745
rect 1397 16711 1455 16717
rect 1397 16677 1409 16711
rect 1443 16708 1455 16711
rect 2317 16711 2375 16717
rect 1443 16680 2176 16708
rect 1443 16677 1455 16680
rect 1397 16671 1455 16677
rect 2148 16640 2176 16680
rect 2317 16677 2329 16711
rect 2363 16677 2375 16711
rect 2317 16671 2375 16677
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 3786 16708 3792 16720
rect 2648 16680 2912 16708
rect 3747 16680 3792 16708
rect 2648 16668 2654 16680
rect 2406 16640 2412 16652
rect 2148 16612 2412 16640
rect 2406 16600 2412 16612
rect 2464 16640 2470 16652
rect 2884 16649 2912 16680
rect 3786 16668 3792 16680
rect 3844 16668 3850 16720
rect 4448 16708 4476 16736
rect 4172 16680 4476 16708
rect 6365 16711 6423 16717
rect 2777 16643 2835 16649
rect 2777 16640 2789 16643
rect 2464 16612 2789 16640
rect 2464 16600 2470 16612
rect 2777 16609 2789 16612
rect 2823 16609 2835 16643
rect 2777 16603 2835 16609
rect 2869 16643 2927 16649
rect 2869 16609 2881 16643
rect 2915 16640 2927 16643
rect 3421 16643 3479 16649
rect 3421 16640 3433 16643
rect 2915 16612 3433 16640
rect 2915 16609 2927 16612
rect 2869 16603 2927 16609
rect 3421 16609 3433 16612
rect 3467 16609 3479 16643
rect 3421 16603 3479 16609
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4172 16640 4200 16680
rect 6365 16677 6377 16711
rect 6411 16708 6423 16711
rect 6914 16708 6920 16720
rect 6411 16680 6920 16708
rect 6411 16677 6423 16680
rect 6365 16671 6423 16677
rect 6914 16668 6920 16680
rect 6972 16668 6978 16720
rect 4430 16640 4436 16652
rect 4120 16612 4200 16640
rect 4343 16612 4436 16640
rect 4120 16600 4126 16612
rect 4430 16600 4436 16612
rect 4488 16640 4494 16652
rect 4798 16640 4804 16652
rect 4488 16612 4804 16640
rect 4488 16600 4494 16612
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 5534 16640 5540 16652
rect 5495 16612 5540 16640
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 6638 16600 6644 16652
rect 6696 16640 6702 16652
rect 6825 16643 6883 16649
rect 6825 16640 6837 16643
rect 6696 16612 6837 16640
rect 6696 16600 6702 16612
rect 6825 16609 6837 16612
rect 6871 16609 6883 16643
rect 7852 16640 7880 16739
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 10229 16779 10287 16785
rect 10229 16745 10241 16779
rect 10275 16776 10287 16779
rect 10686 16776 10692 16788
rect 10275 16748 10692 16776
rect 10275 16745 10287 16748
rect 10229 16739 10287 16745
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 11146 16776 11152 16788
rect 11107 16748 11152 16776
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 8389 16711 8447 16717
rect 8389 16708 8401 16711
rect 8352 16680 8401 16708
rect 8352 16668 8358 16680
rect 8389 16677 8401 16680
rect 8435 16708 8447 16711
rect 9677 16711 9735 16717
rect 9677 16708 9689 16711
rect 8435 16680 9689 16708
rect 8435 16677 8447 16680
rect 8389 16671 8447 16677
rect 9677 16677 9689 16680
rect 9723 16677 9735 16711
rect 9677 16671 9735 16677
rect 10597 16711 10655 16717
rect 10597 16677 10609 16711
rect 10643 16708 10655 16711
rect 11330 16708 11336 16720
rect 10643 16680 11336 16708
rect 10643 16677 10655 16680
rect 10597 16671 10655 16677
rect 11330 16668 11336 16680
rect 11388 16668 11394 16720
rect 7852 16612 8248 16640
rect 6825 16603 6883 16609
rect 2314 16532 2320 16584
rect 2372 16572 2378 16584
rect 2961 16575 3019 16581
rect 2961 16572 2973 16575
rect 2372 16544 2973 16572
rect 2372 16532 2378 16544
rect 2961 16541 2973 16544
rect 3007 16572 3019 16575
rect 3142 16572 3148 16584
rect 3007 16544 3148 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 3142 16532 3148 16544
rect 3200 16532 3206 16584
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 5442 16572 5448 16584
rect 4755 16544 5448 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 5442 16532 5448 16544
rect 5500 16532 5506 16584
rect 6546 16532 6552 16584
rect 6604 16572 6610 16584
rect 6917 16575 6975 16581
rect 6917 16572 6929 16575
rect 6604 16544 6929 16572
rect 6604 16532 6610 16544
rect 6917 16541 6929 16544
rect 6963 16541 6975 16575
rect 6917 16535 6975 16541
rect 7009 16575 7067 16581
rect 7009 16541 7021 16575
rect 7055 16541 7067 16575
rect 8220 16572 8248 16612
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 11514 16640 11520 16652
rect 8536 16612 8581 16640
rect 11475 16612 11520 16640
rect 8536 16600 8542 16612
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 8386 16572 8392 16584
rect 8220 16544 8392 16572
rect 7009 16535 7067 16541
rect 6730 16464 6736 16516
rect 6788 16504 6794 16516
rect 7024 16504 7052 16535
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 8662 16572 8668 16584
rect 8575 16544 8668 16572
rect 8662 16532 8668 16544
rect 8720 16572 8726 16584
rect 11606 16572 11612 16584
rect 8720 16544 9444 16572
rect 11567 16544 11612 16572
rect 8720 16532 8726 16544
rect 6788 16476 7052 16504
rect 6788 16464 6794 16476
rect 7466 16436 7472 16448
rect 7427 16408 7472 16436
rect 7466 16396 7472 16408
rect 7524 16396 7530 16448
rect 9416 16445 9444 16544
rect 11606 16532 11612 16544
rect 11664 16532 11670 16584
rect 11790 16572 11796 16584
rect 11751 16544 11796 16572
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 9401 16439 9459 16445
rect 9401 16405 9413 16439
rect 9447 16436 9459 16439
rect 9582 16436 9588 16448
rect 9447 16408 9588 16436
rect 9447 16405 9459 16408
rect 9401 16399 9459 16405
rect 9582 16396 9588 16408
rect 9640 16436 9646 16448
rect 10594 16436 10600 16448
rect 9640 16408 10600 16436
rect 9640 16396 9646 16408
rect 10594 16396 10600 16408
rect 10652 16396 10658 16448
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 12529 16439 12587 16445
rect 12529 16436 12541 16439
rect 12492 16408 12541 16436
rect 12492 16396 12498 16408
rect 12529 16405 12541 16408
rect 12575 16436 12587 16439
rect 12618 16436 12624 16448
rect 12575 16408 12624 16436
rect 12575 16405 12587 16408
rect 12529 16399 12587 16405
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2406 16232 2412 16244
rect 2367 16204 2412 16232
rect 2406 16192 2412 16204
rect 2464 16192 2470 16244
rect 4430 16192 4436 16244
rect 4488 16232 4494 16244
rect 4617 16235 4675 16241
rect 4617 16232 4629 16235
rect 4488 16204 4629 16232
rect 4488 16192 4494 16204
rect 4617 16201 4629 16204
rect 4663 16201 4675 16235
rect 4617 16195 4675 16201
rect 5077 16235 5135 16241
rect 5077 16201 5089 16235
rect 5123 16232 5135 16235
rect 5442 16232 5448 16244
rect 5123 16204 5448 16232
rect 5123 16201 5135 16204
rect 5077 16195 5135 16201
rect 5442 16192 5448 16204
rect 5500 16192 5506 16244
rect 6822 16232 6828 16244
rect 6783 16204 6828 16232
rect 6822 16192 6828 16204
rect 6880 16192 6886 16244
rect 8294 16232 8300 16244
rect 8255 16204 8300 16232
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 8662 16232 8668 16244
rect 8623 16204 8668 16232
rect 8662 16192 8668 16204
rect 8720 16192 8726 16244
rect 10594 16232 10600 16244
rect 10555 16204 10600 16232
rect 10594 16192 10600 16204
rect 10652 16192 10658 16244
rect 11514 16232 11520 16244
rect 11475 16204 11520 16232
rect 11514 16192 11520 16204
rect 11572 16192 11578 16244
rect 11790 16192 11796 16244
rect 11848 16232 11854 16244
rect 11885 16235 11943 16241
rect 11885 16232 11897 16235
rect 11848 16204 11897 16232
rect 11848 16192 11854 16204
rect 11885 16201 11897 16204
rect 11931 16201 11943 16235
rect 11885 16195 11943 16201
rect 6914 16056 6920 16108
rect 6972 16096 6978 16108
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 6972 16068 7297 16096
rect 6972 16056 6978 16068
rect 7285 16065 7297 16068
rect 7331 16065 7343 16099
rect 7466 16096 7472 16108
rect 7427 16068 7472 16096
rect 7285 16059 7343 16065
rect 7466 16056 7472 16068
rect 7524 16056 7530 16108
rect 9122 16056 9128 16108
rect 9180 16096 9186 16108
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 9180 16068 9229 16096
rect 9180 16056 9186 16068
rect 9217 16065 9229 16068
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1578 16028 1584 16040
rect 1443 16000 1584 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 2685 16031 2743 16037
rect 2685 15997 2697 16031
rect 2731 16028 2743 16031
rect 3418 16028 3424 16040
rect 2731 16000 3424 16028
rect 2731 15997 2743 16000
rect 2685 15991 2743 15997
rect 3418 15988 3424 16000
rect 3476 15988 3482 16040
rect 5169 16031 5227 16037
rect 5169 15997 5181 16031
rect 5215 16028 5227 16031
rect 5534 16028 5540 16040
rect 5215 16000 5540 16028
rect 5215 15997 5227 16000
rect 5169 15991 5227 15997
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 1673 15963 1731 15969
rect 1673 15929 1685 15963
rect 1719 15960 1731 15963
rect 2406 15960 2412 15972
rect 1719 15932 2412 15960
rect 1719 15929 1731 15932
rect 1673 15923 1731 15929
rect 2406 15920 2412 15932
rect 2464 15920 2470 15972
rect 2952 15963 3010 15969
rect 2952 15929 2964 15963
rect 2998 15960 3010 15963
rect 3050 15960 3056 15972
rect 2998 15932 3056 15960
rect 2998 15929 3010 15932
rect 2952 15923 3010 15929
rect 3050 15920 3056 15932
rect 3108 15920 3114 15972
rect 5442 15960 5448 15972
rect 5403 15932 5448 15960
rect 5442 15920 5448 15932
rect 5500 15920 5506 15972
rect 7190 15960 7196 15972
rect 7103 15932 7196 15960
rect 7190 15920 7196 15932
rect 7248 15960 7254 15972
rect 7837 15963 7895 15969
rect 7837 15960 7849 15963
rect 7248 15932 7849 15960
rect 7248 15920 7254 15932
rect 7837 15929 7849 15932
rect 7883 15929 7895 15963
rect 7837 15923 7895 15929
rect 9125 15963 9183 15969
rect 9125 15929 9137 15963
rect 9171 15960 9183 15963
rect 9462 15963 9520 15969
rect 9462 15960 9474 15963
rect 9171 15932 9474 15960
rect 9171 15929 9183 15932
rect 9125 15923 9183 15929
rect 9462 15929 9474 15932
rect 9508 15960 9520 15963
rect 10134 15960 10140 15972
rect 9508 15932 10140 15960
rect 9508 15929 9520 15932
rect 9462 15923 9520 15929
rect 10134 15920 10140 15932
rect 10192 15920 10198 15972
rect 3142 15852 3148 15904
rect 3200 15892 3206 15904
rect 4065 15895 4123 15901
rect 4065 15892 4077 15895
rect 3200 15864 4077 15892
rect 3200 15852 3206 15864
rect 4065 15861 4077 15864
rect 4111 15861 4123 15895
rect 6086 15892 6092 15904
rect 6047 15864 6092 15892
rect 4065 15855 4123 15861
rect 6086 15852 6092 15864
rect 6144 15852 6150 15904
rect 6546 15892 6552 15904
rect 6507 15864 6552 15892
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 11241 15895 11299 15901
rect 11241 15861 11253 15895
rect 11287 15892 11299 15895
rect 11514 15892 11520 15904
rect 11287 15864 11520 15892
rect 11287 15861 11299 15864
rect 11241 15855 11299 15861
rect 11514 15852 11520 15864
rect 11572 15852 11578 15904
rect 11974 15852 11980 15904
rect 12032 15892 12038 15904
rect 12437 15895 12495 15901
rect 12437 15892 12449 15895
rect 12032 15864 12449 15892
rect 12032 15852 12038 15864
rect 12437 15861 12449 15864
rect 12483 15861 12495 15895
rect 12437 15855 12495 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1394 15688 1400 15700
rect 1355 15660 1400 15688
rect 1394 15648 1400 15660
rect 1452 15648 1458 15700
rect 2314 15688 2320 15700
rect 2275 15660 2320 15688
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 2409 15691 2467 15697
rect 2409 15657 2421 15691
rect 2455 15688 2467 15691
rect 2590 15688 2596 15700
rect 2455 15660 2596 15688
rect 2455 15657 2467 15660
rect 2409 15651 2467 15657
rect 2590 15648 2596 15660
rect 2648 15648 2654 15700
rect 3881 15691 3939 15697
rect 3881 15657 3893 15691
rect 3927 15688 3939 15691
rect 4062 15688 4068 15700
rect 3927 15660 4068 15688
rect 3927 15657 3939 15660
rect 3881 15651 3939 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 6549 15691 6607 15697
rect 6549 15657 6561 15691
rect 6595 15688 6607 15691
rect 6730 15688 6736 15700
rect 6595 15660 6736 15688
rect 6595 15657 6607 15660
rect 6549 15651 6607 15657
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7101 15691 7159 15697
rect 7101 15688 7113 15691
rect 6972 15660 7113 15688
rect 6972 15648 6978 15660
rect 7101 15657 7113 15660
rect 7147 15657 7159 15691
rect 7101 15651 7159 15657
rect 8205 15691 8263 15697
rect 8205 15657 8217 15691
rect 8251 15688 8263 15691
rect 8478 15688 8484 15700
rect 8251 15660 8484 15688
rect 8251 15657 8263 15660
rect 8205 15651 8263 15657
rect 8478 15648 8484 15660
rect 8536 15688 8542 15700
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 8536 15660 9689 15688
rect 8536 15648 8542 15660
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 9677 15651 9735 15657
rect 10778 15648 10784 15700
rect 10836 15688 10842 15700
rect 11609 15691 11667 15697
rect 11609 15688 11621 15691
rect 10836 15660 11621 15688
rect 10836 15648 10842 15660
rect 11609 15657 11621 15660
rect 11655 15657 11667 15691
rect 11974 15688 11980 15700
rect 11935 15660 11980 15688
rect 11609 15651 11667 15657
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 12710 15688 12716 15700
rect 12623 15660 12716 15688
rect 12710 15648 12716 15660
rect 12768 15688 12774 15700
rect 13722 15688 13728 15700
rect 12768 15660 13728 15688
rect 12768 15648 12774 15660
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 4246 15580 4252 15632
rect 4304 15629 4310 15632
rect 4304 15623 4368 15629
rect 4304 15589 4322 15623
rect 4356 15589 4368 15623
rect 4304 15583 4368 15589
rect 4304 15580 4310 15583
rect 2774 15552 2780 15564
rect 2735 15524 2780 15552
rect 2774 15512 2780 15524
rect 2832 15512 2838 15564
rect 6181 15555 6239 15561
rect 6181 15521 6193 15555
rect 6227 15552 6239 15555
rect 7009 15555 7067 15561
rect 7009 15552 7021 15555
rect 6227 15524 7021 15552
rect 6227 15521 6239 15524
rect 6181 15515 6239 15521
rect 7009 15521 7021 15524
rect 7055 15521 7067 15555
rect 7009 15515 7067 15521
rect 2866 15484 2872 15496
rect 2827 15456 2872 15484
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 3050 15484 3056 15496
rect 2963 15456 3056 15484
rect 3050 15444 3056 15456
rect 3108 15484 3114 15496
rect 4062 15484 4068 15496
rect 3108 15456 3556 15484
rect 4023 15456 4068 15484
rect 3108 15444 3114 15456
rect 1949 15351 2007 15357
rect 1949 15317 1961 15351
rect 1995 15348 2007 15351
rect 2590 15348 2596 15360
rect 1995 15320 2596 15348
rect 1995 15317 2007 15320
rect 1949 15311 2007 15317
rect 2590 15308 2596 15320
rect 2648 15308 2654 15360
rect 3528 15357 3556 15456
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 7024 15416 7052 15515
rect 7374 15512 7380 15564
rect 7432 15552 7438 15564
rect 7469 15555 7527 15561
rect 7469 15552 7481 15555
rect 7432 15524 7481 15552
rect 7432 15512 7438 15524
rect 7469 15521 7481 15524
rect 7515 15521 7527 15555
rect 7469 15515 7527 15521
rect 9950 15512 9956 15564
rect 10008 15552 10014 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 10008 15524 10057 15552
rect 10008 15512 10014 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 11422 15552 11428 15564
rect 11383 15524 11428 15552
rect 10045 15515 10103 15521
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 7558 15484 7564 15496
rect 7519 15456 7564 15484
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 7742 15484 7748 15496
rect 7703 15456 7748 15484
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 10134 15484 10140 15496
rect 10095 15456 10140 15484
rect 10134 15444 10140 15456
rect 10192 15444 10198 15496
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 12066 15484 12072 15496
rect 10284 15456 10329 15484
rect 12027 15456 12072 15484
rect 10284 15444 10290 15456
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 12250 15484 12256 15496
rect 12211 15456 12256 15484
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 8938 15416 8944 15428
rect 7024 15388 8944 15416
rect 8938 15376 8944 15388
rect 8996 15376 9002 15428
rect 3513 15351 3571 15357
rect 3513 15317 3525 15351
rect 3559 15348 3571 15351
rect 5445 15351 5503 15357
rect 5445 15348 5457 15351
rect 3559 15320 5457 15348
rect 3559 15317 3571 15320
rect 3513 15311 3571 15317
rect 5445 15317 5457 15320
rect 5491 15317 5503 15351
rect 6822 15348 6828 15360
rect 6783 15320 6828 15348
rect 5445 15311 5503 15317
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 8478 15348 8484 15360
rect 8439 15320 8484 15348
rect 8478 15308 8484 15320
rect 8536 15308 8542 15360
rect 9033 15351 9091 15357
rect 9033 15317 9045 15351
rect 9079 15348 9091 15351
rect 9122 15348 9128 15360
rect 9079 15320 9128 15348
rect 9079 15317 9091 15320
rect 9033 15311 9091 15317
rect 9122 15308 9128 15320
rect 9180 15308 9186 15360
rect 9401 15351 9459 15357
rect 9401 15317 9413 15351
rect 9447 15348 9459 15351
rect 9490 15348 9496 15360
rect 9447 15320 9496 15348
rect 9447 15317 9459 15320
rect 9401 15311 9459 15317
rect 9490 15308 9496 15320
rect 9548 15308 9554 15360
rect 11241 15351 11299 15357
rect 11241 15317 11253 15351
rect 11287 15348 11299 15351
rect 12618 15348 12624 15360
rect 11287 15320 12624 15348
rect 11287 15317 11299 15320
rect 11241 15311 11299 15317
rect 12618 15308 12624 15320
rect 12676 15348 12682 15360
rect 12989 15351 13047 15357
rect 12989 15348 13001 15351
rect 12676 15320 13001 15348
rect 12676 15308 12682 15320
rect 12989 15317 13001 15320
rect 13035 15317 13047 15351
rect 12989 15311 13047 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2498 15104 2504 15156
rect 2556 15144 2562 15156
rect 2685 15147 2743 15153
rect 2685 15144 2697 15147
rect 2556 15116 2697 15144
rect 2556 15104 2562 15116
rect 2685 15113 2697 15116
rect 2731 15113 2743 15147
rect 2685 15107 2743 15113
rect 3789 15147 3847 15153
rect 3789 15113 3801 15147
rect 3835 15144 3847 15147
rect 4157 15147 4215 15153
rect 4157 15144 4169 15147
rect 3835 15116 4169 15144
rect 3835 15113 3847 15116
rect 3789 15107 3847 15113
rect 4157 15113 4169 15116
rect 4203 15144 4215 15147
rect 4246 15144 4252 15156
rect 4203 15116 4252 15144
rect 4203 15113 4215 15116
rect 4157 15107 4215 15113
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 2682 15008 2688 15020
rect 1719 14980 2688 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 3329 15011 3387 15017
rect 3329 14977 3341 15011
rect 3375 15008 3387 15011
rect 3804 15008 3832 15107
rect 4246 15104 4252 15116
rect 4304 15144 4310 15156
rect 5629 15147 5687 15153
rect 5629 15144 5641 15147
rect 4304 15116 5641 15144
rect 4304 15104 4310 15116
rect 5629 15113 5641 15116
rect 5675 15113 5687 15147
rect 6270 15144 6276 15156
rect 6231 15116 6276 15144
rect 5629 15107 5687 15113
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 7466 15104 7472 15156
rect 7524 15144 7530 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 7524 15116 8217 15144
rect 7524 15104 7530 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8205 15107 8263 15113
rect 10226 15104 10232 15156
rect 10284 15144 10290 15156
rect 10689 15147 10747 15153
rect 10689 15144 10701 15147
rect 10284 15116 10701 15144
rect 10284 15104 10290 15116
rect 10689 15113 10701 15116
rect 10735 15144 10747 15147
rect 11241 15147 11299 15153
rect 11241 15144 11253 15147
rect 10735 15116 11253 15144
rect 10735 15113 10747 15116
rect 10689 15107 10747 15113
rect 11241 15113 11253 15116
rect 11287 15113 11299 15147
rect 11241 15107 11299 15113
rect 11701 15147 11759 15153
rect 11701 15113 11713 15147
rect 11747 15144 11759 15147
rect 11974 15144 11980 15156
rect 11747 15116 11980 15144
rect 11747 15113 11759 15116
rect 11701 15107 11759 15113
rect 11974 15104 11980 15116
rect 12032 15104 12038 15156
rect 3375 14980 3832 15008
rect 3375 14977 3387 14980
rect 3329 14971 3387 14977
rect 4154 14968 4160 15020
rect 4212 15008 4218 15020
rect 4249 15011 4307 15017
rect 4249 15008 4261 15011
rect 4212 14980 4261 15008
rect 4212 14968 4218 14980
rect 4249 14977 4261 14980
rect 4295 14977 4307 15011
rect 9214 15008 9220 15020
rect 9175 14980 9220 15008
rect 4249 14971 4307 14977
rect 1394 14940 1400 14952
rect 1355 14912 1400 14940
rect 1394 14900 1400 14912
rect 1452 14900 1458 14952
rect 4264 14940 4292 14971
rect 9214 14968 9220 14980
rect 9272 14968 9278 15020
rect 6822 14940 6828 14952
rect 4264 14912 6828 14940
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 12710 14949 12716 14952
rect 9309 14943 9367 14949
rect 9309 14940 9321 14943
rect 9180 14912 9321 14940
rect 9180 14900 9186 14912
rect 9309 14909 9321 14912
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 12704 14940 12716 14949
rect 12671 14912 12716 14940
rect 12437 14903 12495 14909
rect 12704 14903 12716 14912
rect 2774 14832 2780 14884
rect 2832 14872 2838 14884
rect 4522 14881 4528 14884
rect 3145 14875 3203 14881
rect 3145 14872 3157 14875
rect 2832 14844 3157 14872
rect 2832 14832 2838 14844
rect 3145 14841 3157 14844
rect 3191 14841 3203 14875
rect 4516 14872 4528 14881
rect 4483 14844 4528 14872
rect 3145 14835 3203 14841
rect 4516 14835 4528 14844
rect 2498 14804 2504 14816
rect 2459 14776 2504 14804
rect 2498 14764 2504 14776
rect 2556 14764 2562 14816
rect 2958 14764 2964 14816
rect 3016 14804 3022 14816
rect 3053 14807 3111 14813
rect 3053 14804 3065 14807
rect 3016 14776 3065 14804
rect 3016 14764 3022 14776
rect 3053 14773 3065 14776
rect 3099 14773 3111 14807
rect 3160 14804 3188 14835
rect 4522 14832 4528 14835
rect 4580 14832 4586 14884
rect 6730 14832 6736 14884
rect 6788 14872 6794 14884
rect 7092 14875 7150 14881
rect 7092 14872 7104 14875
rect 6788 14844 7104 14872
rect 6788 14832 6794 14844
rect 7092 14841 7104 14844
rect 7138 14872 7150 14875
rect 7742 14872 7748 14884
rect 7138 14844 7748 14872
rect 7138 14841 7150 14844
rect 7092 14835 7150 14841
rect 7742 14832 7748 14844
rect 7800 14832 7806 14884
rect 8386 14832 8392 14884
rect 8444 14872 8450 14884
rect 9490 14872 9496 14884
rect 8444 14844 9496 14872
rect 8444 14832 8450 14844
rect 9490 14832 9496 14844
rect 9548 14881 9554 14884
rect 9548 14875 9612 14881
rect 9548 14841 9566 14875
rect 9600 14841 9612 14875
rect 12452 14872 12480 14903
rect 12710 14900 12716 14903
rect 12768 14900 12774 14952
rect 12618 14872 12624 14884
rect 12452 14844 12624 14872
rect 9548 14835 9612 14841
rect 9548 14832 9554 14835
rect 12618 14832 12624 14844
rect 12676 14832 12682 14884
rect 4890 14804 4896 14816
rect 3160 14776 4896 14804
rect 3053 14767 3111 14773
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 6638 14804 6644 14816
rect 6599 14776 6644 14804
rect 6638 14764 6644 14776
rect 6696 14764 6702 14816
rect 8846 14804 8852 14816
rect 8759 14776 8852 14804
rect 8846 14764 8852 14776
rect 8904 14804 8910 14816
rect 9950 14804 9956 14816
rect 8904 14776 9956 14804
rect 8904 14764 8910 14776
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 12069 14807 12127 14813
rect 12069 14773 12081 14807
rect 12115 14804 12127 14807
rect 12250 14804 12256 14816
rect 12115 14776 12256 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 12250 14764 12256 14776
rect 12308 14804 12314 14816
rect 12802 14804 12808 14816
rect 12308 14776 12808 14804
rect 12308 14764 12314 14776
rect 12802 14764 12808 14776
rect 12860 14804 12866 14816
rect 13817 14807 13875 14813
rect 13817 14804 13829 14807
rect 12860 14776 13829 14804
rect 12860 14764 12866 14776
rect 13817 14773 13829 14776
rect 13863 14773 13875 14807
rect 13817 14767 13875 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1394 14560 1400 14612
rect 1452 14600 1458 14612
rect 1489 14603 1547 14609
rect 1489 14600 1501 14603
rect 1452 14572 1501 14600
rect 1452 14560 1458 14572
rect 1489 14569 1501 14572
rect 1535 14600 1547 14603
rect 4617 14603 4675 14609
rect 4617 14600 4629 14603
rect 1535 14572 4629 14600
rect 1535 14569 1547 14572
rect 1489 14563 1547 14569
rect 4617 14569 4629 14572
rect 4663 14569 4675 14603
rect 4890 14600 4896 14612
rect 4851 14572 4896 14600
rect 4617 14563 4675 14569
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 6273 14603 6331 14609
rect 6273 14569 6285 14603
rect 6319 14600 6331 14603
rect 6641 14603 6699 14609
rect 6641 14600 6653 14603
rect 6319 14572 6653 14600
rect 6319 14569 6331 14572
rect 6273 14563 6331 14569
rect 6641 14569 6653 14572
rect 6687 14600 6699 14603
rect 6730 14600 6736 14612
rect 6687 14572 6736 14600
rect 6687 14569 6699 14572
rect 6641 14563 6699 14569
rect 6730 14560 6736 14572
rect 6788 14560 6794 14612
rect 8478 14560 8484 14612
rect 8536 14600 8542 14612
rect 8665 14603 8723 14609
rect 8665 14600 8677 14603
rect 8536 14572 8677 14600
rect 8536 14560 8542 14572
rect 8665 14569 8677 14572
rect 8711 14569 8723 14603
rect 11146 14600 11152 14612
rect 11107 14572 11152 14600
rect 8665 14563 8723 14569
rect 11146 14560 11152 14572
rect 11204 14560 11210 14612
rect 11793 14603 11851 14609
rect 11793 14569 11805 14603
rect 11839 14600 11851 14603
rect 12066 14600 12072 14612
rect 11839 14572 12072 14600
rect 11839 14569 11851 14572
rect 11793 14563 11851 14569
rect 12066 14560 12072 14572
rect 12124 14560 12130 14612
rect 12618 14560 12624 14612
rect 12676 14560 12682 14612
rect 1946 14532 1952 14544
rect 1907 14504 1952 14532
rect 1946 14492 1952 14504
rect 2004 14492 2010 14544
rect 2314 14492 2320 14544
rect 2372 14532 2378 14544
rect 2501 14535 2559 14541
rect 2501 14532 2513 14535
rect 2372 14504 2513 14532
rect 2372 14492 2378 14504
rect 2501 14501 2513 14504
rect 2547 14501 2559 14535
rect 2501 14495 2559 14501
rect 3050 14492 3056 14544
rect 3108 14532 3114 14544
rect 3237 14535 3295 14541
rect 3237 14532 3249 14535
rect 3108 14504 3249 14532
rect 3108 14492 3114 14504
rect 3237 14501 3249 14504
rect 3283 14501 3295 14535
rect 3237 14495 3295 14501
rect 7000 14535 7058 14541
rect 7000 14501 7012 14535
rect 7046 14532 7058 14535
rect 7466 14532 7472 14544
rect 7046 14504 7472 14532
rect 7046 14501 7058 14504
rect 7000 14495 7058 14501
rect 7466 14492 7472 14504
rect 7524 14492 7530 14544
rect 8938 14492 8944 14544
rect 8996 14532 9002 14544
rect 8996 14504 11468 14532
rect 8996 14492 9002 14504
rect 1670 14424 1676 14476
rect 1728 14464 1734 14476
rect 1857 14467 1915 14473
rect 1857 14464 1869 14467
rect 1728 14436 1869 14464
rect 1728 14424 1734 14436
rect 1857 14433 1869 14436
rect 1903 14433 1915 14467
rect 1964 14464 1992 14492
rect 11440 14476 11468 14504
rect 3605 14467 3663 14473
rect 3605 14464 3617 14467
rect 1964 14436 3617 14464
rect 1857 14427 1915 14433
rect 3605 14433 3617 14436
rect 3651 14433 3663 14467
rect 5258 14464 5264 14476
rect 5219 14436 5264 14464
rect 3605 14427 3663 14433
rect 1872 14328 1900 14427
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14464 6791 14467
rect 6822 14464 6828 14476
rect 6779 14436 6828 14464
rect 6779 14433 6791 14436
rect 6733 14427 6791 14433
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 10042 14473 10048 14476
rect 9401 14467 9459 14473
rect 9401 14464 9413 14467
rect 9088 14436 9413 14464
rect 9088 14424 9094 14436
rect 9401 14433 9413 14436
rect 9447 14433 9459 14467
rect 10036 14464 10048 14473
rect 10003 14436 10048 14464
rect 9401 14427 9459 14433
rect 10036 14427 10048 14436
rect 10042 14424 10048 14427
rect 10100 14424 10106 14476
rect 11422 14424 11428 14476
rect 11480 14464 11486 14476
rect 12069 14467 12127 14473
rect 12069 14464 12081 14467
rect 11480 14436 12081 14464
rect 11480 14424 11486 14436
rect 12069 14433 12081 14436
rect 12115 14433 12127 14467
rect 12069 14427 12127 14433
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 12636 14464 12664 14560
rect 12704 14535 12762 14541
rect 12704 14501 12716 14535
rect 12750 14532 12762 14535
rect 12802 14532 12808 14544
rect 12750 14504 12808 14532
rect 12750 14501 12762 14504
rect 12704 14495 12762 14501
rect 12802 14492 12808 14504
rect 12860 14492 12866 14544
rect 13446 14464 13452 14476
rect 12483 14436 13452 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 3234 14396 3240 14408
rect 2179 14368 3240 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 5350 14396 5356 14408
rect 5311 14368 5356 14396
rect 5350 14356 5356 14368
rect 5408 14356 5414 14408
rect 5537 14399 5595 14405
rect 5537 14365 5549 14399
rect 5583 14396 5595 14399
rect 6178 14396 6184 14408
rect 5583 14368 6184 14396
rect 5583 14365 5595 14368
rect 5537 14359 5595 14365
rect 2406 14328 2412 14340
rect 1872 14300 2412 14328
rect 2406 14288 2412 14300
rect 2464 14288 2470 14340
rect 4341 14331 4399 14337
rect 4341 14297 4353 14331
rect 4387 14328 4399 14331
rect 4522 14328 4528 14340
rect 4387 14300 4528 14328
rect 4387 14297 4399 14300
rect 4341 14291 4399 14297
rect 4522 14288 4528 14300
rect 4580 14328 4586 14340
rect 5552 14328 5580 14359
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 9122 14396 9128 14408
rect 9035 14368 9128 14396
rect 9122 14356 9128 14368
rect 9180 14396 9186 14408
rect 9766 14396 9772 14408
rect 9180 14368 9772 14396
rect 9180 14356 9186 14368
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 4580 14300 5580 14328
rect 4580 14288 4586 14300
rect 8938 14288 8944 14340
rect 8996 14328 9002 14340
rect 9217 14331 9275 14337
rect 9217 14328 9229 14331
rect 8996 14300 9229 14328
rect 8996 14288 9002 14300
rect 9217 14297 9229 14300
rect 9263 14297 9275 14331
rect 9217 14291 9275 14297
rect 1394 14220 1400 14272
rect 1452 14260 1458 14272
rect 2869 14263 2927 14269
rect 2869 14260 2881 14263
rect 1452 14232 2881 14260
rect 1452 14220 1458 14232
rect 2869 14229 2881 14232
rect 2915 14260 2927 14263
rect 2958 14260 2964 14272
rect 2915 14232 2964 14260
rect 2915 14229 2927 14232
rect 2869 14223 2927 14229
rect 2958 14220 2964 14232
rect 3016 14220 3022 14272
rect 7742 14220 7748 14272
rect 7800 14260 7806 14272
rect 8113 14263 8171 14269
rect 8113 14260 8125 14263
rect 7800 14232 8125 14260
rect 7800 14220 7806 14232
rect 8113 14229 8125 14232
rect 8159 14229 8171 14263
rect 8113 14223 8171 14229
rect 13817 14263 13875 14269
rect 13817 14229 13829 14263
rect 13863 14260 13875 14263
rect 13906 14260 13912 14272
rect 13863 14232 13912 14260
rect 13863 14229 13875 14232
rect 13817 14223 13875 14229
rect 13906 14220 13912 14232
rect 13964 14220 13970 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1854 14056 1860 14068
rect 1815 14028 1860 14056
rect 1854 14016 1860 14028
rect 1912 14016 1918 14068
rect 3234 14056 3240 14068
rect 3195 14028 3240 14056
rect 3234 14016 3240 14028
rect 3292 14016 3298 14068
rect 4249 14059 4307 14065
rect 4249 14025 4261 14059
rect 4295 14056 4307 14059
rect 4338 14056 4344 14068
rect 4295 14028 4344 14056
rect 4295 14025 4307 14028
rect 4249 14019 4307 14025
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 6546 14056 6552 14068
rect 6507 14028 6552 14056
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 7006 14056 7012 14068
rect 6967 14028 7012 14056
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7466 14056 7472 14068
rect 7427 14028 7472 14056
rect 7466 14016 7472 14028
rect 7524 14016 7530 14068
rect 7926 14056 7932 14068
rect 7887 14028 7932 14056
rect 7926 14016 7932 14028
rect 7984 14016 7990 14068
rect 9030 14016 9036 14068
rect 9088 14056 9094 14068
rect 10873 14059 10931 14065
rect 10873 14056 10885 14059
rect 9088 14028 10885 14056
rect 9088 14016 9094 14028
rect 10873 14025 10885 14028
rect 10919 14025 10931 14059
rect 10873 14019 10931 14025
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 12437 14059 12495 14065
rect 12437 14056 12449 14059
rect 12124 14028 12449 14056
rect 12124 14016 12130 14028
rect 12437 14025 12449 14028
rect 12483 14025 12495 14059
rect 13446 14056 13452 14068
rect 13407 14028 13452 14056
rect 12437 14019 12495 14025
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 2777 13991 2835 13997
rect 2777 13957 2789 13991
rect 2823 13988 2835 13991
rect 2961 13991 3019 13997
rect 2961 13988 2973 13991
rect 2823 13960 2973 13988
rect 2823 13957 2835 13960
rect 2777 13951 2835 13957
rect 2961 13957 2973 13960
rect 3007 13988 3019 13991
rect 4798 13988 4804 14000
rect 3007 13960 4804 13988
rect 3007 13957 3019 13960
rect 2961 13951 3019 13957
rect 4798 13948 4804 13960
rect 4856 13988 4862 14000
rect 6270 13988 6276 14000
rect 4856 13960 6276 13988
rect 4856 13948 4862 13960
rect 6270 13948 6276 13960
rect 6328 13948 6334 14000
rect 11422 13988 11428 14000
rect 9968 13960 11428 13988
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 2314 13920 2320 13932
rect 1811 13892 2320 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13920 2559 13923
rect 2682 13920 2688 13932
rect 2547 13892 2688 13920
rect 2547 13889 2559 13892
rect 2501 13883 2559 13889
rect 2682 13880 2688 13892
rect 2740 13920 2746 13932
rect 3605 13923 3663 13929
rect 3605 13920 3617 13923
rect 2740 13892 3617 13920
rect 2740 13880 2746 13892
rect 3605 13889 3617 13892
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13920 4215 13923
rect 4893 13923 4951 13929
rect 4893 13920 4905 13923
rect 4203 13892 4905 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 4893 13889 4905 13892
rect 4939 13920 4951 13923
rect 5074 13920 5080 13932
rect 4939 13892 5080 13920
rect 4939 13889 4951 13892
rect 4893 13883 4951 13889
rect 5074 13880 5080 13892
rect 5132 13880 5138 13932
rect 5258 13920 5264 13932
rect 5184 13892 5264 13920
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13821 2835 13855
rect 2777 13815 2835 13821
rect 2225 13787 2283 13793
rect 2225 13753 2237 13787
rect 2271 13784 2283 13787
rect 2792 13784 2820 13815
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 5184 13852 5212 13892
rect 5258 13880 5264 13892
rect 5316 13920 5322 13932
rect 5718 13920 5724 13932
rect 5316 13892 5724 13920
rect 5316 13880 5322 13892
rect 5718 13880 5724 13892
rect 5776 13880 5782 13932
rect 8386 13880 8392 13932
rect 8444 13920 8450 13932
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 8444 13892 8493 13920
rect 8444 13880 8450 13892
rect 8481 13889 8493 13892
rect 8527 13889 8539 13923
rect 8938 13920 8944 13932
rect 8899 13892 8944 13920
rect 8481 13883 8539 13889
rect 8938 13880 8944 13892
rect 8996 13880 9002 13932
rect 9968 13929 9996 13960
rect 11422 13948 11428 13960
rect 11480 13948 11486 14000
rect 11885 13991 11943 13997
rect 11885 13957 11897 13991
rect 11931 13988 11943 13991
rect 12250 13988 12256 14000
rect 11931 13960 12256 13988
rect 11931 13957 11943 13960
rect 11885 13951 11943 13957
rect 12250 13948 12256 13960
rect 12308 13948 12314 14000
rect 24213 13991 24271 13997
rect 24213 13957 24225 13991
rect 24259 13988 24271 13991
rect 24854 13988 24860 14000
rect 24259 13960 24860 13988
rect 24259 13957 24271 13960
rect 24213 13951 24271 13957
rect 24854 13948 24860 13960
rect 24912 13948 24918 14000
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 9953 13923 10011 13929
rect 9953 13920 9965 13923
rect 9447 13892 9965 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 9953 13889 9965 13892
rect 9999 13889 10011 13923
rect 9953 13883 10011 13889
rect 10042 13880 10048 13932
rect 10100 13920 10106 13932
rect 10137 13923 10195 13929
rect 10137 13920 10149 13923
rect 10100 13892 10149 13920
rect 10100 13880 10106 13892
rect 10137 13889 10149 13892
rect 10183 13920 10195 13923
rect 10183 13892 10640 13920
rect 10183 13889 10195 13892
rect 10137 13883 10195 13889
rect 5350 13852 5356 13864
rect 4120 13824 5212 13852
rect 5311 13824 5356 13852
rect 4120 13812 4126 13824
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 6546 13812 6552 13864
rect 6604 13852 6610 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6604 13824 6837 13852
rect 6604 13812 6610 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8956 13852 8984 13880
rect 7883 13824 8340 13852
rect 8956 13824 9628 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 2271 13756 2820 13784
rect 2271 13753 2283 13756
rect 2225 13747 2283 13753
rect 8312 13728 8340 13824
rect 8389 13787 8447 13793
rect 8389 13753 8401 13787
rect 8435 13784 8447 13787
rect 9600 13784 9628 13824
rect 9861 13787 9919 13793
rect 9861 13784 9873 13787
rect 8435 13756 9536 13784
rect 9600 13756 9873 13784
rect 8435 13753 8447 13756
rect 8389 13747 8447 13753
rect 9508 13728 9536 13756
rect 9861 13753 9873 13756
rect 9907 13753 9919 13787
rect 9861 13747 9919 13753
rect 4614 13716 4620 13728
rect 4575 13688 4620 13716
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 4706 13676 4712 13728
rect 4764 13716 4770 13728
rect 6089 13719 6147 13725
rect 4764 13688 4809 13716
rect 4764 13676 4770 13688
rect 6089 13685 6101 13719
rect 6135 13716 6147 13719
rect 6178 13716 6184 13728
rect 6135 13688 6184 13716
rect 6135 13685 6147 13688
rect 6089 13679 6147 13685
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 8294 13716 8300 13728
rect 8255 13688 8300 13716
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 9490 13716 9496 13728
rect 9451 13688 9496 13716
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 10612 13725 10640 13892
rect 12710 13880 12716 13932
rect 12768 13920 12774 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12768 13892 13001 13920
rect 12768 13880 12774 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 12253 13855 12311 13861
rect 12253 13821 12265 13855
rect 12299 13852 12311 13855
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12299 13824 12909 13852
rect 12299 13821 12311 13824
rect 12253 13815 12311 13821
rect 12897 13821 12909 13824
rect 12943 13852 12955 13855
rect 13446 13852 13452 13864
rect 12943 13824 13452 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 24026 13852 24032 13864
rect 23987 13824 24032 13852
rect 24026 13812 24032 13824
rect 24084 13852 24090 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 24084 13824 24593 13852
rect 24084 13812 24090 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 12434 13744 12440 13796
rect 12492 13784 12498 13796
rect 12805 13787 12863 13793
rect 12805 13784 12817 13787
rect 12492 13756 12817 13784
rect 12492 13744 12498 13756
rect 12805 13753 12817 13756
rect 12851 13753 12863 13787
rect 12805 13747 12863 13753
rect 10597 13719 10655 13725
rect 10597 13685 10609 13719
rect 10643 13716 10655 13719
rect 10686 13716 10692 13728
rect 10643 13688 10692 13716
rect 10643 13685 10655 13688
rect 10597 13679 10655 13685
rect 10686 13676 10692 13688
rect 10744 13676 10750 13728
rect 11054 13716 11060 13728
rect 11015 13688 11060 13716
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 14001 13719 14059 13725
rect 14001 13716 14013 13719
rect 13780 13688 14013 13716
rect 13780 13676 13786 13688
rect 14001 13685 14013 13688
rect 14047 13685 14059 13719
rect 14001 13679 14059 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2869 13515 2927 13521
rect 2869 13481 2881 13515
rect 2915 13512 2927 13515
rect 3234 13512 3240 13524
rect 2915 13484 3240 13512
rect 2915 13481 2927 13484
rect 2869 13475 2927 13481
rect 3234 13472 3240 13484
rect 3292 13472 3298 13524
rect 4341 13515 4399 13521
rect 4341 13481 4353 13515
rect 4387 13512 4399 13515
rect 4706 13512 4712 13524
rect 4387 13484 4712 13512
rect 4387 13481 4399 13484
rect 4341 13475 4399 13481
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 6178 13512 6184 13524
rect 6139 13484 6184 13512
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 7282 13512 7288 13524
rect 7243 13484 7288 13512
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 8386 13512 8392 13524
rect 8347 13484 8392 13512
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 9490 13512 9496 13524
rect 8803 13484 9496 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 9953 13515 10011 13521
rect 9953 13481 9965 13515
rect 9999 13512 10011 13515
rect 10686 13512 10692 13524
rect 9999 13484 10692 13512
rect 9999 13481 10011 13484
rect 9953 13475 10011 13481
rect 10686 13472 10692 13484
rect 10744 13512 10750 13524
rect 11425 13515 11483 13521
rect 11425 13512 11437 13515
rect 10744 13484 11437 13512
rect 10744 13472 10750 13484
rect 11425 13481 11437 13484
rect 11471 13481 11483 13515
rect 11425 13475 11483 13481
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12492 13484 12537 13512
rect 12492 13472 12498 13484
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 12768 13484 12817 13512
rect 12768 13472 12774 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 13354 13512 13360 13524
rect 13315 13484 13360 13512
rect 12805 13475 12863 13481
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 1756 13447 1814 13453
rect 1756 13413 1768 13447
rect 1802 13444 1814 13447
rect 2038 13444 2044 13456
rect 1802 13416 2044 13444
rect 1802 13413 1814 13416
rect 1756 13407 1814 13413
rect 2038 13404 2044 13416
rect 2096 13404 2102 13456
rect 2406 13404 2412 13456
rect 2464 13444 2470 13456
rect 3789 13447 3847 13453
rect 3789 13444 3801 13447
rect 2464 13416 3801 13444
rect 2464 13404 2470 13416
rect 3789 13413 3801 13416
rect 3835 13413 3847 13447
rect 3789 13407 3847 13413
rect 2498 13336 2504 13388
rect 2556 13376 2562 13388
rect 3513 13379 3571 13385
rect 3513 13376 3525 13379
rect 2556 13348 3525 13376
rect 2556 13336 2562 13348
rect 3513 13345 3525 13348
rect 3559 13376 3571 13379
rect 4890 13376 4896 13388
rect 3559 13348 4896 13376
rect 3559 13345 3571 13348
rect 3513 13339 3571 13345
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 5074 13385 5080 13388
rect 5068 13376 5080 13385
rect 5035 13348 5080 13376
rect 5068 13339 5080 13348
rect 5074 13336 5080 13339
rect 5132 13336 5138 13388
rect 5350 13336 5356 13388
rect 5408 13376 5414 13388
rect 6546 13376 6552 13388
rect 5408 13348 6552 13376
rect 5408 13336 5414 13348
rect 6546 13336 6552 13348
rect 6604 13376 6610 13388
rect 7653 13379 7711 13385
rect 7653 13376 7665 13379
rect 6604 13348 7665 13376
rect 6604 13336 6610 13348
rect 7653 13345 7665 13348
rect 7699 13376 7711 13379
rect 8202 13376 8208 13388
rect 7699 13348 8208 13376
rect 7699 13345 7711 13348
rect 7653 13339 7711 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 10318 13385 10324 13388
rect 10312 13376 10324 13385
rect 10279 13348 10324 13376
rect 10312 13339 10324 13348
rect 10318 13336 10324 13339
rect 10376 13336 10382 13388
rect 12894 13336 12900 13388
rect 12952 13376 12958 13388
rect 13722 13376 13728 13388
rect 12952 13348 13728 13376
rect 12952 13336 12958 13348
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 15556 13379 15614 13385
rect 15556 13345 15568 13379
rect 15602 13376 15614 13379
rect 15838 13376 15844 13388
rect 15602 13348 15844 13376
rect 15602 13345 15614 13348
rect 15556 13339 15614 13345
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 23382 13376 23388 13388
rect 23343 13348 23388 13376
rect 23382 13336 23388 13348
rect 23440 13336 23446 13388
rect 1486 13308 1492 13320
rect 1447 13280 1492 13308
rect 1486 13268 1492 13280
rect 1544 13268 1550 13320
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 4801 13311 4859 13317
rect 4801 13308 4813 13311
rect 4764 13280 4813 13308
rect 4764 13268 4770 13280
rect 4801 13277 4813 13280
rect 4847 13277 4859 13311
rect 4801 13271 4859 13277
rect 7745 13311 7803 13317
rect 7745 13277 7757 13311
rect 7791 13277 7803 13311
rect 7926 13308 7932 13320
rect 7887 13280 7932 13308
rect 7745 13271 7803 13277
rect 7650 13200 7656 13252
rect 7708 13240 7714 13252
rect 7760 13240 7788 13271
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 9824 13280 10057 13308
rect 9824 13268 9830 13280
rect 10045 13277 10057 13280
rect 10091 13277 10103 13311
rect 13814 13308 13820 13320
rect 13775 13280 13820 13308
rect 10045 13271 10103 13277
rect 7708 13212 7788 13240
rect 7708 13200 7714 13212
rect 4614 13172 4620 13184
rect 4575 13144 4620 13172
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 6972 13144 7017 13172
rect 6972 13132 6978 13144
rect 8570 13132 8576 13184
rect 8628 13172 8634 13184
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8628 13144 9045 13172
rect 8628 13132 8634 13144
rect 9033 13141 9045 13144
rect 9079 13141 9091 13175
rect 9490 13172 9496 13184
rect 9451 13144 9496 13172
rect 9033 13135 9091 13141
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 10060 13172 10088 13271
rect 13814 13268 13820 13280
rect 13872 13268 13878 13320
rect 13998 13308 14004 13320
rect 13959 13280 14004 13308
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 15286 13308 15292 13320
rect 15247 13280 15292 13308
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 16666 13240 16672 13252
rect 16627 13212 16672 13240
rect 16666 13200 16672 13212
rect 16724 13200 16730 13252
rect 11882 13172 11888 13184
rect 10060 13144 11888 13172
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 13170 13172 13176 13184
rect 13131 13144 13176 13172
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 23569 13175 23627 13181
rect 23569 13141 23581 13175
rect 23615 13172 23627 13175
rect 24946 13172 24952 13184
rect 23615 13144 24952 13172
rect 23615 13141 23627 13144
rect 23569 13135 23627 13141
rect 24946 13132 24952 13144
rect 25004 13132 25010 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1854 12968 1860 12980
rect 1815 12940 1860 12968
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 3234 12968 3240 12980
rect 3195 12940 3240 12968
rect 3234 12928 3240 12940
rect 3292 12928 3298 12980
rect 5534 12928 5540 12980
rect 5592 12968 5598 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 5592 12940 6837 12968
rect 5592 12928 5598 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 7926 12928 7932 12980
rect 7984 12968 7990 12980
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 7984 12940 8217 12968
rect 7984 12928 7990 12940
rect 8205 12937 8217 12940
rect 8251 12937 8263 12971
rect 9398 12968 9404 12980
rect 9359 12940 9404 12968
rect 8205 12931 8263 12937
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 11882 12968 11888 12980
rect 11843 12940 11888 12968
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12894 12968 12900 12980
rect 12855 12940 12900 12968
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 13262 12968 13268 12980
rect 13223 12940 13268 12968
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 15657 12971 15715 12977
rect 15657 12968 15669 12971
rect 15344 12940 15669 12968
rect 15344 12928 15350 12940
rect 15657 12937 15669 12940
rect 15703 12937 15715 12971
rect 23382 12968 23388 12980
rect 23343 12940 23388 12968
rect 15657 12931 15715 12937
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 2498 12832 2504 12844
rect 2459 12804 2504 12832
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 3252 12832 3280 12928
rect 4801 12903 4859 12909
rect 4801 12869 4813 12903
rect 4847 12900 4859 12903
rect 4890 12900 4896 12912
rect 4847 12872 4896 12900
rect 4847 12869 4859 12872
rect 4801 12863 4859 12869
rect 4890 12860 4896 12872
rect 4948 12900 4954 12912
rect 7944 12900 7972 12928
rect 4948 12872 7972 12900
rect 23845 12903 23903 12909
rect 4948 12860 4954 12872
rect 23845 12869 23857 12903
rect 23891 12900 23903 12903
rect 25038 12900 25044 12912
rect 23891 12872 25044 12900
rect 23891 12869 23903 12872
rect 23845 12863 23903 12869
rect 25038 12860 25044 12872
rect 25096 12860 25102 12912
rect 6546 12832 6552 12844
rect 3252 12804 3556 12832
rect 6507 12804 6552 12832
rect 1486 12724 1492 12776
rect 1544 12764 1550 12776
rect 3421 12767 3479 12773
rect 3421 12764 3433 12767
rect 1544 12736 3433 12764
rect 1544 12724 1550 12736
rect 3421 12733 3433 12736
rect 3467 12733 3479 12767
rect 3528 12764 3556 12804
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 7248 12804 7389 12832
rect 7248 12792 7254 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 9309 12835 9367 12841
rect 9309 12801 9321 12835
rect 9355 12832 9367 12835
rect 10045 12835 10103 12841
rect 10045 12832 10057 12835
rect 9355 12804 10057 12832
rect 9355 12801 9367 12804
rect 9309 12795 9367 12801
rect 10045 12801 10057 12804
rect 10091 12832 10103 12835
rect 10318 12832 10324 12844
rect 10091 12804 10324 12832
rect 10091 12801 10103 12804
rect 10045 12795 10103 12801
rect 10318 12792 10324 12804
rect 10376 12832 10382 12844
rect 10376 12804 10548 12832
rect 10376 12792 10382 12804
rect 3677 12767 3735 12773
rect 3677 12764 3689 12767
rect 3528 12736 3689 12764
rect 3421 12727 3479 12733
rect 3677 12733 3689 12736
rect 3723 12733 3735 12767
rect 3677 12727 3735 12733
rect 2225 12699 2283 12705
rect 2225 12665 2237 12699
rect 2271 12696 2283 12699
rect 2958 12696 2964 12708
rect 2271 12668 2964 12696
rect 2271 12665 2283 12668
rect 2225 12659 2283 12665
rect 2958 12656 2964 12668
rect 3016 12656 3022 12708
rect 3436 12696 3464 12727
rect 9490 12724 9496 12776
rect 9548 12764 9554 12776
rect 9674 12764 9680 12776
rect 9548 12736 9680 12764
rect 9548 12724 9554 12736
rect 9674 12724 9680 12736
rect 9732 12764 9738 12776
rect 9769 12767 9827 12773
rect 9769 12764 9781 12767
rect 9732 12736 9781 12764
rect 9732 12724 9738 12736
rect 9769 12733 9781 12736
rect 9815 12733 9827 12767
rect 9769 12727 9827 12733
rect 4614 12696 4620 12708
rect 3436 12668 4620 12696
rect 4614 12656 4620 12668
rect 4672 12696 4678 12708
rect 5721 12699 5779 12705
rect 5721 12696 5733 12699
rect 4672 12668 5733 12696
rect 4672 12656 4678 12668
rect 5721 12665 5733 12668
rect 5767 12696 5779 12699
rect 6178 12696 6184 12708
rect 5767 12668 6184 12696
rect 5767 12665 5779 12668
rect 5721 12659 5779 12665
rect 6178 12656 6184 12668
rect 6236 12656 6242 12708
rect 6273 12699 6331 12705
rect 6273 12665 6285 12699
rect 6319 12696 6331 12699
rect 7098 12696 7104 12708
rect 6319 12668 7104 12696
rect 6319 12665 6331 12668
rect 6273 12659 6331 12665
rect 7098 12656 7104 12668
rect 7156 12696 7162 12708
rect 10520 12705 10548 12804
rect 12710 12724 12716 12776
rect 12768 12764 12774 12776
rect 13170 12764 13176 12776
rect 12768 12736 13176 12764
rect 12768 12724 12774 12736
rect 13170 12724 13176 12736
rect 13228 12764 13234 12776
rect 13357 12767 13415 12773
rect 13357 12764 13369 12767
rect 13228 12736 13369 12764
rect 13228 12724 13234 12736
rect 13357 12733 13369 12736
rect 13403 12733 13415 12767
rect 23658 12764 23664 12776
rect 23619 12736 23664 12764
rect 13357 12727 13415 12733
rect 23658 12724 23664 12736
rect 23716 12764 23722 12776
rect 24213 12767 24271 12773
rect 24213 12764 24225 12767
rect 23716 12736 24225 12764
rect 23716 12724 23722 12736
rect 24213 12733 24225 12736
rect 24259 12733 24271 12767
rect 24213 12727 24271 12733
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 7156 12668 7205 12696
rect 7156 12656 7162 12668
rect 7193 12665 7205 12668
rect 7239 12665 7251 12699
rect 7193 12659 7251 12665
rect 10505 12699 10563 12705
rect 10505 12665 10517 12699
rect 10551 12696 10563 12699
rect 10962 12696 10968 12708
rect 10551 12668 10968 12696
rect 10551 12665 10563 12668
rect 10505 12659 10563 12665
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 13630 12705 13636 12708
rect 13624 12659 13636 12705
rect 13688 12696 13694 12708
rect 15381 12699 15439 12705
rect 15381 12696 15393 12699
rect 13688 12668 13724 12696
rect 14752 12668 15393 12696
rect 13630 12656 13636 12659
rect 13688 12656 13694 12668
rect 1765 12631 1823 12637
rect 1765 12597 1777 12631
rect 1811 12628 1823 12631
rect 2317 12631 2375 12637
rect 2317 12628 2329 12631
rect 1811 12600 2329 12628
rect 1811 12597 1823 12600
rect 1765 12591 1823 12597
rect 2317 12597 2329 12600
rect 2363 12628 2375 12631
rect 4154 12628 4160 12640
rect 2363 12600 4160 12628
rect 2363 12597 2375 12600
rect 2317 12591 2375 12597
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 5074 12588 5080 12640
rect 5132 12628 5138 12640
rect 5445 12631 5503 12637
rect 5445 12628 5457 12631
rect 5132 12600 5457 12628
rect 5132 12588 5138 12600
rect 5445 12597 5457 12600
rect 5491 12628 5503 12631
rect 5534 12628 5540 12640
rect 5491 12600 5540 12628
rect 5491 12597 5503 12600
rect 5445 12591 5503 12597
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7285 12631 7343 12637
rect 7285 12628 7297 12631
rect 6972 12600 7297 12628
rect 6972 12588 6978 12600
rect 7285 12597 7297 12600
rect 7331 12597 7343 12631
rect 7285 12591 7343 12597
rect 7650 12588 7656 12640
rect 7708 12628 7714 12640
rect 7837 12631 7895 12637
rect 7837 12628 7849 12631
rect 7708 12600 7849 12628
rect 7708 12588 7714 12600
rect 7837 12597 7849 12600
rect 7883 12597 7895 12631
rect 8386 12628 8392 12640
rect 8347 12600 8392 12628
rect 7837 12591 7895 12597
rect 8386 12588 8392 12600
rect 8444 12588 8450 12640
rect 8570 12588 8576 12640
rect 8628 12628 8634 12640
rect 8849 12631 8907 12637
rect 8849 12628 8861 12631
rect 8628 12600 8861 12628
rect 8628 12588 8634 12600
rect 8849 12597 8861 12600
rect 8895 12597 8907 12631
rect 9858 12628 9864 12640
rect 9819 12600 9864 12628
rect 8849 12591 8907 12597
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 10778 12628 10784 12640
rect 10739 12600 10784 12628
rect 10778 12588 10784 12600
rect 10836 12628 10842 12640
rect 11149 12631 11207 12637
rect 11149 12628 11161 12631
rect 10836 12600 11161 12628
rect 10836 12588 10842 12600
rect 11149 12597 11161 12600
rect 11195 12597 11207 12631
rect 11330 12628 11336 12640
rect 11291 12600 11336 12628
rect 11149 12591 11207 12597
rect 11330 12588 11336 12600
rect 11388 12588 11394 12640
rect 14752 12637 14780 12668
rect 15381 12665 15393 12668
rect 15427 12696 15439 12699
rect 15838 12696 15844 12708
rect 15427 12668 15844 12696
rect 15427 12665 15439 12668
rect 15381 12659 15439 12665
rect 15838 12656 15844 12668
rect 15896 12656 15902 12708
rect 14737 12631 14795 12637
rect 14737 12597 14749 12631
rect 14783 12597 14795 12631
rect 14737 12591 14795 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2038 12384 2044 12436
rect 2096 12424 2102 12436
rect 2869 12427 2927 12433
rect 2869 12424 2881 12427
rect 2096 12396 2881 12424
rect 2096 12384 2102 12396
rect 2869 12393 2881 12396
rect 2915 12424 2927 12427
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 2915 12396 3433 12424
rect 2915 12393 2927 12396
rect 2869 12387 2927 12393
rect 3421 12393 3433 12396
rect 3467 12393 3479 12427
rect 3421 12387 3479 12393
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 5997 12427 6055 12433
rect 5997 12424 6009 12427
rect 5592 12396 6009 12424
rect 5592 12384 5598 12396
rect 5997 12393 6009 12396
rect 6043 12393 6055 12427
rect 7098 12424 7104 12436
rect 7059 12396 7104 12424
rect 5997 12387 6055 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11701 12427 11759 12433
rect 11701 12424 11713 12427
rect 11112 12396 11713 12424
rect 11112 12384 11118 12396
rect 11701 12393 11713 12396
rect 11747 12393 11759 12427
rect 11701 12387 11759 12393
rect 12805 12427 12863 12433
rect 12805 12393 12817 12427
rect 12851 12424 12863 12427
rect 12986 12424 12992 12436
rect 12851 12396 12992 12424
rect 12851 12393 12863 12396
rect 12805 12387 12863 12393
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 4890 12365 4896 12368
rect 4884 12356 4896 12365
rect 4851 12328 4896 12356
rect 4884 12319 4896 12328
rect 4890 12316 4896 12319
rect 4948 12316 4954 12368
rect 10778 12356 10784 12368
rect 10336 12328 10784 12356
rect 1756 12291 1814 12297
rect 1756 12257 1768 12291
rect 1802 12288 1814 12291
rect 2590 12288 2596 12300
rect 1802 12260 2596 12288
rect 1802 12257 1814 12260
rect 1756 12251 1814 12257
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 4614 12288 4620 12300
rect 4575 12260 4620 12288
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 6362 12248 6368 12300
rect 6420 12288 6426 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 6420 12260 7481 12288
rect 6420 12248 6426 12260
rect 7469 12257 7481 12260
rect 7515 12288 7527 12291
rect 8202 12288 8208 12300
rect 7515 12260 8208 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 8849 12291 8907 12297
rect 8849 12257 8861 12291
rect 8895 12288 8907 12291
rect 9030 12288 9036 12300
rect 8895 12260 9036 12288
rect 8895 12257 8907 12260
rect 8849 12251 8907 12257
rect 9030 12248 9036 12260
rect 9088 12248 9094 12300
rect 10336 12232 10364 12328
rect 10778 12316 10784 12328
rect 10836 12356 10842 12368
rect 12253 12359 12311 12365
rect 12253 12356 12265 12359
rect 10836 12328 12265 12356
rect 10836 12316 10842 12328
rect 12253 12325 12265 12328
rect 12299 12356 12311 12359
rect 12710 12356 12716 12368
rect 12299 12328 12716 12356
rect 12299 12325 12311 12328
rect 12253 12319 12311 12325
rect 12710 12316 12716 12328
rect 12768 12316 12774 12368
rect 10588 12291 10646 12297
rect 10588 12257 10600 12291
rect 10634 12288 10646 12291
rect 11146 12288 11152 12300
rect 10634 12260 11152 12288
rect 10634 12257 10646 12260
rect 10588 12251 10646 12257
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 13173 12291 13231 12297
rect 13173 12288 13185 12291
rect 12216 12260 13185 12288
rect 12216 12248 12222 12260
rect 13173 12257 13185 12260
rect 13219 12257 13231 12291
rect 13630 12288 13636 12300
rect 13173 12251 13231 12257
rect 13372 12260 13636 12288
rect 13372 12232 13400 12260
rect 13630 12248 13636 12260
rect 13688 12288 13694 12300
rect 13909 12291 13967 12297
rect 13909 12288 13921 12291
rect 13688 12260 13921 12288
rect 13688 12248 13694 12260
rect 13909 12257 13921 12260
rect 13955 12257 13967 12291
rect 13909 12251 13967 12257
rect 14366 12248 14372 12300
rect 14424 12288 14430 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 14424 12260 15669 12288
rect 14424 12248 14430 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 22278 12288 22284 12300
rect 22239 12260 22284 12288
rect 15657 12251 15715 12257
rect 22278 12248 22284 12260
rect 22336 12248 22342 12300
rect 1486 12220 1492 12232
rect 1399 12192 1492 12220
rect 1486 12180 1492 12192
rect 1544 12180 1550 12232
rect 7006 12180 7012 12232
rect 7064 12220 7070 12232
rect 7561 12223 7619 12229
rect 7561 12220 7573 12223
rect 7064 12192 7573 12220
rect 7064 12180 7070 12192
rect 7561 12189 7573 12192
rect 7607 12189 7619 12223
rect 7561 12183 7619 12189
rect 7653 12223 7711 12229
rect 7653 12189 7665 12223
rect 7699 12189 7711 12223
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 7653 12183 7711 12189
rect 1504 12084 1532 12180
rect 6917 12155 6975 12161
rect 6917 12121 6929 12155
rect 6963 12152 6975 12155
rect 7190 12152 7196 12164
rect 6963 12124 7196 12152
rect 6963 12121 6975 12124
rect 6917 12115 6975 12121
rect 7190 12112 7196 12124
rect 7248 12112 7254 12164
rect 7466 12112 7472 12164
rect 7524 12152 7530 12164
rect 7668 12152 7696 12183
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 12713 12223 12771 12229
rect 12713 12189 12725 12223
rect 12759 12220 12771 12223
rect 12802 12220 12808 12232
rect 12759 12192 12808 12220
rect 12759 12189 12771 12192
rect 12713 12183 12771 12189
rect 12802 12180 12808 12192
rect 12860 12220 12866 12232
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 12860 12192 13277 12220
rect 12860 12180 12866 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 13412 12192 13457 12220
rect 13412 12180 13418 12192
rect 13814 12180 13820 12232
rect 13872 12180 13878 12232
rect 15470 12180 15476 12232
rect 15528 12220 15534 12232
rect 15749 12223 15807 12229
rect 15749 12220 15761 12223
rect 15528 12192 15761 12220
rect 15528 12180 15534 12192
rect 15749 12189 15761 12192
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 15896 12192 15941 12220
rect 15896 12180 15902 12192
rect 7524 12124 7696 12152
rect 8205 12155 8263 12161
rect 7524 12112 7530 12124
rect 8205 12121 8217 12155
rect 8251 12152 8263 12155
rect 8570 12152 8576 12164
rect 8251 12124 8576 12152
rect 8251 12121 8263 12124
rect 8205 12115 8263 12121
rect 1762 12084 1768 12096
rect 1504 12056 1768 12084
rect 1762 12044 1768 12056
rect 1820 12044 1826 12096
rect 3878 12084 3884 12096
rect 3839 12056 3884 12084
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 4338 12084 4344 12096
rect 4299 12056 4344 12084
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 8220 12084 8248 12115
rect 8570 12112 8576 12124
rect 8628 12112 8634 12164
rect 9582 12152 9588 12164
rect 8680 12124 9588 12152
rect 8680 12096 8708 12124
rect 9582 12112 9588 12124
rect 9640 12152 9646 12164
rect 9861 12155 9919 12161
rect 9861 12152 9873 12155
rect 9640 12124 9873 12152
rect 9640 12112 9646 12124
rect 9861 12121 9873 12124
rect 9907 12121 9919 12155
rect 13832 12152 13860 12180
rect 14277 12155 14335 12161
rect 14277 12152 14289 12155
rect 13832 12124 14289 12152
rect 9861 12115 9919 12121
rect 14277 12121 14289 12124
rect 14323 12152 14335 12155
rect 15289 12155 15347 12161
rect 15289 12152 15301 12155
rect 14323 12124 15301 12152
rect 14323 12121 14335 12124
rect 14277 12115 14335 12121
rect 15289 12121 15301 12124
rect 15335 12121 15347 12155
rect 15289 12115 15347 12121
rect 8662 12084 8668 12096
rect 6788 12056 8248 12084
rect 8623 12056 8668 12084
rect 6788 12044 6794 12056
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 9490 12084 9496 12096
rect 9451 12056 9496 12084
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 22462 12084 22468 12096
rect 22423 12056 22468 12084
rect 22462 12044 22468 12056
rect 22520 12044 22526 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2590 11880 2596 11892
rect 2551 11852 2596 11880
rect 2590 11840 2596 11852
rect 2648 11880 2654 11892
rect 2958 11880 2964 11892
rect 2648 11852 2964 11880
rect 2648 11840 2654 11852
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 4890 11880 4896 11892
rect 4851 11852 4896 11880
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 5534 11880 5540 11892
rect 5495 11852 5540 11880
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 6362 11880 6368 11892
rect 6323 11852 6368 11880
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 10318 11880 10324 11892
rect 9692 11852 10324 11880
rect 3418 11772 3424 11824
rect 3476 11812 3482 11824
rect 4062 11812 4068 11824
rect 3476 11784 4068 11812
rect 3476 11772 3482 11784
rect 4062 11772 4068 11784
rect 4120 11772 4126 11824
rect 6178 11772 6184 11824
rect 6236 11812 6242 11824
rect 6457 11815 6515 11821
rect 6457 11812 6469 11815
rect 6236 11784 6469 11812
rect 6236 11772 6242 11784
rect 6457 11781 6469 11784
rect 6503 11812 6515 11815
rect 6730 11812 6736 11824
rect 6503 11784 6736 11812
rect 6503 11781 6515 11784
rect 6457 11775 6515 11781
rect 6730 11772 6736 11784
rect 6788 11772 6794 11824
rect 2130 11744 2136 11756
rect 2091 11716 2136 11744
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 3878 11704 3884 11756
rect 3936 11744 3942 11756
rect 4341 11747 4399 11753
rect 4341 11744 4353 11747
rect 3936 11716 4353 11744
rect 3936 11704 3942 11716
rect 4341 11713 4353 11716
rect 4387 11744 4399 11747
rect 4614 11744 4620 11756
rect 4387 11716 4620 11744
rect 4387 11713 4399 11716
rect 4341 11707 4399 11713
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 9692 11753 9720 11852
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 12158 11880 12164 11892
rect 11388 11852 12164 11880
rect 11388 11840 11394 11852
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 14093 11883 14151 11889
rect 14093 11880 14105 11883
rect 13412 11852 14105 11880
rect 13412 11840 13418 11852
rect 14093 11849 14105 11852
rect 14139 11849 14151 11883
rect 14093 11843 14151 11849
rect 15197 11883 15255 11889
rect 15197 11849 15209 11883
rect 15243 11880 15255 11883
rect 15378 11880 15384 11892
rect 15243 11852 15384 11880
rect 15243 11849 15255 11852
rect 15197 11843 15255 11849
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 22278 11880 22284 11892
rect 22239 11852 22284 11880
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11744 5319 11747
rect 9677 11747 9735 11753
rect 9677 11744 9689 11747
rect 5307 11716 6684 11744
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 6656 11688 6684 11716
rect 9232 11716 9689 11744
rect 1946 11676 1952 11688
rect 1907 11648 1952 11676
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 3970 11636 3976 11688
rect 4028 11676 4034 11688
rect 4157 11679 4215 11685
rect 4157 11676 4169 11679
rect 4028 11648 4169 11676
rect 4028 11636 4034 11648
rect 4157 11645 4169 11648
rect 4203 11676 4215 11679
rect 5166 11676 5172 11688
rect 4203 11648 5172 11676
rect 4203 11645 4215 11648
rect 4157 11639 4215 11645
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 5353 11679 5411 11685
rect 5353 11645 5365 11679
rect 5399 11676 5411 11679
rect 5442 11676 5448 11688
rect 5399 11648 5448 11676
rect 5399 11645 5411 11648
rect 5353 11639 5411 11645
rect 5442 11636 5448 11648
rect 5500 11676 5506 11688
rect 5905 11679 5963 11685
rect 5905 11676 5917 11679
rect 5500 11648 5917 11676
rect 5500 11636 5506 11648
rect 5905 11645 5917 11648
rect 5951 11645 5963 11679
rect 6638 11676 6644 11688
rect 6599 11648 6644 11676
rect 5905 11639 5963 11645
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 6822 11676 6828 11688
rect 6783 11648 6828 11676
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 7098 11617 7104 11620
rect 3697 11611 3755 11617
rect 3697 11577 3709 11611
rect 3743 11608 3755 11611
rect 7092 11608 7104 11617
rect 3743 11580 4292 11608
rect 7059 11580 7104 11608
rect 3743 11577 3755 11580
rect 3697 11571 3755 11577
rect 1486 11500 1492 11552
rect 1544 11540 1550 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 1544 11512 1593 11540
rect 1544 11500 1550 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 1581 11503 1639 11509
rect 2041 11543 2099 11549
rect 2041 11509 2053 11543
rect 2087 11540 2099 11543
rect 2498 11540 2504 11552
rect 2087 11512 2504 11540
rect 2087 11509 2099 11512
rect 2041 11503 2099 11509
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 3786 11540 3792 11552
rect 3747 11512 3792 11540
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 4264 11549 4292 11580
rect 7092 11571 7104 11580
rect 7098 11568 7104 11571
rect 7156 11568 7162 11620
rect 7466 11568 7472 11620
rect 7524 11608 7530 11620
rect 8757 11611 8815 11617
rect 8757 11608 8769 11611
rect 7524 11580 8769 11608
rect 7524 11568 7530 11580
rect 8757 11577 8769 11580
rect 8803 11577 8815 11611
rect 8757 11571 8815 11577
rect 4249 11543 4307 11549
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 4982 11540 4988 11552
rect 4295 11512 4988 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 8076 11512 8217 11540
rect 8076 11500 8082 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 8205 11503 8263 11509
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 9232 11540 9260 11716
rect 9677 11713 9689 11716
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11744 11943 11747
rect 15746 11744 15752 11756
rect 11931 11716 12848 11744
rect 15707 11716 15752 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 9582 11676 9588 11688
rect 9543 11648 9588 11676
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 12710 11676 12716 11688
rect 12623 11648 12716 11676
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 12820 11676 12848 11716
rect 15746 11704 15752 11716
rect 15804 11744 15810 11756
rect 16209 11747 16267 11753
rect 16209 11744 16221 11747
rect 15804 11716 16221 11744
rect 15804 11704 15810 11716
rect 16209 11713 16221 11716
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 12980 11679 13038 11685
rect 12980 11676 12992 11679
rect 12820 11648 12992 11676
rect 12980 11645 12992 11648
rect 13026 11676 13038 11679
rect 13722 11676 13728 11688
rect 13026 11648 13728 11676
rect 13026 11645 13038 11648
rect 12980 11639 13038 11645
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 15562 11676 15568 11688
rect 15523 11648 15568 11676
rect 15562 11636 15568 11648
rect 15620 11636 15626 11688
rect 9950 11617 9956 11620
rect 9309 11611 9367 11617
rect 9309 11577 9321 11611
rect 9355 11608 9367 11611
rect 9944 11608 9956 11617
rect 9355 11580 9956 11608
rect 9355 11577 9367 11580
rect 9309 11571 9367 11577
rect 9944 11571 9956 11580
rect 9950 11568 9956 11571
rect 10008 11568 10014 11620
rect 12728 11608 12756 11636
rect 14458 11608 14464 11620
rect 12728 11580 14464 11608
rect 14458 11568 14464 11580
rect 14516 11568 14522 11620
rect 14550 11568 14556 11620
rect 14608 11608 14614 11620
rect 15013 11611 15071 11617
rect 15013 11608 15025 11611
rect 14608 11580 15025 11608
rect 14608 11568 14614 11580
rect 15013 11577 15025 11580
rect 15059 11608 15071 11611
rect 15470 11608 15476 11620
rect 15059 11580 15476 11608
rect 15059 11577 15071 11580
rect 15013 11571 15071 11577
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 9401 11543 9459 11549
rect 9401 11540 9413 11543
rect 8536 11512 9413 11540
rect 8536 11500 8542 11512
rect 9401 11509 9413 11512
rect 9447 11509 9459 11543
rect 9401 11503 9459 11509
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 11146 11540 11152 11552
rect 11103 11512 11152 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14645 11543 14703 11549
rect 14645 11540 14657 11543
rect 14424 11512 14657 11540
rect 14424 11500 14430 11512
rect 14645 11509 14657 11512
rect 14691 11509 14703 11543
rect 15654 11540 15660 11552
rect 15615 11512 15660 11540
rect 14645 11503 14703 11509
rect 15654 11500 15660 11512
rect 15712 11540 15718 11552
rect 16577 11543 16635 11549
rect 16577 11540 16589 11543
rect 15712 11512 16589 11540
rect 15712 11500 15718 11512
rect 16577 11509 16589 11512
rect 16623 11509 16635 11543
rect 16577 11503 16635 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1394 11336 1400 11348
rect 1355 11308 1400 11336
rect 1394 11296 1400 11308
rect 1452 11296 1458 11348
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2130 11336 2136 11348
rect 1995 11308 2136 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 2409 11339 2467 11345
rect 2409 11336 2421 11339
rect 2280 11308 2421 11336
rect 2280 11296 2286 11308
rect 2409 11305 2421 11308
rect 2455 11305 2467 11339
rect 2409 11299 2467 11305
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 2556 11308 3433 11336
rect 2556 11296 2562 11308
rect 3421 11305 3433 11308
rect 3467 11336 3479 11339
rect 4062 11336 4068 11348
rect 3467 11308 4068 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4430 11296 4436 11348
rect 4488 11336 4494 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4488 11308 4537 11336
rect 4488 11296 4494 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 5810 11336 5816 11348
rect 5771 11308 5816 11336
rect 4525 11299 4583 11305
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 9674 11336 9680 11348
rect 9635 11308 9680 11336
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 11054 11336 11060 11348
rect 11015 11308 11060 11336
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 11238 11336 11244 11348
rect 11199 11308 11244 11336
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 12802 11336 12808 11348
rect 12763 11308 12808 11336
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 13998 11336 14004 11348
rect 13959 11308 14004 11336
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 14458 11336 14464 11348
rect 14419 11308 14464 11336
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 15562 11336 15568 11348
rect 15523 11308 15568 11336
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 15838 11336 15844 11348
rect 15799 11308 15844 11336
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 3881 11271 3939 11277
rect 3881 11237 3893 11271
rect 3927 11268 3939 11271
rect 3970 11268 3976 11280
rect 3927 11240 3976 11268
rect 3927 11237 3939 11240
rect 3881 11231 3939 11237
rect 3970 11228 3976 11240
rect 4028 11228 4034 11280
rect 6917 11271 6975 11277
rect 6917 11237 6929 11271
rect 6963 11268 6975 11271
rect 7098 11268 7104 11280
rect 6963 11240 7104 11268
rect 6963 11237 6975 11240
rect 6917 11231 6975 11237
rect 7098 11228 7104 11240
rect 7156 11228 7162 11280
rect 7368 11271 7426 11277
rect 7368 11237 7380 11271
rect 7414 11268 7426 11271
rect 8018 11268 8024 11280
rect 7414 11240 8024 11268
rect 7414 11237 7426 11240
rect 7368 11231 7426 11237
rect 8018 11228 8024 11240
rect 8076 11228 8082 11280
rect 12713 11271 12771 11277
rect 12713 11237 12725 11271
rect 12759 11268 12771 11271
rect 13354 11268 13360 11280
rect 12759 11240 13360 11268
rect 12759 11237 12771 11240
rect 12713 11231 12771 11237
rect 13354 11228 13360 11240
rect 13412 11228 13418 11280
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 3418 11200 3424 11212
rect 2823 11172 3424 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 3418 11160 3424 11172
rect 3476 11160 3482 11212
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4212 11172 4445 11200
rect 4212 11160 4218 11172
rect 4433 11169 4445 11172
rect 4479 11200 4491 11203
rect 5350 11200 5356 11212
rect 4479 11172 5356 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 5350 11160 5356 11172
rect 5408 11160 5414 11212
rect 5629 11203 5687 11209
rect 5629 11169 5641 11203
rect 5675 11200 5687 11203
rect 5994 11200 6000 11212
rect 5675 11172 6000 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 8478 11200 8484 11212
rect 6880 11172 8484 11200
rect 6880 11160 6886 11172
rect 2866 11132 2872 11144
rect 2827 11104 2872 11132
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 2958 11092 2964 11144
rect 3016 11132 3022 11144
rect 4614 11132 4620 11144
rect 3016 11104 3061 11132
rect 4575 11104 4620 11132
rect 3016 11092 3022 11104
rect 4614 11092 4620 11104
rect 4672 11132 4678 11144
rect 5442 11132 5448 11144
rect 4672 11104 5448 11132
rect 4672 11092 4678 11104
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 7116 11141 7144 11172
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 10045 11203 10103 11209
rect 10045 11169 10057 11203
rect 10091 11200 10103 11203
rect 10778 11200 10784 11212
rect 10091 11172 10784 11200
rect 10091 11169 10103 11172
rect 10045 11163 10103 11169
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 11606 11200 11612 11212
rect 11567 11172 11612 11200
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 13173 11203 13231 11209
rect 13173 11200 13185 11203
rect 12492 11172 13185 11200
rect 12492 11160 12498 11172
rect 13173 11169 13185 11172
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11101 7159 11135
rect 10134 11132 10140 11144
rect 10095 11104 10140 11132
rect 7101 11095 7159 11101
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11101 10379 11135
rect 11698 11132 11704 11144
rect 11659 11104 11704 11132
rect 10321 11095 10379 11101
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11033 4123 11067
rect 4065 11027 4123 11033
rect 6549 11067 6607 11073
rect 6549 11033 6561 11067
rect 6595 11064 6607 11067
rect 7006 11064 7012 11076
rect 6595 11036 7012 11064
rect 6595 11033 6607 11036
rect 6549 11027 6607 11033
rect 2038 10956 2044 11008
rect 2096 10996 2102 11008
rect 2225 10999 2283 11005
rect 2225 10996 2237 10999
rect 2096 10968 2237 10996
rect 2096 10956 2102 10968
rect 2225 10965 2237 10968
rect 2271 10965 2283 10999
rect 4080 10996 4108 11027
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 9030 11064 9036 11076
rect 8991 11036 9036 11064
rect 9030 11024 9036 11036
rect 9088 11024 9094 11076
rect 9493 11067 9551 11073
rect 9493 11033 9505 11067
rect 9539 11064 9551 11067
rect 10336 11064 10364 11095
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11132 13323 11135
rect 13354 11132 13360 11144
rect 13311 11104 13360 11132
rect 13311 11101 13323 11104
rect 13265 11095 13323 11101
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 9539 11036 10793 11064
rect 9539 11033 9551 11036
rect 9493 11027 9551 11033
rect 10781 11033 10793 11036
rect 10827 11064 10839 11067
rect 11146 11064 11152 11076
rect 10827 11036 11152 11064
rect 10827 11033 10839 11036
rect 10781 11027 10839 11033
rect 11146 11024 11152 11036
rect 11204 11064 11210 11076
rect 11808 11064 11836 11095
rect 13354 11092 13360 11104
rect 13412 11092 13418 11144
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11132 13507 11135
rect 13722 11132 13728 11144
rect 13495 11104 13728 11132
rect 13495 11101 13507 11104
rect 13449 11095 13507 11101
rect 11204 11036 11836 11064
rect 12345 11067 12403 11073
rect 11204 11024 11210 11036
rect 12345 11033 12357 11067
rect 12391 11064 12403 11067
rect 13464 11064 13492 11095
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13906 11064 13912 11076
rect 12391 11036 13492 11064
rect 13867 11036 13912 11064
rect 12391 11033 12403 11036
rect 12345 11027 12403 11033
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 4706 10996 4712 11008
rect 4080 10968 4712 10996
rect 2225 10959 2283 10965
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 5074 10996 5080 11008
rect 5035 10968 5080 10996
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 5442 10996 5448 11008
rect 5403 10968 5448 10996
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 8481 10999 8539 11005
rect 8481 10965 8493 10999
rect 8527 10996 8539 10999
rect 8754 10996 8760 11008
rect 8527 10968 8760 10996
rect 8527 10965 8539 10968
rect 8481 10959 8539 10965
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1673 10795 1731 10801
rect 1673 10761 1685 10795
rect 1719 10792 1731 10795
rect 2682 10792 2688 10804
rect 1719 10764 2688 10792
rect 1719 10761 1731 10764
rect 1673 10755 1731 10761
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 3145 10795 3203 10801
rect 3145 10792 3157 10795
rect 3016 10764 3157 10792
rect 3016 10752 3022 10764
rect 3145 10761 3157 10764
rect 3191 10761 3203 10795
rect 3145 10755 3203 10761
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 3476 10764 3709 10792
rect 3476 10752 3482 10764
rect 3697 10761 3709 10764
rect 3743 10761 3755 10795
rect 3697 10755 3755 10761
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5592 10764 5641 10792
rect 5592 10752 5598 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5629 10755 5687 10761
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 9861 10795 9919 10801
rect 6972 10764 7017 10792
rect 6972 10752 6978 10764
rect 9861 10761 9873 10795
rect 9907 10792 9919 10795
rect 9950 10792 9956 10804
rect 9907 10764 9956 10792
rect 9907 10761 9919 10764
rect 9861 10755 9919 10761
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 10192 10764 10425 10792
rect 10192 10752 10198 10764
rect 10413 10761 10425 10764
rect 10459 10761 10471 10795
rect 10778 10792 10784 10804
rect 10739 10764 10784 10792
rect 10413 10755 10471 10761
rect 10778 10752 10784 10764
rect 10836 10792 10842 10804
rect 10836 10764 11008 10792
rect 10836 10752 10842 10764
rect 4249 10727 4307 10733
rect 4249 10693 4261 10727
rect 4295 10724 4307 10727
rect 5258 10724 5264 10736
rect 4295 10696 5264 10724
rect 4295 10693 4307 10696
rect 4249 10687 4307 10693
rect 5258 10684 5264 10696
rect 5316 10684 5322 10736
rect 4893 10659 4951 10665
rect 4893 10625 4905 10659
rect 4939 10656 4951 10659
rect 5074 10656 5080 10668
rect 4939 10628 5080 10656
rect 4939 10625 4951 10628
rect 4893 10619 4951 10625
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 7466 10656 7472 10668
rect 6687 10628 7472 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 10980 10665 11008 10764
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 11664 10764 11805 10792
rect 11664 10752 11670 10764
rect 11793 10761 11805 10764
rect 11839 10761 11851 10795
rect 11793 10755 11851 10761
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 1762 10588 1768 10600
rect 1675 10560 1768 10588
rect 1762 10548 1768 10560
rect 1820 10588 1826 10600
rect 2314 10588 2320 10600
rect 1820 10560 2320 10588
rect 1820 10548 1826 10560
rect 2314 10548 2320 10560
rect 2372 10548 2378 10600
rect 4706 10588 4712 10600
rect 4619 10560 4712 10588
rect 4706 10548 4712 10560
rect 4764 10588 4770 10600
rect 5442 10588 5448 10600
rect 4764 10560 5448 10588
rect 4764 10548 4770 10560
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 8478 10588 8484 10600
rect 8439 10560 8484 10588
rect 8478 10548 8484 10560
rect 8536 10548 8542 10600
rect 13173 10591 13231 10597
rect 13173 10557 13185 10591
rect 13219 10588 13231 10591
rect 13722 10588 13728 10600
rect 13219 10560 13728 10588
rect 13219 10557 13231 10560
rect 13173 10551 13231 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 2038 10529 2044 10532
rect 2032 10520 2044 10529
rect 1999 10492 2044 10520
rect 2032 10483 2044 10492
rect 2038 10480 2044 10483
rect 2096 10480 2102 10532
rect 7098 10480 7104 10532
rect 7156 10520 7162 10532
rect 7377 10523 7435 10529
rect 7377 10520 7389 10523
rect 7156 10492 7389 10520
rect 7156 10480 7162 10492
rect 7377 10489 7389 10492
rect 7423 10489 7435 10523
rect 8018 10520 8024 10532
rect 7979 10492 8024 10520
rect 7377 10483 7435 10489
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 8754 10529 8760 10532
rect 8389 10523 8447 10529
rect 8389 10489 8401 10523
rect 8435 10520 8447 10523
rect 8748 10520 8760 10529
rect 8435 10492 8760 10520
rect 8435 10489 8447 10492
rect 8389 10483 8447 10489
rect 8748 10483 8760 10492
rect 8754 10480 8760 10483
rect 8812 10480 8818 10532
rect 11606 10480 11612 10532
rect 11664 10520 11670 10532
rect 12161 10523 12219 10529
rect 12161 10520 12173 10523
rect 11664 10492 12173 10520
rect 11664 10480 11670 10492
rect 12161 10489 12173 10492
rect 12207 10520 12219 10523
rect 12434 10520 12440 10532
rect 12207 10492 12440 10520
rect 12207 10489 12219 10492
rect 12161 10483 12219 10489
rect 12434 10480 12440 10492
rect 12492 10480 12498 10532
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10452 4215 10455
rect 4430 10452 4436 10464
rect 4203 10424 4436 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 4617 10455 4675 10461
rect 4617 10421 4629 10455
rect 4663 10452 4675 10455
rect 5166 10452 5172 10464
rect 4663 10424 5172 10452
rect 4663 10421 4675 10424
rect 4617 10415 4675 10421
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 5350 10452 5356 10464
rect 5311 10424 5356 10452
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 6273 10455 6331 10461
rect 6273 10421 6285 10455
rect 6319 10452 6331 10455
rect 7282 10452 7288 10464
rect 6319 10424 7288 10452
rect 6319 10421 6331 10424
rect 6273 10415 6331 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11425 10455 11483 10461
rect 11425 10452 11437 10455
rect 11112 10424 11437 10452
rect 11112 10412 11118 10424
rect 11425 10421 11437 10424
rect 11471 10452 11483 10455
rect 11698 10452 11704 10464
rect 11471 10424 11704 10452
rect 11471 10421 11483 10424
rect 11425 10415 11483 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13354 10452 13360 10464
rect 12943 10424 13360 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13354 10412 13360 10424
rect 13412 10412 13418 10464
rect 14458 10452 14464 10464
rect 14419 10424 14464 10452
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 2096 10220 2789 10248
rect 2096 10208 2102 10220
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 4062 10248 4068 10260
rect 4023 10220 4068 10248
rect 2777 10211 2835 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 5997 10251 6055 10257
rect 5997 10217 6009 10251
rect 6043 10248 6055 10251
rect 6086 10248 6092 10260
rect 6043 10220 6092 10248
rect 6043 10217 6055 10220
rect 5997 10211 6055 10217
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7064 10220 7941 10248
rect 7064 10208 7070 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 8386 10248 8392 10260
rect 8347 10220 8392 10248
rect 7929 10211 7987 10217
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 9674 10248 9680 10260
rect 9635 10220 9680 10248
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 10042 10248 10048 10260
rect 10003 10220 10048 10248
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 11146 10248 11152 10260
rect 11107 10220 11152 10248
rect 11146 10208 11152 10220
rect 11204 10208 11210 10260
rect 11241 10251 11299 10257
rect 11241 10217 11253 10251
rect 11287 10248 11299 10251
rect 12437 10251 12495 10257
rect 11287 10220 12388 10248
rect 11287 10217 11299 10220
rect 11241 10211 11299 10217
rect 4338 10140 4344 10192
rect 4396 10180 4402 10192
rect 4396 10152 4660 10180
rect 4396 10140 4402 10152
rect 1670 10121 1676 10124
rect 1664 10075 1676 10121
rect 1728 10112 1734 10124
rect 3881 10115 3939 10121
rect 1728 10084 1764 10112
rect 1670 10072 1676 10075
rect 1728 10072 1734 10084
rect 3881 10081 3893 10115
rect 3927 10112 3939 10115
rect 4062 10112 4068 10124
rect 3927 10084 4068 10112
rect 3927 10081 3939 10084
rect 3881 10075 3939 10081
rect 4062 10072 4068 10084
rect 4120 10112 4126 10124
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 4120 10084 4445 10112
rect 4120 10072 4126 10084
rect 4433 10081 4445 10084
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10013 1455 10047
rect 4522 10044 4528 10056
rect 4483 10016 4528 10044
rect 1397 10007 1455 10013
rect 1412 9908 1440 10007
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 4632 10053 4660 10152
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 5592 10152 6132 10180
rect 5592 10140 5598 10152
rect 5626 10112 5632 10124
rect 5552 10084 5632 10112
rect 4617 10047 4675 10053
rect 4617 10013 4629 10047
rect 4663 10013 4675 10047
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 4617 10007 4675 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 5552 10053 5580 10084
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 6104 10112 6132 10152
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 8297 10183 8355 10189
rect 8297 10180 8309 10183
rect 8260 10152 8309 10180
rect 8260 10140 8266 10152
rect 8297 10149 8309 10152
rect 8343 10180 8355 10183
rect 10134 10180 10140 10192
rect 8343 10152 10140 10180
rect 8343 10149 8355 10152
rect 8297 10143 8355 10149
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 11701 10183 11759 10189
rect 11701 10149 11713 10183
rect 11747 10180 11759 10183
rect 11790 10180 11796 10192
rect 11747 10152 11796 10180
rect 11747 10149 11759 10152
rect 11701 10143 11759 10149
rect 11790 10140 11796 10152
rect 11848 10140 11854 10192
rect 12360 10180 12388 10220
rect 12437 10217 12449 10251
rect 12483 10248 12495 10251
rect 12618 10248 12624 10260
rect 12483 10220 12624 10248
rect 12483 10217 12495 10220
rect 12437 10211 12495 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13262 10248 13268 10260
rect 13223 10220 13268 10248
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13722 10180 13728 10192
rect 12360 10152 12940 10180
rect 13683 10152 13728 10180
rect 6104 10084 6224 10112
rect 6196 10053 6224 10084
rect 9858 10072 9864 10124
rect 9916 10112 9922 10124
rect 10502 10112 10508 10124
rect 9916 10084 10508 10112
rect 9916 10072 9922 10084
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10013 6147 10047
rect 6089 10007 6147 10013
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 8846 10044 8852 10056
rect 8619 10016 8852 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 2682 9936 2688 9988
rect 2740 9976 2746 9988
rect 3421 9979 3479 9985
rect 3421 9976 3433 9979
rect 2740 9948 3433 9976
rect 2740 9936 2746 9948
rect 3421 9945 3433 9948
rect 3467 9976 3479 9979
rect 5629 9979 5687 9985
rect 5629 9976 5641 9979
rect 3467 9948 5641 9976
rect 3467 9945 3479 9948
rect 3421 9939 3479 9945
rect 5629 9945 5641 9948
rect 5675 9945 5687 9979
rect 6104 9976 6132 10007
rect 8846 10004 8852 10016
rect 8904 10044 8910 10056
rect 10152 10053 10180 10084
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 11606 10112 11612 10124
rect 11567 10084 11612 10112
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 12912 10121 12940 10152
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 12805 10115 12863 10121
rect 12805 10112 12817 10115
rect 12492 10084 12817 10112
rect 12492 10072 12498 10084
rect 12805 10081 12817 10084
rect 12851 10081 12863 10115
rect 12805 10075 12863 10081
rect 12897 10115 12955 10121
rect 12897 10081 12909 10115
rect 12943 10112 12955 10115
rect 13078 10112 13084 10124
rect 12943 10084 13084 10112
rect 12943 10081 12955 10084
rect 12897 10075 12955 10081
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 13633 10115 13691 10121
rect 13633 10081 13645 10115
rect 13679 10112 13691 10115
rect 14366 10112 14372 10124
rect 13679 10084 14372 10112
rect 13679 10081 13691 10084
rect 13633 10075 13691 10081
rect 14366 10072 14372 10084
rect 14424 10072 14430 10124
rect 10137 10047 10195 10053
rect 8904 10016 9168 10044
rect 8904 10004 8910 10016
rect 6454 9976 6460 9988
rect 6104 9948 6460 9976
rect 5629 9939 5687 9945
rect 6454 9936 6460 9948
rect 6512 9936 6518 9988
rect 7006 9936 7012 9988
rect 7064 9976 7070 9988
rect 9140 9985 9168 10016
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 10226 10004 10232 10056
rect 10284 10044 10290 10056
rect 11882 10044 11888 10056
rect 10284 10016 10329 10044
rect 11843 10016 11888 10044
rect 10284 10004 10290 10016
rect 11882 10004 11888 10016
rect 11940 10004 11946 10056
rect 12250 10004 12256 10056
rect 12308 10044 12314 10056
rect 12989 10047 13047 10053
rect 12989 10044 13001 10047
rect 12308 10016 13001 10044
rect 12308 10004 12314 10016
rect 12989 10013 13001 10016
rect 13035 10013 13047 10047
rect 13814 10044 13820 10056
rect 13775 10016 13820 10044
rect 12989 10007 13047 10013
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 15286 10044 15292 10056
rect 15247 10016 15292 10044
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 7377 9979 7435 9985
rect 7377 9976 7389 9979
rect 7064 9948 7389 9976
rect 7064 9936 7070 9948
rect 7377 9945 7389 9948
rect 7423 9976 7435 9979
rect 7653 9979 7711 9985
rect 7653 9976 7665 9979
rect 7423 9948 7665 9976
rect 7423 9945 7435 9948
rect 7377 9939 7435 9945
rect 7653 9945 7665 9948
rect 7699 9945 7711 9979
rect 7653 9939 7711 9945
rect 9125 9979 9183 9985
rect 9125 9945 9137 9979
rect 9171 9976 9183 9979
rect 9493 9979 9551 9985
rect 9493 9976 9505 9979
rect 9171 9948 9505 9976
rect 9171 9945 9183 9948
rect 9125 9939 9183 9945
rect 9493 9945 9505 9948
rect 9539 9976 9551 9979
rect 10244 9976 10272 10004
rect 9539 9948 10272 9976
rect 9539 9945 9551 9948
rect 9493 9939 9551 9945
rect 2314 9908 2320 9920
rect 1412 9880 2320 9908
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 6917 9911 6975 9917
rect 6917 9877 6929 9911
rect 6963 9908 6975 9911
rect 7098 9908 7104 9920
rect 6963 9880 7104 9908
rect 6963 9877 6975 9880
rect 6917 9871 6975 9877
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 10689 9911 10747 9917
rect 10689 9908 10701 9911
rect 8536 9880 10701 9908
rect 8536 9868 8542 9880
rect 10689 9877 10701 9880
rect 10735 9877 10747 9911
rect 12342 9908 12348 9920
rect 12303 9880 12348 9908
rect 10689 9871 10747 9877
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 13998 9868 14004 9920
rect 14056 9908 14062 9920
rect 14277 9911 14335 9917
rect 14277 9908 14289 9911
rect 14056 9880 14289 9908
rect 14056 9868 14062 9880
rect 14277 9877 14289 9880
rect 14323 9908 14335 9911
rect 14642 9908 14648 9920
rect 14323 9880 14648 9908
rect 14323 9877 14335 9880
rect 14277 9871 14335 9877
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1670 9704 1676 9716
rect 1631 9676 1676 9704
rect 1670 9664 1676 9676
rect 1728 9704 1734 9716
rect 2041 9707 2099 9713
rect 2041 9704 2053 9707
rect 1728 9676 2053 9704
rect 1728 9664 1734 9676
rect 2041 9673 2053 9676
rect 2087 9673 2099 9707
rect 4522 9704 4528 9716
rect 2041 9667 2099 9673
rect 3804 9676 4528 9704
rect 2056 9568 2084 9667
rect 2590 9596 2596 9648
rect 2648 9636 2654 9648
rect 3329 9639 3387 9645
rect 3329 9636 3341 9639
rect 2648 9608 3341 9636
rect 2648 9596 2654 9608
rect 3329 9605 3341 9608
rect 3375 9636 3387 9639
rect 3804 9636 3832 9676
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 5074 9664 5080 9716
rect 5132 9704 5138 9716
rect 5169 9707 5227 9713
rect 5169 9704 5181 9707
rect 5132 9676 5181 9704
rect 5132 9664 5138 9676
rect 5169 9673 5181 9676
rect 5215 9673 5227 9707
rect 5169 9667 5227 9673
rect 5813 9707 5871 9713
rect 5813 9673 5825 9707
rect 5859 9704 5871 9707
rect 6454 9704 6460 9716
rect 5859 9676 6460 9704
rect 5859 9673 5871 9676
rect 5813 9667 5871 9673
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 7156 9676 8340 9704
rect 7156 9664 7162 9676
rect 3375 9608 3832 9636
rect 8312 9636 8340 9676
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 8757 9707 8815 9713
rect 8757 9704 8769 9707
rect 8444 9676 8769 9704
rect 8444 9664 8450 9676
rect 8757 9673 8769 9676
rect 8803 9704 8815 9707
rect 11149 9707 11207 9713
rect 11149 9704 11161 9707
rect 8803 9676 11161 9704
rect 8803 9673 8815 9676
rect 8757 9667 8815 9673
rect 11149 9673 11161 9676
rect 11195 9704 11207 9707
rect 11606 9704 11612 9716
rect 11195 9676 11612 9704
rect 11195 9673 11207 9676
rect 11149 9667 11207 9673
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 13136 9676 13952 9704
rect 13136 9664 13142 9676
rect 9493 9639 9551 9645
rect 9493 9636 9505 9639
rect 8312 9608 9505 9636
rect 3375 9605 3387 9608
rect 3329 9599 3387 9605
rect 9493 9605 9505 9608
rect 9539 9605 9551 9639
rect 10502 9636 10508 9648
rect 10463 9608 10508 9636
rect 9493 9599 9551 9605
rect 10502 9596 10508 9608
rect 10560 9596 10566 9648
rect 13814 9636 13820 9648
rect 13775 9608 13820 9636
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 13924 9636 13952 9676
rect 14642 9664 14648 9716
rect 14700 9704 14706 9716
rect 14700 9676 15148 9704
rect 14700 9664 14706 9676
rect 14737 9639 14795 9645
rect 14737 9636 14749 9639
rect 13924 9608 14749 9636
rect 14737 9605 14749 9608
rect 14783 9605 14795 9639
rect 15120 9636 15148 9676
rect 15378 9636 15384 9648
rect 15120 9608 15384 9636
rect 14737 9599 14795 9605
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 2056 9540 2881 9568
rect 2869 9537 2881 9540
rect 2915 9568 2927 9571
rect 6641 9571 6699 9577
rect 2915 9540 3924 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 2593 9503 2651 9509
rect 2593 9469 2605 9503
rect 2639 9500 2651 9503
rect 2682 9500 2688 9512
rect 2639 9472 2688 9500
rect 2639 9469 2651 9472
rect 2593 9463 2651 9469
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 3510 9460 3516 9512
rect 3568 9500 3574 9512
rect 3789 9503 3847 9509
rect 3789 9500 3801 9503
rect 3568 9472 3801 9500
rect 3568 9460 3574 9472
rect 3789 9469 3801 9472
rect 3835 9469 3847 9503
rect 3896 9500 3924 9540
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 10134 9568 10140 9580
rect 6687 9540 6960 9568
rect 10095 9540 10140 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 5074 9500 5080 9512
rect 3896 9472 5080 9500
rect 3789 9463 3847 9469
rect 5074 9460 5080 9472
rect 5132 9460 5138 9512
rect 6730 9460 6736 9512
rect 6788 9500 6794 9512
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6788 9472 6837 9500
rect 6788 9460 6794 9472
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 6932 9500 6960 9540
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 7092 9503 7150 9509
rect 7092 9500 7104 9503
rect 6932 9472 7104 9500
rect 6825 9463 6883 9469
rect 7092 9469 7104 9472
rect 7138 9500 7150 9503
rect 7466 9500 7472 9512
rect 7138 9472 7472 9500
rect 7138 9469 7150 9472
rect 7092 9463 7150 9469
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9824 9472 9873 9500
rect 9824 9460 9830 9472
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 11698 9460 11704 9512
rect 11756 9500 11762 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 11756 9472 12449 9500
rect 11756 9460 11762 9472
rect 12437 9469 12449 9472
rect 12483 9500 12495 9503
rect 13998 9500 14004 9512
rect 12483 9472 14004 9500
rect 12483 9469 12495 9472
rect 12437 9463 12495 9469
rect 13998 9460 14004 9472
rect 14056 9460 14062 9512
rect 3878 9392 3884 9444
rect 3936 9432 3942 9444
rect 4056 9435 4114 9441
rect 4056 9432 4068 9435
rect 3936 9404 4068 9432
rect 3936 9392 3942 9404
rect 4056 9401 4068 9404
rect 4102 9432 4114 9435
rect 4614 9432 4620 9444
rect 4102 9404 4620 9432
rect 4102 9401 4114 9404
rect 4056 9395 4114 9401
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 6454 9392 6460 9444
rect 6512 9432 6518 9444
rect 6914 9432 6920 9444
rect 6512 9404 6920 9432
rect 6512 9392 6518 9404
rect 6914 9392 6920 9404
rect 6972 9432 6978 9444
rect 9401 9435 9459 9441
rect 6972 9404 7065 9432
rect 6972 9392 6978 9404
rect 9401 9401 9413 9435
rect 9447 9432 9459 9435
rect 9953 9435 10011 9441
rect 9953 9432 9965 9435
rect 9447 9404 9965 9432
rect 9447 9401 9459 9404
rect 9401 9395 9459 9401
rect 9953 9401 9965 9404
rect 9999 9432 10011 9435
rect 10686 9432 10692 9444
rect 9999 9404 10692 9432
rect 9999 9401 10011 9404
rect 9953 9395 10011 9401
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 12342 9392 12348 9444
rect 12400 9432 12406 9444
rect 12682 9435 12740 9441
rect 12682 9432 12694 9435
rect 12400 9404 12694 9432
rect 12400 9392 12406 9404
rect 12682 9401 12694 9404
rect 12728 9401 12740 9435
rect 12682 9395 12740 9401
rect 2225 9367 2283 9373
rect 2225 9333 2237 9367
rect 2271 9364 2283 9367
rect 2314 9364 2320 9376
rect 2271 9336 2320 9364
rect 2271 9333 2283 9336
rect 2225 9327 2283 9333
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 2682 9364 2688 9376
rect 2643 9336 2688 9364
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 3697 9367 3755 9373
rect 3697 9333 3709 9367
rect 3743 9364 3755 9367
rect 4338 9364 4344 9376
rect 3743 9336 4344 9364
rect 3743 9333 3755 9336
rect 3697 9327 3755 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 6089 9367 6147 9373
rect 6089 9364 6101 9367
rect 6052 9336 6101 9364
rect 6052 9324 6058 9336
rect 6089 9333 6101 9336
rect 6135 9333 6147 9367
rect 6932 9364 6960 9392
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 6932 9336 8217 9364
rect 6089 9327 6147 9333
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 11330 9364 11336 9376
rect 11291 9336 11336 9364
rect 8205 9327 8263 9333
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 11790 9364 11796 9376
rect 11751 9336 11796 9364
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 12158 9364 12164 9376
rect 12119 9336 12164 9364
rect 12158 9324 12164 9336
rect 12216 9364 12222 9376
rect 12434 9364 12440 9376
rect 12216 9336 12440 9364
rect 12216 9324 12222 9336
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 14366 9364 14372 9376
rect 14327 9336 14372 9364
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 14826 9324 14832 9376
rect 14884 9364 14890 9376
rect 14921 9367 14979 9373
rect 14921 9364 14933 9367
rect 14884 9336 14933 9364
rect 14884 9324 14890 9336
rect 14921 9333 14933 9336
rect 14967 9333 14979 9367
rect 14921 9327 14979 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1578 9120 1584 9172
rect 1636 9160 1642 9172
rect 1857 9163 1915 9169
rect 1857 9160 1869 9163
rect 1636 9132 1869 9160
rect 1636 9120 1642 9132
rect 1857 9129 1869 9132
rect 1903 9129 1915 9163
rect 3878 9160 3884 9172
rect 3839 9132 3884 9160
rect 1857 9123 1915 9129
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 4062 9160 4068 9172
rect 4023 9132 4068 9160
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 4525 9163 4583 9169
rect 4525 9160 4537 9163
rect 4304 9132 4537 9160
rect 4304 9120 4310 9132
rect 4525 9129 4537 9132
rect 4571 9129 4583 9163
rect 4525 9123 4583 9129
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 4672 9132 5641 9160
rect 4672 9120 4678 9132
rect 5629 9129 5641 9132
rect 5675 9129 5687 9163
rect 8294 9160 8300 9172
rect 8255 9132 8300 9160
rect 5629 9123 5687 9129
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 8846 9160 8852 9172
rect 8807 9132 8852 9160
rect 8846 9120 8852 9132
rect 8904 9120 8910 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 9766 9160 9772 9172
rect 9539 9132 9772 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 9953 9163 10011 9169
rect 9953 9129 9965 9163
rect 9999 9160 10011 9163
rect 10042 9160 10048 9172
rect 9999 9132 10048 9160
rect 9999 9129 10011 9132
rect 9953 9123 10011 9129
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 11701 9163 11759 9169
rect 11701 9129 11713 9163
rect 11747 9160 11759 9163
rect 12250 9160 12256 9172
rect 11747 9132 12256 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 12986 9160 12992 9172
rect 12400 9132 12992 9160
rect 12400 9120 12406 9132
rect 12986 9120 12992 9132
rect 13044 9160 13050 9172
rect 13173 9163 13231 9169
rect 13173 9160 13185 9163
rect 13044 9132 13185 9160
rect 13044 9120 13050 9132
rect 13173 9129 13185 9132
rect 13219 9129 13231 9163
rect 13173 9123 13231 9129
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 14093 9163 14151 9169
rect 14093 9160 14105 9163
rect 13964 9132 14105 9160
rect 13964 9120 13970 9132
rect 14093 9129 14105 9132
rect 14139 9129 14151 9163
rect 14093 9123 14151 9129
rect 2314 9092 2320 9104
rect 2275 9064 2320 9092
rect 2314 9052 2320 9064
rect 2372 9092 2378 9104
rect 5077 9095 5135 9101
rect 5077 9092 5089 9095
rect 2372 9064 5089 9092
rect 2372 9052 2378 9064
rect 5077 9061 5089 9064
rect 5123 9061 5135 9095
rect 6362 9092 6368 9104
rect 5077 9055 5135 9061
rect 5828 9064 6368 9092
rect 2222 9024 2228 9036
rect 2183 8996 2228 9024
rect 2222 8984 2228 8996
rect 2280 8984 2286 9036
rect 2682 8984 2688 9036
rect 2740 9024 2746 9036
rect 3329 9027 3387 9033
rect 3329 9024 3341 9027
rect 2740 8996 3341 9024
rect 2740 8984 2746 8996
rect 3329 8993 3341 8996
rect 3375 9024 3387 9027
rect 3786 9024 3792 9036
rect 3375 8996 3792 9024
rect 3375 8993 3387 8996
rect 3329 8987 3387 8993
rect 3786 8984 3792 8996
rect 3844 8984 3850 9036
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4798 9024 4804 9036
rect 4479 8996 4804 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4798 8984 4804 8996
rect 4856 8984 4862 9036
rect 5828 9033 5856 9064
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 8021 9095 8079 9101
rect 8021 9061 8033 9095
rect 8067 9092 8079 9095
rect 8202 9092 8208 9104
rect 8067 9064 8208 9092
rect 8067 9061 8079 9064
rect 8021 9055 8079 9061
rect 8202 9052 8208 9064
rect 8260 9052 8266 9104
rect 11333 9095 11391 9101
rect 11333 9061 11345 9095
rect 11379 9092 11391 9095
rect 11882 9092 11888 9104
rect 11379 9064 11888 9092
rect 11379 9061 11391 9064
rect 11333 9055 11391 9061
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 13814 9092 13820 9104
rect 13775 9064 13820 9092
rect 13814 9052 13820 9064
rect 13872 9052 13878 9104
rect 6086 9033 6092 9036
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 8993 5871 9027
rect 6080 9024 6092 9033
rect 5999 8996 6092 9024
rect 5813 8987 5871 8993
rect 6080 8987 6092 8996
rect 6144 9024 6150 9036
rect 6454 9024 6460 9036
rect 6144 8996 6460 9024
rect 6086 8984 6092 8987
rect 6144 8984 6150 8996
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 10594 9024 10600 9036
rect 10555 8996 10600 9024
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 12060 9027 12118 9033
rect 12060 9024 12072 9027
rect 10888 8996 12072 9024
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 2038 8956 2044 8968
rect 1811 8928 2044 8956
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 2038 8916 2044 8928
rect 2096 8956 2102 8968
rect 2409 8959 2467 8965
rect 2409 8956 2421 8959
rect 2096 8928 2421 8956
rect 2096 8916 2102 8928
rect 2409 8925 2421 8928
rect 2455 8925 2467 8959
rect 2409 8919 2467 8925
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 10686 8956 10692 8968
rect 4755 8928 5212 8956
rect 10647 8928 10692 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 1486 8848 1492 8900
rect 1544 8888 1550 8900
rect 2869 8891 2927 8897
rect 2869 8888 2881 8891
rect 1544 8860 2881 8888
rect 1544 8848 1550 8860
rect 2869 8857 2881 8860
rect 2915 8857 2927 8891
rect 2869 8851 2927 8857
rect 5184 8832 5212 8928
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 10888 8965 10916 8996
rect 12060 8993 12072 8996
rect 12106 9024 12118 9027
rect 13538 9024 13544 9036
rect 12106 8996 13544 9024
rect 12106 8993 12118 8996
rect 12060 8987 12118 8993
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 15378 9024 15384 9036
rect 15339 8996 15384 9024
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 15654 9033 15660 9036
rect 15648 9024 15660 9033
rect 15615 8996 15660 9024
rect 15648 8987 15660 8996
rect 15654 8984 15660 8987
rect 15712 8984 15718 9036
rect 10873 8959 10931 8965
rect 10873 8925 10885 8959
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 9582 8848 9588 8900
rect 9640 8888 9646 8900
rect 10888 8888 10916 8919
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11698 8956 11704 8968
rect 11296 8928 11704 8956
rect 11296 8916 11302 8928
rect 11698 8916 11704 8928
rect 11756 8956 11762 8968
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 11756 8928 11805 8956
rect 11756 8916 11762 8928
rect 11793 8925 11805 8928
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 14458 8888 14464 8900
rect 9640 8860 10916 8888
rect 14419 8860 14464 8888
rect 9640 8848 9646 8860
rect 14458 8848 14464 8860
rect 14516 8848 14522 8900
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 5224 8792 7205 8820
rect 5224 8780 5230 8792
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 10226 8820 10232 8832
rect 10187 8792 10232 8820
rect 7193 8783 7251 8789
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 14734 8780 14740 8832
rect 14792 8820 14798 8832
rect 14829 8823 14887 8829
rect 14829 8820 14841 8823
rect 14792 8792 14841 8820
rect 14792 8780 14798 8792
rect 14829 8789 14841 8792
rect 14875 8789 14887 8823
rect 16758 8820 16764 8832
rect 16719 8792 16764 8820
rect 14829 8783 14887 8789
rect 16758 8780 16764 8792
rect 16816 8780 16822 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 2593 8619 2651 8625
rect 2593 8616 2605 8619
rect 2188 8588 2605 8616
rect 2188 8576 2194 8588
rect 2593 8585 2605 8588
rect 2639 8585 2651 8619
rect 2593 8579 2651 8585
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 1762 8480 1768 8492
rect 1719 8452 1768 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 1762 8440 1768 8452
rect 1820 8440 1826 8492
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1486 8412 1492 8424
rect 1443 8384 1492 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1486 8372 1492 8384
rect 1544 8372 1550 8424
rect 2608 8344 2636 8579
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 4157 8619 4215 8625
rect 4157 8616 4169 8619
rect 3936 8588 4169 8616
rect 3936 8576 3942 8588
rect 4157 8585 4169 8588
rect 4203 8585 4215 8619
rect 4157 8579 4215 8585
rect 4246 8576 4252 8628
rect 4304 8616 4310 8628
rect 4709 8619 4767 8625
rect 4709 8616 4721 8619
rect 4304 8588 4721 8616
rect 4304 8576 4310 8588
rect 4709 8585 4721 8588
rect 4755 8585 4767 8619
rect 5166 8616 5172 8628
rect 5127 8588 5172 8616
rect 4709 8579 4767 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 6086 8616 6092 8628
rect 5675 8588 6092 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 7929 8619 7987 8625
rect 7929 8585 7941 8619
rect 7975 8616 7987 8619
rect 9030 8616 9036 8628
rect 7975 8588 9036 8616
rect 7975 8585 7987 8588
rect 7929 8579 7987 8585
rect 5442 8508 5448 8560
rect 5500 8548 5506 8560
rect 6825 8551 6883 8557
rect 6825 8548 6837 8551
rect 5500 8520 6837 8548
rect 5500 8508 5506 8520
rect 6825 8517 6837 8520
rect 6871 8517 6883 8551
rect 8386 8548 8392 8560
rect 8347 8520 8392 8548
rect 6825 8511 6883 8517
rect 8386 8508 8392 8520
rect 8444 8508 8450 8560
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 6914 8480 6920 8492
rect 6687 8452 6920 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 6914 8440 6920 8452
rect 6972 8480 6978 8492
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 6972 8452 7297 8480
rect 6972 8440 6978 8452
rect 7285 8449 7297 8452
rect 7331 8449 7343 8483
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 7285 8443 7343 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 2774 8412 2780 8424
rect 2735 8384 2780 8412
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 3418 8372 3424 8424
rect 3476 8412 3482 8424
rect 8202 8412 8208 8424
rect 3476 8384 8208 8412
rect 3476 8372 3482 8384
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 8588 8421 8616 8588
rect 9030 8576 9036 8588
rect 9088 8616 9094 8628
rect 9088 8588 9628 8616
rect 9088 8576 9094 8588
rect 9600 8548 9628 8588
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 9732 8588 10057 8616
rect 9732 8576 9738 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10686 8616 10692 8628
rect 10647 8588 10692 8616
rect 10045 8579 10103 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 11330 8576 11336 8628
rect 11388 8616 11394 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 11388 8588 12173 8616
rect 11388 8576 11394 8588
rect 12161 8585 12173 8588
rect 12207 8616 12219 8619
rect 12207 8588 12664 8616
rect 12207 8585 12219 8588
rect 12161 8579 12219 8585
rect 9600 8520 9904 8548
rect 9876 8480 9904 8520
rect 10594 8508 10600 8560
rect 10652 8548 10658 8560
rect 10965 8551 11023 8557
rect 10965 8548 10977 8551
rect 10652 8520 10977 8548
rect 10652 8508 10658 8520
rect 10965 8517 10977 8520
rect 11011 8517 11023 8551
rect 10965 8511 11023 8517
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 12492 8520 12537 8548
rect 12492 8508 12498 8520
rect 11606 8480 11612 8492
rect 9876 8452 11612 8480
rect 11606 8440 11612 8452
rect 11664 8480 11670 8492
rect 11790 8480 11796 8492
rect 11664 8452 11796 8480
rect 11664 8440 11670 8452
rect 11790 8440 11796 8452
rect 11848 8440 11854 8492
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12342 8480 12348 8492
rect 11931 8452 12348 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8412 8723 8415
rect 9674 8412 9680 8424
rect 8711 8384 9680 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 2866 8344 2872 8356
rect 2608 8316 2872 8344
rect 2866 8304 2872 8316
rect 2924 8344 2930 8356
rect 3022 8347 3080 8353
rect 3022 8344 3034 8347
rect 2924 8316 3034 8344
rect 2924 8304 2930 8316
rect 3022 8313 3034 8316
rect 3068 8313 3080 8347
rect 5166 8344 5172 8356
rect 3022 8307 3080 8313
rect 4080 8316 5172 8344
rect 2038 8236 2044 8288
rect 2096 8276 2102 8288
rect 2133 8279 2191 8285
rect 2133 8276 2145 8279
rect 2096 8248 2145 8276
rect 2096 8236 2102 8248
rect 2133 8245 2145 8248
rect 2179 8245 2191 8279
rect 2133 8239 2191 8245
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 4080 8276 4108 8316
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 5718 8344 5724 8356
rect 5679 8316 5724 8344
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 6273 8347 6331 8353
rect 6273 8313 6285 8347
rect 6319 8344 6331 8347
rect 7190 8344 7196 8356
rect 6319 8316 7196 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 7190 8304 7196 8316
rect 7248 8304 7254 8356
rect 8297 8347 8355 8353
rect 8297 8313 8309 8347
rect 8343 8344 8355 8347
rect 8846 8344 8852 8356
rect 8343 8316 8852 8344
rect 8343 8313 8355 8316
rect 8297 8307 8355 8313
rect 8846 8304 8852 8316
rect 8904 8353 8910 8356
rect 8904 8347 8968 8353
rect 8904 8313 8922 8347
rect 8956 8313 8968 8347
rect 12636 8344 12664 8588
rect 15378 8576 15384 8628
rect 15436 8616 15442 8628
rect 17129 8619 17187 8625
rect 17129 8616 17141 8619
rect 15436 8588 17141 8616
rect 15436 8576 15442 8588
rect 17129 8585 17141 8588
rect 17175 8616 17187 8619
rect 17218 8616 17224 8628
rect 17175 8588 17224 8616
rect 17175 8585 17187 8588
rect 17129 8579 17187 8585
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 13538 8548 13544 8560
rect 13499 8520 13544 8548
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 14734 8508 14740 8560
rect 14792 8548 14798 8560
rect 15841 8551 15899 8557
rect 15841 8548 15853 8551
rect 14792 8520 15853 8548
rect 14792 8508 14798 8520
rect 15841 8517 15853 8520
rect 15887 8517 15899 8551
rect 15841 8511 15899 8517
rect 12986 8480 12992 8492
rect 12947 8452 12992 8480
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8480 14059 8483
rect 15102 8480 15108 8492
rect 14047 8452 15108 8480
rect 14047 8449 14059 8452
rect 14001 8443 14059 8449
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 16298 8480 16304 8492
rect 16259 8452 16304 8480
rect 16298 8440 16304 8452
rect 16356 8440 16362 8492
rect 12894 8412 12900 8424
rect 12855 8384 12900 8412
rect 12894 8372 12900 8384
rect 12952 8372 12958 8424
rect 14458 8372 14464 8424
rect 14516 8412 14522 8424
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 14516 8384 14841 8412
rect 14516 8372 14522 8384
rect 14829 8381 14841 8384
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 15930 8372 15936 8424
rect 15988 8412 15994 8424
rect 16025 8415 16083 8421
rect 16025 8412 16037 8415
rect 15988 8384 16037 8412
rect 15988 8372 15994 8384
rect 16025 8381 16037 8384
rect 16071 8412 16083 8415
rect 16761 8415 16819 8421
rect 16761 8412 16773 8415
rect 16071 8384 16773 8412
rect 16071 8381 16083 8384
rect 16025 8375 16083 8381
rect 16761 8381 16773 8384
rect 16807 8381 16819 8415
rect 20898 8412 20904 8424
rect 20859 8384 20904 8412
rect 16761 8375 16819 8381
rect 20898 8372 20904 8384
rect 20956 8412 20962 8424
rect 21637 8415 21695 8421
rect 21637 8412 21649 8415
rect 20956 8384 21649 8412
rect 20956 8372 20962 8384
rect 21637 8381 21649 8384
rect 21683 8381 21695 8415
rect 21637 8375 21695 8381
rect 12805 8347 12863 8353
rect 12805 8344 12817 8347
rect 12636 8316 12817 8344
rect 8904 8307 8968 8313
rect 12805 8313 12817 8316
rect 12851 8313 12863 8347
rect 12805 8307 12863 8313
rect 8904 8304 8910 8307
rect 13906 8304 13912 8356
rect 13964 8344 13970 8356
rect 14277 8347 14335 8353
rect 14277 8344 14289 8347
rect 13964 8316 14289 8344
rect 13964 8304 13970 8316
rect 14277 8313 14289 8316
rect 14323 8344 14335 8347
rect 14921 8347 14979 8353
rect 14921 8344 14933 8347
rect 14323 8316 14933 8344
rect 14323 8313 14335 8316
rect 14277 8307 14335 8313
rect 14921 8313 14933 8316
rect 14967 8313 14979 8347
rect 14921 8307 14979 8313
rect 15565 8347 15623 8353
rect 15565 8313 15577 8347
rect 15611 8344 15623 8347
rect 15654 8344 15660 8356
rect 15611 8316 15660 8344
rect 15611 8313 15623 8316
rect 15565 8307 15623 8313
rect 15654 8304 15660 8316
rect 15712 8344 15718 8356
rect 21177 8347 21235 8353
rect 15712 8316 16620 8344
rect 15712 8304 15718 8316
rect 3200 8248 4108 8276
rect 3200 8236 3206 8248
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 11333 8279 11391 8285
rect 11333 8276 11345 8279
rect 11204 8248 11345 8276
rect 11204 8236 11210 8248
rect 11333 8245 11345 8248
rect 11379 8245 11391 8279
rect 14458 8276 14464 8288
rect 14419 8248 14464 8276
rect 11333 8239 11391 8245
rect 14458 8236 14464 8248
rect 14516 8236 14522 8288
rect 16592 8276 16620 8316
rect 21177 8313 21189 8347
rect 21223 8344 21235 8347
rect 22002 8344 22008 8356
rect 21223 8316 22008 8344
rect 21223 8313 21235 8316
rect 21177 8307 21235 8313
rect 22002 8304 22008 8316
rect 22060 8304 22066 8356
rect 16666 8276 16672 8288
rect 16592 8248 16672 8276
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1394 8072 1400 8084
rect 1355 8044 1400 8072
rect 1394 8032 1400 8044
rect 1452 8032 1458 8084
rect 2409 8075 2467 8081
rect 2409 8041 2421 8075
rect 2455 8072 2467 8075
rect 2590 8072 2596 8084
rect 2455 8044 2596 8072
rect 2455 8041 2467 8044
rect 2409 8035 2467 8041
rect 2590 8032 2596 8044
rect 2648 8032 2654 8084
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 2958 8072 2964 8084
rect 2823 8044 2964 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 2958 8032 2964 8044
rect 3016 8072 3022 8084
rect 3510 8072 3516 8084
rect 3016 8044 3516 8072
rect 3016 8032 3022 8044
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 3927 8044 5089 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 5077 8041 5089 8044
rect 5123 8072 5135 8075
rect 5442 8072 5448 8084
rect 5123 8044 5448 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6604 8044 6653 8072
rect 6604 8032 6610 8044
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 7834 8072 7840 8084
rect 7795 8044 7840 8072
rect 6641 8035 6699 8041
rect 4341 8007 4399 8013
rect 4341 7973 4353 8007
rect 4387 8004 4399 8007
rect 4798 8004 4804 8016
rect 4387 7976 4804 8004
rect 4387 7973 4399 7976
rect 4341 7967 4399 7973
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 5258 7964 5264 8016
rect 5316 8004 5322 8016
rect 5721 8007 5779 8013
rect 5721 8004 5733 8007
rect 5316 7976 5733 8004
rect 5316 7964 5322 7976
rect 5721 7973 5733 7976
rect 5767 7973 5779 8007
rect 6656 8004 6684 8035
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 8202 8072 8208 8084
rect 8163 8044 8208 8072
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 8478 8032 8484 8084
rect 8536 8072 8542 8084
rect 8849 8075 8907 8081
rect 8849 8072 8861 8075
rect 8536 8044 8861 8072
rect 8536 8032 8542 8044
rect 8849 8041 8861 8044
rect 8895 8041 8907 8075
rect 8849 8035 8907 8041
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9582 8072 9588 8084
rect 9539 8044 9588 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10321 8075 10379 8081
rect 10321 8072 10333 8075
rect 10008 8044 10333 8072
rect 10008 8032 10014 8044
rect 10321 8041 10333 8044
rect 10367 8072 10379 8075
rect 10686 8072 10692 8084
rect 10367 8044 10692 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 7006 8004 7012 8016
rect 6656 7976 7012 8004
rect 5721 7967 5779 7973
rect 7006 7964 7012 7976
rect 7064 7964 7070 8016
rect 10134 7964 10140 8016
rect 10192 8004 10198 8016
rect 10229 8007 10287 8013
rect 10229 8004 10241 8007
rect 10192 7976 10241 8004
rect 10192 7964 10198 7976
rect 10229 7973 10241 7976
rect 10275 7973 10287 8007
rect 11054 8004 11060 8016
rect 10229 7967 10287 7973
rect 10336 7976 11060 8004
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7936 5227 7939
rect 5350 7936 5356 7948
rect 5215 7908 5356 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 7282 7896 7288 7948
rect 7340 7936 7346 7948
rect 8297 7939 8355 7945
rect 8297 7936 8309 7939
rect 7340 7908 8309 7936
rect 7340 7896 7346 7908
rect 8297 7905 8309 7908
rect 8343 7936 8355 7939
rect 10336 7936 10364 7976
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 11698 7945 11704 7948
rect 8343 7908 10364 7936
rect 10965 7939 11023 7945
rect 8343 7905 8355 7908
rect 8297 7899 8355 7905
rect 10965 7905 10977 7939
rect 11011 7936 11023 7939
rect 11692 7936 11704 7945
rect 11011 7908 11704 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 11692 7899 11704 7908
rect 11698 7896 11704 7899
rect 11756 7896 11762 7948
rect 15102 7896 15108 7948
rect 15160 7936 15166 7948
rect 15562 7945 15568 7948
rect 15556 7936 15568 7945
rect 15160 7908 15568 7936
rect 15160 7896 15166 7908
rect 15556 7899 15568 7908
rect 15562 7896 15568 7899
rect 15620 7896 15626 7948
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2556 7840 2881 7868
rect 2556 7828 2562 7840
rect 2869 7837 2881 7840
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3142 7868 3148 7880
rect 3099 7840 3148 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3234 7828 3240 7880
rect 3292 7868 3298 7880
rect 3292 7840 4936 7868
rect 3292 7828 3298 7840
rect 1762 7760 1768 7812
rect 1820 7800 1826 7812
rect 2225 7803 2283 7809
rect 2225 7800 2237 7803
rect 1820 7772 2237 7800
rect 1820 7760 1826 7772
rect 2225 7769 2237 7772
rect 2271 7769 2283 7803
rect 2225 7763 2283 7769
rect 1854 7732 1860 7744
rect 1815 7704 1860 7732
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 3234 7692 3240 7744
rect 3292 7732 3298 7744
rect 3421 7735 3479 7741
rect 3421 7732 3433 7735
rect 3292 7704 3433 7732
rect 3292 7692 3298 7704
rect 3421 7701 3433 7704
rect 3467 7701 3479 7735
rect 4706 7732 4712 7744
rect 4667 7704 4712 7732
rect 3421 7695 3479 7701
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 4908 7732 4936 7840
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 6730 7868 6736 7880
rect 5316 7840 5361 7868
rect 6691 7840 6736 7868
rect 5316 7828 5322 7840
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7868 10563 7871
rect 11054 7868 11060 7880
rect 10551 7840 11060 7868
rect 10551 7837 10563 7840
rect 10505 7831 10563 7837
rect 6178 7800 6184 7812
rect 6139 7772 6184 7800
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 6932 7800 6960 7831
rect 7742 7800 7748 7812
rect 6932 7772 7748 7800
rect 7742 7760 7748 7772
rect 7800 7760 7806 7812
rect 7926 7760 7932 7812
rect 7984 7800 7990 7812
rect 8404 7800 8432 7831
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11330 7828 11336 7880
rect 11388 7868 11394 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11388 7840 11437 7868
rect 11388 7828 11394 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 14182 7868 14188 7880
rect 14143 7840 14188 7868
rect 11425 7831 11483 7837
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 15286 7868 15292 7880
rect 15247 7840 15292 7868
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 7984 7772 8432 7800
rect 9861 7803 9919 7809
rect 7984 7760 7990 7772
rect 9861 7769 9873 7803
rect 9907 7800 9919 7803
rect 11238 7800 11244 7812
rect 9907 7772 11244 7800
rect 9907 7769 9919 7772
rect 9861 7763 9919 7769
rect 11238 7760 11244 7772
rect 11296 7760 11302 7812
rect 12802 7800 12808 7812
rect 12763 7772 12808 7800
rect 12802 7760 12808 7772
rect 12860 7760 12866 7812
rect 6086 7732 6092 7744
rect 4908 7704 6092 7732
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6270 7732 6276 7744
rect 6231 7704 6276 7732
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 7377 7735 7435 7741
rect 7377 7701 7389 7735
rect 7423 7732 7435 7735
rect 7466 7732 7472 7744
rect 7423 7704 7472 7732
rect 7423 7701 7435 7704
rect 7377 7695 7435 7701
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 13449 7735 13507 7741
rect 13449 7701 13461 7735
rect 13495 7732 13507 7735
rect 13630 7732 13636 7744
rect 13495 7704 13636 7732
rect 13495 7701 13507 7704
rect 13449 7695 13507 7701
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 13817 7735 13875 7741
rect 13817 7701 13829 7735
rect 13863 7732 13875 7735
rect 13998 7732 14004 7744
rect 13863 7704 14004 7732
rect 13863 7701 13875 7704
rect 13817 7695 13875 7701
rect 13998 7692 14004 7704
rect 14056 7732 14062 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 14056 7704 14657 7732
rect 14056 7692 14062 7704
rect 14645 7701 14657 7704
rect 14691 7732 14703 7735
rect 14734 7732 14740 7744
rect 14691 7704 14740 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 14734 7692 14740 7704
rect 14792 7732 14798 7744
rect 15013 7735 15071 7741
rect 15013 7732 15025 7735
rect 14792 7704 15025 7732
rect 14792 7692 14798 7704
rect 15013 7701 15025 7704
rect 15059 7701 15071 7735
rect 16666 7732 16672 7744
rect 16627 7704 16672 7732
rect 15013 7695 15071 7701
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1397 7531 1455 7537
rect 1397 7497 1409 7531
rect 1443 7528 1455 7531
rect 3234 7528 3240 7540
rect 1443 7500 3240 7528
rect 1443 7497 1455 7500
rect 1397 7491 1455 7497
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 4985 7531 5043 7537
rect 4985 7497 4997 7531
rect 5031 7528 5043 7531
rect 5258 7528 5264 7540
rect 5031 7500 5264 7528
rect 5031 7497 5043 7500
rect 4985 7491 5043 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 6365 7531 6423 7537
rect 6365 7497 6377 7531
rect 6411 7528 6423 7531
rect 6454 7528 6460 7540
rect 6411 7500 6460 7528
rect 6411 7497 6423 7500
rect 6365 7491 6423 7497
rect 6454 7488 6460 7500
rect 6512 7528 6518 7540
rect 6730 7528 6736 7540
rect 6512 7500 6736 7528
rect 6512 7488 6518 7500
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7006 7528 7012 7540
rect 6967 7500 7012 7528
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7469 7531 7527 7537
rect 7469 7528 7481 7531
rect 7340 7500 7481 7528
rect 7340 7488 7346 7500
rect 7469 7497 7481 7500
rect 7515 7497 7527 7531
rect 9950 7528 9956 7540
rect 9911 7500 9956 7528
rect 7469 7491 7527 7497
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10229 7531 10287 7537
rect 10229 7528 10241 7531
rect 10192 7500 10241 7528
rect 10192 7488 10198 7500
rect 10229 7497 10241 7500
rect 10275 7497 10287 7531
rect 10229 7491 10287 7497
rect 10686 7488 10692 7540
rect 10744 7528 10750 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 10744 7500 12173 7528
rect 10744 7488 10750 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12161 7491 12219 7497
rect 12713 7531 12771 7537
rect 12713 7497 12725 7531
rect 12759 7528 12771 7531
rect 12894 7528 12900 7540
rect 12759 7500 12900 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 14461 7531 14519 7537
rect 14461 7497 14473 7531
rect 14507 7528 14519 7531
rect 15562 7528 15568 7540
rect 14507 7500 15568 7528
rect 14507 7497 14519 7500
rect 14461 7491 14519 7497
rect 15562 7488 15568 7500
rect 15620 7488 15626 7540
rect 17218 7528 17224 7540
rect 17179 7500 17224 7528
rect 17218 7488 17224 7500
rect 17276 7528 17282 7540
rect 17589 7531 17647 7537
rect 17589 7528 17601 7531
rect 17276 7500 17601 7528
rect 17276 7488 17282 7500
rect 17589 7497 17601 7500
rect 17635 7497 17647 7531
rect 17589 7491 17647 7497
rect 2869 7463 2927 7469
rect 2869 7429 2881 7463
rect 2915 7460 2927 7463
rect 2958 7460 2964 7472
rect 2915 7432 2964 7460
rect 2915 7429 2927 7432
rect 2869 7423 2927 7429
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 3970 7420 3976 7472
rect 4028 7460 4034 7472
rect 4338 7460 4344 7472
rect 4028 7432 4344 7460
rect 4028 7420 4034 7432
rect 4338 7420 4344 7432
rect 4396 7420 4402 7472
rect 5445 7463 5503 7469
rect 5445 7429 5457 7463
rect 5491 7460 5503 7463
rect 5626 7460 5632 7472
rect 5491 7432 5632 7460
rect 5491 7429 5503 7432
rect 5445 7423 5503 7429
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2682 7284 2688 7336
rect 2740 7324 2746 7336
rect 2961 7327 3019 7333
rect 2961 7324 2973 7327
rect 2740 7296 2973 7324
rect 2740 7284 2746 7296
rect 2961 7293 2973 7296
rect 3007 7324 3019 7327
rect 5460 7324 5488 7423
rect 5626 7420 5632 7432
rect 5684 7420 5690 7472
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 10505 7463 10563 7469
rect 10505 7460 10517 7463
rect 9732 7432 10517 7460
rect 9732 7420 9738 7432
rect 10505 7429 10517 7432
rect 10551 7460 10563 7463
rect 11330 7460 11336 7472
rect 10551 7432 11336 7460
rect 10551 7429 10563 7432
rect 10505 7423 10563 7429
rect 11330 7420 11336 7432
rect 11388 7420 11394 7472
rect 11238 7392 11244 7404
rect 11199 7364 11244 7392
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 11425 7395 11483 7401
rect 11425 7361 11437 7395
rect 11471 7392 11483 7395
rect 11698 7392 11704 7404
rect 11471 7364 11704 7392
rect 11471 7361 11483 7364
rect 11425 7355 11483 7361
rect 11698 7352 11704 7364
rect 11756 7392 11762 7404
rect 11756 7364 11928 7392
rect 11756 7352 11762 7364
rect 3007 7296 5488 7324
rect 5629 7327 5687 7333
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 5629 7293 5641 7327
rect 5675 7324 5687 7327
rect 6178 7324 6184 7336
rect 5675 7296 6184 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 7653 7327 7711 7333
rect 7653 7324 7665 7327
rect 7616 7296 7665 7324
rect 7616 7284 7622 7296
rect 7653 7293 7665 7296
rect 7699 7293 7711 7327
rect 7653 7287 7711 7293
rect 7742 7284 7748 7336
rect 7800 7324 7806 7336
rect 7909 7327 7967 7333
rect 7909 7324 7921 7327
rect 7800 7296 7921 7324
rect 7800 7284 7806 7296
rect 7909 7293 7921 7296
rect 7955 7293 7967 7327
rect 10686 7324 10692 7336
rect 10647 7296 10692 7324
rect 7909 7287 7967 7293
rect 10686 7284 10692 7296
rect 10744 7284 10750 7336
rect 11146 7324 11152 7336
rect 11107 7296 11152 7324
rect 11146 7284 11152 7296
rect 11204 7284 11210 7336
rect 1762 7256 1768 7268
rect 1723 7228 1768 7256
rect 1762 7216 1768 7228
rect 1820 7216 1826 7268
rect 3142 7216 3148 7268
rect 3200 7265 3206 7268
rect 3200 7259 3264 7265
rect 3200 7225 3218 7259
rect 3252 7225 3264 7259
rect 5350 7256 5356 7268
rect 5263 7228 5356 7256
rect 3200 7219 3264 7225
rect 3200 7216 3206 7219
rect 5350 7216 5356 7228
rect 5408 7256 5414 7268
rect 6086 7256 6092 7268
rect 5408 7228 6092 7256
rect 5408 7216 5414 7228
rect 6086 7216 6092 7228
rect 6144 7216 6150 7268
rect 1854 7188 1860 7200
rect 1815 7160 1860 7188
rect 1854 7148 1860 7160
rect 1912 7148 1918 7200
rect 2498 7188 2504 7200
rect 2459 7160 2504 7188
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 5718 7188 5724 7200
rect 5679 7160 5724 7188
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 8846 7148 8852 7200
rect 8904 7188 8910 7200
rect 9033 7191 9091 7197
rect 9033 7188 9045 7191
rect 8904 7160 9045 7188
rect 8904 7148 8910 7160
rect 9033 7157 9045 7160
rect 9079 7157 9091 7191
rect 10778 7188 10784 7200
rect 10739 7160 10784 7188
rect 9033 7151 9091 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11900 7197 11928 7364
rect 13630 7352 13636 7404
rect 13688 7392 13694 7404
rect 13814 7392 13820 7404
rect 13688 7364 13820 7392
rect 13688 7352 13694 7364
rect 13814 7352 13820 7364
rect 13872 7392 13878 7404
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13872 7364 13921 7392
rect 13872 7352 13878 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 13354 7284 13360 7336
rect 13412 7324 13418 7336
rect 13725 7327 13783 7333
rect 13725 7324 13737 7327
rect 13412 7296 13737 7324
rect 13412 7284 13418 7296
rect 13725 7293 13737 7296
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 15010 7324 15016 7336
rect 14967 7296 15016 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 18046 7324 18052 7336
rect 18007 7296 18052 7324
rect 18046 7284 18052 7296
rect 18104 7324 18110 7336
rect 18785 7327 18843 7333
rect 18785 7324 18797 7327
rect 18104 7296 18797 7324
rect 18104 7284 18110 7296
rect 18785 7293 18797 7296
rect 18831 7293 18843 7327
rect 18785 7287 18843 7293
rect 13817 7259 13875 7265
rect 13817 7256 13829 7259
rect 13188 7228 13829 7256
rect 11885 7191 11943 7197
rect 11885 7157 11897 7191
rect 11931 7188 11943 7191
rect 12342 7188 12348 7200
rect 11931 7160 12348 7188
rect 11931 7157 11943 7160
rect 11885 7151 11943 7157
rect 12342 7148 12348 7160
rect 12400 7148 12406 7200
rect 12894 7148 12900 7200
rect 12952 7188 12958 7200
rect 13188 7197 13216 7228
rect 13817 7225 13829 7228
rect 13863 7256 13875 7259
rect 13906 7256 13912 7268
rect 13863 7228 13912 7256
rect 13863 7225 13875 7228
rect 13817 7219 13875 7225
rect 13906 7216 13912 7228
rect 13964 7216 13970 7268
rect 14829 7259 14887 7265
rect 14829 7225 14841 7259
rect 14875 7256 14887 7259
rect 15188 7259 15246 7265
rect 15188 7256 15200 7259
rect 14875 7228 15200 7256
rect 14875 7225 14887 7228
rect 14829 7219 14887 7225
rect 15188 7225 15200 7228
rect 15234 7256 15246 7259
rect 15838 7256 15844 7268
rect 15234 7228 15844 7256
rect 15234 7225 15246 7228
rect 15188 7219 15246 7225
rect 15838 7216 15844 7228
rect 15896 7216 15902 7268
rect 18322 7256 18328 7268
rect 18283 7228 18328 7256
rect 18322 7216 18328 7228
rect 18380 7216 18386 7268
rect 13173 7191 13231 7197
rect 13173 7188 13185 7191
rect 12952 7160 13185 7188
rect 12952 7148 12958 7160
rect 13173 7157 13185 7160
rect 13219 7157 13231 7191
rect 13173 7151 13231 7157
rect 13357 7191 13415 7197
rect 13357 7157 13369 7191
rect 13403 7188 13415 7191
rect 13722 7188 13728 7200
rect 13403 7160 13728 7188
rect 13403 7157 13415 7160
rect 13357 7151 13415 7157
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 16298 7188 16304 7200
rect 16259 7160 16304 7188
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 16850 7188 16856 7200
rect 16811 7160 16856 7188
rect 16850 7148 16856 7160
rect 16908 7148 16914 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 3142 6944 3148 6996
rect 3200 6984 3206 6996
rect 3421 6987 3479 6993
rect 3421 6984 3433 6987
rect 3200 6956 3433 6984
rect 3200 6944 3206 6956
rect 3421 6953 3433 6956
rect 3467 6953 3479 6987
rect 3421 6947 3479 6953
rect 4430 6944 4436 6996
rect 4488 6984 4494 6996
rect 4798 6984 4804 6996
rect 4488 6956 4804 6984
rect 4488 6944 4494 6956
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 4982 6944 4988 6996
rect 5040 6984 5046 6996
rect 5442 6984 5448 6996
rect 5040 6956 5448 6984
rect 5040 6944 5046 6956
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 6365 6987 6423 6993
rect 6365 6953 6377 6987
rect 6411 6984 6423 6987
rect 7742 6984 7748 6996
rect 6411 6956 7748 6984
rect 6411 6953 6423 6956
rect 6365 6947 6423 6953
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 13354 6984 13360 6996
rect 13315 6956 13360 6984
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 14182 6944 14188 6996
rect 14240 6984 14246 6996
rect 15749 6987 15807 6993
rect 15749 6984 15761 6987
rect 14240 6956 15761 6984
rect 14240 6944 14246 6956
rect 15749 6953 15761 6956
rect 15795 6984 15807 6987
rect 16298 6984 16304 6996
rect 15795 6956 16304 6984
rect 15795 6953 15807 6956
rect 15749 6947 15807 6953
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 17218 6984 17224 6996
rect 17179 6956 17224 6984
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 19150 6984 19156 6996
rect 19111 6956 19156 6984
rect 19150 6944 19156 6956
rect 19208 6944 19214 6996
rect 5261 6919 5319 6925
rect 5261 6885 5273 6919
rect 5307 6916 5319 6919
rect 5350 6916 5356 6928
rect 5307 6888 5356 6916
rect 5307 6885 5319 6888
rect 5261 6879 5319 6885
rect 5350 6876 5356 6888
rect 5408 6876 5414 6928
rect 10042 6916 10048 6928
rect 10003 6888 10048 6916
rect 10042 6876 10048 6888
rect 10100 6876 10106 6928
rect 11146 6916 11152 6928
rect 11072 6888 11152 6916
rect 1756 6851 1814 6857
rect 1756 6817 1768 6851
rect 1802 6848 1814 6851
rect 2590 6848 2596 6860
rect 1802 6820 2596 6848
rect 1802 6817 1814 6820
rect 1756 6811 1814 6817
rect 2590 6808 2596 6820
rect 2648 6848 2654 6860
rect 3970 6848 3976 6860
rect 2648 6820 3976 6848
rect 2648 6808 2654 6820
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 6362 6848 6368 6860
rect 5684 6820 6368 6848
rect 5684 6808 5690 6820
rect 6362 6808 6368 6820
rect 6420 6848 6426 6860
rect 6730 6857 6736 6860
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 6420 6820 6469 6848
rect 6420 6808 6426 6820
rect 6457 6817 6469 6820
rect 6503 6817 6515 6851
rect 6724 6848 6736 6857
rect 6691 6820 6736 6848
rect 6457 6811 6515 6817
rect 6724 6811 6736 6820
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6749 1547 6783
rect 1489 6743 1547 6749
rect 1504 6644 1532 6743
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 5350 6780 5356 6792
rect 4212 6752 5356 6780
rect 4212 6740 4218 6752
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 2866 6712 2872 6724
rect 2827 6684 2872 6712
rect 2866 6672 2872 6684
rect 2924 6672 2930 6724
rect 3050 6672 3056 6724
rect 3108 6712 3114 6724
rect 3418 6712 3424 6724
rect 3108 6684 3424 6712
rect 3108 6672 3114 6684
rect 3418 6672 3424 6684
rect 3476 6672 3482 6724
rect 5166 6672 5172 6724
rect 5224 6712 5230 6724
rect 5460 6712 5488 6743
rect 5224 6684 5488 6712
rect 5224 6672 5230 6684
rect 2682 6644 2688 6656
rect 1504 6616 2688 6644
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 2832 6616 3801 6644
rect 2832 6604 2838 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 4246 6644 4252 6656
rect 4207 6616 4252 6644
rect 3789 6607 3847 6613
rect 4246 6604 4252 6616
rect 4304 6604 4310 6656
rect 4614 6604 4620 6656
rect 4672 6644 4678 6656
rect 4709 6647 4767 6653
rect 4709 6644 4721 6647
rect 4672 6616 4721 6644
rect 4672 6604 4678 6616
rect 4709 6613 4721 6616
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 4893 6647 4951 6653
rect 4893 6613 4905 6647
rect 4939 6644 4951 6647
rect 5994 6644 6000 6656
rect 4939 6616 6000 6644
rect 4939 6613 4951 6616
rect 4893 6607 4951 6613
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 6472 6644 6500 6811
rect 6730 6808 6736 6811
rect 6788 6808 6794 6860
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 8389 6851 8447 6857
rect 8389 6848 8401 6851
rect 8352 6820 8401 6848
rect 8352 6808 8358 6820
rect 8389 6817 8401 6820
rect 8435 6817 8447 6851
rect 9490 6848 9496 6860
rect 9451 6820 9496 6848
rect 8389 6811 8447 6817
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 9858 6848 9864 6860
rect 9732 6820 9864 6848
rect 9732 6808 9738 6820
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 10873 6851 10931 6857
rect 10873 6817 10885 6851
rect 10919 6848 10931 6851
rect 11072 6848 11100 6888
rect 11146 6876 11152 6888
rect 11204 6876 11210 6928
rect 13998 6876 14004 6928
rect 14056 6916 14062 6928
rect 14921 6919 14979 6925
rect 14921 6916 14933 6919
rect 14056 6888 14933 6916
rect 14056 6876 14062 6888
rect 14921 6885 14933 6888
rect 14967 6916 14979 6919
rect 15013 6919 15071 6925
rect 15013 6916 15025 6919
rect 14967 6888 15025 6916
rect 14967 6885 14979 6888
rect 14921 6879 14979 6885
rect 15013 6885 15025 6888
rect 15059 6885 15071 6919
rect 15013 6879 15071 6885
rect 24118 6876 24124 6928
rect 24176 6916 24182 6928
rect 24670 6916 24676 6928
rect 24176 6888 24676 6916
rect 24176 6876 24182 6888
rect 24670 6876 24676 6888
rect 24728 6876 24734 6928
rect 11514 6857 11520 6860
rect 11508 6848 11520 6857
rect 10919 6820 11100 6848
rect 11475 6820 11520 6848
rect 10919 6817 10931 6820
rect 10873 6811 10931 6817
rect 11508 6811 11520 6820
rect 11514 6808 11520 6811
rect 11572 6808 11578 6860
rect 13906 6848 13912 6860
rect 13867 6820 13912 6848
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 14458 6808 14464 6860
rect 14516 6848 14522 6860
rect 15841 6851 15899 6857
rect 15841 6848 15853 6851
rect 14516 6820 15853 6848
rect 14516 6808 14522 6820
rect 15841 6817 15853 6820
rect 15887 6817 15899 6851
rect 15841 6811 15899 6817
rect 18040 6851 18098 6857
rect 18040 6817 18052 6851
rect 18086 6848 18098 6851
rect 19058 6848 19064 6860
rect 18086 6820 19064 6848
rect 18086 6817 18098 6820
rect 18040 6811 18098 6817
rect 19058 6808 19064 6820
rect 19116 6808 19122 6860
rect 20898 6848 20904 6860
rect 20859 6820 20904 6848
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 9876 6752 10149 6780
rect 9876 6724 9904 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6749 11299 6783
rect 14182 6780 14188 6792
rect 14143 6752 14188 6780
rect 11241 6743 11299 6749
rect 7558 6712 7564 6724
rect 7392 6684 7564 6712
rect 7098 6644 7104 6656
rect 6472 6616 7104 6644
rect 7098 6604 7104 6616
rect 7156 6644 7162 6656
rect 7392 6644 7420 6684
rect 7558 6672 7564 6684
rect 7616 6672 7622 6724
rect 9858 6672 9864 6724
rect 9916 6672 9922 6724
rect 9950 6672 9956 6724
rect 10008 6712 10014 6724
rect 10244 6712 10272 6743
rect 10008 6684 10272 6712
rect 10008 6672 10014 6684
rect 7156 6616 7420 6644
rect 7156 6604 7162 6616
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 7524 6616 7849 6644
rect 7524 6604 7530 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 7837 6607 7895 6613
rect 8849 6647 8907 6653
rect 8849 6613 8861 6647
rect 8895 6644 8907 6647
rect 9306 6644 9312 6656
rect 8895 6616 9312 6644
rect 8895 6613 8907 6616
rect 8849 6607 8907 6613
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 9677 6647 9735 6653
rect 9677 6613 9689 6647
rect 9723 6644 9735 6647
rect 10778 6644 10784 6656
rect 9723 6616 10784 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 11256 6644 11284 6743
rect 14182 6740 14188 6752
rect 14240 6740 14246 6792
rect 16022 6780 16028 6792
rect 15983 6752 16028 6780
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 17773 6783 17831 6789
rect 17773 6780 17785 6783
rect 17604 6752 17785 6780
rect 12434 6672 12440 6724
rect 12492 6712 12498 6724
rect 12621 6715 12679 6721
rect 12621 6712 12633 6715
rect 12492 6684 12633 6712
rect 12492 6672 12498 6684
rect 12621 6681 12633 6684
rect 12667 6681 12679 6715
rect 15378 6712 15384 6724
rect 15339 6684 15384 6712
rect 12621 6675 12679 6681
rect 15378 6672 15384 6684
rect 15436 6672 15442 6724
rect 11882 6644 11888 6656
rect 11256 6616 11888 6644
rect 11882 6604 11888 6616
rect 11940 6644 11946 6656
rect 12342 6644 12348 6656
rect 11940 6616 12348 6644
rect 11940 6604 11946 6616
rect 12342 6604 12348 6616
rect 12400 6644 12406 6656
rect 13817 6647 13875 6653
rect 13817 6644 13829 6647
rect 12400 6616 13829 6644
rect 12400 6604 12406 6616
rect 13817 6613 13829 6616
rect 13863 6644 13875 6647
rect 14366 6644 14372 6656
rect 13863 6616 14372 6644
rect 13863 6613 13875 6616
rect 13817 6607 13875 6613
rect 14366 6604 14372 6616
rect 14424 6644 14430 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 14424 6616 14657 6644
rect 14424 6604 14430 6616
rect 14645 6613 14657 6616
rect 14691 6613 14703 6647
rect 14645 6607 14703 6613
rect 14921 6647 14979 6653
rect 14921 6613 14933 6647
rect 14967 6644 14979 6647
rect 16393 6647 16451 6653
rect 16393 6644 16405 6647
rect 14967 6616 16405 6644
rect 14967 6613 14979 6616
rect 14921 6607 14979 6613
rect 16393 6613 16405 6616
rect 16439 6644 16451 6647
rect 16761 6647 16819 6653
rect 16761 6644 16773 6647
rect 16439 6616 16773 6644
rect 16439 6613 16451 6616
rect 16393 6607 16451 6613
rect 16761 6613 16773 6616
rect 16807 6644 16819 6647
rect 16850 6644 16856 6656
rect 16807 6616 16856 6644
rect 16807 6613 16819 6616
rect 16761 6607 16819 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17604 6653 17632 6752
rect 17773 6749 17785 6752
rect 17819 6749 17831 6783
rect 21174 6780 21180 6792
rect 21135 6752 21180 6780
rect 17773 6743 17831 6749
rect 21174 6740 21180 6752
rect 21232 6740 21238 6792
rect 17589 6647 17647 6653
rect 17589 6644 17601 6647
rect 17276 6616 17601 6644
rect 17276 6604 17282 6616
rect 17589 6613 17601 6616
rect 17635 6613 17647 6647
rect 17589 6607 17647 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2685 6443 2743 6449
rect 2685 6409 2697 6443
rect 2731 6440 2743 6443
rect 3142 6440 3148 6452
rect 2731 6412 3148 6440
rect 2731 6409 2743 6412
rect 2685 6403 2743 6409
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 5350 6400 5356 6452
rect 5408 6440 5414 6452
rect 5721 6443 5779 6449
rect 5721 6440 5733 6443
rect 5408 6412 5733 6440
rect 5408 6400 5414 6412
rect 5721 6409 5733 6412
rect 5767 6409 5779 6443
rect 7926 6440 7932 6452
rect 7887 6412 7932 6440
rect 5721 6403 5779 6409
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 10100 6412 10517 6440
rect 10100 6400 10106 6412
rect 10505 6409 10517 6412
rect 10551 6409 10563 6443
rect 10505 6403 10563 6409
rect 11514 6400 11520 6452
rect 11572 6440 11578 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11572 6412 11805 6440
rect 11572 6400 11578 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14185 6443 14243 6449
rect 14185 6440 14197 6443
rect 13872 6412 14197 6440
rect 13872 6400 13878 6412
rect 14185 6409 14197 6412
rect 14231 6409 14243 6443
rect 14185 6403 14243 6409
rect 3510 6332 3516 6384
rect 3568 6372 3574 6384
rect 3786 6372 3792 6384
rect 3568 6344 3792 6372
rect 3568 6332 3574 6344
rect 3786 6332 3792 6344
rect 3844 6332 3850 6384
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 4709 6375 4767 6381
rect 4709 6372 4721 6375
rect 4120 6344 4721 6372
rect 4120 6332 4126 6344
rect 4709 6341 4721 6344
rect 4755 6341 4767 6375
rect 4709 6335 4767 6341
rect 9858 6332 9864 6384
rect 9916 6372 9922 6384
rect 10873 6375 10931 6381
rect 10873 6372 10885 6375
rect 9916 6344 10885 6372
rect 9916 6332 9922 6344
rect 10873 6341 10885 6344
rect 10919 6341 10931 6375
rect 10873 6335 10931 6341
rect 12434 6332 12440 6384
rect 12492 6372 12498 6384
rect 12492 6344 12537 6372
rect 12492 6332 12498 6344
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 2038 6304 2044 6316
rect 1636 6276 2044 6304
rect 1636 6264 1642 6276
rect 2038 6264 2044 6276
rect 2096 6304 2102 6316
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 2096 6276 2145 6304
rect 2096 6264 2102 6276
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 3142 6304 3148 6316
rect 3099 6276 3148 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3142 6264 3148 6276
rect 3200 6304 3206 6316
rect 3697 6307 3755 6313
rect 3697 6304 3709 6307
rect 3200 6276 3709 6304
rect 3200 6264 3206 6276
rect 3697 6273 3709 6276
rect 3743 6273 3755 6307
rect 3697 6267 3755 6273
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 4580 6276 5365 6304
rect 4580 6264 4586 6276
rect 5353 6273 5365 6276
rect 5399 6304 5411 6307
rect 6089 6307 6147 6313
rect 6089 6304 6101 6307
rect 5399 6276 6101 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 6089 6273 6101 6276
rect 6135 6273 6147 6307
rect 7282 6304 7288 6316
rect 7243 6276 7288 6304
rect 6089 6267 6147 6273
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 8481 6307 8539 6313
rect 8481 6273 8493 6307
rect 8527 6304 8539 6307
rect 12986 6304 12992 6316
rect 8527 6276 8708 6304
rect 12947 6276 12992 6304
rect 8527 6273 8539 6276
rect 8481 6267 8539 6273
rect 1946 6236 1952 6248
rect 1907 6208 1952 6236
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 2774 6236 2780 6248
rect 2455 6208 2780 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 3513 6239 3571 6245
rect 3513 6236 3525 6239
rect 3292 6208 3525 6236
rect 3292 6196 3298 6208
rect 3513 6205 3525 6208
rect 3559 6205 3571 6239
rect 3513 6199 3571 6205
rect 4154 6196 4160 6248
rect 4212 6236 4218 6248
rect 4430 6236 4436 6248
rect 4212 6208 4436 6236
rect 4212 6196 4218 6208
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 4614 6196 4620 6248
rect 4672 6236 4678 6248
rect 5077 6239 5135 6245
rect 5077 6236 5089 6239
rect 4672 6208 5089 6236
rect 4672 6196 4678 6208
rect 5077 6205 5089 6208
rect 5123 6205 5135 6239
rect 5077 6199 5135 6205
rect 5994 6196 6000 6248
rect 6052 6236 6058 6248
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 6052 6208 7205 6236
rect 6052 6196 6058 6208
rect 7193 6205 7205 6208
rect 7239 6205 7251 6239
rect 8570 6236 8576 6248
rect 8531 6208 8576 6236
rect 7193 6199 7251 6205
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 8680 6236 8708 6276
rect 12986 6264 12992 6276
rect 13044 6304 13050 6316
rect 13449 6307 13507 6313
rect 13449 6304 13461 6307
rect 13044 6276 13461 6304
rect 13044 6264 13050 6276
rect 13449 6273 13461 6276
rect 13495 6273 13507 6307
rect 13449 6267 13507 6273
rect 8846 6245 8852 6248
rect 8840 6236 8852 6245
rect 8680 6208 8852 6236
rect 8840 6199 8852 6208
rect 8904 6236 8910 6248
rect 9950 6236 9956 6248
rect 8904 6208 9956 6236
rect 8846 6196 8852 6199
rect 8904 6196 8910 6208
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 14200 6236 14228 6403
rect 16022 6400 16028 6452
rect 16080 6440 16086 6452
rect 16666 6440 16672 6452
rect 16080 6412 16672 6440
rect 16080 6400 16086 6412
rect 16666 6400 16672 6412
rect 16724 6400 16730 6452
rect 19058 6440 19064 6452
rect 19019 6412 19064 6440
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 20898 6440 20904 6452
rect 20859 6412 20904 6440
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 16298 6372 16304 6384
rect 16259 6344 16304 6372
rect 16298 6332 16304 6344
rect 16356 6332 16362 6384
rect 17037 6375 17095 6381
rect 17037 6341 17049 6375
rect 17083 6372 17095 6375
rect 18138 6372 18144 6384
rect 17083 6344 18144 6372
rect 17083 6341 17095 6344
rect 17037 6335 17095 6341
rect 18138 6332 18144 6344
rect 18196 6332 18202 6384
rect 14366 6304 14372 6316
rect 14327 6276 14372 6304
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 18690 6304 18696 6316
rect 18603 6276 18696 6304
rect 18690 6264 18696 6276
rect 18748 6304 18754 6316
rect 19429 6307 19487 6313
rect 19429 6304 19441 6307
rect 18748 6276 19441 6304
rect 18748 6264 18754 6276
rect 19429 6273 19441 6276
rect 19475 6273 19487 6307
rect 19429 6267 19487 6273
rect 14642 6245 14648 6248
rect 14625 6239 14648 6245
rect 14625 6236 14637 6239
rect 14200 6208 14637 6236
rect 14625 6205 14637 6208
rect 14700 6236 14706 6248
rect 16850 6236 16856 6248
rect 14700 6208 14773 6236
rect 16811 6208 16856 6236
rect 14625 6199 14648 6205
rect 14642 6196 14648 6199
rect 14700 6196 14706 6208
rect 16850 6196 16856 6208
rect 16908 6196 16914 6248
rect 17770 6236 17776 6248
rect 17731 6208 17776 6236
rect 17770 6196 17776 6208
rect 17828 6236 17834 6248
rect 18509 6239 18567 6245
rect 18509 6236 18521 6239
rect 17828 6208 18521 6236
rect 17828 6196 17834 6208
rect 18509 6205 18521 6208
rect 18555 6205 18567 6239
rect 18509 6199 18567 6205
rect 3418 6168 3424 6180
rect 1596 6140 3424 6168
rect 1596 6109 1624 6140
rect 3418 6128 3424 6140
rect 3476 6168 3482 6180
rect 3605 6171 3663 6177
rect 3605 6168 3617 6171
rect 3476 6140 3617 6168
rect 3476 6128 3482 6140
rect 3605 6137 3617 6140
rect 3651 6137 3663 6171
rect 3605 6131 3663 6137
rect 4249 6171 4307 6177
rect 4249 6137 4261 6171
rect 4295 6168 4307 6171
rect 5350 6168 5356 6180
rect 4295 6140 5356 6168
rect 4295 6137 4307 6140
rect 4249 6131 4307 6137
rect 5350 6128 5356 6140
rect 5408 6128 5414 6180
rect 6641 6171 6699 6177
rect 6641 6137 6653 6171
rect 6687 6168 6699 6171
rect 7466 6168 7472 6180
rect 6687 6140 7472 6168
rect 6687 6137 6699 6140
rect 6641 6131 6699 6137
rect 7466 6128 7472 6140
rect 7524 6128 7530 6180
rect 12897 6171 12955 6177
rect 12897 6137 12909 6171
rect 12943 6168 12955 6171
rect 13078 6168 13084 6180
rect 12943 6140 13084 6168
rect 12943 6137 12955 6140
rect 12897 6131 12955 6137
rect 13078 6128 13084 6140
rect 13136 6168 13142 6180
rect 13817 6171 13875 6177
rect 13817 6168 13829 6171
rect 13136 6140 13829 6168
rect 13136 6128 13142 6140
rect 13817 6137 13829 6140
rect 13863 6137 13875 6171
rect 13817 6131 13875 6137
rect 17497 6171 17555 6177
rect 17497 6137 17509 6171
rect 17543 6168 17555 6171
rect 18417 6171 18475 6177
rect 18417 6168 18429 6171
rect 17543 6140 18429 6168
rect 17543 6137 17555 6140
rect 17497 6131 17555 6137
rect 18417 6137 18429 6140
rect 18463 6168 18475 6171
rect 19613 6171 19671 6177
rect 19613 6168 19625 6171
rect 18463 6140 19625 6168
rect 18463 6137 18475 6140
rect 18417 6131 18475 6137
rect 19613 6137 19625 6140
rect 19659 6137 19671 6171
rect 19613 6131 19671 6137
rect 1581 6103 1639 6109
rect 1581 6069 1593 6103
rect 1627 6069 1639 6103
rect 1581 6063 1639 6069
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 2041 6103 2099 6109
rect 2041 6100 2053 6103
rect 1728 6072 2053 6100
rect 1728 6060 1734 6072
rect 2041 6069 2053 6072
rect 2087 6100 2099 6103
rect 2409 6103 2467 6109
rect 2409 6100 2421 6103
rect 2087 6072 2421 6100
rect 2087 6069 2099 6072
rect 2041 6063 2099 6069
rect 2409 6069 2421 6072
rect 2455 6069 2467 6103
rect 2409 6063 2467 6069
rect 3145 6103 3203 6109
rect 3145 6069 3157 6103
rect 3191 6100 3203 6103
rect 3510 6100 3516 6112
rect 3191 6072 3516 6100
rect 3191 6069 3203 6072
rect 3145 6063 3203 6069
rect 3510 6060 3516 6072
rect 3568 6060 3574 6112
rect 4430 6060 4436 6112
rect 4488 6100 4494 6112
rect 4525 6103 4583 6109
rect 4525 6100 4537 6103
rect 4488 6072 4537 6100
rect 4488 6060 4494 6072
rect 4525 6069 4537 6072
rect 4571 6100 4583 6103
rect 5169 6103 5227 6109
rect 5169 6100 5181 6103
rect 4571 6072 5181 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 5169 6069 5181 6072
rect 5215 6069 5227 6103
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 5169 6063 5227 6069
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 9953 6103 10011 6109
rect 9953 6100 9965 6103
rect 9916 6072 9965 6100
rect 9916 6060 9922 6072
rect 9953 6069 9965 6072
rect 9999 6069 10011 6103
rect 11330 6100 11336 6112
rect 11291 6072 11336 6100
rect 9953 6063 10011 6069
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 12158 6100 12164 6112
rect 12119 6072 12164 6100
rect 12158 6060 12164 6072
rect 12216 6100 12222 6112
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 12216 6072 12817 6100
rect 12216 6060 12222 6072
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 12805 6063 12863 6069
rect 15749 6103 15807 6109
rect 15749 6069 15761 6103
rect 15795 6100 15807 6103
rect 15838 6100 15844 6112
rect 15795 6072 15844 6100
rect 15795 6069 15807 6072
rect 15749 6063 15807 6069
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 18046 6100 18052 6112
rect 18007 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1946 5856 1952 5908
rect 2004 5896 2010 5908
rect 2133 5899 2191 5905
rect 2133 5896 2145 5899
rect 2004 5868 2145 5896
rect 2004 5856 2010 5868
rect 2133 5865 2145 5868
rect 2179 5865 2191 5899
rect 3142 5896 3148 5908
rect 3103 5868 3148 5896
rect 2133 5859 2191 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 4525 5899 4583 5905
rect 4525 5865 4537 5899
rect 4571 5896 4583 5899
rect 5166 5896 5172 5908
rect 4571 5868 5172 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 5166 5856 5172 5868
rect 5224 5896 5230 5908
rect 5997 5899 6055 5905
rect 5997 5896 6009 5899
rect 5224 5868 6009 5896
rect 5224 5856 5230 5868
rect 5997 5865 6009 5868
rect 6043 5896 6055 5899
rect 6549 5899 6607 5905
rect 6549 5896 6561 5899
rect 6043 5868 6561 5896
rect 6043 5865 6055 5868
rect 5997 5859 6055 5865
rect 6549 5865 6561 5868
rect 6595 5896 6607 5899
rect 6730 5896 6736 5908
rect 6595 5868 6736 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7009 5899 7067 5905
rect 7009 5865 7021 5899
rect 7055 5896 7067 5899
rect 7282 5896 7288 5908
rect 7055 5868 7288 5896
rect 7055 5865 7067 5868
rect 7009 5859 7067 5865
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 9950 5896 9956 5908
rect 9911 5868 9956 5896
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 10321 5899 10379 5905
rect 10321 5865 10333 5899
rect 10367 5896 10379 5899
rect 10962 5896 10968 5908
rect 10367 5868 10968 5896
rect 10367 5865 10379 5868
rect 10321 5859 10379 5865
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 11790 5896 11796 5908
rect 11751 5868 11796 5896
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 14366 5896 14372 5908
rect 14327 5868 14372 5896
rect 14366 5856 14372 5868
rect 14424 5856 14430 5908
rect 14826 5856 14832 5908
rect 14884 5896 14890 5908
rect 15286 5896 15292 5908
rect 14884 5868 15292 5896
rect 14884 5856 14890 5868
rect 15286 5856 15292 5868
rect 15344 5896 15350 5908
rect 15657 5899 15715 5905
rect 15657 5896 15669 5899
rect 15344 5868 15669 5896
rect 15344 5856 15350 5868
rect 15657 5865 15669 5868
rect 15703 5865 15715 5899
rect 15657 5859 15715 5865
rect 15746 5856 15752 5908
rect 15804 5896 15810 5908
rect 16298 5896 16304 5908
rect 15804 5868 15849 5896
rect 16259 5868 16304 5896
rect 15804 5856 15810 5868
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 18877 5899 18935 5905
rect 18877 5865 18889 5899
rect 18923 5896 18935 5899
rect 19058 5896 19064 5908
rect 18923 5868 19064 5896
rect 18923 5865 18935 5868
rect 18877 5859 18935 5865
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 2501 5831 2559 5837
rect 2501 5797 2513 5831
rect 2547 5828 2559 5831
rect 2590 5828 2596 5840
rect 2547 5800 2596 5828
rect 2547 5797 2559 5800
rect 2501 5791 2559 5797
rect 2590 5788 2596 5800
rect 2648 5788 2654 5840
rect 2682 5788 2688 5840
rect 2740 5828 2746 5840
rect 3513 5831 3571 5837
rect 3513 5828 3525 5831
rect 2740 5800 3525 5828
rect 2740 5788 2746 5800
rect 3513 5797 3525 5800
rect 3559 5797 3571 5831
rect 7098 5828 7104 5840
rect 3513 5791 3571 5797
rect 4632 5800 7104 5828
rect 4632 5769 4660 5800
rect 7098 5788 7104 5800
rect 7156 5788 7162 5840
rect 7368 5831 7426 5837
rect 7368 5797 7380 5831
rect 7414 5828 7426 5831
rect 7466 5828 7472 5840
rect 7414 5800 7472 5828
rect 7414 5797 7426 5800
rect 7368 5791 7426 5797
rect 7466 5788 7472 5800
rect 7524 5788 7530 5840
rect 14458 5788 14464 5840
rect 14516 5828 14522 5840
rect 15013 5831 15071 5837
rect 15013 5828 15025 5831
rect 14516 5800 15025 5828
rect 14516 5788 14522 5800
rect 15013 5797 15025 5800
rect 15059 5797 15071 5831
rect 15013 5791 15071 5797
rect 17494 5788 17500 5840
rect 17552 5828 17558 5840
rect 17764 5831 17822 5837
rect 17764 5828 17776 5831
rect 17552 5800 17776 5828
rect 17552 5788 17558 5800
rect 17764 5797 17776 5800
rect 17810 5828 17822 5831
rect 18690 5828 18696 5840
rect 17810 5800 18696 5828
rect 17810 5797 17822 5800
rect 17764 5791 17822 5797
rect 18690 5788 18696 5800
rect 18748 5788 18754 5840
rect 4890 5769 4896 5772
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5729 4675 5763
rect 4884 5760 4896 5769
rect 4851 5732 4896 5760
rect 4617 5723 4675 5729
rect 4884 5723 4896 5732
rect 4890 5720 4896 5723
rect 4948 5720 4954 5772
rect 10686 5760 10692 5772
rect 10647 5732 10692 5760
rect 10686 5720 10692 5732
rect 10744 5760 10750 5772
rect 10962 5760 10968 5772
rect 10744 5732 10968 5760
rect 10744 5720 10750 5732
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 12141 5763 12199 5769
rect 12141 5760 12153 5763
rect 11716 5732 12153 5760
rect 2406 5652 2412 5704
rect 2464 5692 2470 5704
rect 2593 5695 2651 5701
rect 2593 5692 2605 5695
rect 2464 5664 2605 5692
rect 2464 5652 2470 5664
rect 2593 5661 2605 5664
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5661 2743 5695
rect 7098 5692 7104 5704
rect 7059 5664 7104 5692
rect 2685 5655 2743 5661
rect 2041 5627 2099 5633
rect 2041 5593 2053 5627
rect 2087 5624 2099 5627
rect 2222 5624 2228 5636
rect 2087 5596 2228 5624
rect 2087 5593 2099 5596
rect 2041 5587 2099 5593
rect 2222 5584 2228 5596
rect 2280 5624 2286 5636
rect 2700 5624 2728 5655
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 9950 5652 9956 5704
rect 10008 5692 10014 5704
rect 10781 5695 10839 5701
rect 10781 5692 10793 5695
rect 10008 5664 10793 5692
rect 10008 5652 10014 5664
rect 10781 5661 10793 5664
rect 10827 5661 10839 5695
rect 10781 5655 10839 5661
rect 10873 5695 10931 5701
rect 10873 5661 10885 5695
rect 10919 5661 10931 5695
rect 10873 5655 10931 5661
rect 2280 5596 2728 5624
rect 8481 5627 8539 5633
rect 2280 5584 2286 5596
rect 8481 5593 8493 5627
rect 8527 5624 8539 5627
rect 10888 5624 10916 5655
rect 11716 5636 11744 5732
rect 12141 5729 12153 5732
rect 12187 5729 12199 5763
rect 20898 5760 20904 5772
rect 20859 5732 20904 5760
rect 12141 5723 12199 5729
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 11882 5692 11888 5704
rect 11843 5664 11888 5692
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 13906 5692 13912 5704
rect 13867 5664 13912 5692
rect 13906 5652 13912 5664
rect 13964 5652 13970 5704
rect 15838 5652 15844 5704
rect 15896 5692 15902 5704
rect 16482 5692 16488 5704
rect 15896 5664 16488 5692
rect 15896 5652 15902 5664
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 17497 5695 17555 5701
rect 17497 5692 17509 5695
rect 17236 5664 17509 5692
rect 11698 5624 11704 5636
rect 8527 5596 11704 5624
rect 8527 5593 8539 5596
rect 8481 5587 8539 5593
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 15289 5627 15347 5633
rect 15289 5593 15301 5627
rect 15335 5624 15347 5627
rect 15930 5624 15936 5636
rect 15335 5596 15936 5624
rect 15335 5593 15347 5596
rect 15289 5587 15347 5593
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 16850 5624 16856 5636
rect 16811 5596 16856 5624
rect 16850 5584 16856 5596
rect 16908 5584 16914 5636
rect 17236 5568 17264 5664
rect 17497 5661 17509 5664
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 9125 5559 9183 5565
rect 9125 5525 9137 5559
rect 9171 5556 9183 5559
rect 9306 5556 9312 5568
rect 9171 5528 9312 5556
rect 9171 5525 9183 5528
rect 9125 5519 9183 5525
rect 9306 5516 9312 5528
rect 9364 5556 9370 5568
rect 9401 5559 9459 5565
rect 9401 5556 9413 5559
rect 9364 5528 9413 5556
rect 9364 5516 9370 5528
rect 9401 5525 9413 5528
rect 9447 5525 9459 5559
rect 9401 5519 9459 5525
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 11204 5528 11345 5556
rect 11204 5516 11210 5528
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 11333 5519 11391 5525
rect 13265 5559 13323 5565
rect 13265 5525 13277 5559
rect 13311 5556 13323 5559
rect 13630 5556 13636 5568
rect 13311 5528 13636 5556
rect 13311 5525 13323 5528
rect 13265 5519 13323 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 17218 5556 17224 5568
rect 17179 5528 17224 5556
rect 17218 5516 17224 5528
rect 17276 5516 17282 5568
rect 21082 5556 21088 5568
rect 21043 5528 21088 5556
rect 21082 5516 21088 5528
rect 21140 5516 21146 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 4522 5352 4528 5364
rect 4295 5324 4528 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 7466 5352 7472 5364
rect 7427 5324 7472 5352
rect 7466 5312 7472 5324
rect 7524 5312 7530 5364
rect 10778 5312 10784 5364
rect 10836 5352 10842 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10836 5324 10885 5352
rect 10836 5312 10842 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 11425 5355 11483 5361
rect 11425 5352 11437 5355
rect 11112 5324 11437 5352
rect 11112 5312 11118 5324
rect 11425 5321 11437 5324
rect 11471 5321 11483 5355
rect 11425 5315 11483 5321
rect 11698 5312 11704 5364
rect 11756 5352 11762 5364
rect 11793 5355 11851 5361
rect 11793 5352 11805 5355
rect 11756 5324 11805 5352
rect 11756 5312 11762 5324
rect 11793 5321 11805 5324
rect 11839 5352 11851 5355
rect 12621 5355 12679 5361
rect 12621 5352 12633 5355
rect 11839 5324 12633 5352
rect 11839 5321 11851 5324
rect 11793 5315 11851 5321
rect 12621 5321 12633 5324
rect 12667 5321 12679 5355
rect 12621 5315 12679 5321
rect 14642 5312 14648 5364
rect 14700 5352 14706 5364
rect 14737 5355 14795 5361
rect 14737 5352 14749 5355
rect 14700 5324 14749 5352
rect 14700 5312 14706 5324
rect 14737 5321 14749 5324
rect 14783 5321 14795 5355
rect 15286 5352 15292 5364
rect 15247 5324 15292 5352
rect 14737 5315 14795 5321
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 16482 5312 16488 5364
rect 16540 5352 16546 5364
rect 16853 5355 16911 5361
rect 16853 5352 16865 5355
rect 16540 5324 16865 5352
rect 16540 5312 16546 5324
rect 16853 5321 16865 5324
rect 16899 5321 16911 5355
rect 17494 5352 17500 5364
rect 17455 5324 17500 5352
rect 16853 5315 16911 5321
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 17865 5355 17923 5361
rect 17865 5321 17877 5355
rect 17911 5352 17923 5355
rect 20898 5352 20904 5364
rect 17911 5324 18736 5352
rect 17911 5321 17923 5324
rect 17865 5315 17923 5321
rect 9033 5287 9091 5293
rect 9033 5284 9045 5287
rect 8404 5256 9045 5284
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5216 1455 5219
rect 1762 5216 1768 5228
rect 1443 5188 1768 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 5350 5176 5356 5228
rect 5408 5216 5414 5228
rect 8404 5225 8432 5256
rect 9033 5253 9045 5256
rect 9079 5284 9091 5287
rect 9490 5284 9496 5296
rect 9079 5256 9496 5284
rect 9079 5253 9091 5256
rect 9033 5247 9091 5253
rect 9490 5244 9496 5256
rect 9548 5244 9554 5296
rect 18049 5287 18107 5293
rect 18049 5253 18061 5287
rect 18095 5253 18107 5287
rect 18049 5247 18107 5253
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5408 5188 5733 5216
rect 5408 5176 5414 5188
rect 5721 5185 5733 5188
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5185 8539 5219
rect 15654 5216 15660 5228
rect 15615 5188 15660 5216
rect 8481 5179 8539 5185
rect 1486 5108 1492 5160
rect 1544 5148 1550 5160
rect 3142 5157 3148 5160
rect 2869 5151 2927 5157
rect 2869 5148 2881 5151
rect 1544 5120 2881 5148
rect 1544 5108 1550 5120
rect 2869 5117 2881 5120
rect 2915 5117 2927 5151
rect 3136 5148 3148 5157
rect 3103 5120 3148 5148
rect 2869 5111 2927 5117
rect 3136 5111 3148 5120
rect 2884 5080 2912 5111
rect 3142 5108 3148 5111
rect 3200 5108 3206 5160
rect 4890 5148 4896 5160
rect 4803 5120 4896 5148
rect 4890 5108 4896 5120
rect 4948 5148 4954 5160
rect 6178 5148 6184 5160
rect 4948 5120 6184 5148
rect 4948 5108 4954 5120
rect 6178 5108 6184 5120
rect 6236 5108 6242 5160
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5148 7895 5151
rect 8202 5148 8208 5160
rect 7883 5120 8208 5148
rect 7883 5117 7895 5120
rect 7837 5111 7895 5117
rect 8202 5108 8208 5120
rect 8260 5148 8266 5160
rect 8496 5148 8524 5179
rect 15654 5176 15660 5188
rect 15712 5216 15718 5228
rect 16390 5216 16396 5228
rect 15712 5188 16252 5216
rect 16351 5188 16396 5216
rect 15712 5176 15718 5188
rect 8260 5120 8524 5148
rect 8260 5108 8266 5120
rect 9306 5108 9312 5160
rect 9364 5148 9370 5160
rect 9493 5151 9551 5157
rect 9493 5148 9505 5151
rect 9364 5120 9505 5148
rect 9364 5108 9370 5120
rect 9493 5117 9505 5120
rect 9539 5117 9551 5151
rect 9493 5111 9551 5117
rect 11790 5108 11796 5160
rect 11848 5148 11854 5160
rect 12161 5151 12219 5157
rect 12161 5148 12173 5151
rect 11848 5120 12173 5148
rect 11848 5108 11854 5120
rect 12161 5117 12173 5120
rect 12207 5117 12219 5151
rect 12161 5111 12219 5117
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 16224 5157 16252 5188
rect 16390 5176 16396 5188
rect 16448 5176 16454 5228
rect 13357 5151 13415 5157
rect 13357 5148 13369 5151
rect 12492 5120 13369 5148
rect 12492 5108 12498 5120
rect 13357 5117 13369 5120
rect 13403 5148 13415 5151
rect 16209 5151 16267 5157
rect 13403 5120 13768 5148
rect 13403 5117 13415 5120
rect 13357 5111 13415 5117
rect 13740 5092 13768 5120
rect 16209 5117 16221 5151
rect 16255 5117 16267 5151
rect 16209 5111 16267 5117
rect 16298 5108 16304 5160
rect 16356 5148 16362 5160
rect 18064 5148 18092 5247
rect 18708 5225 18736 5324
rect 20088 5324 20904 5352
rect 18693 5219 18751 5225
rect 18693 5185 18705 5219
rect 18739 5216 18751 5219
rect 19058 5216 19064 5228
rect 18739 5188 19064 5216
rect 18739 5185 18751 5188
rect 18693 5179 18751 5185
rect 19058 5176 19064 5188
rect 19116 5176 19122 5228
rect 20088 5225 20116 5324
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 20073 5219 20131 5225
rect 20073 5185 20085 5219
rect 20119 5185 20131 5219
rect 20073 5179 20131 5185
rect 19797 5151 19855 5157
rect 19797 5148 19809 5151
rect 16356 5120 16401 5148
rect 18064 5120 19809 5148
rect 16356 5108 16362 5120
rect 19797 5117 19809 5120
rect 19843 5148 19855 5151
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 19843 5120 20545 5148
rect 19843 5117 19855 5120
rect 19797 5111 19855 5117
rect 20533 5117 20545 5120
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 21085 5151 21143 5157
rect 21085 5117 21097 5151
rect 21131 5148 21143 5151
rect 21131 5120 21680 5148
rect 21131 5117 21143 5120
rect 21085 5111 21143 5117
rect 5169 5083 5227 5089
rect 5169 5080 5181 5083
rect 2884 5052 5181 5080
rect 5169 5049 5181 5052
rect 5215 5080 5227 5083
rect 5350 5080 5356 5092
rect 5215 5052 5356 5080
rect 5215 5049 5227 5052
rect 5169 5043 5227 5049
rect 5350 5040 5356 5052
rect 5408 5080 5414 5092
rect 5537 5083 5595 5089
rect 5537 5080 5549 5083
rect 5408 5052 5549 5080
rect 5408 5040 5414 5052
rect 5537 5049 5549 5052
rect 5583 5080 5595 5083
rect 6273 5083 6331 5089
rect 6273 5080 6285 5083
rect 5583 5052 6285 5080
rect 5583 5049 5595 5052
rect 5537 5043 5595 5049
rect 6273 5049 6285 5052
rect 6319 5080 6331 5083
rect 6549 5083 6607 5089
rect 6549 5080 6561 5083
rect 6319 5052 6561 5080
rect 6319 5049 6331 5052
rect 6273 5043 6331 5049
rect 6549 5049 6561 5052
rect 6595 5080 6607 5083
rect 7282 5080 7288 5092
rect 6595 5052 7288 5080
rect 6595 5049 6607 5052
rect 6549 5043 6607 5049
rect 7282 5040 7288 5052
rect 7340 5040 7346 5092
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 8297 5083 8355 5089
rect 8297 5080 8309 5083
rect 7616 5052 8309 5080
rect 7616 5040 7622 5052
rect 8297 5049 8309 5052
rect 8343 5080 8355 5083
rect 9398 5080 9404 5092
rect 8343 5052 9404 5080
rect 8343 5049 8355 5052
rect 8297 5043 8355 5049
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 9760 5083 9818 5089
rect 9760 5080 9772 5083
rect 9692 5052 9772 5080
rect 2225 5015 2283 5021
rect 2225 4981 2237 5015
rect 2271 5012 2283 5015
rect 2406 5012 2412 5024
rect 2271 4984 2412 5012
rect 2271 4981 2283 4984
rect 2225 4975 2283 4981
rect 2406 4972 2412 4984
rect 2464 4972 2470 5024
rect 2590 5012 2596 5024
rect 2551 4984 2596 5012
rect 2590 4972 2596 4984
rect 2648 4972 2654 5024
rect 6917 5015 6975 5021
rect 6917 4981 6929 5015
rect 6963 5012 6975 5015
rect 7466 5012 7472 5024
rect 6963 4984 7472 5012
rect 6963 4981 6975 4984
rect 6917 4975 6975 4981
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 7926 5012 7932 5024
rect 7887 4984 7932 5012
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 9309 5015 9367 5021
rect 9309 4981 9321 5015
rect 9355 5012 9367 5015
rect 9692 5012 9720 5052
rect 9760 5049 9772 5052
rect 9806 5080 9818 5083
rect 9858 5080 9864 5092
rect 9806 5052 9864 5080
rect 9806 5049 9818 5052
rect 9760 5043 9818 5049
rect 9858 5040 9864 5052
rect 9916 5080 9922 5092
rect 10686 5080 10692 5092
rect 9916 5052 10692 5080
rect 9916 5040 9922 5052
rect 10686 5040 10692 5052
rect 10744 5040 10750 5092
rect 13630 5089 13636 5092
rect 13265 5083 13323 5089
rect 13265 5049 13277 5083
rect 13311 5080 13323 5083
rect 13624 5080 13636 5089
rect 13311 5052 13636 5080
rect 13311 5049 13323 5052
rect 13265 5043 13323 5049
rect 13624 5043 13636 5052
rect 13630 5040 13636 5043
rect 13688 5040 13694 5092
rect 13722 5040 13728 5092
rect 13780 5040 13786 5092
rect 18046 5040 18052 5092
rect 18104 5080 18110 5092
rect 18417 5083 18475 5089
rect 18417 5080 18429 5083
rect 18104 5052 18429 5080
rect 18104 5040 18110 5052
rect 18417 5049 18429 5052
rect 18463 5080 18475 5083
rect 19429 5083 19487 5089
rect 19429 5080 19441 5083
rect 18463 5052 19441 5080
rect 18463 5049 18475 5052
rect 18417 5043 18475 5049
rect 19429 5049 19441 5052
rect 19475 5049 19487 5083
rect 19429 5043 19487 5049
rect 21652 5024 21680 5120
rect 9355 4984 9720 5012
rect 9355 4981 9367 4984
rect 9309 4975 9367 4981
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 11977 5015 12035 5021
rect 11977 5012 11989 5015
rect 11940 4984 11989 5012
rect 11940 4972 11946 4984
rect 11977 4981 11989 4984
rect 12023 4981 12035 5015
rect 11977 4975 12035 4981
rect 14826 4972 14832 5024
rect 14884 5012 14890 5024
rect 15841 5015 15899 5021
rect 15841 5012 15853 5015
rect 14884 4984 15853 5012
rect 14884 4972 14890 4984
rect 15841 4981 15853 4984
rect 15887 4981 15899 5015
rect 15841 4975 15899 4981
rect 18506 4972 18512 5024
rect 18564 5012 18570 5024
rect 19061 5015 19119 5021
rect 19061 5012 19073 5015
rect 18564 4984 19073 5012
rect 18564 4972 18570 4984
rect 19061 4981 19073 4984
rect 19107 4981 19119 5015
rect 19061 4975 19119 4981
rect 21269 5015 21327 5021
rect 21269 4981 21281 5015
rect 21315 5012 21327 5015
rect 21542 5012 21548 5024
rect 21315 4984 21548 5012
rect 21315 4981 21327 4984
rect 21269 4975 21327 4981
rect 21542 4972 21548 4984
rect 21600 4972 21606 5024
rect 21634 4972 21640 5024
rect 21692 5012 21698 5024
rect 21692 4984 21737 5012
rect 21692 4972 21698 4984
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 3142 4808 3148 4820
rect 2915 4780 3148 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 3418 4808 3424 4820
rect 3379 4780 3424 4808
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 3602 4768 3608 4820
rect 3660 4808 3666 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3660 4780 3801 4808
rect 3660 4768 3666 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4808 5871 4811
rect 6086 4808 6092 4820
rect 5859 4780 6092 4808
rect 5859 4777 5871 4780
rect 5813 4771 5871 4777
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 7558 4808 7564 4820
rect 7519 4780 7564 4808
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 8294 4808 8300 4820
rect 8255 4780 8300 4808
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 12618 4808 12624 4820
rect 12579 4780 12624 4808
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 13078 4808 13084 4820
rect 13039 4780 13084 4808
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 14734 4768 14740 4820
rect 14792 4808 14798 4820
rect 15013 4811 15071 4817
rect 15013 4808 15025 4811
rect 14792 4780 15025 4808
rect 14792 4768 14798 4780
rect 15013 4777 15025 4780
rect 15059 4777 15071 4811
rect 15746 4808 15752 4820
rect 15707 4780 15752 4808
rect 15013 4771 15071 4777
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 16390 4808 16396 4820
rect 16351 4780 16396 4808
rect 16390 4768 16396 4780
rect 16448 4768 16454 4820
rect 18417 4811 18475 4817
rect 18417 4777 18429 4811
rect 18463 4808 18475 4811
rect 18690 4808 18696 4820
rect 18463 4780 18696 4808
rect 18463 4777 18475 4780
rect 18417 4771 18475 4777
rect 18690 4768 18696 4780
rect 18748 4768 18754 4820
rect 10778 4700 10784 4752
rect 10836 4749 10842 4752
rect 10836 4743 10900 4749
rect 10836 4709 10854 4743
rect 10888 4709 10900 4743
rect 10836 4703 10900 4709
rect 10836 4700 10842 4703
rect 10962 4700 10968 4752
rect 11020 4700 11026 4752
rect 12989 4743 13047 4749
rect 12989 4709 13001 4743
rect 13035 4740 13047 4743
rect 13722 4740 13728 4752
rect 13035 4712 13728 4740
rect 13035 4709 13047 4712
rect 12989 4703 13047 4709
rect 13722 4700 13728 4712
rect 13780 4700 13786 4752
rect 24210 4749 24216 4752
rect 24204 4740 24216 4749
rect 24171 4712 24216 4740
rect 24204 4703 24216 4712
rect 24210 4700 24216 4703
rect 24268 4700 24274 4752
rect 1578 4632 1584 4684
rect 1636 4672 1642 4684
rect 1756 4675 1814 4681
rect 1756 4672 1768 4675
rect 1636 4644 1768 4672
rect 1636 4632 1642 4644
rect 1756 4641 1768 4644
rect 1802 4672 1814 4675
rect 2590 4672 2596 4684
rect 1802 4644 2596 4672
rect 1802 4641 1814 4644
rect 1756 4635 1814 4641
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 4614 4672 4620 4684
rect 4575 4644 4620 4672
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 4709 4675 4767 4681
rect 4709 4641 4721 4675
rect 4755 4672 4767 4675
rect 4890 4672 4896 4684
rect 4755 4644 4896 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 6086 4632 6092 4684
rect 6144 4672 6150 4684
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 6144 4644 6193 4672
rect 6144 4632 6150 4644
rect 6181 4641 6193 4644
rect 6227 4672 6239 4675
rect 6454 4672 6460 4684
rect 6227 4644 6460 4672
rect 6227 4641 6239 4644
rect 6181 4635 6239 4641
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 7193 4675 7251 4681
rect 7193 4641 7205 4675
rect 7239 4672 7251 4675
rect 7834 4672 7840 4684
rect 7239 4644 7840 4672
rect 7239 4641 7251 4644
rect 7193 4635 7251 4641
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 7944 4644 8953 4672
rect 1486 4604 1492 4616
rect 1447 4576 1492 4604
rect 1486 4564 1492 4576
rect 1544 4564 1550 4616
rect 4798 4604 4804 4616
rect 4759 4576 4804 4604
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 6270 4604 6276 4616
rect 6231 4576 6276 4604
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 7944 4604 7972 4644
rect 8941 4641 8953 4644
rect 8987 4672 8999 4675
rect 9306 4672 9312 4684
rect 8987 4644 9312 4672
rect 8987 4641 8999 4644
rect 8941 4635 8999 4641
rect 9306 4632 9312 4644
rect 9364 4672 9370 4684
rect 10597 4675 10655 4681
rect 10597 4672 10609 4675
rect 9364 4644 10609 4672
rect 9364 4632 9370 4644
rect 10597 4641 10609 4644
rect 10643 4672 10655 4675
rect 10980 4672 11008 4700
rect 10643 4644 11008 4672
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 13262 4632 13268 4684
rect 13320 4672 13326 4684
rect 13449 4675 13507 4681
rect 13449 4672 13461 4675
rect 13320 4644 13461 4672
rect 13320 4632 13326 4644
rect 13449 4641 13461 4644
rect 13495 4641 13507 4675
rect 14090 4672 14096 4684
rect 14051 4644 14096 4672
rect 13449 4635 13507 4641
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 15654 4672 15660 4684
rect 15615 4644 15660 4672
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 17126 4632 17132 4684
rect 17184 4672 17190 4684
rect 17293 4675 17351 4681
rect 17293 4672 17305 4675
rect 17184 4644 17305 4672
rect 17184 4632 17190 4644
rect 17293 4641 17305 4644
rect 17339 4641 17351 4675
rect 17293 4635 17351 4641
rect 19426 4632 19432 4684
rect 19484 4672 19490 4684
rect 19521 4675 19579 4681
rect 19521 4672 19533 4675
rect 19484 4644 19533 4672
rect 19484 4632 19490 4644
rect 19521 4641 19533 4644
rect 19567 4641 19579 4675
rect 20898 4672 20904 4684
rect 20859 4644 20904 4672
rect 19521 4635 19579 4641
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 21174 4632 21180 4684
rect 21232 4672 21238 4684
rect 21818 4672 21824 4684
rect 21232 4644 21824 4672
rect 21232 4632 21238 4644
rect 21818 4632 21824 4644
rect 21876 4672 21882 4684
rect 22005 4675 22063 4681
rect 22005 4672 22017 4675
rect 21876 4644 22017 4672
rect 21876 4632 21882 4644
rect 22005 4641 22017 4644
rect 22051 4641 22063 4675
rect 22005 4635 22063 4641
rect 6365 4567 6423 4573
rect 7668 4576 7972 4604
rect 4430 4496 4436 4548
rect 4488 4536 4494 4548
rect 5994 4536 6000 4548
rect 4488 4508 6000 4536
rect 4488 4496 4494 4508
rect 5994 4496 6000 4508
rect 6052 4496 6058 4548
rect 6178 4496 6184 4548
rect 6236 4536 6242 4548
rect 6380 4536 6408 4567
rect 6236 4508 6408 4536
rect 6236 4496 6242 4508
rect 7282 4496 7288 4548
rect 7340 4536 7346 4548
rect 7668 4545 7696 4576
rect 8018 4564 8024 4616
rect 8076 4604 8082 4616
rect 8386 4604 8392 4616
rect 8076 4576 8392 4604
rect 8076 4564 8082 4576
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 8570 4604 8576 4616
rect 8531 4576 8576 4604
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 13412 4576 13553 4604
rect 13412 4564 13418 4576
rect 13541 4573 13553 4576
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 13630 4564 13636 4616
rect 13688 4604 13694 4616
rect 13688 4576 13733 4604
rect 13688 4564 13694 4576
rect 15838 4564 15844 4616
rect 15896 4604 15902 4616
rect 17037 4607 17095 4613
rect 15896 4576 15941 4604
rect 15896 4564 15902 4576
rect 17037 4573 17049 4607
rect 17083 4573 17095 4607
rect 17037 4567 17095 4573
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4604 19855 4607
rect 20622 4604 20628 4616
rect 19843 4576 20628 4604
rect 19843 4573 19855 4576
rect 19797 4567 19855 4573
rect 7653 4539 7711 4545
rect 7653 4536 7665 4539
rect 7340 4508 7665 4536
rect 7340 4496 7346 4508
rect 7653 4505 7665 4508
rect 7699 4505 7711 4539
rect 7653 4499 7711 4505
rect 7929 4539 7987 4545
rect 7929 4505 7941 4539
rect 7975 4536 7987 4539
rect 9953 4539 10011 4545
rect 9953 4536 9965 4539
rect 7975 4508 9965 4536
rect 7975 4505 7987 4508
rect 7929 4499 7987 4505
rect 9953 4505 9965 4508
rect 9999 4536 10011 4539
rect 10502 4536 10508 4548
rect 9999 4508 10508 4536
rect 9999 4505 10011 4508
rect 9953 4499 10011 4505
rect 10502 4496 10508 4508
rect 10560 4496 10566 4548
rect 4246 4468 4252 4480
rect 4207 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 5074 4428 5080 4480
rect 5132 4468 5138 4480
rect 5261 4471 5319 4477
rect 5261 4468 5273 4471
rect 5132 4440 5273 4468
rect 5132 4428 5138 4440
rect 5261 4437 5273 4440
rect 5307 4437 5319 4471
rect 5261 4431 5319 4437
rect 5350 4428 5356 4480
rect 5408 4468 5414 4480
rect 5629 4471 5687 4477
rect 5629 4468 5641 4471
rect 5408 4440 5641 4468
rect 5408 4428 5414 4440
rect 5629 4437 5641 4440
rect 5675 4437 5687 4471
rect 5629 4431 5687 4437
rect 10042 4428 10048 4480
rect 10100 4468 10106 4480
rect 10413 4471 10471 4477
rect 10413 4468 10425 4471
rect 10100 4440 10425 4468
rect 10100 4428 10106 4440
rect 10413 4437 10425 4440
rect 10459 4468 10471 4471
rect 10962 4468 10968 4480
rect 10459 4440 10968 4468
rect 10459 4437 10471 4440
rect 10413 4431 10471 4437
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11698 4428 11704 4480
rect 11756 4468 11762 4480
rect 11977 4471 12035 4477
rect 11977 4468 11989 4471
rect 11756 4440 11989 4468
rect 11756 4428 11762 4440
rect 11977 4437 11989 4440
rect 12023 4437 12035 4471
rect 11977 4431 12035 4437
rect 14553 4471 14611 4477
rect 14553 4437 14565 4471
rect 14599 4468 14611 4471
rect 14642 4468 14648 4480
rect 14599 4440 14648 4468
rect 14599 4437 14611 4440
rect 14553 4431 14611 4437
rect 14642 4428 14648 4440
rect 14700 4428 14706 4480
rect 15286 4468 15292 4480
rect 15247 4440 15292 4468
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 16761 4471 16819 4477
rect 16761 4437 16773 4471
rect 16807 4468 16819 4471
rect 17052 4468 17080 4567
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 23934 4604 23940 4616
rect 23895 4576 23940 4604
rect 23934 4564 23940 4576
rect 23992 4564 23998 4616
rect 25314 4536 25320 4548
rect 25275 4508 25320 4536
rect 25314 4496 25320 4508
rect 25372 4496 25378 4548
rect 17218 4468 17224 4480
rect 16807 4440 17224 4468
rect 16807 4437 16819 4440
rect 16761 4431 16819 4437
rect 17218 4428 17224 4440
rect 17276 4468 17282 4480
rect 17678 4468 17684 4480
rect 17276 4440 17684 4468
rect 17276 4428 17282 4440
rect 17678 4428 17684 4440
rect 17736 4468 17742 4480
rect 19061 4471 19119 4477
rect 19061 4468 19073 4471
rect 17736 4440 19073 4468
rect 17736 4428 17742 4440
rect 19061 4437 19073 4440
rect 19107 4468 19119 4471
rect 19242 4468 19248 4480
rect 19107 4440 19248 4468
rect 19107 4437 19119 4440
rect 19061 4431 19119 4437
rect 19242 4428 19248 4440
rect 19300 4428 19306 4480
rect 20346 4428 20352 4480
rect 20404 4468 20410 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 20404 4440 21097 4468
rect 20404 4428 20410 4440
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 22189 4471 22247 4477
rect 22189 4437 22201 4471
rect 22235 4468 22247 4471
rect 23198 4468 23204 4480
rect 22235 4440 23204 4468
rect 22235 4437 22247 4440
rect 22189 4431 22247 4437
rect 23198 4428 23204 4440
rect 23256 4428 23262 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1670 4264 1676 4276
rect 1631 4236 1676 4264
rect 1670 4224 1676 4236
rect 1728 4224 1734 4276
rect 4154 4224 4160 4276
rect 4212 4264 4218 4276
rect 4249 4267 4307 4273
rect 4249 4264 4261 4267
rect 4212 4236 4261 4264
rect 4212 4224 4218 4236
rect 4249 4233 4261 4236
rect 4295 4264 4307 4267
rect 4798 4264 4804 4276
rect 4295 4236 4804 4264
rect 4295 4233 4307 4236
rect 4249 4227 4307 4233
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 6178 4224 6184 4276
rect 6236 4264 6242 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6236 4236 6561 4264
rect 6236 4224 6242 4236
rect 6549 4233 6561 4236
rect 6595 4264 6607 4267
rect 6730 4264 6736 4276
rect 6595 4236 6736 4264
rect 6595 4233 6607 4236
rect 6549 4227 6607 4233
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 10229 4267 10287 4273
rect 10229 4233 10241 4267
rect 10275 4264 10287 4267
rect 10778 4264 10784 4276
rect 10275 4236 10784 4264
rect 10275 4233 10287 4236
rect 10229 4227 10287 4233
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 13722 4264 13728 4276
rect 13004 4236 13728 4264
rect 4617 4199 4675 4205
rect 4617 4165 4629 4199
rect 4663 4196 4675 4199
rect 4663 4168 5304 4196
rect 4663 4165 4675 4168
rect 4617 4159 4675 4165
rect 5276 4140 5304 4168
rect 5994 4156 6000 4208
rect 6052 4196 6058 4208
rect 7929 4199 7987 4205
rect 7929 4196 7941 4199
rect 6052 4168 7941 4196
rect 6052 4156 6058 4168
rect 7929 4165 7941 4168
rect 7975 4196 7987 4199
rect 8018 4196 8024 4208
rect 7975 4168 8024 4196
rect 7975 4165 7987 4168
rect 7929 4159 7987 4165
rect 8018 4156 8024 4168
rect 8076 4156 8082 4208
rect 9398 4156 9404 4208
rect 9456 4196 9462 4208
rect 13004 4196 13032 4236
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 15654 4224 15660 4276
rect 15712 4264 15718 4276
rect 16393 4267 16451 4273
rect 16393 4264 16405 4267
rect 15712 4236 16405 4264
rect 15712 4224 15718 4236
rect 16393 4233 16405 4236
rect 16439 4233 16451 4267
rect 16393 4227 16451 4233
rect 18049 4267 18107 4273
rect 18049 4233 18061 4267
rect 18095 4264 18107 4267
rect 18506 4264 18512 4276
rect 18095 4236 18512 4264
rect 18095 4233 18107 4236
rect 18049 4227 18107 4233
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 18690 4224 18696 4276
rect 18748 4264 18754 4276
rect 19061 4267 19119 4273
rect 19061 4264 19073 4267
rect 18748 4236 19073 4264
rect 18748 4224 18754 4236
rect 19061 4233 19073 4236
rect 19107 4233 19119 4267
rect 19061 4227 19119 4233
rect 20809 4267 20867 4273
rect 20809 4233 20821 4267
rect 20855 4264 20867 4267
rect 20898 4264 20904 4276
rect 20855 4236 20904 4264
rect 20855 4233 20867 4236
rect 20809 4227 20867 4233
rect 9456 4168 9628 4196
rect 9456 4156 9462 4168
rect 2222 4128 2228 4140
rect 2183 4100 2228 4128
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2961 4131 3019 4137
rect 2961 4128 2973 4131
rect 2332 4100 2973 4128
rect 1394 4020 1400 4072
rect 1452 4060 1458 4072
rect 2041 4063 2099 4069
rect 2041 4060 2053 4063
rect 1452 4032 2053 4060
rect 1452 4020 1458 4032
rect 2041 4029 2053 4032
rect 2087 4060 2099 4063
rect 2332 4060 2360 4100
rect 2961 4097 2973 4100
rect 3007 4128 3019 4131
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 3007 4100 3065 4128
rect 3007 4097 3019 4100
rect 2961 4091 3019 4097
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4128 3295 4131
rect 3326 4128 3332 4140
rect 3283 4100 3332 4128
rect 3283 4097 3295 4100
rect 3237 4091 3295 4097
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 4246 4088 4252 4140
rect 4304 4128 4310 4140
rect 5166 4128 5172 4140
rect 4304 4100 5172 4128
rect 4304 4088 4310 4100
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 7006 4128 7012 4140
rect 5316 4100 5409 4128
rect 6967 4100 7012 4128
rect 5316 4088 5322 4100
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7282 4088 7288 4140
rect 7340 4128 7346 4140
rect 8205 4131 8263 4137
rect 8205 4128 8217 4131
rect 7340 4100 8217 4128
rect 7340 4088 7346 4100
rect 8205 4097 8217 4100
rect 8251 4097 8263 4131
rect 9600 4128 9628 4168
rect 12360 4168 13032 4196
rect 9600 4100 9720 4128
rect 8205 4091 8263 4097
rect 5813 4063 5871 4069
rect 5813 4060 5825 4063
rect 2087 4032 2360 4060
rect 2700 4032 5825 4060
rect 2087 4029 2099 4032
rect 2041 4023 2099 4029
rect 290 3952 296 4004
rect 348 3992 354 4004
rect 2700 4001 2728 4032
rect 5813 4029 5825 4032
rect 5859 4060 5871 4063
rect 6270 4060 6276 4072
rect 5859 4032 6276 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 9692 4060 9720 4100
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 11149 4131 11207 4137
rect 11149 4128 11161 4131
rect 10560 4100 11161 4128
rect 10560 4088 10566 4100
rect 11149 4097 11161 4100
rect 11195 4097 11207 4131
rect 11149 4091 11207 4097
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 11885 4131 11943 4137
rect 11296 4100 11341 4128
rect 11296 4088 11302 4100
rect 11885 4097 11897 4131
rect 11931 4128 11943 4131
rect 12360 4128 12388 4168
rect 13004 4137 13032 4168
rect 13262 4156 13268 4208
rect 13320 4196 13326 4208
rect 13320 4168 13768 4196
rect 13320 4156 13326 4168
rect 11931 4100 12388 4128
rect 12989 4131 13047 4137
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 13740 4128 13768 4168
rect 18708 4137 18736 4224
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13740 4100 13829 4128
rect 12989 4091 13047 4097
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 18693 4131 18751 4137
rect 18693 4097 18705 4131
rect 18739 4097 18751 4131
rect 18693 4091 18751 4097
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4128 19947 4131
rect 20824 4128 20852 4227
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 21818 4264 21824 4276
rect 21779 4236 21824 4264
rect 21818 4224 21824 4236
rect 21876 4224 21882 4276
rect 24029 4267 24087 4273
rect 24029 4233 24041 4267
rect 24075 4264 24087 4267
rect 24210 4264 24216 4276
rect 24075 4236 24216 4264
rect 24075 4233 24087 4236
rect 24029 4227 24087 4233
rect 24210 4224 24216 4236
rect 24268 4224 24274 4276
rect 23934 4156 23940 4208
rect 23992 4196 23998 4208
rect 24305 4199 24363 4205
rect 24305 4196 24317 4199
rect 23992 4168 24317 4196
rect 23992 4156 23998 4168
rect 24305 4165 24317 4168
rect 24351 4165 24363 4199
rect 24305 4159 24363 4165
rect 19935 4100 20852 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 11054 4060 11060 4072
rect 9692 4032 10732 4060
rect 11015 4032 11060 4060
rect 2133 3995 2191 4001
rect 2133 3992 2145 3995
rect 348 3964 2145 3992
rect 348 3952 354 3964
rect 2133 3961 2145 3964
rect 2179 3992 2191 3995
rect 2685 3995 2743 4001
rect 2685 3992 2697 3995
rect 2179 3964 2697 3992
rect 2179 3961 2191 3964
rect 2133 3955 2191 3961
rect 2685 3961 2697 3964
rect 2731 3961 2743 3995
rect 2685 3955 2743 3961
rect 2866 3952 2872 4004
rect 2924 3992 2930 4004
rect 3697 3995 3755 4001
rect 3697 3992 3709 3995
rect 2924 3964 3709 3992
rect 2924 3952 2930 3964
rect 3697 3961 3709 3964
rect 3743 3961 3755 3995
rect 6086 3992 6092 4004
rect 3697 3955 3755 3961
rect 4080 3964 6092 3992
rect 2961 3927 3019 3933
rect 2961 3893 2973 3927
rect 3007 3924 3019 3927
rect 4080 3924 4108 3964
rect 6086 3952 6092 3964
rect 6144 3992 6150 4004
rect 6181 3995 6239 4001
rect 6181 3992 6193 3995
rect 6144 3964 6193 3992
rect 6144 3952 6150 3964
rect 6181 3961 6193 3964
rect 6227 3961 6239 3995
rect 6181 3955 6239 3961
rect 8472 3995 8530 4001
rect 8472 3961 8484 3995
rect 8518 3992 8530 3995
rect 8570 3992 8576 4004
rect 8518 3964 8576 3992
rect 8518 3961 8530 3964
rect 8472 3955 8530 3961
rect 8570 3952 8576 3964
rect 8628 3952 8634 4004
rect 10502 3992 10508 4004
rect 10463 3964 10508 3992
rect 10502 3952 10508 3964
rect 10560 3952 10566 4004
rect 3007 3896 4108 3924
rect 4709 3927 4767 3933
rect 3007 3893 3019 3896
rect 2961 3887 3019 3893
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 4982 3924 4988 3936
rect 4755 3896 4988 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5074 3884 5080 3936
rect 5132 3924 5138 3936
rect 7190 3924 7196 3936
rect 5132 3896 5177 3924
rect 7151 3896 7196 3924
rect 5132 3884 5138 3896
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 9585 3927 9643 3933
rect 9585 3924 9597 3927
rect 8352 3896 9597 3924
rect 8352 3884 8358 3896
rect 9585 3893 9597 3896
rect 9631 3924 9643 3927
rect 10042 3924 10048 3936
rect 9631 3896 10048 3924
rect 9631 3893 9643 3896
rect 9585 3887 9643 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10704 3933 10732 4032
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 12618 4020 12624 4072
rect 12676 4060 12682 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12676 4032 12817 4060
rect 12676 4020 12682 4032
rect 12805 4029 12817 4032
rect 12851 4029 12863 4063
rect 12805 4023 12863 4029
rect 14090 4020 14096 4072
rect 14148 4060 14154 4072
rect 14185 4063 14243 4069
rect 14185 4060 14197 4063
rect 14148 4032 14197 4060
rect 14148 4020 14154 4032
rect 14185 4029 14197 4032
rect 14231 4029 14243 4063
rect 14185 4023 14243 4029
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4060 14519 4063
rect 14507 4032 14964 4060
rect 14507 4029 14519 4032
rect 14461 4023 14519 4029
rect 12897 3995 12955 4001
rect 12897 3992 12909 3995
rect 12176 3964 12909 3992
rect 10689 3927 10747 3933
rect 10689 3893 10701 3927
rect 10735 3893 10747 3927
rect 10689 3887 10747 3893
rect 12066 3884 12072 3936
rect 12124 3924 12130 3936
rect 12176 3933 12204 3964
rect 12897 3961 12909 3964
rect 12943 3961 12955 3995
rect 12897 3955 12955 3961
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 12124 3896 12173 3924
rect 12124 3884 12130 3896
rect 12161 3893 12173 3896
rect 12207 3893 12219 3927
rect 12161 3887 12219 3893
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12492 3896 12537 3924
rect 12492 3884 12498 3896
rect 13354 3884 13360 3936
rect 13412 3924 13418 3936
rect 13449 3927 13507 3933
rect 13449 3924 13461 3927
rect 13412 3896 13461 3924
rect 13412 3884 13418 3896
rect 13449 3893 13461 3896
rect 13495 3893 13507 3927
rect 13449 3887 13507 3893
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 14001 3927 14059 3933
rect 14001 3924 14013 3927
rect 13872 3896 14013 3924
rect 13872 3884 13878 3896
rect 14001 3893 14013 3896
rect 14047 3924 14059 3927
rect 14476 3924 14504 4023
rect 14936 4004 14964 4032
rect 19518 4020 19524 4072
rect 19576 4060 19582 4072
rect 19613 4063 19671 4069
rect 19613 4060 19625 4063
rect 19576 4032 19625 4060
rect 19576 4020 19582 4032
rect 19613 4029 19625 4032
rect 19659 4060 19671 4063
rect 20349 4063 20407 4069
rect 20349 4060 20361 4063
rect 19659 4032 20361 4060
rect 19659 4029 19671 4032
rect 19613 4023 19671 4029
rect 20349 4029 20361 4032
rect 20395 4029 20407 4063
rect 20898 4060 20904 4072
rect 20859 4032 20904 4060
rect 20349 4023 20407 4029
rect 20898 4020 20904 4032
rect 20956 4060 20962 4072
rect 21453 4063 21511 4069
rect 21453 4060 21465 4063
rect 20956 4032 21465 4060
rect 20956 4020 20962 4032
rect 21453 4029 21465 4032
rect 21499 4029 21511 4063
rect 21453 4023 21511 4029
rect 22005 4063 22063 4069
rect 22005 4029 22017 4063
rect 22051 4060 22063 4063
rect 22557 4063 22615 4069
rect 22557 4060 22569 4063
rect 22051 4032 22569 4060
rect 22051 4029 22063 4032
rect 22005 4023 22063 4029
rect 22557 4029 22569 4032
rect 22603 4029 22615 4063
rect 22557 4023 22615 4029
rect 14642 3952 14648 4004
rect 14700 4001 14706 4004
rect 14700 3995 14764 4001
rect 14700 3961 14718 3995
rect 14752 3961 14764 3995
rect 14700 3955 14764 3961
rect 14700 3952 14706 3955
rect 14918 3952 14924 4004
rect 14976 3952 14982 4004
rect 17954 3952 17960 4004
rect 18012 3992 18018 4004
rect 18506 3992 18512 4004
rect 18012 3964 18512 3992
rect 18012 3952 18018 3964
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 20714 3952 20720 4004
rect 20772 3992 20778 4004
rect 22020 3992 22048 4023
rect 20772 3964 22048 3992
rect 20772 3952 20778 3964
rect 15838 3924 15844 3936
rect 14047 3896 14504 3924
rect 15799 3896 15844 3924
rect 14047 3893 14059 3896
rect 14001 3887 14059 3893
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 16850 3924 16856 3936
rect 16811 3896 16856 3924
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 16942 3884 16948 3936
rect 17000 3924 17006 3936
rect 17000 3896 17045 3924
rect 17000 3884 17006 3896
rect 17126 3884 17132 3936
rect 17184 3924 17190 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 17184 3896 17417 3924
rect 17184 3884 17190 3896
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 17770 3924 17776 3936
rect 17731 3896 17776 3924
rect 17405 3887 17463 3893
rect 17770 3884 17776 3896
rect 17828 3924 17834 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 17828 3896 18429 3924
rect 17828 3884 17834 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 19426 3924 19432 3936
rect 19387 3896 19432 3924
rect 18417 3887 18475 3893
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 21082 3924 21088 3936
rect 21043 3896 21088 3924
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 22186 3924 22192 3936
rect 22147 3896 22192 3924
rect 22186 3884 22192 3896
rect 22244 3884 22250 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 2866 3720 2872 3732
rect 2648 3692 2872 3720
rect 2648 3680 2654 3692
rect 2866 3680 2872 3692
rect 2924 3680 2930 3732
rect 3142 3680 3148 3732
rect 3200 3720 3206 3732
rect 3513 3723 3571 3729
rect 3513 3720 3525 3723
rect 3200 3692 3525 3720
rect 3200 3680 3206 3692
rect 3513 3689 3525 3692
rect 3559 3720 3571 3723
rect 4062 3720 4068 3732
rect 3559 3692 4068 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 5166 3720 5172 3732
rect 5127 3692 5172 3720
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 6730 3720 6736 3732
rect 6691 3692 6736 3720
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 7745 3723 7803 3729
rect 7745 3689 7757 3723
rect 7791 3720 7803 3723
rect 8570 3720 8576 3732
rect 7791 3692 8576 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10100 3692 10701 3720
rect 10100 3680 10106 3692
rect 10689 3689 10701 3692
rect 10735 3720 10747 3723
rect 11057 3723 11115 3729
rect 11057 3720 11069 3723
rect 10735 3692 11069 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 11057 3689 11069 3692
rect 11103 3720 11115 3723
rect 11146 3720 11152 3732
rect 11103 3692 11152 3720
rect 11103 3689 11115 3692
rect 11057 3683 11115 3689
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 13265 3723 13323 3729
rect 13265 3689 13277 3723
rect 13311 3720 13323 3723
rect 13630 3720 13636 3732
rect 13311 3692 13636 3720
rect 13311 3689 13323 3692
rect 13265 3683 13323 3689
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 14737 3723 14795 3729
rect 14737 3689 14749 3723
rect 14783 3720 14795 3723
rect 14826 3720 14832 3732
rect 14783 3692 14832 3720
rect 14783 3689 14795 3692
rect 14737 3683 14795 3689
rect 1756 3655 1814 3661
rect 1756 3621 1768 3655
rect 1802 3652 1814 3655
rect 2222 3652 2228 3664
rect 1802 3624 2228 3652
rect 1802 3621 1814 3624
rect 1756 3615 1814 3621
rect 2222 3612 2228 3624
rect 2280 3612 2286 3664
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 5598 3655 5656 3661
rect 5598 3652 5610 3655
rect 5316 3624 5610 3652
rect 5316 3612 5322 3624
rect 5598 3621 5610 3624
rect 5644 3621 5656 3655
rect 5598 3615 5656 3621
rect 7282 3612 7288 3664
rect 7340 3652 7346 3664
rect 8297 3655 8355 3661
rect 8297 3652 8309 3655
rect 7340 3624 8309 3652
rect 7340 3612 7346 3624
rect 8297 3621 8309 3624
rect 8343 3652 8355 3655
rect 10137 3655 10195 3661
rect 10137 3652 10149 3655
rect 8343 3624 10149 3652
rect 8343 3621 8355 3624
rect 8297 3615 8355 3621
rect 10137 3621 10149 3624
rect 10183 3652 10195 3655
rect 10226 3652 10232 3664
rect 10183 3624 10232 3652
rect 10183 3621 10195 3624
rect 10137 3615 10195 3621
rect 10226 3612 10232 3624
rect 10284 3652 10290 3664
rect 10778 3652 10784 3664
rect 10284 3624 10784 3652
rect 10284 3612 10290 3624
rect 10778 3612 10784 3624
rect 10836 3612 10842 3664
rect 11508 3655 11566 3661
rect 11508 3621 11520 3655
rect 11554 3652 11566 3655
rect 11698 3652 11704 3664
rect 11554 3624 11704 3652
rect 11554 3621 11566 3624
rect 11508 3615 11566 3621
rect 11698 3612 11704 3624
rect 11756 3612 11762 3664
rect 14182 3652 14188 3664
rect 14143 3624 14188 3652
rect 14182 3612 14188 3624
rect 14240 3612 14246 3664
rect 5350 3584 5356 3596
rect 5311 3556 5356 3584
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 8251 3556 10057 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 10045 3553 10057 3556
rect 10091 3584 10103 3587
rect 10410 3584 10416 3596
rect 10091 3556 10416 3584
rect 10091 3553 10103 3556
rect 10045 3547 10103 3553
rect 1486 3516 1492 3528
rect 1447 3488 1492 3516
rect 1486 3476 1492 3488
rect 1544 3476 1550 3528
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 4341 3519 4399 3525
rect 4341 3516 4353 3519
rect 3108 3488 4353 3516
rect 3108 3476 3114 3488
rect 4341 3485 4353 3488
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3516 7435 3519
rect 7466 3516 7472 3528
rect 7423 3488 7472 3516
rect 7423 3485 7435 3488
rect 7377 3479 7435 3485
rect 7466 3476 7472 3488
rect 7524 3516 7530 3528
rect 7524 3488 7972 3516
rect 7524 3476 7530 3488
rect 3878 3448 3884 3460
rect 3839 3420 3884 3448
rect 3878 3408 3884 3420
rect 3936 3408 3942 3460
rect 7834 3448 7840 3460
rect 7795 3420 7840 3448
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 7944 3448 7972 3488
rect 8018 3476 8024 3528
rect 8076 3516 8082 3528
rect 8220 3516 8248 3547
rect 10410 3544 10416 3556
rect 10468 3584 10474 3596
rect 12066 3584 12072 3596
rect 10468 3556 12072 3584
rect 10468 3544 10474 3556
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 13814 3544 13820 3596
rect 13872 3544 13878 3596
rect 13909 3587 13967 3593
rect 13909 3553 13921 3587
rect 13955 3584 13967 3587
rect 14752 3584 14780 3683
rect 14826 3680 14832 3692
rect 14884 3680 14890 3732
rect 15565 3723 15623 3729
rect 15565 3689 15577 3723
rect 15611 3720 15623 3723
rect 15746 3720 15752 3732
rect 15611 3692 15752 3720
rect 15611 3689 15623 3692
rect 15565 3683 15623 3689
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 16942 3680 16948 3732
rect 17000 3720 17006 3732
rect 18601 3723 18659 3729
rect 18601 3720 18613 3723
rect 17000 3692 18613 3720
rect 17000 3680 17006 3692
rect 18601 3689 18613 3692
rect 18647 3720 18659 3723
rect 19058 3720 19064 3732
rect 18647 3692 19064 3720
rect 18647 3689 18659 3692
rect 18601 3683 18659 3689
rect 19058 3680 19064 3692
rect 19116 3680 19122 3732
rect 19242 3680 19248 3732
rect 19300 3720 19306 3732
rect 19337 3723 19395 3729
rect 19337 3720 19349 3723
rect 19300 3692 19349 3720
rect 19300 3680 19306 3692
rect 19337 3689 19349 3692
rect 19383 3720 19395 3723
rect 20070 3720 20076 3732
rect 19383 3692 20076 3720
rect 19383 3689 19395 3692
rect 19337 3683 19395 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20898 3680 20904 3732
rect 20956 3720 20962 3732
rect 22186 3720 22192 3732
rect 20956 3692 22192 3720
rect 20956 3680 20962 3692
rect 22186 3680 22192 3692
rect 22244 3680 22250 3732
rect 15838 3612 15844 3664
rect 15896 3652 15902 3664
rect 16016 3655 16074 3661
rect 16016 3652 16028 3655
rect 15896 3624 16028 3652
rect 15896 3612 15902 3624
rect 16016 3621 16028 3624
rect 16062 3652 16074 3655
rect 16850 3652 16856 3664
rect 16062 3624 16856 3652
rect 16062 3621 16074 3624
rect 16016 3615 16074 3621
rect 16850 3612 16856 3624
rect 16908 3612 16914 3664
rect 17678 3652 17684 3664
rect 16960 3624 17684 3652
rect 16960 3596 16988 3624
rect 17678 3612 17684 3624
rect 17736 3612 17742 3664
rect 17954 3612 17960 3664
rect 18012 3652 18018 3664
rect 18049 3655 18107 3661
rect 18049 3652 18061 3655
rect 18012 3624 18061 3652
rect 18012 3612 18018 3624
rect 18049 3621 18061 3624
rect 18095 3621 18107 3655
rect 18690 3652 18696 3664
rect 18651 3624 18696 3652
rect 18049 3615 18107 3621
rect 18690 3612 18696 3624
rect 18748 3652 18754 3664
rect 18966 3652 18972 3664
rect 18748 3624 18972 3652
rect 18748 3612 18754 3624
rect 18966 3612 18972 3624
rect 19024 3612 19030 3664
rect 22094 3612 22100 3664
rect 22152 3652 22158 3664
rect 22152 3624 23336 3652
rect 22152 3612 22158 3624
rect 23308 3596 23336 3624
rect 24854 3612 24860 3664
rect 24912 3652 24918 3664
rect 25958 3652 25964 3664
rect 24912 3624 25964 3652
rect 24912 3612 24918 3624
rect 25958 3612 25964 3624
rect 26016 3612 26022 3664
rect 13955 3556 14780 3584
rect 13955 3553 13967 3556
rect 13909 3547 13967 3553
rect 14826 3544 14832 3596
rect 14884 3584 14890 3596
rect 15105 3587 15163 3593
rect 15105 3584 15117 3587
rect 14884 3556 15117 3584
rect 14884 3544 14890 3556
rect 15105 3553 15117 3556
rect 15151 3584 15163 3587
rect 15749 3587 15807 3593
rect 15749 3584 15761 3587
rect 15151 3556 15761 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15749 3553 15761 3556
rect 15795 3584 15807 3587
rect 16942 3584 16948 3596
rect 15795 3556 16948 3584
rect 15795 3553 15807 3556
rect 15749 3547 15807 3553
rect 16942 3544 16948 3556
rect 17000 3544 17006 3596
rect 20901 3587 20959 3593
rect 20901 3553 20913 3587
rect 20947 3553 20959 3587
rect 22186 3584 22192 3596
rect 22147 3556 22192 3584
rect 20901 3547 20959 3553
rect 8076 3488 8248 3516
rect 8389 3519 8447 3525
rect 8076 3476 8082 3488
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8404 3448 8432 3479
rect 8570 3476 8576 3528
rect 8628 3516 8634 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8628 3488 8953 3516
rect 8628 3476 8634 3488
rect 8941 3485 8953 3488
rect 8987 3516 8999 3519
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 8987 3488 9505 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 9493 3485 9505 3488
rect 9539 3516 9551 3519
rect 10321 3519 10379 3525
rect 10321 3516 10333 3519
rect 9539 3488 10333 3516
rect 9539 3485 9551 3488
rect 9493 3479 9551 3485
rect 10321 3485 10333 3488
rect 10367 3516 10379 3519
rect 10686 3516 10692 3528
rect 10367 3488 10692 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 11241 3519 11299 3525
rect 11241 3485 11253 3519
rect 11287 3485 11299 3519
rect 11241 3479 11299 3485
rect 7944 3420 8432 3448
rect 9677 3451 9735 3457
rect 9677 3417 9689 3451
rect 9723 3448 9735 3451
rect 10778 3448 10784 3460
rect 9723 3420 10784 3448
rect 9723 3417 9735 3420
rect 9677 3411 9735 3417
rect 10778 3408 10784 3420
rect 10836 3408 10842 3460
rect 4890 3380 4896 3392
rect 4851 3352 4896 3380
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 11256 3380 11284 3479
rect 13832 3448 13860 3544
rect 18782 3516 18788 3528
rect 18743 3488 18788 3516
rect 18782 3476 18788 3488
rect 18840 3476 18846 3528
rect 12452 3420 13860 3448
rect 18233 3451 18291 3457
rect 12342 3380 12348 3392
rect 11256 3352 12348 3380
rect 12342 3340 12348 3352
rect 12400 3380 12406 3392
rect 12452 3380 12480 3420
rect 18233 3417 18245 3451
rect 18279 3448 18291 3451
rect 20714 3448 20720 3460
rect 18279 3420 20720 3448
rect 18279 3417 18291 3420
rect 18233 3411 18291 3417
rect 20714 3408 20720 3420
rect 20772 3448 20778 3460
rect 20916 3448 20944 3547
rect 22186 3544 22192 3556
rect 22244 3544 22250 3596
rect 23290 3584 23296 3596
rect 23203 3556 23296 3584
rect 23290 3544 23296 3556
rect 23348 3544 23354 3596
rect 24946 3544 24952 3596
rect 25004 3584 25010 3596
rect 25406 3584 25412 3596
rect 25004 3556 25412 3584
rect 25004 3544 25010 3556
rect 25406 3544 25412 3556
rect 25464 3544 25470 3596
rect 21174 3516 21180 3528
rect 21135 3488 21180 3516
rect 21174 3476 21180 3488
rect 21232 3476 21238 3528
rect 20772 3420 20944 3448
rect 20772 3408 20778 3420
rect 12618 3380 12624 3392
rect 12400 3352 12480 3380
rect 12579 3352 12624 3380
rect 12400 3340 12406 3352
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 13633 3383 13691 3389
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 13722 3380 13728 3392
rect 13679 3352 13728 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 17126 3380 17132 3392
rect 17087 3352 17132 3380
rect 17126 3340 17132 3352
rect 17184 3340 17190 3392
rect 22370 3380 22376 3392
rect 22331 3352 22376 3380
rect 22370 3340 22376 3352
rect 22428 3340 22434 3392
rect 23477 3383 23535 3389
rect 23477 3349 23489 3383
rect 23523 3380 23535 3383
rect 23750 3380 23756 3392
rect 23523 3352 23756 3380
rect 23523 3349 23535 3352
rect 23477 3343 23535 3349
rect 23750 3340 23756 3352
rect 23808 3340 23814 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2041 3179 2099 3185
rect 2041 3145 2053 3179
rect 2087 3176 2099 3179
rect 2222 3176 2228 3188
rect 2087 3148 2228 3176
rect 2087 3145 2099 3148
rect 2041 3139 2099 3145
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 2682 3176 2688 3188
rect 2643 3148 2688 3176
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 4154 3176 4160 3188
rect 4115 3148 4160 3176
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 5629 3179 5687 3185
rect 5629 3176 5641 3179
rect 5224 3148 5641 3176
rect 5224 3136 5230 3148
rect 5629 3145 5641 3148
rect 5675 3176 5687 3179
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 5675 3148 6193 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 6181 3145 6193 3148
rect 6227 3145 6239 3179
rect 6546 3176 6552 3188
rect 6507 3148 6552 3176
rect 6181 3139 6239 3145
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7282 3176 7288 3188
rect 6972 3148 7288 3176
rect 6972 3136 6978 3148
rect 7282 3136 7288 3148
rect 7340 3176 7346 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7340 3148 7849 3176
rect 7340 3136 7346 3148
rect 7837 3145 7849 3148
rect 7883 3145 7895 3179
rect 7837 3139 7895 3145
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 9548 3148 10609 3176
rect 9548 3136 9554 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 14366 3176 14372 3188
rect 12492 3148 14372 3176
rect 12492 3136 12498 3148
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 16850 3176 16856 3188
rect 16811 3148 16856 3176
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 17184 3148 17509 3176
rect 17184 3136 17190 3148
rect 17497 3145 17509 3148
rect 17543 3176 17555 3179
rect 18782 3176 18788 3188
rect 17543 3148 18788 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 18782 3136 18788 3148
rect 18840 3136 18846 3188
rect 19058 3176 19064 3188
rect 19019 3148 19064 3176
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 20714 3176 20720 3188
rect 20675 3148 20720 3176
rect 20714 3136 20720 3148
rect 20772 3136 20778 3188
rect 22097 3179 22155 3185
rect 22097 3145 22109 3179
rect 22143 3176 22155 3179
rect 22186 3176 22192 3188
rect 22143 3148 22192 3176
rect 22143 3145 22155 3148
rect 22097 3139 22155 3145
rect 2240 3108 2268 3136
rect 2866 3108 2872 3120
rect 2240 3080 2872 3108
rect 2866 3068 2872 3080
rect 2924 3108 2930 3120
rect 3697 3111 3755 3117
rect 3697 3108 3709 3111
rect 2924 3080 3709 3108
rect 2924 3068 2930 3080
rect 3697 3077 3709 3080
rect 3743 3077 3755 3111
rect 3697 3071 3755 3077
rect 3142 3040 3148 3052
rect 3103 3012 3148 3040
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3040 3387 3043
rect 3510 3040 3516 3052
rect 3375 3012 3516 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 3510 3000 3516 3012
rect 3568 3040 3574 3052
rect 4172 3040 4200 3136
rect 10137 3111 10195 3117
rect 10137 3077 10149 3111
rect 10183 3108 10195 3111
rect 10226 3108 10232 3120
rect 10183 3080 10232 3108
rect 10183 3077 10195 3080
rect 10137 3071 10195 3077
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 10410 3108 10416 3120
rect 10371 3080 10416 3108
rect 10410 3068 10416 3080
rect 10468 3068 10474 3120
rect 13814 3108 13820 3120
rect 13775 3080 13820 3108
rect 13814 3068 13820 3080
rect 13872 3108 13878 3120
rect 14737 3111 14795 3117
rect 14737 3108 14749 3111
rect 13872 3080 14749 3108
rect 13872 3068 13878 3080
rect 14737 3077 14749 3080
rect 14783 3077 14795 3111
rect 14737 3071 14795 3077
rect 18049 3111 18107 3117
rect 18049 3077 18061 3111
rect 18095 3108 18107 3111
rect 19426 3108 19432 3120
rect 18095 3080 19432 3108
rect 18095 3077 18107 3080
rect 18049 3071 18107 3077
rect 3568 3012 4384 3040
rect 3568 3000 3574 3012
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2972 2651 2975
rect 3050 2972 3056 2984
rect 2639 2944 3056 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 3050 2932 3056 2944
rect 3108 2932 3114 2984
rect 4062 2932 4068 2984
rect 4120 2972 4126 2984
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 4120 2944 4261 2972
rect 4120 2932 4126 2944
rect 4249 2941 4261 2944
rect 4295 2941 4307 2975
rect 4356 2972 4384 3012
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 7156 3012 8125 3040
rect 7156 3000 7162 3012
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 11146 3040 11152 3052
rect 11107 3012 11152 3040
rect 8113 3003 8171 3009
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 12342 3000 12348 3052
rect 12400 3040 12406 3052
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 12400 3012 12449 3040
rect 12400 3000 12406 3012
rect 12437 3009 12449 3012
rect 12483 3009 12495 3043
rect 14752 3040 14780 3071
rect 19426 3068 19432 3080
rect 19484 3068 19490 3120
rect 18598 3040 18604 3052
rect 14752 3012 15056 3040
rect 18559 3012 18604 3040
rect 12437 3003 12495 3009
rect 4505 2975 4563 2981
rect 4505 2972 4517 2975
rect 4356 2944 4517 2972
rect 4249 2935 4307 2941
rect 4505 2941 4517 2944
rect 4551 2941 4563 2975
rect 4505 2935 4563 2941
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11057 2975 11115 2981
rect 11057 2972 11069 2975
rect 11020 2944 11069 2972
rect 11020 2932 11026 2944
rect 11057 2941 11069 2944
rect 11103 2941 11115 2975
rect 11057 2935 11115 2941
rect 14826 2932 14832 2984
rect 14884 2972 14890 2984
rect 14921 2975 14979 2981
rect 14921 2972 14933 2975
rect 14884 2944 14933 2972
rect 14884 2932 14890 2944
rect 14921 2941 14933 2944
rect 14967 2941 14979 2975
rect 15028 2972 15056 3012
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 20349 3043 20407 3049
rect 20349 3040 20361 3043
rect 19392 3012 20361 3040
rect 19392 3000 19398 3012
rect 15177 2975 15235 2981
rect 15177 2972 15189 2975
rect 15028 2944 15189 2972
rect 14921 2935 14979 2941
rect 15177 2941 15189 2944
rect 15223 2941 15235 2975
rect 18506 2972 18512 2984
rect 18467 2944 18512 2972
rect 15177 2935 15235 2941
rect 18506 2932 18512 2944
rect 18564 2972 18570 2984
rect 19628 2981 19656 3012
rect 20349 3009 20361 3012
rect 20395 3009 20407 3043
rect 20349 3003 20407 3009
rect 21177 3043 21235 3049
rect 21177 3009 21189 3043
rect 21223 3040 21235 3043
rect 22112 3040 22140 3139
rect 22186 3136 22192 3148
rect 22244 3136 22250 3188
rect 22373 3179 22431 3185
rect 22373 3145 22385 3179
rect 22419 3176 22431 3179
rect 22462 3176 22468 3188
rect 22419 3148 22468 3176
rect 22419 3145 22431 3148
rect 22373 3139 22431 3145
rect 22462 3136 22468 3148
rect 22520 3136 22526 3188
rect 23290 3176 23296 3188
rect 23251 3148 23296 3176
rect 23290 3136 23296 3148
rect 23348 3136 23354 3188
rect 24949 3111 25007 3117
rect 24949 3077 24961 3111
rect 24995 3108 25007 3111
rect 26510 3108 26516 3120
rect 24995 3080 26516 3108
rect 24995 3077 25007 3080
rect 24949 3071 25007 3077
rect 26510 3068 26516 3080
rect 26568 3068 26574 3120
rect 21223 3012 22140 3040
rect 21223 3009 21235 3012
rect 21177 3003 21235 3009
rect 19429 2975 19487 2981
rect 19429 2972 19441 2975
rect 18564 2944 19441 2972
rect 18564 2932 18570 2944
rect 19429 2941 19441 2944
rect 19475 2941 19487 2975
rect 19429 2935 19487 2941
rect 19613 2975 19671 2981
rect 19613 2941 19625 2975
rect 19659 2941 19671 2975
rect 19613 2935 19671 2941
rect 20806 2932 20812 2984
rect 20864 2972 20870 2984
rect 20901 2975 20959 2981
rect 20901 2972 20913 2975
rect 20864 2944 20913 2972
rect 20864 2932 20870 2944
rect 20901 2941 20913 2944
rect 20947 2972 20959 2975
rect 21637 2975 21695 2981
rect 21637 2972 21649 2975
rect 20947 2944 21649 2972
rect 20947 2941 20959 2944
rect 20901 2935 20959 2941
rect 21637 2941 21649 2944
rect 21683 2941 21695 2975
rect 21637 2935 21695 2941
rect 22189 2975 22247 2981
rect 22189 2941 22201 2975
rect 22235 2972 22247 2975
rect 22278 2972 22284 2984
rect 22235 2944 22284 2972
rect 22235 2941 22247 2944
rect 22189 2935 22247 2941
rect 22278 2932 22284 2944
rect 22336 2972 22342 2984
rect 22741 2975 22799 2981
rect 22741 2972 22753 2975
rect 22336 2944 22753 2972
rect 22336 2932 22342 2944
rect 22741 2941 22753 2944
rect 22787 2941 22799 2975
rect 23658 2972 23664 2984
rect 23619 2944 23664 2972
rect 22741 2935 22799 2941
rect 23658 2932 23664 2944
rect 23716 2972 23722 2984
rect 24213 2975 24271 2981
rect 24213 2972 24225 2975
rect 23716 2944 24225 2972
rect 23716 2932 23722 2944
rect 24213 2941 24225 2944
rect 24259 2941 24271 2975
rect 24213 2935 24271 2941
rect 24670 2932 24676 2984
rect 24728 2972 24734 2984
rect 24765 2975 24823 2981
rect 24765 2972 24777 2975
rect 24728 2944 24777 2972
rect 24728 2932 24734 2944
rect 24765 2941 24777 2944
rect 24811 2972 24823 2975
rect 25317 2975 25375 2981
rect 25317 2972 25329 2975
rect 24811 2944 25329 2972
rect 24811 2941 24823 2944
rect 24765 2935 24823 2941
rect 25317 2941 25329 2944
rect 25363 2941 25375 2975
rect 25317 2935 25375 2941
rect 1670 2904 1676 2916
rect 1631 2876 1676 2904
rect 1670 2864 1676 2876
rect 1728 2864 1734 2916
rect 7098 2904 7104 2916
rect 7059 2876 7104 2904
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 8386 2913 8392 2916
rect 8380 2904 8392 2913
rect 8347 2876 8392 2904
rect 8380 2867 8392 2876
rect 8386 2864 8392 2867
rect 8444 2864 8450 2916
rect 12253 2907 12311 2913
rect 12253 2873 12265 2907
rect 12299 2904 12311 2907
rect 12618 2904 12624 2916
rect 12299 2876 12624 2904
rect 12299 2873 12311 2876
rect 12253 2867 12311 2873
rect 12618 2864 12624 2876
rect 12676 2913 12682 2916
rect 12676 2907 12740 2913
rect 12676 2873 12694 2907
rect 12728 2904 12740 2907
rect 12728 2876 12769 2904
rect 12728 2873 12740 2876
rect 12676 2867 12740 2873
rect 12676 2864 12682 2867
rect 14642 2864 14648 2916
rect 14700 2904 14706 2916
rect 17770 2904 17776 2916
rect 14700 2876 14872 2904
rect 17731 2876 17776 2904
rect 14700 2864 14706 2876
rect 6546 2796 6552 2848
rect 6604 2836 6610 2848
rect 7466 2836 7472 2848
rect 6604 2808 7472 2836
rect 6604 2796 6610 2808
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 9490 2836 9496 2848
rect 9451 2808 9496 2836
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 10778 2796 10784 2848
rect 10836 2836 10842 2848
rect 10965 2839 11023 2845
rect 10965 2836 10977 2839
rect 10836 2808 10977 2836
rect 10836 2796 10842 2808
rect 10965 2805 10977 2808
rect 11011 2805 11023 2839
rect 11698 2836 11704 2848
rect 11659 2808 11704 2836
rect 10965 2799 11023 2805
rect 11698 2796 11704 2808
rect 11756 2796 11762 2848
rect 14844 2836 14872 2876
rect 17770 2864 17776 2876
rect 17828 2904 17834 2916
rect 18417 2907 18475 2913
rect 18417 2904 18429 2907
rect 17828 2876 18429 2904
rect 17828 2864 17834 2876
rect 18417 2873 18429 2876
rect 18463 2873 18475 2907
rect 18417 2867 18475 2873
rect 19334 2864 19340 2916
rect 19392 2904 19398 2916
rect 19889 2907 19947 2913
rect 19889 2904 19901 2907
rect 19392 2876 19901 2904
rect 19392 2864 19398 2876
rect 19889 2873 19901 2876
rect 19935 2873 19947 2907
rect 19889 2867 19947 2873
rect 22094 2864 22100 2916
rect 22152 2904 22158 2916
rect 22152 2876 23888 2904
rect 22152 2864 22158 2876
rect 16301 2839 16359 2845
rect 16301 2836 16313 2839
rect 14844 2808 16313 2836
rect 16301 2805 16313 2808
rect 16347 2805 16359 2839
rect 16301 2799 16359 2805
rect 18046 2796 18052 2848
rect 18104 2836 18110 2848
rect 18598 2836 18604 2848
rect 18104 2808 18604 2836
rect 18104 2796 18110 2808
rect 18598 2796 18604 2808
rect 18656 2796 18662 2848
rect 23860 2845 23888 2876
rect 23845 2839 23903 2845
rect 23845 2805 23857 2839
rect 23891 2805 23903 2839
rect 23845 2799 23903 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2866 2632 2872 2644
rect 2827 2604 2872 2632
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 6914 2632 6920 2644
rect 6875 2604 6920 2632
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 8386 2632 8392 2644
rect 8347 2604 8392 2632
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 10686 2592 10692 2644
rect 10744 2632 10750 2644
rect 10781 2635 10839 2641
rect 10781 2632 10793 2635
rect 10744 2604 10793 2632
rect 10744 2592 10750 2604
rect 10781 2601 10793 2604
rect 10827 2601 10839 2635
rect 11606 2632 11612 2644
rect 11567 2604 11612 2632
rect 10781 2595 10839 2601
rect 11606 2592 11612 2604
rect 11664 2592 11670 2644
rect 12894 2632 12900 2644
rect 12855 2604 12900 2632
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 14366 2632 14372 2644
rect 14323 2604 14372 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 15473 2635 15531 2641
rect 15473 2601 15485 2635
rect 15519 2632 15531 2635
rect 15654 2632 15660 2644
rect 15519 2604 15660 2632
rect 15519 2601 15531 2604
rect 15473 2595 15531 2601
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 16942 2632 16948 2644
rect 16903 2604 16948 2632
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 17678 2632 17684 2644
rect 17639 2604 17684 2632
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 18966 2592 18972 2644
rect 19024 2632 19030 2644
rect 19061 2635 19119 2641
rect 19061 2632 19073 2635
rect 19024 2604 19073 2632
rect 19024 2592 19030 2604
rect 19061 2601 19073 2604
rect 19107 2601 19119 2635
rect 22646 2632 22652 2644
rect 22607 2604 22652 2632
rect 19061 2595 19119 2601
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 24762 2632 24768 2644
rect 24723 2604 24768 2632
rect 24762 2592 24768 2604
rect 24820 2592 24826 2644
rect 1670 2524 1676 2576
rect 1728 2573 1734 2576
rect 1728 2567 1792 2573
rect 1728 2533 1746 2567
rect 1780 2533 1792 2567
rect 1728 2527 1792 2533
rect 3881 2567 3939 2573
rect 3881 2533 3893 2567
rect 3927 2564 3939 2567
rect 4332 2567 4390 2573
rect 4332 2564 4344 2567
rect 3927 2536 4344 2564
rect 3927 2533 3939 2536
rect 3881 2527 3939 2533
rect 4332 2533 4344 2536
rect 4378 2564 4390 2567
rect 4522 2564 4528 2576
rect 4378 2536 4528 2564
rect 4378 2533 4390 2536
rect 4332 2527 4390 2533
rect 1728 2524 1734 2527
rect 4522 2524 4528 2536
rect 4580 2524 4586 2576
rect 9493 2567 9551 2573
rect 9493 2564 9505 2567
rect 7300 2536 9505 2564
rect 1486 2496 1492 2508
rect 1447 2468 1492 2496
rect 1486 2456 1492 2468
rect 1544 2496 1550 2508
rect 4062 2496 4068 2508
rect 1544 2468 4068 2496
rect 1544 2456 1550 2468
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 6638 2496 6644 2508
rect 6599 2468 6644 2496
rect 6638 2456 6644 2468
rect 6696 2496 6702 2508
rect 7300 2505 7328 2536
rect 9493 2533 9505 2536
rect 9539 2564 9551 2567
rect 9674 2564 9680 2576
rect 9539 2536 9680 2564
rect 9539 2533 9551 2536
rect 9493 2527 9551 2533
rect 9674 2524 9680 2536
rect 9732 2564 9738 2576
rect 10137 2567 10195 2573
rect 10137 2564 10149 2567
rect 9732 2536 10149 2564
rect 9732 2524 9738 2536
rect 10137 2533 10149 2536
rect 10183 2533 10195 2567
rect 10137 2527 10195 2533
rect 13357 2567 13415 2573
rect 13357 2533 13369 2567
rect 13403 2564 13415 2567
rect 13403 2536 14504 2564
rect 13403 2533 13415 2536
rect 13357 2527 13415 2533
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6696 2468 7297 2496
rect 6696 2456 6702 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 7285 2459 7343 2465
rect 7392 2468 9137 2496
rect 7392 2437 7420 2468
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 12066 2496 12072 2508
rect 11471 2468 12072 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 6411 2400 7389 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 8662 2428 8668 2440
rect 7524 2400 7569 2428
rect 8623 2400 8668 2428
rect 7524 2388 7530 2400
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 9140 2428 9168 2459
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 12437 2499 12495 2505
rect 12437 2465 12449 2499
rect 12483 2496 12495 2499
rect 12710 2496 12716 2508
rect 12483 2468 12716 2496
rect 12483 2465 12495 2468
rect 12437 2459 12495 2465
rect 12710 2456 12716 2468
rect 12768 2456 12774 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13648 2468 14197 2496
rect 9858 2428 9864 2440
rect 9140 2400 9864 2428
rect 9858 2388 9864 2400
rect 9916 2428 9922 2440
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 9916 2400 10241 2428
rect 9916 2388 9922 2400
rect 10229 2397 10241 2400
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10686 2428 10692 2440
rect 10459 2400 10692 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 10836 2400 11989 2428
rect 10836 2388 10842 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 9769 2363 9827 2369
rect 9769 2329 9781 2363
rect 9815 2360 9827 2363
rect 10962 2360 10968 2372
rect 9815 2332 10968 2360
rect 9815 2329 9827 2332
rect 9769 2323 9827 2329
rect 10962 2320 10968 2332
rect 11020 2360 11026 2372
rect 11149 2363 11207 2369
rect 11149 2360 11161 2363
rect 11020 2332 11161 2360
rect 11020 2320 11026 2332
rect 11149 2329 11161 2332
rect 11195 2329 11207 2363
rect 11149 2323 11207 2329
rect 13538 2320 13544 2372
rect 13596 2360 13602 2372
rect 13648 2369 13676 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 14476 2437 14504 2536
rect 15286 2524 15292 2576
rect 15344 2564 15350 2576
rect 15933 2567 15991 2573
rect 15933 2564 15945 2567
rect 15344 2536 15945 2564
rect 15344 2524 15350 2536
rect 15933 2533 15945 2536
rect 15979 2533 15991 2567
rect 15933 2527 15991 2533
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 14844 2468 15853 2496
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 14642 2428 14648 2440
rect 14507 2400 14648 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 14642 2388 14648 2400
rect 14700 2388 14706 2440
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 13596 2332 13645 2360
rect 13596 2320 13602 2332
rect 13633 2329 13645 2332
rect 13679 2329 13691 2363
rect 13814 2360 13820 2372
rect 13775 2332 13820 2360
rect 13633 2323 13691 2329
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 3510 2292 3516 2304
rect 3423 2264 3516 2292
rect 3510 2252 3516 2264
rect 3568 2292 3574 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 3568 2264 5457 2292
rect 3568 2252 3574 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 14550 2252 14556 2304
rect 14608 2292 14614 2304
rect 14844 2301 14872 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2496 17095 2499
rect 17696 2496 17724 2592
rect 21453 2567 21511 2573
rect 21453 2533 21465 2567
rect 21499 2564 21511 2567
rect 21634 2564 21640 2576
rect 21499 2536 21640 2564
rect 21499 2533 21511 2536
rect 21453 2527 21511 2533
rect 21634 2524 21640 2536
rect 21692 2524 21698 2576
rect 18322 2496 18328 2508
rect 17083 2468 17724 2496
rect 18283 2468 18328 2496
rect 17083 2465 17095 2468
rect 17037 2459 17095 2465
rect 18322 2456 18328 2468
rect 18380 2496 18386 2508
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 18380 2468 19441 2496
rect 18380 2456 18386 2468
rect 19429 2465 19441 2468
rect 19475 2465 19487 2499
rect 19610 2496 19616 2508
rect 19571 2468 19616 2496
rect 19429 2459 19487 2465
rect 19610 2456 19616 2468
rect 19668 2496 19674 2508
rect 20349 2499 20407 2505
rect 20349 2496 20361 2499
rect 19668 2468 20361 2496
rect 19668 2456 19674 2468
rect 20349 2465 20361 2468
rect 20395 2465 20407 2499
rect 21174 2496 21180 2508
rect 21135 2468 21180 2496
rect 20349 2459 20407 2465
rect 21174 2456 21180 2468
rect 21232 2496 21238 2508
rect 21913 2499 21971 2505
rect 21913 2496 21925 2499
rect 21232 2468 21925 2496
rect 21232 2456 21238 2468
rect 21913 2465 21925 2468
rect 21959 2465 21971 2499
rect 22462 2496 22468 2508
rect 22423 2468 22468 2496
rect 21913 2459 21971 2465
rect 22462 2456 22468 2468
rect 22520 2496 22526 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22520 2468 23029 2496
rect 22520 2456 22526 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 23017 2459 23075 2465
rect 24118 2456 24124 2508
rect 24176 2496 24182 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 24176 2468 24593 2496
rect 24176 2456 24182 2468
rect 24581 2465 24593 2468
rect 24627 2496 24639 2499
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24627 2468 25145 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 16022 2428 16028 2440
rect 15983 2400 16028 2428
rect 16022 2388 16028 2400
rect 16080 2428 16086 2440
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 16080 2400 16497 2428
rect 16080 2388 16086 2400
rect 16485 2397 16497 2400
rect 16531 2397 16543 2431
rect 18506 2428 18512 2440
rect 18467 2400 18512 2428
rect 16485 2391 16543 2397
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 19794 2428 19800 2440
rect 19755 2400 19800 2428
rect 19794 2388 19800 2400
rect 19852 2388 19858 2440
rect 14829 2295 14887 2301
rect 14829 2292 14841 2295
rect 14608 2264 14841 2292
rect 14608 2252 14614 2264
rect 14829 2261 14841 2264
rect 14875 2261 14887 2295
rect 15286 2292 15292 2304
rect 15247 2264 15292 2292
rect 14829 2255 14887 2261
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 16574 2252 16580 2304
rect 16632 2292 16638 2304
rect 17221 2295 17279 2301
rect 17221 2292 17233 2295
rect 16632 2264 17233 2292
rect 16632 2252 16638 2264
rect 17221 2261 17233 2264
rect 17267 2261 17279 2295
rect 17221 2255 17279 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 8662 1368 8668 1420
rect 8720 1408 8726 1420
rect 9582 1408 9588 1420
rect 8720 1380 9588 1408
rect 8720 1368 8726 1380
rect 9582 1368 9588 1380
rect 9640 1368 9646 1420
rect 11790 552 11796 604
rect 11848 592 11854 604
rect 13078 592 13084 604
rect 11848 564 13084 592
rect 11848 552 11854 564
rect 13078 552 13084 564
rect 13136 552 13142 604
<< via1 >>
rect 3332 26664 3384 26716
rect 5448 26664 5500 26716
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 2780 25440 2832 25492
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 1584 24939 1636 24948
rect 1584 24905 1593 24939
rect 1593 24905 1627 24939
rect 1627 24905 1636 24939
rect 1584 24896 1636 24905
rect 2136 24556 2188 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1492 24352 1544 24404
rect 2688 24395 2740 24404
rect 2688 24361 2697 24395
rect 2697 24361 2731 24395
rect 2731 24361 2740 24395
rect 2688 24352 2740 24361
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 2504 24259 2556 24268
rect 2504 24225 2513 24259
rect 2513 24225 2547 24259
rect 2547 24225 2556 24259
rect 2504 24216 2556 24225
rect 2044 24123 2096 24132
rect 2044 24089 2053 24123
rect 2053 24089 2087 24123
rect 2087 24089 2096 24123
rect 2044 24080 2096 24089
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2504 23851 2556 23860
rect 2504 23817 2513 23851
rect 2513 23817 2547 23851
rect 2547 23817 2556 23851
rect 2504 23808 2556 23817
rect 3240 23851 3292 23860
rect 3240 23817 3249 23851
rect 3249 23817 3283 23851
rect 3283 23817 3292 23851
rect 3240 23808 3292 23817
rect 24768 23851 24820 23860
rect 24768 23817 24777 23851
rect 24777 23817 24811 23851
rect 24811 23817 24820 23851
rect 24768 23808 24820 23817
rect 3700 23715 3752 23724
rect 1952 23604 2004 23656
rect 3700 23681 3709 23715
rect 3709 23681 3743 23715
rect 3743 23681 3752 23715
rect 3700 23672 3752 23681
rect 1400 23468 1452 23520
rect 1952 23468 2004 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2136 23196 2188 23248
rect 12716 23239 12768 23248
rect 12716 23205 12725 23239
rect 12725 23205 12759 23239
rect 12759 23205 12768 23239
rect 12716 23196 12768 23205
rect 1676 23128 1728 23180
rect 12440 23171 12492 23180
rect 12440 23137 12449 23171
rect 12449 23137 12483 23171
rect 12483 23137 12492 23171
rect 12440 23128 12492 23137
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2964 22720 3016 22772
rect 1952 22627 2004 22636
rect 1952 22593 1961 22627
rect 1961 22593 1995 22627
rect 1995 22593 2004 22627
rect 1952 22584 2004 22593
rect 1676 22559 1728 22568
rect 1676 22525 1685 22559
rect 1685 22525 1719 22559
rect 1719 22525 1728 22559
rect 1676 22516 1728 22525
rect 2596 22423 2648 22432
rect 2596 22389 2605 22423
rect 2605 22389 2639 22423
rect 2639 22389 2648 22423
rect 2596 22380 2648 22389
rect 3700 22423 3752 22432
rect 3700 22389 3709 22423
rect 3709 22389 3743 22423
rect 3743 22389 3752 22423
rect 3700 22380 3752 22389
rect 12440 22380 12492 22432
rect 13360 22380 13412 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1400 22083 1452 22092
rect 1400 22049 1409 22083
rect 1409 22049 1443 22083
rect 1443 22049 1452 22083
rect 1400 22040 1452 22049
rect 2412 22040 2464 22092
rect 2688 21947 2740 21956
rect 2688 21913 2697 21947
rect 2697 21913 2731 21947
rect 2731 21913 2740 21947
rect 2688 21904 2740 21913
rect 1584 21879 1636 21888
rect 1584 21845 1593 21879
rect 1593 21845 1627 21879
rect 1627 21845 1636 21879
rect 1584 21836 1636 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1492 21632 1544 21684
rect 8576 21675 8628 21684
rect 8576 21641 8585 21675
rect 8585 21641 8619 21675
rect 8619 21641 8628 21675
rect 8576 21632 8628 21641
rect 2688 21607 2740 21616
rect 2688 21573 2697 21607
rect 2697 21573 2731 21607
rect 2731 21573 2740 21607
rect 2688 21564 2740 21573
rect 7288 21539 7340 21548
rect 7288 21505 7297 21539
rect 7297 21505 7331 21539
rect 7331 21505 7340 21539
rect 7288 21496 7340 21505
rect 1676 21428 1728 21480
rect 2044 21428 2096 21480
rect 2412 21403 2464 21412
rect 2412 21369 2421 21403
rect 2421 21369 2455 21403
rect 2455 21369 2464 21403
rect 2412 21360 2464 21369
rect 8760 21428 8812 21480
rect 1400 21292 1452 21344
rect 2504 21292 2556 21344
rect 7840 21335 7892 21344
rect 7840 21301 7849 21335
rect 7849 21301 7883 21335
rect 7883 21301 7892 21335
rect 7840 21292 7892 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1768 20995 1820 21004
rect 1768 20961 1777 20995
rect 1777 20961 1811 20995
rect 1811 20961 1820 20995
rect 1768 20952 1820 20961
rect 7932 20995 7984 21004
rect 7932 20961 7941 20995
rect 7941 20961 7975 20995
rect 7975 20961 7984 20995
rect 7932 20952 7984 20961
rect 1676 20927 1728 20936
rect 1676 20893 1685 20927
rect 1685 20893 1719 20927
rect 1719 20893 1728 20927
rect 1676 20884 1728 20893
rect 2688 20884 2740 20936
rect 8116 20927 8168 20936
rect 8116 20893 8125 20927
rect 8125 20893 8159 20927
rect 8159 20893 8168 20927
rect 8116 20884 8168 20893
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2596 20587 2648 20596
rect 2596 20553 2605 20587
rect 2605 20553 2639 20587
rect 2639 20553 2648 20587
rect 2596 20544 2648 20553
rect 4160 20544 4212 20596
rect 2044 20451 2096 20460
rect 2044 20417 2053 20451
rect 2053 20417 2087 20451
rect 2087 20417 2096 20451
rect 2044 20408 2096 20417
rect 8760 20451 8812 20460
rect 8760 20417 8769 20451
rect 8769 20417 8803 20451
rect 8803 20417 8812 20451
rect 8760 20408 8812 20417
rect 2596 20340 2648 20392
rect 2780 20340 2832 20392
rect 4160 20383 4212 20392
rect 4160 20349 4169 20383
rect 4169 20349 4203 20383
rect 4203 20349 4212 20383
rect 4160 20340 4212 20349
rect 1768 20204 1820 20256
rect 3240 20247 3292 20256
rect 3240 20213 3249 20247
rect 3249 20213 3283 20247
rect 3283 20213 3292 20247
rect 3240 20204 3292 20213
rect 7932 20247 7984 20256
rect 7932 20213 7941 20247
rect 7941 20213 7975 20247
rect 7975 20213 7984 20247
rect 7932 20204 7984 20213
rect 9404 20247 9456 20256
rect 9404 20213 9413 20247
rect 9413 20213 9447 20247
rect 9447 20213 9456 20247
rect 9404 20204 9456 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 4252 20043 4304 20052
rect 4252 20009 4261 20043
rect 4261 20009 4295 20043
rect 4295 20009 4304 20043
rect 4252 20000 4304 20009
rect 7380 19932 7432 19984
rect 1676 19864 1728 19916
rect 2964 19864 3016 19916
rect 4068 19907 4120 19916
rect 4068 19873 4077 19907
rect 4077 19873 4111 19907
rect 4111 19873 4120 19907
rect 4068 19864 4120 19873
rect 7656 19907 7708 19916
rect 7656 19873 7665 19907
rect 7665 19873 7699 19907
rect 7699 19873 7708 19907
rect 7656 19864 7708 19873
rect 4804 19796 4856 19848
rect 2872 19660 2924 19712
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 4068 19499 4120 19508
rect 4068 19465 4077 19499
rect 4077 19465 4111 19499
rect 4111 19465 4120 19499
rect 4068 19456 4120 19465
rect 2504 19320 2556 19372
rect 6920 19320 6972 19372
rect 7380 19363 7432 19372
rect 7380 19329 7389 19363
rect 7389 19329 7423 19363
rect 7423 19329 7432 19363
rect 7380 19320 7432 19329
rect 2688 19252 2740 19304
rect 1676 19159 1728 19168
rect 1676 19125 1685 19159
rect 1685 19125 1719 19159
rect 1719 19125 1728 19159
rect 1676 19116 1728 19125
rect 2688 19159 2740 19168
rect 2688 19125 2697 19159
rect 2697 19125 2731 19159
rect 2731 19125 2740 19159
rect 2688 19116 2740 19125
rect 4160 19252 4212 19304
rect 6460 19252 6512 19304
rect 11980 19252 12032 19304
rect 12992 19252 13044 19304
rect 3240 19116 3292 19168
rect 4620 19159 4672 19168
rect 4620 19125 4629 19159
rect 4629 19125 4663 19159
rect 4663 19125 4672 19159
rect 4620 19116 4672 19125
rect 6460 19116 6512 19168
rect 6828 19159 6880 19168
rect 6828 19125 6837 19159
rect 6837 19125 6871 19159
rect 6871 19125 6880 19159
rect 6828 19116 6880 19125
rect 7656 19116 7708 19168
rect 12164 19116 12216 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1492 18912 1544 18964
rect 4344 18912 4396 18964
rect 5540 18844 5592 18896
rect 10600 18844 10652 18896
rect 2596 18776 2648 18828
rect 3148 18776 3200 18828
rect 3700 18708 3752 18760
rect 1768 18640 1820 18692
rect 2964 18640 3016 18692
rect 4252 18683 4304 18692
rect 4252 18649 4261 18683
rect 4261 18649 4295 18683
rect 4295 18649 4304 18683
rect 4252 18640 4304 18649
rect 2320 18615 2372 18624
rect 2320 18581 2329 18615
rect 2329 18581 2363 18615
rect 2363 18581 2372 18615
rect 2320 18572 2372 18581
rect 3056 18615 3108 18624
rect 3056 18581 3065 18615
rect 3065 18581 3099 18615
rect 3099 18581 3108 18615
rect 3056 18572 3108 18581
rect 3884 18615 3936 18624
rect 3884 18581 3893 18615
rect 3893 18581 3927 18615
rect 3927 18581 3936 18615
rect 8024 18708 8076 18760
rect 3884 18572 3936 18581
rect 6736 18615 6788 18624
rect 6736 18581 6745 18615
rect 6745 18581 6779 18615
rect 6779 18581 6788 18615
rect 6736 18572 6788 18581
rect 8208 18572 8260 18624
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9312 18572 9364 18581
rect 11796 18615 11848 18624
rect 11796 18581 11805 18615
rect 11805 18581 11839 18615
rect 11839 18581 11848 18615
rect 11796 18572 11848 18581
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 3700 18411 3752 18420
rect 3700 18377 3709 18411
rect 3709 18377 3743 18411
rect 3743 18377 3752 18411
rect 3700 18368 3752 18377
rect 7656 18411 7708 18420
rect 7656 18377 7665 18411
rect 7665 18377 7699 18411
rect 7699 18377 7708 18411
rect 7656 18368 7708 18377
rect 12164 18411 12216 18420
rect 12164 18377 12173 18411
rect 12173 18377 12207 18411
rect 12207 18377 12216 18411
rect 12164 18368 12216 18377
rect 10600 18343 10652 18352
rect 10600 18309 10609 18343
rect 10609 18309 10643 18343
rect 10643 18309 10652 18343
rect 10600 18300 10652 18309
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 2596 18232 2648 18284
rect 4160 18232 4212 18284
rect 8208 18275 8260 18284
rect 8208 18241 8217 18275
rect 8217 18241 8251 18275
rect 8251 18241 8260 18275
rect 8208 18232 8260 18241
rect 12532 18232 12584 18284
rect 1492 18207 1544 18216
rect 1492 18173 1501 18207
rect 1501 18173 1535 18207
rect 1535 18173 1544 18207
rect 1492 18164 1544 18173
rect 3884 18164 3936 18216
rect 4252 18207 4304 18216
rect 4252 18173 4261 18207
rect 4261 18173 4295 18207
rect 4295 18173 4304 18207
rect 4252 18164 4304 18173
rect 8024 18207 8076 18216
rect 8024 18173 8033 18207
rect 8033 18173 8067 18207
rect 8067 18173 8076 18207
rect 8024 18164 8076 18173
rect 9312 18164 9364 18216
rect 12164 18164 12216 18216
rect 4988 18096 5040 18148
rect 9772 18096 9824 18148
rect 2688 18071 2740 18080
rect 2688 18037 2697 18071
rect 2697 18037 2731 18071
rect 2731 18037 2740 18071
rect 2688 18028 2740 18037
rect 5540 18028 5592 18080
rect 8116 18071 8168 18080
rect 8116 18037 8125 18071
rect 8125 18037 8159 18071
rect 8159 18037 8168 18071
rect 8116 18028 8168 18037
rect 11152 18028 11204 18080
rect 12440 18071 12492 18080
rect 12440 18037 12449 18071
rect 12449 18037 12483 18071
rect 12483 18037 12492 18071
rect 12440 18028 12492 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1860 17824 1912 17876
rect 2320 17824 2372 17876
rect 7380 17824 7432 17876
rect 7840 17824 7892 17876
rect 8024 17824 8076 17876
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 12532 17824 12584 17876
rect 6736 17756 6788 17808
rect 9772 17756 9824 17808
rect 2504 17688 2556 17740
rect 4620 17688 4672 17740
rect 5356 17688 5408 17740
rect 8760 17688 8812 17740
rect 2136 17620 2188 17672
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 10140 17663 10192 17672
rect 6000 17552 6052 17604
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 11796 17756 11848 17808
rect 10692 17620 10744 17672
rect 11336 17663 11388 17672
rect 9312 17552 9364 17604
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 1952 17484 2004 17536
rect 2688 17484 2740 17536
rect 3148 17484 3200 17536
rect 3424 17484 3476 17536
rect 4252 17527 4304 17536
rect 4252 17493 4261 17527
rect 4261 17493 4295 17527
rect 4295 17493 4304 17527
rect 4252 17484 4304 17493
rect 4436 17527 4488 17536
rect 4436 17493 4445 17527
rect 4445 17493 4479 17527
rect 4479 17493 4488 17527
rect 4436 17484 4488 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 4988 17280 5040 17332
rect 6736 17280 6788 17332
rect 10048 17280 10100 17332
rect 10692 17323 10744 17332
rect 10692 17289 10701 17323
rect 10701 17289 10735 17323
rect 10735 17289 10744 17323
rect 10692 17280 10744 17289
rect 11796 17280 11848 17332
rect 12440 17280 12492 17332
rect 3332 17212 3384 17264
rect 2136 17144 2188 17196
rect 6000 17144 6052 17196
rect 6828 17187 6880 17196
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 9312 17187 9364 17196
rect 9312 17153 9321 17187
rect 9321 17153 9355 17187
rect 9355 17153 9364 17187
rect 9312 17144 9364 17153
rect 3424 17076 3476 17128
rect 11336 17076 11388 17128
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 7380 17008 7432 17060
rect 9588 17051 9640 17060
rect 9588 17017 9622 17051
rect 9622 17017 9640 17051
rect 9588 17008 9640 17017
rect 12532 17008 12584 17060
rect 1676 16983 1728 16992
rect 1676 16949 1685 16983
rect 1685 16949 1719 16983
rect 1719 16949 1728 16983
rect 1676 16940 1728 16949
rect 1768 16940 1820 16992
rect 2136 16983 2188 16992
rect 2136 16949 2145 16983
rect 2145 16949 2179 16983
rect 2179 16949 2188 16983
rect 2136 16940 2188 16949
rect 2320 16940 2372 16992
rect 2504 16940 2556 16992
rect 3148 16983 3200 16992
rect 3148 16949 3157 16983
rect 3157 16949 3191 16983
rect 3191 16949 3200 16983
rect 3148 16940 3200 16949
rect 5356 16983 5408 16992
rect 5356 16949 5365 16983
rect 5365 16949 5399 16983
rect 5399 16949 5408 16983
rect 5356 16940 5408 16949
rect 7748 16940 7800 16992
rect 8760 16983 8812 16992
rect 8760 16949 8769 16983
rect 8769 16949 8803 16983
rect 8803 16949 8812 16983
rect 8760 16940 8812 16949
rect 13820 16983 13872 16992
rect 13820 16949 13829 16983
rect 13829 16949 13863 16983
rect 13863 16949 13872 16983
rect 13820 16940 13872 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1768 16736 1820 16788
rect 2044 16736 2096 16788
rect 2780 16736 2832 16788
rect 4068 16779 4120 16788
rect 4068 16745 4077 16779
rect 4077 16745 4111 16779
rect 4111 16745 4120 16779
rect 4068 16736 4120 16745
rect 4436 16736 4488 16788
rect 4620 16736 4672 16788
rect 5264 16736 5316 16788
rect 6000 16736 6052 16788
rect 6460 16779 6512 16788
rect 6460 16745 6469 16779
rect 6469 16745 6503 16779
rect 6503 16745 6512 16779
rect 6460 16736 6512 16745
rect 6828 16736 6880 16788
rect 8024 16779 8076 16788
rect 2596 16668 2648 16720
rect 3792 16711 3844 16720
rect 2412 16600 2464 16652
rect 3792 16677 3801 16711
rect 3801 16677 3835 16711
rect 3835 16677 3844 16711
rect 3792 16668 3844 16677
rect 4068 16600 4120 16652
rect 6920 16668 6972 16720
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 4804 16600 4856 16652
rect 5540 16643 5592 16652
rect 5540 16609 5549 16643
rect 5549 16609 5583 16643
rect 5583 16609 5592 16643
rect 5540 16600 5592 16609
rect 6644 16600 6696 16652
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 10692 16736 10744 16788
rect 11152 16779 11204 16788
rect 11152 16745 11161 16779
rect 11161 16745 11195 16779
rect 11195 16745 11204 16779
rect 11152 16736 11204 16745
rect 8300 16668 8352 16720
rect 11336 16668 11388 16720
rect 2320 16532 2372 16584
rect 3148 16532 3200 16584
rect 5448 16532 5500 16584
rect 6552 16532 6604 16584
rect 8484 16643 8536 16652
rect 8484 16609 8493 16643
rect 8493 16609 8527 16643
rect 8527 16609 8536 16643
rect 11520 16643 11572 16652
rect 8484 16600 8536 16609
rect 11520 16609 11529 16643
rect 11529 16609 11563 16643
rect 11563 16609 11572 16643
rect 11520 16600 11572 16609
rect 6736 16464 6788 16516
rect 8392 16532 8444 16584
rect 8668 16575 8720 16584
rect 8668 16541 8677 16575
rect 8677 16541 8711 16575
rect 8711 16541 8720 16575
rect 11612 16575 11664 16584
rect 8668 16532 8720 16541
rect 7472 16439 7524 16448
rect 7472 16405 7481 16439
rect 7481 16405 7515 16439
rect 7515 16405 7524 16439
rect 7472 16396 7524 16405
rect 11612 16541 11621 16575
rect 11621 16541 11655 16575
rect 11655 16541 11664 16575
rect 11612 16532 11664 16541
rect 11796 16575 11848 16584
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 9588 16396 9640 16448
rect 10600 16396 10652 16448
rect 12440 16396 12492 16448
rect 12624 16396 12676 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2412 16235 2464 16244
rect 2412 16201 2421 16235
rect 2421 16201 2455 16235
rect 2455 16201 2464 16235
rect 2412 16192 2464 16201
rect 4436 16192 4488 16244
rect 5448 16192 5500 16244
rect 6828 16235 6880 16244
rect 6828 16201 6837 16235
rect 6837 16201 6871 16235
rect 6871 16201 6880 16235
rect 6828 16192 6880 16201
rect 8300 16235 8352 16244
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 8300 16192 8352 16201
rect 8668 16235 8720 16244
rect 8668 16201 8677 16235
rect 8677 16201 8711 16235
rect 8711 16201 8720 16235
rect 8668 16192 8720 16201
rect 10600 16235 10652 16244
rect 10600 16201 10609 16235
rect 10609 16201 10643 16235
rect 10643 16201 10652 16235
rect 10600 16192 10652 16201
rect 11520 16235 11572 16244
rect 11520 16201 11529 16235
rect 11529 16201 11563 16235
rect 11563 16201 11572 16235
rect 11520 16192 11572 16201
rect 11796 16192 11848 16244
rect 6920 16056 6972 16108
rect 7472 16099 7524 16108
rect 7472 16065 7481 16099
rect 7481 16065 7515 16099
rect 7515 16065 7524 16099
rect 7472 16056 7524 16065
rect 9128 16056 9180 16108
rect 1584 15988 1636 16040
rect 3424 15988 3476 16040
rect 5540 15988 5592 16040
rect 2412 15920 2464 15972
rect 3056 15920 3108 15972
rect 5448 15963 5500 15972
rect 5448 15929 5457 15963
rect 5457 15929 5491 15963
rect 5491 15929 5500 15963
rect 5448 15920 5500 15929
rect 7196 15963 7248 15972
rect 7196 15929 7205 15963
rect 7205 15929 7239 15963
rect 7239 15929 7248 15963
rect 7196 15920 7248 15929
rect 10140 15920 10192 15972
rect 3148 15852 3200 15904
rect 6092 15895 6144 15904
rect 6092 15861 6101 15895
rect 6101 15861 6135 15895
rect 6135 15861 6144 15895
rect 6092 15852 6144 15861
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 11520 15852 11572 15904
rect 11980 15852 12032 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1400 15691 1452 15700
rect 1400 15657 1409 15691
rect 1409 15657 1443 15691
rect 1443 15657 1452 15691
rect 1400 15648 1452 15657
rect 2320 15691 2372 15700
rect 2320 15657 2329 15691
rect 2329 15657 2363 15691
rect 2363 15657 2372 15691
rect 2320 15648 2372 15657
rect 2596 15648 2648 15700
rect 4068 15648 4120 15700
rect 6736 15648 6788 15700
rect 6920 15648 6972 15700
rect 8484 15648 8536 15700
rect 10784 15648 10836 15700
rect 11980 15691 12032 15700
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 12716 15691 12768 15700
rect 12716 15657 12725 15691
rect 12725 15657 12759 15691
rect 12759 15657 12768 15691
rect 12716 15648 12768 15657
rect 13728 15648 13780 15700
rect 4252 15580 4304 15632
rect 2780 15555 2832 15564
rect 2780 15521 2789 15555
rect 2789 15521 2823 15555
rect 2823 15521 2832 15555
rect 2780 15512 2832 15521
rect 2872 15487 2924 15496
rect 2872 15453 2881 15487
rect 2881 15453 2915 15487
rect 2915 15453 2924 15487
rect 2872 15444 2924 15453
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 4068 15487 4120 15496
rect 3056 15444 3108 15453
rect 2596 15308 2648 15360
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 7380 15512 7432 15564
rect 9956 15512 10008 15564
rect 11428 15555 11480 15564
rect 11428 15521 11437 15555
rect 11437 15521 11471 15555
rect 11471 15521 11480 15555
rect 11428 15512 11480 15521
rect 7564 15487 7616 15496
rect 7564 15453 7573 15487
rect 7573 15453 7607 15487
rect 7607 15453 7616 15487
rect 7564 15444 7616 15453
rect 7748 15487 7800 15496
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 12072 15487 12124 15496
rect 10232 15444 10284 15453
rect 12072 15453 12081 15487
rect 12081 15453 12115 15487
rect 12115 15453 12124 15487
rect 12072 15444 12124 15453
rect 12256 15487 12308 15496
rect 12256 15453 12265 15487
rect 12265 15453 12299 15487
rect 12299 15453 12308 15487
rect 12256 15444 12308 15453
rect 8944 15376 8996 15428
rect 6828 15351 6880 15360
rect 6828 15317 6837 15351
rect 6837 15317 6871 15351
rect 6871 15317 6880 15351
rect 6828 15308 6880 15317
rect 8484 15351 8536 15360
rect 8484 15317 8493 15351
rect 8493 15317 8527 15351
rect 8527 15317 8536 15351
rect 8484 15308 8536 15317
rect 9128 15308 9180 15360
rect 9496 15308 9548 15360
rect 12624 15308 12676 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2504 15104 2556 15156
rect 2688 14968 2740 15020
rect 4252 15104 4304 15156
rect 6276 15147 6328 15156
rect 6276 15113 6285 15147
rect 6285 15113 6319 15147
rect 6319 15113 6328 15147
rect 6276 15104 6328 15113
rect 7472 15104 7524 15156
rect 10232 15104 10284 15156
rect 11980 15104 12032 15156
rect 4160 14968 4212 15020
rect 9220 15011 9272 15020
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 9220 14977 9229 15011
rect 9229 14977 9263 15011
rect 9263 14977 9272 15011
rect 9220 14968 9272 14977
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 9128 14900 9180 14952
rect 12716 14943 12768 14952
rect 12716 14909 12750 14943
rect 12750 14909 12768 14943
rect 2780 14832 2832 14884
rect 4528 14875 4580 14884
rect 4528 14841 4562 14875
rect 4562 14841 4580 14875
rect 2504 14807 2556 14816
rect 2504 14773 2513 14807
rect 2513 14773 2547 14807
rect 2547 14773 2556 14807
rect 2504 14764 2556 14773
rect 2964 14764 3016 14816
rect 4528 14832 4580 14841
rect 6736 14832 6788 14884
rect 7748 14832 7800 14884
rect 8392 14832 8444 14884
rect 9496 14832 9548 14884
rect 12716 14900 12768 14909
rect 12624 14832 12676 14884
rect 4896 14764 4948 14816
rect 6644 14807 6696 14816
rect 6644 14773 6653 14807
rect 6653 14773 6687 14807
rect 6687 14773 6696 14807
rect 6644 14764 6696 14773
rect 8852 14807 8904 14816
rect 8852 14773 8861 14807
rect 8861 14773 8895 14807
rect 8895 14773 8904 14807
rect 8852 14764 8904 14773
rect 9956 14764 10008 14816
rect 12256 14764 12308 14816
rect 12808 14764 12860 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1400 14560 1452 14612
rect 4896 14603 4948 14612
rect 4896 14569 4905 14603
rect 4905 14569 4939 14603
rect 4939 14569 4948 14603
rect 4896 14560 4948 14569
rect 6736 14560 6788 14612
rect 8484 14560 8536 14612
rect 11152 14603 11204 14612
rect 11152 14569 11161 14603
rect 11161 14569 11195 14603
rect 11195 14569 11204 14603
rect 11152 14560 11204 14569
rect 12072 14560 12124 14612
rect 12624 14560 12676 14612
rect 1952 14535 2004 14544
rect 1952 14501 1961 14535
rect 1961 14501 1995 14535
rect 1995 14501 2004 14535
rect 1952 14492 2004 14501
rect 2320 14492 2372 14544
rect 3056 14492 3108 14544
rect 7472 14492 7524 14544
rect 8944 14492 8996 14544
rect 1676 14424 1728 14476
rect 5264 14467 5316 14476
rect 5264 14433 5273 14467
rect 5273 14433 5307 14467
rect 5307 14433 5316 14467
rect 5264 14424 5316 14433
rect 6828 14424 6880 14476
rect 9036 14424 9088 14476
rect 10048 14467 10100 14476
rect 10048 14433 10082 14467
rect 10082 14433 10100 14467
rect 10048 14424 10100 14433
rect 11428 14424 11480 14476
rect 12808 14492 12860 14544
rect 13452 14424 13504 14476
rect 3240 14356 3292 14408
rect 5356 14399 5408 14408
rect 5356 14365 5365 14399
rect 5365 14365 5399 14399
rect 5399 14365 5408 14399
rect 5356 14356 5408 14365
rect 2412 14288 2464 14340
rect 4528 14288 4580 14340
rect 6184 14356 6236 14408
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9772 14399 9824 14408
rect 9128 14356 9180 14365
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 8944 14288 8996 14340
rect 1400 14220 1452 14272
rect 2964 14220 3016 14272
rect 7748 14220 7800 14272
rect 13912 14220 13964 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1860 14059 1912 14068
rect 1860 14025 1869 14059
rect 1869 14025 1903 14059
rect 1903 14025 1912 14059
rect 1860 14016 1912 14025
rect 3240 14059 3292 14068
rect 3240 14025 3249 14059
rect 3249 14025 3283 14059
rect 3283 14025 3292 14059
rect 3240 14016 3292 14025
rect 4344 14016 4396 14068
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 7012 14059 7064 14068
rect 7012 14025 7021 14059
rect 7021 14025 7055 14059
rect 7055 14025 7064 14059
rect 7012 14016 7064 14025
rect 7472 14059 7524 14068
rect 7472 14025 7481 14059
rect 7481 14025 7515 14059
rect 7515 14025 7524 14059
rect 7472 14016 7524 14025
rect 7932 14059 7984 14068
rect 7932 14025 7941 14059
rect 7941 14025 7975 14059
rect 7975 14025 7984 14059
rect 7932 14016 7984 14025
rect 9036 14016 9088 14068
rect 12072 14016 12124 14068
rect 13452 14059 13504 14068
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 4804 13948 4856 14000
rect 6276 13948 6328 14000
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 2688 13880 2740 13932
rect 5080 13880 5132 13932
rect 4068 13812 4120 13864
rect 5264 13880 5316 13932
rect 5724 13923 5776 13932
rect 5724 13889 5733 13923
rect 5733 13889 5767 13923
rect 5767 13889 5776 13923
rect 5724 13880 5776 13889
rect 8392 13880 8444 13932
rect 8944 13923 8996 13932
rect 8944 13889 8953 13923
rect 8953 13889 8987 13923
rect 8987 13889 8996 13923
rect 8944 13880 8996 13889
rect 11428 13948 11480 14000
rect 12256 13948 12308 14000
rect 24860 13948 24912 14000
rect 10048 13880 10100 13932
rect 5356 13855 5408 13864
rect 5356 13821 5365 13855
rect 5365 13821 5399 13855
rect 5399 13821 5408 13855
rect 5356 13812 5408 13821
rect 6552 13812 6604 13864
rect 4620 13719 4672 13728
rect 4620 13685 4629 13719
rect 4629 13685 4663 13719
rect 4663 13685 4672 13719
rect 4620 13676 4672 13685
rect 4712 13719 4764 13728
rect 4712 13685 4721 13719
rect 4721 13685 4755 13719
rect 4755 13685 4764 13719
rect 4712 13676 4764 13685
rect 6184 13676 6236 13728
rect 8300 13719 8352 13728
rect 8300 13685 8309 13719
rect 8309 13685 8343 13719
rect 8343 13685 8352 13719
rect 8300 13676 8352 13685
rect 9496 13719 9548 13728
rect 9496 13685 9505 13719
rect 9505 13685 9539 13719
rect 9539 13685 9548 13719
rect 9496 13676 9548 13685
rect 12716 13880 12768 13932
rect 13452 13812 13504 13864
rect 24032 13855 24084 13864
rect 24032 13821 24041 13855
rect 24041 13821 24075 13855
rect 24075 13821 24084 13855
rect 24032 13812 24084 13821
rect 12440 13744 12492 13796
rect 10692 13676 10744 13728
rect 11060 13719 11112 13728
rect 11060 13685 11069 13719
rect 11069 13685 11103 13719
rect 11103 13685 11112 13719
rect 11060 13676 11112 13685
rect 13728 13676 13780 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 3240 13472 3292 13524
rect 4712 13472 4764 13524
rect 6184 13515 6236 13524
rect 6184 13481 6193 13515
rect 6193 13481 6227 13515
rect 6227 13481 6236 13515
rect 6184 13472 6236 13481
rect 7288 13515 7340 13524
rect 7288 13481 7297 13515
rect 7297 13481 7331 13515
rect 7331 13481 7340 13515
rect 7288 13472 7340 13481
rect 8392 13515 8444 13524
rect 8392 13481 8401 13515
rect 8401 13481 8435 13515
rect 8435 13481 8444 13515
rect 8392 13472 8444 13481
rect 9496 13472 9548 13524
rect 10692 13472 10744 13524
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 12716 13472 12768 13524
rect 13360 13515 13412 13524
rect 13360 13481 13369 13515
rect 13369 13481 13403 13515
rect 13403 13481 13412 13515
rect 13360 13472 13412 13481
rect 2044 13404 2096 13456
rect 2412 13404 2464 13456
rect 2504 13336 2556 13388
rect 4896 13336 4948 13388
rect 5080 13379 5132 13388
rect 5080 13345 5114 13379
rect 5114 13345 5132 13379
rect 5080 13336 5132 13345
rect 5356 13336 5408 13388
rect 6552 13336 6604 13388
rect 8208 13336 8260 13388
rect 10324 13379 10376 13388
rect 10324 13345 10358 13379
rect 10358 13345 10376 13379
rect 10324 13336 10376 13345
rect 12900 13336 12952 13388
rect 13728 13379 13780 13388
rect 13728 13345 13737 13379
rect 13737 13345 13771 13379
rect 13771 13345 13780 13379
rect 13728 13336 13780 13345
rect 15844 13336 15896 13388
rect 23388 13379 23440 13388
rect 23388 13345 23397 13379
rect 23397 13345 23431 13379
rect 23431 13345 23440 13379
rect 23388 13336 23440 13345
rect 1492 13311 1544 13320
rect 1492 13277 1501 13311
rect 1501 13277 1535 13311
rect 1535 13277 1544 13311
rect 1492 13268 1544 13277
rect 4712 13268 4764 13320
rect 7932 13311 7984 13320
rect 7656 13200 7708 13252
rect 7932 13277 7941 13311
rect 7941 13277 7975 13311
rect 7975 13277 7984 13311
rect 7932 13268 7984 13277
rect 9772 13268 9824 13320
rect 13820 13311 13872 13320
rect 4620 13175 4672 13184
rect 4620 13141 4629 13175
rect 4629 13141 4663 13175
rect 4663 13141 4672 13175
rect 4620 13132 4672 13141
rect 6920 13175 6972 13184
rect 6920 13141 6929 13175
rect 6929 13141 6963 13175
rect 6963 13141 6972 13175
rect 6920 13132 6972 13141
rect 8576 13132 8628 13184
rect 9496 13175 9548 13184
rect 9496 13141 9505 13175
rect 9505 13141 9539 13175
rect 9539 13141 9548 13175
rect 9496 13132 9548 13141
rect 13820 13277 13829 13311
rect 13829 13277 13863 13311
rect 13863 13277 13872 13311
rect 13820 13268 13872 13277
rect 14004 13311 14056 13320
rect 14004 13277 14013 13311
rect 14013 13277 14047 13311
rect 14047 13277 14056 13311
rect 14004 13268 14056 13277
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 16672 13243 16724 13252
rect 16672 13209 16681 13243
rect 16681 13209 16715 13243
rect 16715 13209 16724 13243
rect 16672 13200 16724 13209
rect 11888 13132 11940 13184
rect 13176 13175 13228 13184
rect 13176 13141 13185 13175
rect 13185 13141 13219 13175
rect 13219 13141 13228 13175
rect 13176 13132 13228 13141
rect 24952 13132 25004 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1860 12971 1912 12980
rect 1860 12937 1869 12971
rect 1869 12937 1903 12971
rect 1903 12937 1912 12971
rect 1860 12928 1912 12937
rect 3240 12971 3292 12980
rect 3240 12937 3249 12971
rect 3249 12937 3283 12971
rect 3283 12937 3292 12971
rect 3240 12928 3292 12937
rect 5540 12928 5592 12980
rect 7932 12928 7984 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 12900 12971 12952 12980
rect 12900 12937 12909 12971
rect 12909 12937 12943 12971
rect 12943 12937 12952 12971
rect 12900 12928 12952 12937
rect 13268 12971 13320 12980
rect 13268 12937 13277 12971
rect 13277 12937 13311 12971
rect 13311 12937 13320 12971
rect 13268 12928 13320 12937
rect 15292 12928 15344 12980
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 4896 12860 4948 12912
rect 25044 12860 25096 12912
rect 6552 12835 6604 12844
rect 1492 12724 1544 12776
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 7196 12792 7248 12844
rect 10324 12792 10376 12844
rect 2964 12699 3016 12708
rect 2964 12665 2973 12699
rect 2973 12665 3007 12699
rect 3007 12665 3016 12699
rect 2964 12656 3016 12665
rect 9496 12724 9548 12776
rect 9680 12724 9732 12776
rect 4620 12656 4672 12708
rect 6184 12656 6236 12708
rect 7104 12656 7156 12708
rect 12716 12724 12768 12776
rect 13176 12724 13228 12776
rect 23664 12767 23716 12776
rect 23664 12733 23673 12767
rect 23673 12733 23707 12767
rect 23707 12733 23716 12767
rect 23664 12724 23716 12733
rect 10968 12656 11020 12708
rect 13636 12699 13688 12708
rect 13636 12665 13670 12699
rect 13670 12665 13688 12699
rect 13636 12656 13688 12665
rect 4160 12588 4212 12640
rect 5080 12588 5132 12640
rect 5540 12588 5592 12640
rect 6920 12588 6972 12640
rect 7656 12588 7708 12640
rect 8392 12631 8444 12640
rect 8392 12597 8401 12631
rect 8401 12597 8435 12631
rect 8435 12597 8444 12631
rect 8392 12588 8444 12597
rect 8576 12588 8628 12640
rect 9864 12631 9916 12640
rect 9864 12597 9873 12631
rect 9873 12597 9907 12631
rect 9907 12597 9916 12631
rect 9864 12588 9916 12597
rect 10784 12631 10836 12640
rect 10784 12597 10793 12631
rect 10793 12597 10827 12631
rect 10827 12597 10836 12631
rect 10784 12588 10836 12597
rect 11336 12631 11388 12640
rect 11336 12597 11345 12631
rect 11345 12597 11379 12631
rect 11379 12597 11388 12631
rect 11336 12588 11388 12597
rect 15844 12656 15896 12708
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2044 12384 2096 12436
rect 5540 12384 5592 12436
rect 7104 12427 7156 12436
rect 7104 12393 7113 12427
rect 7113 12393 7147 12427
rect 7147 12393 7156 12427
rect 7104 12384 7156 12393
rect 11060 12384 11112 12436
rect 12992 12384 13044 12436
rect 4896 12359 4948 12368
rect 4896 12325 4930 12359
rect 4930 12325 4948 12359
rect 4896 12316 4948 12325
rect 2596 12248 2648 12300
rect 4620 12291 4672 12300
rect 4620 12257 4629 12291
rect 4629 12257 4663 12291
rect 4663 12257 4672 12291
rect 4620 12248 4672 12257
rect 6368 12248 6420 12300
rect 8208 12248 8260 12300
rect 9036 12248 9088 12300
rect 10784 12316 10836 12368
rect 12716 12316 12768 12368
rect 11152 12248 11204 12300
rect 12164 12248 12216 12300
rect 13636 12248 13688 12300
rect 14372 12248 14424 12300
rect 22284 12291 22336 12300
rect 22284 12257 22293 12291
rect 22293 12257 22327 12291
rect 22327 12257 22336 12291
rect 22284 12248 22336 12257
rect 1492 12223 1544 12232
rect 1492 12189 1501 12223
rect 1501 12189 1535 12223
rect 1535 12189 1544 12223
rect 1492 12180 1544 12189
rect 7012 12180 7064 12232
rect 10324 12223 10376 12232
rect 7196 12112 7248 12164
rect 7472 12112 7524 12164
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 12808 12180 12860 12232
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 13820 12180 13872 12232
rect 15476 12180 15528 12232
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 8576 12155 8628 12164
rect 1768 12044 1820 12096
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 4344 12087 4396 12096
rect 4344 12053 4353 12087
rect 4353 12053 4387 12087
rect 4387 12053 4396 12087
rect 4344 12044 4396 12053
rect 6736 12044 6788 12096
rect 8576 12121 8585 12155
rect 8585 12121 8619 12155
rect 8619 12121 8628 12155
rect 8576 12112 8628 12121
rect 9588 12112 9640 12164
rect 8668 12087 8720 12096
rect 8668 12053 8677 12087
rect 8677 12053 8711 12087
rect 8711 12053 8720 12087
rect 8668 12044 8720 12053
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 22468 12087 22520 12096
rect 22468 12053 22477 12087
rect 22477 12053 22511 12087
rect 22511 12053 22520 12087
rect 22468 12044 22520 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2596 11883 2648 11892
rect 2596 11849 2605 11883
rect 2605 11849 2639 11883
rect 2639 11849 2648 11883
rect 2964 11883 3016 11892
rect 2596 11840 2648 11849
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 4896 11883 4948 11892
rect 4896 11849 4905 11883
rect 4905 11849 4939 11883
rect 4939 11849 4948 11883
rect 4896 11840 4948 11849
rect 5540 11883 5592 11892
rect 5540 11849 5549 11883
rect 5549 11849 5583 11883
rect 5583 11849 5592 11883
rect 5540 11840 5592 11849
rect 6368 11883 6420 11892
rect 6368 11849 6377 11883
rect 6377 11849 6411 11883
rect 6411 11849 6420 11883
rect 6368 11840 6420 11849
rect 3424 11772 3476 11824
rect 4068 11772 4120 11824
rect 6184 11772 6236 11824
rect 6736 11772 6788 11824
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 3884 11704 3936 11756
rect 4620 11704 4672 11756
rect 10324 11840 10376 11892
rect 11336 11840 11388 11892
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 13360 11840 13412 11892
rect 15384 11840 15436 11892
rect 22284 11883 22336 11892
rect 22284 11849 22293 11883
rect 22293 11849 22327 11883
rect 22327 11849 22336 11883
rect 22284 11840 22336 11849
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 1952 11636 2004 11645
rect 3976 11636 4028 11688
rect 5172 11636 5224 11688
rect 5448 11636 5500 11688
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 7104 11611 7156 11620
rect 1492 11500 1544 11552
rect 2504 11500 2556 11552
rect 3792 11543 3844 11552
rect 3792 11509 3801 11543
rect 3801 11509 3835 11543
rect 3835 11509 3844 11543
rect 3792 11500 3844 11509
rect 7104 11577 7138 11611
rect 7138 11577 7156 11611
rect 7104 11568 7156 11577
rect 7472 11568 7524 11620
rect 4988 11500 5040 11552
rect 8024 11500 8076 11552
rect 8484 11500 8536 11552
rect 15752 11747 15804 11756
rect 9588 11679 9640 11688
rect 9588 11645 9597 11679
rect 9597 11645 9631 11679
rect 9631 11645 9640 11679
rect 9588 11636 9640 11645
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 13728 11636 13780 11688
rect 15568 11679 15620 11688
rect 15568 11645 15577 11679
rect 15577 11645 15611 11679
rect 15611 11645 15620 11679
rect 15568 11636 15620 11645
rect 9956 11611 10008 11620
rect 9956 11577 9990 11611
rect 9990 11577 10008 11611
rect 9956 11568 10008 11577
rect 14464 11568 14516 11620
rect 14556 11568 14608 11620
rect 15476 11568 15528 11620
rect 11152 11500 11204 11552
rect 14372 11500 14424 11552
rect 15660 11543 15712 11552
rect 15660 11509 15669 11543
rect 15669 11509 15703 11543
rect 15703 11509 15712 11543
rect 15660 11500 15712 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 2136 11296 2188 11348
rect 2228 11296 2280 11348
rect 2504 11296 2556 11348
rect 4068 11296 4120 11348
rect 4436 11296 4488 11348
rect 5816 11339 5868 11348
rect 5816 11305 5825 11339
rect 5825 11305 5859 11339
rect 5859 11305 5868 11339
rect 5816 11296 5868 11305
rect 9680 11339 9732 11348
rect 9680 11305 9689 11339
rect 9689 11305 9723 11339
rect 9723 11305 9732 11339
rect 9680 11296 9732 11305
rect 11060 11339 11112 11348
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 12808 11339 12860 11348
rect 12808 11305 12817 11339
rect 12817 11305 12851 11339
rect 12851 11305 12860 11339
rect 12808 11296 12860 11305
rect 14004 11339 14056 11348
rect 14004 11305 14013 11339
rect 14013 11305 14047 11339
rect 14047 11305 14056 11339
rect 14004 11296 14056 11305
rect 14464 11339 14516 11348
rect 14464 11305 14473 11339
rect 14473 11305 14507 11339
rect 14507 11305 14516 11339
rect 14464 11296 14516 11305
rect 15568 11339 15620 11348
rect 15568 11305 15577 11339
rect 15577 11305 15611 11339
rect 15611 11305 15620 11339
rect 15568 11296 15620 11305
rect 15844 11339 15896 11348
rect 15844 11305 15853 11339
rect 15853 11305 15887 11339
rect 15887 11305 15896 11339
rect 15844 11296 15896 11305
rect 3976 11228 4028 11280
rect 7104 11228 7156 11280
rect 8024 11228 8076 11280
rect 13360 11228 13412 11280
rect 3424 11160 3476 11212
rect 4160 11160 4212 11212
rect 5356 11160 5408 11212
rect 6000 11160 6052 11212
rect 6828 11160 6880 11212
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 4620 11135 4672 11144
rect 2964 11092 3016 11101
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 5448 11092 5500 11144
rect 8484 11160 8536 11212
rect 10784 11160 10836 11212
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 12440 11160 12492 11212
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 11704 11135 11756 11144
rect 2044 10956 2096 11008
rect 7012 11024 7064 11076
rect 9036 11067 9088 11076
rect 9036 11033 9045 11067
rect 9045 11033 9079 11067
rect 9079 11033 9088 11067
rect 9036 11024 9088 11033
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 11704 11092 11756 11101
rect 11152 11024 11204 11076
rect 13360 11092 13412 11144
rect 13728 11092 13780 11144
rect 13912 11067 13964 11076
rect 13912 11033 13921 11067
rect 13921 11033 13955 11067
rect 13955 11033 13964 11067
rect 13912 11024 13964 11033
rect 4712 10956 4764 11008
rect 5080 10999 5132 11008
rect 5080 10965 5089 10999
rect 5089 10965 5123 10999
rect 5123 10965 5132 10999
rect 5080 10956 5132 10965
rect 5448 10999 5500 11008
rect 5448 10965 5457 10999
rect 5457 10965 5491 10999
rect 5491 10965 5500 10999
rect 5448 10956 5500 10965
rect 8760 10956 8812 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2688 10752 2740 10804
rect 2964 10752 3016 10804
rect 3424 10752 3476 10804
rect 5540 10752 5592 10804
rect 6920 10795 6972 10804
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 6920 10752 6972 10761
rect 9956 10752 10008 10804
rect 10140 10752 10192 10804
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 5264 10684 5316 10736
rect 5080 10616 5132 10668
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 11612 10752 11664 10804
rect 1768 10591 1820 10600
rect 1768 10557 1777 10591
rect 1777 10557 1811 10591
rect 1811 10557 1820 10591
rect 1768 10548 1820 10557
rect 2320 10548 2372 10600
rect 4712 10591 4764 10600
rect 4712 10557 4721 10591
rect 4721 10557 4755 10591
rect 4755 10557 4764 10591
rect 4712 10548 4764 10557
rect 5448 10548 5500 10600
rect 8484 10591 8536 10600
rect 8484 10557 8493 10591
rect 8493 10557 8527 10591
rect 8527 10557 8536 10591
rect 8484 10548 8536 10557
rect 13728 10548 13780 10600
rect 2044 10523 2096 10532
rect 2044 10489 2078 10523
rect 2078 10489 2096 10523
rect 2044 10480 2096 10489
rect 7104 10480 7156 10532
rect 8024 10523 8076 10532
rect 8024 10489 8033 10523
rect 8033 10489 8067 10523
rect 8067 10489 8076 10523
rect 8024 10480 8076 10489
rect 8760 10523 8812 10532
rect 8760 10489 8794 10523
rect 8794 10489 8812 10523
rect 8760 10480 8812 10489
rect 11612 10480 11664 10532
rect 12440 10480 12492 10532
rect 4436 10412 4488 10464
rect 5172 10412 5224 10464
rect 5356 10455 5408 10464
rect 5356 10421 5365 10455
rect 5365 10421 5399 10455
rect 5399 10421 5408 10455
rect 5356 10412 5408 10421
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 7288 10412 7340 10421
rect 11060 10412 11112 10464
rect 11704 10412 11756 10464
rect 13360 10412 13412 10464
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2044 10208 2096 10260
rect 4068 10251 4120 10260
rect 4068 10217 4077 10251
rect 4077 10217 4111 10251
rect 4111 10217 4120 10251
rect 4068 10208 4120 10217
rect 6092 10208 6144 10260
rect 7012 10208 7064 10260
rect 8392 10251 8444 10260
rect 8392 10217 8401 10251
rect 8401 10217 8435 10251
rect 8435 10217 8444 10251
rect 8392 10208 8444 10217
rect 9680 10251 9732 10260
rect 9680 10217 9689 10251
rect 9689 10217 9723 10251
rect 9723 10217 9732 10251
rect 9680 10208 9732 10217
rect 10048 10251 10100 10260
rect 10048 10217 10057 10251
rect 10057 10217 10091 10251
rect 10091 10217 10100 10251
rect 10048 10208 10100 10217
rect 11152 10251 11204 10260
rect 11152 10217 11161 10251
rect 11161 10217 11195 10251
rect 11195 10217 11204 10251
rect 11152 10208 11204 10217
rect 4344 10140 4396 10192
rect 1676 10115 1728 10124
rect 1676 10081 1710 10115
rect 1710 10081 1728 10115
rect 1676 10072 1728 10081
rect 4068 10072 4120 10124
rect 4528 10047 4580 10056
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 5540 10140 5592 10192
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 5632 10072 5684 10124
rect 8208 10140 8260 10192
rect 10140 10140 10192 10192
rect 11796 10140 11848 10192
rect 12624 10208 12676 10260
rect 13268 10251 13320 10260
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 13728 10183 13780 10192
rect 9864 10072 9916 10124
rect 2688 9936 2740 9988
rect 8852 10004 8904 10056
rect 10508 10072 10560 10124
rect 11612 10115 11664 10124
rect 11612 10081 11621 10115
rect 11621 10081 11655 10115
rect 11655 10081 11664 10115
rect 11612 10072 11664 10081
rect 12440 10072 12492 10124
rect 13728 10149 13737 10183
rect 13737 10149 13771 10183
rect 13771 10149 13780 10183
rect 13728 10140 13780 10149
rect 13084 10072 13136 10124
rect 14372 10072 14424 10124
rect 6460 9936 6512 9988
rect 7012 9936 7064 9988
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 11888 10047 11940 10056
rect 10232 10004 10284 10013
rect 11888 10013 11897 10047
rect 11897 10013 11931 10047
rect 11931 10013 11940 10047
rect 11888 10004 11940 10013
rect 12256 10004 12308 10056
rect 13820 10047 13872 10056
rect 13820 10013 13829 10047
rect 13829 10013 13863 10047
rect 13863 10013 13872 10047
rect 13820 10004 13872 10013
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 2320 9868 2372 9920
rect 7104 9868 7156 9920
rect 8484 9868 8536 9920
rect 12348 9911 12400 9920
rect 12348 9877 12357 9911
rect 12357 9877 12391 9911
rect 12391 9877 12400 9911
rect 12348 9868 12400 9877
rect 14004 9868 14056 9920
rect 14648 9911 14700 9920
rect 14648 9877 14657 9911
rect 14657 9877 14691 9911
rect 14691 9877 14700 9911
rect 14648 9868 14700 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1676 9707 1728 9716
rect 1676 9673 1685 9707
rect 1685 9673 1719 9707
rect 1719 9673 1728 9707
rect 1676 9664 1728 9673
rect 2596 9596 2648 9648
rect 4528 9664 4580 9716
rect 5080 9664 5132 9716
rect 6460 9664 6512 9716
rect 7104 9664 7156 9716
rect 8392 9664 8444 9716
rect 11612 9664 11664 9716
rect 13084 9664 13136 9716
rect 10508 9639 10560 9648
rect 10508 9605 10517 9639
rect 10517 9605 10551 9639
rect 10551 9605 10560 9639
rect 10508 9596 10560 9605
rect 13820 9639 13872 9648
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 14648 9664 14700 9716
rect 15384 9639 15436 9648
rect 15384 9605 15393 9639
rect 15393 9605 15427 9639
rect 15427 9605 15436 9639
rect 15384 9596 15436 9605
rect 2688 9460 2740 9512
rect 3516 9460 3568 9512
rect 10140 9571 10192 9580
rect 5080 9460 5132 9512
rect 6736 9460 6788 9512
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 7472 9460 7524 9512
rect 9772 9460 9824 9512
rect 11704 9460 11756 9512
rect 14004 9460 14056 9512
rect 3884 9392 3936 9444
rect 4620 9392 4672 9444
rect 6460 9392 6512 9444
rect 6920 9392 6972 9444
rect 10692 9392 10744 9444
rect 12348 9392 12400 9444
rect 2320 9324 2372 9376
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 4344 9324 4396 9376
rect 6000 9324 6052 9376
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 11796 9367 11848 9376
rect 11796 9333 11805 9367
rect 11805 9333 11839 9367
rect 11839 9333 11848 9367
rect 11796 9324 11848 9333
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 12440 9324 12492 9376
rect 14372 9367 14424 9376
rect 14372 9333 14381 9367
rect 14381 9333 14415 9367
rect 14415 9333 14424 9367
rect 14372 9324 14424 9333
rect 14832 9324 14884 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1584 9120 1636 9172
rect 3884 9163 3936 9172
rect 3884 9129 3893 9163
rect 3893 9129 3927 9163
rect 3927 9129 3936 9163
rect 3884 9120 3936 9129
rect 4068 9163 4120 9172
rect 4068 9129 4077 9163
rect 4077 9129 4111 9163
rect 4111 9129 4120 9163
rect 4068 9120 4120 9129
rect 4252 9120 4304 9172
rect 4620 9120 4672 9172
rect 8300 9163 8352 9172
rect 8300 9129 8309 9163
rect 8309 9129 8343 9163
rect 8343 9129 8352 9163
rect 8300 9120 8352 9129
rect 8852 9163 8904 9172
rect 8852 9129 8861 9163
rect 8861 9129 8895 9163
rect 8895 9129 8904 9163
rect 8852 9120 8904 9129
rect 9772 9120 9824 9172
rect 10048 9120 10100 9172
rect 12256 9120 12308 9172
rect 12348 9120 12400 9172
rect 12992 9120 13044 9172
rect 13912 9120 13964 9172
rect 2320 9095 2372 9104
rect 2320 9061 2329 9095
rect 2329 9061 2363 9095
rect 2363 9061 2372 9095
rect 2320 9052 2372 9061
rect 2228 9027 2280 9036
rect 2228 8993 2237 9027
rect 2237 8993 2271 9027
rect 2271 8993 2280 9027
rect 2228 8984 2280 8993
rect 2688 8984 2740 9036
rect 3792 8984 3844 9036
rect 4804 8984 4856 9036
rect 6368 9052 6420 9104
rect 8208 9052 8260 9104
rect 11888 9052 11940 9104
rect 13820 9095 13872 9104
rect 13820 9061 13829 9095
rect 13829 9061 13863 9095
rect 13863 9061 13872 9095
rect 13820 9052 13872 9061
rect 6092 9027 6144 9036
rect 6092 8993 6126 9027
rect 6126 8993 6144 9027
rect 6092 8984 6144 8993
rect 6460 8984 6512 9036
rect 10600 9027 10652 9036
rect 10600 8993 10609 9027
rect 10609 8993 10643 9027
rect 10643 8993 10652 9027
rect 10600 8984 10652 8993
rect 2044 8916 2096 8968
rect 10692 8959 10744 8968
rect 1492 8848 1544 8900
rect 10692 8925 10701 8959
rect 10701 8925 10735 8959
rect 10735 8925 10744 8959
rect 10692 8916 10744 8925
rect 13544 8984 13596 9036
rect 15384 9027 15436 9036
rect 15384 8993 15393 9027
rect 15393 8993 15427 9027
rect 15427 8993 15436 9027
rect 15384 8984 15436 8993
rect 15660 9027 15712 9036
rect 15660 8993 15694 9027
rect 15694 8993 15712 9027
rect 15660 8984 15712 8993
rect 9588 8848 9640 8900
rect 11244 8916 11296 8968
rect 11704 8916 11756 8968
rect 14464 8891 14516 8900
rect 14464 8857 14473 8891
rect 14473 8857 14507 8891
rect 14507 8857 14516 8891
rect 14464 8848 14516 8857
rect 5172 8780 5224 8832
rect 10232 8823 10284 8832
rect 10232 8789 10241 8823
rect 10241 8789 10275 8823
rect 10275 8789 10284 8823
rect 10232 8780 10284 8789
rect 14740 8780 14792 8832
rect 16764 8823 16816 8832
rect 16764 8789 16773 8823
rect 16773 8789 16807 8823
rect 16807 8789 16816 8823
rect 16764 8780 16816 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2136 8576 2188 8628
rect 1768 8440 1820 8492
rect 1492 8372 1544 8424
rect 3884 8576 3936 8628
rect 4252 8576 4304 8628
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 6092 8576 6144 8628
rect 5448 8508 5500 8560
rect 8392 8551 8444 8560
rect 8392 8517 8401 8551
rect 8401 8517 8435 8551
rect 8435 8517 8444 8551
rect 8392 8508 8444 8517
rect 6920 8440 6972 8492
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 3424 8372 3476 8424
rect 8208 8372 8260 8424
rect 9036 8576 9088 8628
rect 9680 8576 9732 8628
rect 10692 8619 10744 8628
rect 10692 8585 10701 8619
rect 10701 8585 10735 8619
rect 10735 8585 10744 8619
rect 10692 8576 10744 8585
rect 11336 8576 11388 8628
rect 10600 8508 10652 8560
rect 12440 8551 12492 8560
rect 12440 8517 12449 8551
rect 12449 8517 12483 8551
rect 12483 8517 12492 8551
rect 12440 8508 12492 8517
rect 11612 8440 11664 8492
rect 11796 8440 11848 8492
rect 12348 8440 12400 8492
rect 9680 8372 9732 8424
rect 2872 8304 2924 8356
rect 2044 8236 2096 8288
rect 3148 8236 3200 8288
rect 5172 8304 5224 8356
rect 5724 8347 5776 8356
rect 5724 8313 5733 8347
rect 5733 8313 5767 8347
rect 5767 8313 5776 8347
rect 5724 8304 5776 8313
rect 7196 8347 7248 8356
rect 7196 8313 7205 8347
rect 7205 8313 7239 8347
rect 7239 8313 7248 8347
rect 7196 8304 7248 8313
rect 8852 8304 8904 8356
rect 15384 8576 15436 8628
rect 17224 8576 17276 8628
rect 13544 8551 13596 8560
rect 13544 8517 13553 8551
rect 13553 8517 13587 8551
rect 13587 8517 13596 8551
rect 13544 8508 13596 8517
rect 14740 8508 14792 8560
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 16304 8483 16356 8492
rect 16304 8449 16313 8483
rect 16313 8449 16347 8483
rect 16347 8449 16356 8483
rect 16304 8440 16356 8449
rect 12900 8415 12952 8424
rect 12900 8381 12909 8415
rect 12909 8381 12943 8415
rect 12943 8381 12952 8415
rect 12900 8372 12952 8381
rect 14464 8372 14516 8424
rect 15936 8372 15988 8424
rect 20904 8415 20956 8424
rect 20904 8381 20913 8415
rect 20913 8381 20947 8415
rect 20947 8381 20956 8415
rect 20904 8372 20956 8381
rect 13912 8304 13964 8356
rect 15660 8304 15712 8356
rect 11152 8236 11204 8288
rect 14464 8279 14516 8288
rect 14464 8245 14473 8279
rect 14473 8245 14507 8279
rect 14507 8245 14516 8279
rect 14464 8236 14516 8245
rect 22008 8304 22060 8356
rect 16672 8236 16724 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1400 8075 1452 8084
rect 1400 8041 1409 8075
rect 1409 8041 1443 8075
rect 1443 8041 1452 8075
rect 1400 8032 1452 8041
rect 2596 8032 2648 8084
rect 2964 8032 3016 8084
rect 3516 8032 3568 8084
rect 5448 8032 5500 8084
rect 6552 8032 6604 8084
rect 7840 8075 7892 8084
rect 4804 7964 4856 8016
rect 5264 7964 5316 8016
rect 7840 8041 7849 8075
rect 7849 8041 7883 8075
rect 7883 8041 7892 8075
rect 7840 8032 7892 8041
rect 8208 8075 8260 8084
rect 8208 8041 8217 8075
rect 8217 8041 8251 8075
rect 8251 8041 8260 8075
rect 8208 8032 8260 8041
rect 8484 8032 8536 8084
rect 9588 8032 9640 8084
rect 9956 8032 10008 8084
rect 10692 8032 10744 8084
rect 7012 7964 7064 8016
rect 10140 7964 10192 8016
rect 5356 7896 5408 7948
rect 7288 7896 7340 7948
rect 11060 7964 11112 8016
rect 11704 7939 11756 7948
rect 11704 7905 11738 7939
rect 11738 7905 11756 7939
rect 11704 7896 11756 7905
rect 15108 7896 15160 7948
rect 15568 7939 15620 7948
rect 15568 7905 15602 7939
rect 15602 7905 15620 7939
rect 15568 7896 15620 7905
rect 2504 7828 2556 7880
rect 3148 7828 3200 7880
rect 3240 7828 3292 7880
rect 1768 7760 1820 7812
rect 1860 7735 1912 7744
rect 1860 7701 1869 7735
rect 1869 7701 1903 7735
rect 1903 7701 1912 7735
rect 1860 7692 1912 7701
rect 3240 7692 3292 7744
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 6736 7871 6788 7880
rect 5264 7828 5316 7837
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 6184 7803 6236 7812
rect 6184 7769 6193 7803
rect 6193 7769 6227 7803
rect 6227 7769 6236 7803
rect 6184 7760 6236 7769
rect 7748 7803 7800 7812
rect 7748 7769 7757 7803
rect 7757 7769 7791 7803
rect 7791 7769 7800 7803
rect 7748 7760 7800 7769
rect 7932 7760 7984 7812
rect 11060 7828 11112 7880
rect 11336 7828 11388 7880
rect 14188 7871 14240 7880
rect 14188 7837 14197 7871
rect 14197 7837 14231 7871
rect 14231 7837 14240 7871
rect 14188 7828 14240 7837
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 11244 7803 11296 7812
rect 11244 7769 11253 7803
rect 11253 7769 11287 7803
rect 11287 7769 11296 7803
rect 11244 7760 11296 7769
rect 12808 7803 12860 7812
rect 12808 7769 12817 7803
rect 12817 7769 12851 7803
rect 12851 7769 12860 7803
rect 12808 7760 12860 7769
rect 6092 7692 6144 7744
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6276 7692 6328 7701
rect 7472 7692 7524 7744
rect 13636 7692 13688 7744
rect 14004 7692 14056 7744
rect 14740 7692 14792 7744
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 3240 7488 3292 7540
rect 5264 7488 5316 7540
rect 6460 7488 6512 7540
rect 6736 7488 6788 7540
rect 7012 7531 7064 7540
rect 7012 7497 7021 7531
rect 7021 7497 7055 7531
rect 7055 7497 7064 7531
rect 7012 7488 7064 7497
rect 7288 7488 7340 7540
rect 9956 7531 10008 7540
rect 9956 7497 9965 7531
rect 9965 7497 9999 7531
rect 9999 7497 10008 7531
rect 9956 7488 10008 7497
rect 10140 7488 10192 7540
rect 10692 7488 10744 7540
rect 12900 7488 12952 7540
rect 15568 7488 15620 7540
rect 17224 7531 17276 7540
rect 17224 7497 17233 7531
rect 17233 7497 17267 7531
rect 17267 7497 17276 7531
rect 17224 7488 17276 7497
rect 2964 7420 3016 7472
rect 3976 7420 4028 7472
rect 4344 7463 4396 7472
rect 4344 7429 4353 7463
rect 4353 7429 4387 7463
rect 4387 7429 4396 7463
rect 4344 7420 4396 7429
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 2688 7284 2740 7336
rect 5632 7420 5684 7472
rect 9680 7420 9732 7472
rect 11336 7420 11388 7472
rect 11244 7395 11296 7404
rect 11244 7361 11253 7395
rect 11253 7361 11287 7395
rect 11287 7361 11296 7395
rect 11244 7352 11296 7361
rect 11704 7352 11756 7404
rect 6184 7284 6236 7336
rect 7564 7284 7616 7336
rect 7748 7284 7800 7336
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 11152 7327 11204 7336
rect 11152 7293 11161 7327
rect 11161 7293 11195 7327
rect 11195 7293 11204 7327
rect 11152 7284 11204 7293
rect 1768 7259 1820 7268
rect 1768 7225 1777 7259
rect 1777 7225 1811 7259
rect 1811 7225 1820 7259
rect 1768 7216 1820 7225
rect 3148 7216 3200 7268
rect 5356 7259 5408 7268
rect 5356 7225 5365 7259
rect 5365 7225 5399 7259
rect 5399 7225 5408 7259
rect 5356 7216 5408 7225
rect 6092 7216 6144 7268
rect 1860 7191 1912 7200
rect 1860 7157 1869 7191
rect 1869 7157 1903 7191
rect 1903 7157 1912 7191
rect 1860 7148 1912 7157
rect 2504 7191 2556 7200
rect 2504 7157 2513 7191
rect 2513 7157 2547 7191
rect 2547 7157 2556 7191
rect 2504 7148 2556 7157
rect 5724 7191 5776 7200
rect 5724 7157 5733 7191
rect 5733 7157 5767 7191
rect 5767 7157 5776 7191
rect 5724 7148 5776 7157
rect 8852 7148 8904 7200
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 13636 7352 13688 7404
rect 13820 7352 13872 7404
rect 13360 7284 13412 7336
rect 15016 7284 15068 7336
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 12348 7148 12400 7200
rect 12900 7148 12952 7200
rect 13912 7216 13964 7268
rect 15844 7216 15896 7268
rect 18328 7259 18380 7268
rect 18328 7225 18337 7259
rect 18337 7225 18371 7259
rect 18371 7225 18380 7259
rect 18328 7216 18380 7225
rect 13728 7148 13780 7200
rect 16304 7191 16356 7200
rect 16304 7157 16313 7191
rect 16313 7157 16347 7191
rect 16347 7157 16356 7191
rect 16304 7148 16356 7157
rect 16856 7191 16908 7200
rect 16856 7157 16865 7191
rect 16865 7157 16899 7191
rect 16899 7157 16908 7191
rect 16856 7148 16908 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 3148 6944 3200 6996
rect 4436 6944 4488 6996
rect 4804 6944 4856 6996
rect 4988 6944 5040 6996
rect 5448 6944 5500 6996
rect 7748 6944 7800 6996
rect 13360 6987 13412 6996
rect 13360 6953 13369 6987
rect 13369 6953 13403 6987
rect 13403 6953 13412 6987
rect 13360 6944 13412 6953
rect 14188 6944 14240 6996
rect 16304 6944 16356 6996
rect 17224 6987 17276 6996
rect 17224 6953 17233 6987
rect 17233 6953 17267 6987
rect 17267 6953 17276 6987
rect 17224 6944 17276 6953
rect 19156 6987 19208 6996
rect 19156 6953 19165 6987
rect 19165 6953 19199 6987
rect 19199 6953 19208 6987
rect 19156 6944 19208 6953
rect 5356 6876 5408 6928
rect 10048 6919 10100 6928
rect 10048 6885 10057 6919
rect 10057 6885 10091 6919
rect 10091 6885 10100 6919
rect 10048 6876 10100 6885
rect 2596 6808 2648 6860
rect 3976 6808 4028 6860
rect 5632 6808 5684 6860
rect 6368 6808 6420 6860
rect 6736 6851 6788 6860
rect 6736 6817 6770 6851
rect 6770 6817 6788 6851
rect 4160 6740 4212 6792
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 2872 6715 2924 6724
rect 2872 6681 2881 6715
rect 2881 6681 2915 6715
rect 2915 6681 2924 6715
rect 2872 6672 2924 6681
rect 3056 6672 3108 6724
rect 3424 6672 3476 6724
rect 5172 6672 5224 6724
rect 2688 6604 2740 6656
rect 2780 6604 2832 6656
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 4252 6604 4304 6613
rect 4620 6604 4672 6656
rect 6000 6647 6052 6656
rect 6000 6613 6009 6647
rect 6009 6613 6043 6647
rect 6043 6613 6052 6647
rect 6000 6604 6052 6613
rect 6736 6808 6788 6817
rect 8300 6808 8352 6860
rect 9496 6851 9548 6860
rect 9496 6817 9505 6851
rect 9505 6817 9539 6851
rect 9539 6817 9548 6851
rect 9496 6808 9548 6817
rect 9680 6808 9732 6860
rect 9864 6808 9916 6860
rect 11152 6876 11204 6928
rect 14004 6876 14056 6928
rect 24124 6876 24176 6928
rect 24676 6876 24728 6928
rect 11520 6851 11572 6860
rect 11520 6817 11554 6851
rect 11554 6817 11572 6851
rect 11520 6808 11572 6817
rect 13912 6851 13964 6860
rect 13912 6817 13921 6851
rect 13921 6817 13955 6851
rect 13955 6817 13964 6851
rect 13912 6808 13964 6817
rect 14464 6808 14516 6860
rect 19064 6808 19116 6860
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 14188 6783 14240 6792
rect 7104 6604 7156 6656
rect 7564 6672 7616 6724
rect 9864 6672 9916 6724
rect 9956 6672 10008 6724
rect 7472 6604 7524 6656
rect 9312 6604 9364 6656
rect 10784 6604 10836 6656
rect 14188 6749 14197 6783
rect 14197 6749 14231 6783
rect 14231 6749 14240 6783
rect 14188 6740 14240 6749
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 12440 6672 12492 6724
rect 15384 6715 15436 6724
rect 15384 6681 15393 6715
rect 15393 6681 15427 6715
rect 15427 6681 15436 6715
rect 15384 6672 15436 6681
rect 11888 6604 11940 6656
rect 12348 6604 12400 6656
rect 14372 6604 14424 6656
rect 16856 6604 16908 6656
rect 17224 6604 17276 6656
rect 21180 6783 21232 6792
rect 21180 6749 21189 6783
rect 21189 6749 21223 6783
rect 21223 6749 21232 6783
rect 21180 6740 21232 6749
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 3148 6400 3200 6452
rect 5356 6400 5408 6452
rect 7932 6443 7984 6452
rect 7932 6409 7941 6443
rect 7941 6409 7975 6443
rect 7975 6409 7984 6443
rect 7932 6400 7984 6409
rect 10048 6400 10100 6452
rect 11520 6400 11572 6452
rect 13820 6400 13872 6452
rect 3516 6332 3568 6384
rect 3792 6332 3844 6384
rect 4068 6332 4120 6384
rect 9864 6332 9916 6384
rect 12440 6375 12492 6384
rect 12440 6341 12449 6375
rect 12449 6341 12483 6375
rect 12483 6341 12492 6375
rect 12440 6332 12492 6341
rect 1584 6264 1636 6316
rect 2044 6264 2096 6316
rect 3148 6264 3200 6316
rect 4528 6264 4580 6316
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 12992 6307 13044 6316
rect 1952 6239 2004 6248
rect 1952 6205 1961 6239
rect 1961 6205 1995 6239
rect 1995 6205 2004 6239
rect 1952 6196 2004 6205
rect 2780 6196 2832 6248
rect 3240 6196 3292 6248
rect 4160 6196 4212 6248
rect 4436 6196 4488 6248
rect 4620 6196 4672 6248
rect 6000 6196 6052 6248
rect 8576 6239 8628 6248
rect 8576 6205 8585 6239
rect 8585 6205 8619 6239
rect 8619 6205 8628 6239
rect 8576 6196 8628 6205
rect 12992 6273 13001 6307
rect 13001 6273 13035 6307
rect 13035 6273 13044 6307
rect 12992 6264 13044 6273
rect 8852 6239 8904 6248
rect 8852 6205 8886 6239
rect 8886 6205 8904 6239
rect 8852 6196 8904 6205
rect 9956 6196 10008 6248
rect 16028 6400 16080 6452
rect 16672 6443 16724 6452
rect 16672 6409 16681 6443
rect 16681 6409 16715 6443
rect 16715 6409 16724 6443
rect 16672 6400 16724 6409
rect 19064 6443 19116 6452
rect 19064 6409 19073 6443
rect 19073 6409 19107 6443
rect 19107 6409 19116 6443
rect 19064 6400 19116 6409
rect 20904 6443 20956 6452
rect 20904 6409 20913 6443
rect 20913 6409 20947 6443
rect 20947 6409 20956 6443
rect 20904 6400 20956 6409
rect 16304 6375 16356 6384
rect 16304 6341 16313 6375
rect 16313 6341 16347 6375
rect 16347 6341 16356 6375
rect 16304 6332 16356 6341
rect 18144 6332 18196 6384
rect 14372 6307 14424 6316
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 18696 6307 18748 6316
rect 18696 6273 18705 6307
rect 18705 6273 18739 6307
rect 18739 6273 18748 6307
rect 18696 6264 18748 6273
rect 14648 6239 14700 6248
rect 14648 6205 14671 6239
rect 14671 6205 14700 6239
rect 16856 6239 16908 6248
rect 14648 6196 14700 6205
rect 16856 6205 16865 6239
rect 16865 6205 16899 6239
rect 16899 6205 16908 6239
rect 16856 6196 16908 6205
rect 17776 6239 17828 6248
rect 17776 6205 17785 6239
rect 17785 6205 17819 6239
rect 17819 6205 17828 6239
rect 17776 6196 17828 6205
rect 3424 6128 3476 6180
rect 5356 6128 5408 6180
rect 7472 6128 7524 6180
rect 13084 6128 13136 6180
rect 1676 6060 1728 6112
rect 3516 6060 3568 6112
rect 4436 6060 4488 6112
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 9864 6060 9916 6112
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 11336 6060 11388 6069
rect 12164 6103 12216 6112
rect 12164 6069 12173 6103
rect 12173 6069 12207 6103
rect 12207 6069 12216 6103
rect 12164 6060 12216 6069
rect 15844 6060 15896 6112
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1952 5856 2004 5908
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 5172 5856 5224 5908
rect 6736 5856 6788 5908
rect 7288 5856 7340 5908
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 10968 5856 11020 5908
rect 11796 5899 11848 5908
rect 11796 5865 11805 5899
rect 11805 5865 11839 5899
rect 11839 5865 11848 5899
rect 11796 5856 11848 5865
rect 14372 5899 14424 5908
rect 14372 5865 14381 5899
rect 14381 5865 14415 5899
rect 14415 5865 14424 5899
rect 14372 5856 14424 5865
rect 14832 5856 14884 5908
rect 15292 5856 15344 5908
rect 15752 5899 15804 5908
rect 15752 5865 15761 5899
rect 15761 5865 15795 5899
rect 15795 5865 15804 5899
rect 16304 5899 16356 5908
rect 15752 5856 15804 5865
rect 16304 5865 16313 5899
rect 16313 5865 16347 5899
rect 16347 5865 16356 5899
rect 16304 5856 16356 5865
rect 19064 5856 19116 5908
rect 2596 5788 2648 5840
rect 2688 5788 2740 5840
rect 7104 5788 7156 5840
rect 7472 5788 7524 5840
rect 14464 5788 14516 5840
rect 17500 5788 17552 5840
rect 18696 5788 18748 5840
rect 4896 5763 4948 5772
rect 4896 5729 4930 5763
rect 4930 5729 4948 5763
rect 4896 5720 4948 5729
rect 10692 5763 10744 5772
rect 10692 5729 10701 5763
rect 10701 5729 10735 5763
rect 10735 5729 10744 5763
rect 10692 5720 10744 5729
rect 10968 5720 11020 5772
rect 2412 5652 2464 5704
rect 7104 5695 7156 5704
rect 2228 5584 2280 5636
rect 7104 5661 7113 5695
rect 7113 5661 7147 5695
rect 7147 5661 7156 5695
rect 7104 5652 7156 5661
rect 9956 5652 10008 5704
rect 20904 5763 20956 5772
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 11888 5695 11940 5704
rect 11888 5661 11897 5695
rect 11897 5661 11931 5695
rect 11931 5661 11940 5695
rect 11888 5652 11940 5661
rect 13912 5695 13964 5704
rect 13912 5661 13921 5695
rect 13921 5661 13955 5695
rect 13955 5661 13964 5695
rect 13912 5652 13964 5661
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 16488 5652 16540 5704
rect 11704 5584 11756 5636
rect 15936 5584 15988 5636
rect 16856 5627 16908 5636
rect 16856 5593 16865 5627
rect 16865 5593 16899 5627
rect 16899 5593 16908 5627
rect 16856 5584 16908 5593
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 9312 5516 9364 5568
rect 11152 5516 11204 5568
rect 13636 5516 13688 5568
rect 17224 5559 17276 5568
rect 17224 5525 17233 5559
rect 17233 5525 17267 5559
rect 17267 5525 17276 5559
rect 17224 5516 17276 5525
rect 21088 5559 21140 5568
rect 21088 5525 21097 5559
rect 21097 5525 21131 5559
rect 21131 5525 21140 5559
rect 21088 5516 21140 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 4528 5312 4580 5364
rect 7472 5355 7524 5364
rect 7472 5321 7481 5355
rect 7481 5321 7515 5355
rect 7515 5321 7524 5355
rect 7472 5312 7524 5321
rect 10784 5312 10836 5364
rect 11060 5312 11112 5364
rect 11704 5312 11756 5364
rect 14648 5312 14700 5364
rect 15292 5355 15344 5364
rect 15292 5321 15301 5355
rect 15301 5321 15335 5355
rect 15335 5321 15344 5355
rect 15292 5312 15344 5321
rect 16488 5312 16540 5364
rect 17500 5355 17552 5364
rect 17500 5321 17509 5355
rect 17509 5321 17543 5355
rect 17543 5321 17552 5355
rect 17500 5312 17552 5321
rect 20904 5355 20956 5364
rect 1768 5176 1820 5228
rect 5356 5176 5408 5228
rect 9496 5244 9548 5296
rect 15660 5219 15712 5228
rect 1492 5108 1544 5160
rect 3148 5151 3200 5160
rect 3148 5117 3182 5151
rect 3182 5117 3200 5151
rect 3148 5108 3200 5117
rect 4896 5151 4948 5160
rect 4896 5117 4905 5151
rect 4905 5117 4939 5151
rect 4939 5117 4948 5151
rect 4896 5108 4948 5117
rect 6184 5108 6236 5160
rect 8208 5108 8260 5160
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 16396 5219 16448 5228
rect 15660 5176 15712 5185
rect 9312 5108 9364 5160
rect 11796 5108 11848 5160
rect 12440 5108 12492 5160
rect 16396 5185 16405 5219
rect 16405 5185 16439 5219
rect 16439 5185 16448 5219
rect 16396 5176 16448 5185
rect 16304 5151 16356 5160
rect 16304 5117 16313 5151
rect 16313 5117 16347 5151
rect 16347 5117 16356 5151
rect 19064 5176 19116 5228
rect 20904 5321 20913 5355
rect 20913 5321 20947 5355
rect 20947 5321 20956 5355
rect 20904 5312 20956 5321
rect 16304 5108 16356 5117
rect 5356 5040 5408 5092
rect 7288 5040 7340 5092
rect 7564 5040 7616 5092
rect 9404 5040 9456 5092
rect 2412 4972 2464 5024
rect 2596 5015 2648 5024
rect 2596 4981 2605 5015
rect 2605 4981 2639 5015
rect 2639 4981 2648 5015
rect 2596 4972 2648 4981
rect 7472 4972 7524 5024
rect 7932 5015 7984 5024
rect 7932 4981 7941 5015
rect 7941 4981 7975 5015
rect 7975 4981 7984 5015
rect 7932 4972 7984 4981
rect 9864 5040 9916 5092
rect 10692 5040 10744 5092
rect 13636 5083 13688 5092
rect 13636 5049 13670 5083
rect 13670 5049 13688 5083
rect 13636 5040 13688 5049
rect 13728 5040 13780 5092
rect 18052 5040 18104 5092
rect 11888 4972 11940 5024
rect 14832 4972 14884 5024
rect 18512 5015 18564 5024
rect 18512 4981 18521 5015
rect 18521 4981 18555 5015
rect 18555 4981 18564 5015
rect 18512 4972 18564 4981
rect 21548 4972 21600 5024
rect 21640 5015 21692 5024
rect 21640 4981 21649 5015
rect 21649 4981 21683 5015
rect 21683 4981 21692 5015
rect 21640 4972 21692 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 3148 4768 3200 4820
rect 3424 4811 3476 4820
rect 3424 4777 3433 4811
rect 3433 4777 3467 4811
rect 3467 4777 3476 4811
rect 3424 4768 3476 4777
rect 3608 4768 3660 4820
rect 6092 4768 6144 4820
rect 7564 4811 7616 4820
rect 7564 4777 7573 4811
rect 7573 4777 7607 4811
rect 7607 4777 7616 4811
rect 7564 4768 7616 4777
rect 8300 4811 8352 4820
rect 8300 4777 8309 4811
rect 8309 4777 8343 4811
rect 8343 4777 8352 4811
rect 8300 4768 8352 4777
rect 12624 4811 12676 4820
rect 12624 4777 12633 4811
rect 12633 4777 12667 4811
rect 12667 4777 12676 4811
rect 12624 4768 12676 4777
rect 13084 4811 13136 4820
rect 13084 4777 13093 4811
rect 13093 4777 13127 4811
rect 13127 4777 13136 4811
rect 13084 4768 13136 4777
rect 14740 4768 14792 4820
rect 15752 4811 15804 4820
rect 15752 4777 15761 4811
rect 15761 4777 15795 4811
rect 15795 4777 15804 4811
rect 15752 4768 15804 4777
rect 16396 4811 16448 4820
rect 16396 4777 16405 4811
rect 16405 4777 16439 4811
rect 16439 4777 16448 4811
rect 16396 4768 16448 4777
rect 18696 4768 18748 4820
rect 10784 4700 10836 4752
rect 10968 4700 11020 4752
rect 13728 4700 13780 4752
rect 24216 4743 24268 4752
rect 24216 4709 24250 4743
rect 24250 4709 24268 4743
rect 24216 4700 24268 4709
rect 1584 4632 1636 4684
rect 2596 4632 2648 4684
rect 4620 4675 4672 4684
rect 4620 4641 4629 4675
rect 4629 4641 4663 4675
rect 4663 4641 4672 4675
rect 4620 4632 4672 4641
rect 4896 4632 4948 4684
rect 6092 4632 6144 4684
rect 6460 4632 6512 4684
rect 7840 4675 7892 4684
rect 7840 4641 7849 4675
rect 7849 4641 7883 4675
rect 7883 4641 7892 4675
rect 7840 4632 7892 4641
rect 1492 4607 1544 4616
rect 1492 4573 1501 4607
rect 1501 4573 1535 4607
rect 1535 4573 1544 4607
rect 1492 4564 1544 4573
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 13268 4632 13320 4684
rect 14096 4675 14148 4684
rect 14096 4641 14105 4675
rect 14105 4641 14139 4675
rect 14139 4641 14148 4675
rect 14096 4632 14148 4641
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 17132 4632 17184 4684
rect 19432 4632 19484 4684
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 21180 4632 21232 4684
rect 21824 4632 21876 4684
rect 4436 4496 4488 4548
rect 6000 4496 6052 4548
rect 6184 4496 6236 4548
rect 7288 4496 7340 4548
rect 8024 4564 8076 4616
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 13360 4564 13412 4616
rect 13636 4607 13688 4616
rect 13636 4573 13645 4607
rect 13645 4573 13679 4607
rect 13679 4573 13688 4607
rect 13636 4564 13688 4573
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 10508 4496 10560 4548
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 5080 4428 5132 4480
rect 5356 4428 5408 4480
rect 10048 4428 10100 4480
rect 10968 4428 11020 4480
rect 11704 4428 11756 4480
rect 14648 4428 14700 4480
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 20628 4564 20680 4616
rect 23940 4607 23992 4616
rect 23940 4573 23949 4607
rect 23949 4573 23983 4607
rect 23983 4573 23992 4607
rect 23940 4564 23992 4573
rect 25320 4539 25372 4548
rect 25320 4505 25329 4539
rect 25329 4505 25363 4539
rect 25363 4505 25372 4539
rect 25320 4496 25372 4505
rect 17224 4428 17276 4480
rect 17684 4428 17736 4480
rect 19248 4428 19300 4480
rect 20352 4428 20404 4480
rect 23204 4428 23256 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 4160 4224 4212 4276
rect 4804 4224 4856 4276
rect 6184 4224 6236 4276
rect 6736 4224 6788 4276
rect 10784 4224 10836 4276
rect 6000 4156 6052 4208
rect 8024 4156 8076 4208
rect 9404 4156 9456 4208
rect 13728 4224 13780 4276
rect 15660 4224 15712 4276
rect 18512 4224 18564 4276
rect 18696 4224 18748 4276
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 1400 4020 1452 4072
rect 3332 4088 3384 4140
rect 4252 4088 4304 4140
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 7012 4131 7064 4140
rect 5264 4088 5316 4097
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7012 4088 7064 4097
rect 7288 4088 7340 4140
rect 296 3952 348 4004
rect 6276 4020 6328 4072
rect 10508 4088 10560 4140
rect 11244 4131 11296 4140
rect 11244 4097 11253 4131
rect 11253 4097 11287 4131
rect 11287 4097 11296 4131
rect 11244 4088 11296 4097
rect 13268 4156 13320 4208
rect 20904 4224 20956 4276
rect 21824 4267 21876 4276
rect 21824 4233 21833 4267
rect 21833 4233 21867 4267
rect 21867 4233 21876 4267
rect 21824 4224 21876 4233
rect 24216 4224 24268 4276
rect 23940 4156 23992 4208
rect 11060 4063 11112 4072
rect 2872 3952 2924 4004
rect 6092 3952 6144 4004
rect 8576 3952 8628 4004
rect 10508 3995 10560 4004
rect 10508 3961 10517 3995
rect 10517 3961 10551 3995
rect 10551 3961 10560 3995
rect 10508 3952 10560 3961
rect 4988 3884 5040 3936
rect 5080 3927 5132 3936
rect 5080 3893 5089 3927
rect 5089 3893 5123 3927
rect 5123 3893 5132 3927
rect 7196 3927 7248 3936
rect 5080 3884 5132 3893
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 8300 3884 8352 3936
rect 10048 3884 10100 3936
rect 11060 4029 11069 4063
rect 11069 4029 11103 4063
rect 11103 4029 11112 4063
rect 11060 4020 11112 4029
rect 12624 4020 12676 4072
rect 14096 4020 14148 4072
rect 12072 3884 12124 3936
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 13360 3884 13412 3936
rect 13820 3884 13872 3936
rect 19524 4020 19576 4072
rect 20904 4063 20956 4072
rect 20904 4029 20913 4063
rect 20913 4029 20947 4063
rect 20947 4029 20956 4063
rect 20904 4020 20956 4029
rect 14648 3952 14700 4004
rect 14924 3952 14976 4004
rect 17960 3952 18012 4004
rect 18512 3995 18564 4004
rect 18512 3961 18521 3995
rect 18521 3961 18555 3995
rect 18555 3961 18564 3995
rect 18512 3952 18564 3961
rect 20720 3952 20772 4004
rect 15844 3927 15896 3936
rect 15844 3893 15853 3927
rect 15853 3893 15887 3927
rect 15887 3893 15896 3927
rect 15844 3884 15896 3893
rect 16856 3927 16908 3936
rect 16856 3893 16865 3927
rect 16865 3893 16899 3927
rect 16899 3893 16908 3927
rect 16856 3884 16908 3893
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 17132 3884 17184 3936
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 19432 3927 19484 3936
rect 19432 3893 19441 3927
rect 19441 3893 19475 3927
rect 19475 3893 19484 3927
rect 19432 3884 19484 3893
rect 21088 3927 21140 3936
rect 21088 3893 21097 3927
rect 21097 3893 21131 3927
rect 21131 3893 21140 3927
rect 21088 3884 21140 3893
rect 22192 3927 22244 3936
rect 22192 3893 22201 3927
rect 22201 3893 22235 3927
rect 22235 3893 22244 3927
rect 22192 3884 22244 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2596 3680 2648 3732
rect 2872 3723 2924 3732
rect 2872 3689 2881 3723
rect 2881 3689 2915 3723
rect 2915 3689 2924 3723
rect 2872 3680 2924 3689
rect 3148 3680 3200 3732
rect 4068 3680 4120 3732
rect 5172 3723 5224 3732
rect 5172 3689 5181 3723
rect 5181 3689 5215 3723
rect 5215 3689 5224 3723
rect 5172 3680 5224 3689
rect 6736 3723 6788 3732
rect 6736 3689 6745 3723
rect 6745 3689 6779 3723
rect 6779 3689 6788 3723
rect 6736 3680 6788 3689
rect 8576 3680 8628 3732
rect 10048 3680 10100 3732
rect 11152 3680 11204 3732
rect 13636 3680 13688 3732
rect 2228 3612 2280 3664
rect 5264 3612 5316 3664
rect 7288 3612 7340 3664
rect 10232 3612 10284 3664
rect 10784 3612 10836 3664
rect 11704 3612 11756 3664
rect 14188 3655 14240 3664
rect 14188 3621 14197 3655
rect 14197 3621 14231 3655
rect 14231 3621 14240 3655
rect 14188 3612 14240 3621
rect 5356 3587 5408 3596
rect 5356 3553 5365 3587
rect 5365 3553 5399 3587
rect 5399 3553 5408 3587
rect 5356 3544 5408 3553
rect 1492 3519 1544 3528
rect 1492 3485 1501 3519
rect 1501 3485 1535 3519
rect 1535 3485 1544 3519
rect 1492 3476 1544 3485
rect 3056 3476 3108 3528
rect 7472 3476 7524 3528
rect 3884 3451 3936 3460
rect 3884 3417 3893 3451
rect 3893 3417 3927 3451
rect 3927 3417 3936 3451
rect 3884 3408 3936 3417
rect 7840 3451 7892 3460
rect 7840 3417 7849 3451
rect 7849 3417 7883 3451
rect 7883 3417 7892 3451
rect 7840 3408 7892 3417
rect 8024 3476 8076 3528
rect 10416 3544 10468 3596
rect 12072 3544 12124 3596
rect 13820 3544 13872 3596
rect 14832 3680 14884 3732
rect 15752 3680 15804 3732
rect 16948 3680 17000 3732
rect 19064 3680 19116 3732
rect 19248 3680 19300 3732
rect 20076 3680 20128 3732
rect 20904 3680 20956 3732
rect 22192 3680 22244 3732
rect 15844 3612 15896 3664
rect 16856 3612 16908 3664
rect 17684 3655 17736 3664
rect 17684 3621 17693 3655
rect 17693 3621 17727 3655
rect 17727 3621 17736 3655
rect 17684 3612 17736 3621
rect 17960 3612 18012 3664
rect 18696 3655 18748 3664
rect 18696 3621 18705 3655
rect 18705 3621 18739 3655
rect 18739 3621 18748 3655
rect 18696 3612 18748 3621
rect 18972 3612 19024 3664
rect 22100 3612 22152 3664
rect 24860 3612 24912 3664
rect 25964 3612 26016 3664
rect 14832 3544 14884 3596
rect 16948 3544 17000 3596
rect 22192 3587 22244 3596
rect 8576 3476 8628 3528
rect 10692 3476 10744 3528
rect 10784 3408 10836 3460
rect 4896 3383 4948 3392
rect 4896 3349 4905 3383
rect 4905 3349 4939 3383
rect 4939 3349 4948 3383
rect 4896 3340 4948 3349
rect 18788 3519 18840 3528
rect 18788 3485 18797 3519
rect 18797 3485 18831 3519
rect 18831 3485 18840 3519
rect 18788 3476 18840 3485
rect 12348 3340 12400 3392
rect 20720 3408 20772 3460
rect 22192 3553 22201 3587
rect 22201 3553 22235 3587
rect 22235 3553 22244 3587
rect 22192 3544 22244 3553
rect 23296 3587 23348 3596
rect 23296 3553 23305 3587
rect 23305 3553 23339 3587
rect 23339 3553 23348 3587
rect 23296 3544 23348 3553
rect 24952 3544 25004 3596
rect 25412 3544 25464 3596
rect 21180 3519 21232 3528
rect 21180 3485 21189 3519
rect 21189 3485 21223 3519
rect 21223 3485 21232 3519
rect 21180 3476 21232 3485
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 13728 3340 13780 3392
rect 17132 3383 17184 3392
rect 17132 3349 17141 3383
rect 17141 3349 17175 3383
rect 17175 3349 17184 3383
rect 17132 3340 17184 3349
rect 22376 3383 22428 3392
rect 22376 3349 22385 3383
rect 22385 3349 22419 3383
rect 22419 3349 22428 3383
rect 22376 3340 22428 3349
rect 23756 3340 23808 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 2228 3136 2280 3188
rect 2688 3179 2740 3188
rect 2688 3145 2697 3179
rect 2697 3145 2731 3179
rect 2731 3145 2740 3179
rect 2688 3136 2740 3145
rect 4160 3179 4212 3188
rect 4160 3145 4169 3179
rect 4169 3145 4203 3179
rect 4203 3145 4212 3179
rect 4160 3136 4212 3145
rect 5172 3136 5224 3188
rect 6552 3179 6604 3188
rect 6552 3145 6561 3179
rect 6561 3145 6595 3179
rect 6595 3145 6604 3179
rect 6552 3136 6604 3145
rect 6920 3136 6972 3188
rect 7288 3136 7340 3188
rect 9496 3136 9548 3188
rect 12440 3136 12492 3188
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 16856 3179 16908 3188
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 17132 3136 17184 3188
rect 18788 3136 18840 3188
rect 19064 3179 19116 3188
rect 19064 3145 19073 3179
rect 19073 3145 19107 3179
rect 19107 3145 19116 3179
rect 19064 3136 19116 3145
rect 20720 3179 20772 3188
rect 20720 3145 20729 3179
rect 20729 3145 20763 3179
rect 20763 3145 20772 3179
rect 20720 3136 20772 3145
rect 2872 3068 2924 3120
rect 3148 3043 3200 3052
rect 3148 3009 3157 3043
rect 3157 3009 3191 3043
rect 3191 3009 3200 3043
rect 3148 3000 3200 3009
rect 3516 3000 3568 3052
rect 10232 3068 10284 3120
rect 10416 3111 10468 3120
rect 10416 3077 10425 3111
rect 10425 3077 10459 3111
rect 10459 3077 10468 3111
rect 10416 3068 10468 3077
rect 13820 3111 13872 3120
rect 13820 3077 13829 3111
rect 13829 3077 13863 3111
rect 13863 3077 13872 3111
rect 13820 3068 13872 3077
rect 3056 2975 3108 2984
rect 3056 2941 3065 2975
rect 3065 2941 3099 2975
rect 3099 2941 3108 2975
rect 3056 2932 3108 2941
rect 4068 2932 4120 2984
rect 7104 3000 7156 3052
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 12348 3000 12400 3052
rect 19432 3068 19484 3120
rect 18604 3043 18656 3052
rect 10968 2932 11020 2984
rect 14832 2932 14884 2984
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 19340 3000 19392 3052
rect 18512 2975 18564 2984
rect 18512 2941 18521 2975
rect 18521 2941 18555 2975
rect 18555 2941 18564 2975
rect 22192 3136 22244 3188
rect 22468 3136 22520 3188
rect 23296 3179 23348 3188
rect 23296 3145 23305 3179
rect 23305 3145 23339 3179
rect 23339 3145 23348 3179
rect 23296 3136 23348 3145
rect 26516 3068 26568 3120
rect 18512 2932 18564 2941
rect 20812 2932 20864 2984
rect 22284 2932 22336 2984
rect 23664 2975 23716 2984
rect 23664 2941 23673 2975
rect 23673 2941 23707 2975
rect 23707 2941 23716 2975
rect 23664 2932 23716 2941
rect 24676 2932 24728 2984
rect 1676 2907 1728 2916
rect 1676 2873 1685 2907
rect 1685 2873 1719 2907
rect 1719 2873 1728 2907
rect 1676 2864 1728 2873
rect 7104 2907 7156 2916
rect 7104 2873 7113 2907
rect 7113 2873 7147 2907
rect 7147 2873 7156 2907
rect 7104 2864 7156 2873
rect 8392 2907 8444 2916
rect 8392 2873 8426 2907
rect 8426 2873 8444 2907
rect 8392 2864 8444 2873
rect 12624 2864 12676 2916
rect 14648 2864 14700 2916
rect 17776 2907 17828 2916
rect 6552 2796 6604 2848
rect 7472 2796 7524 2848
rect 9496 2839 9548 2848
rect 9496 2805 9505 2839
rect 9505 2805 9539 2839
rect 9539 2805 9548 2839
rect 9496 2796 9548 2805
rect 10784 2796 10836 2848
rect 11704 2839 11756 2848
rect 11704 2805 11713 2839
rect 11713 2805 11747 2839
rect 11747 2805 11756 2839
rect 11704 2796 11756 2805
rect 17776 2873 17785 2907
rect 17785 2873 17819 2907
rect 17819 2873 17828 2907
rect 17776 2864 17828 2873
rect 19340 2864 19392 2916
rect 22100 2864 22152 2916
rect 18052 2796 18104 2848
rect 18604 2796 18656 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 10692 2592 10744 2644
rect 11612 2635 11664 2644
rect 11612 2601 11621 2635
rect 11621 2601 11655 2635
rect 11655 2601 11664 2635
rect 11612 2592 11664 2601
rect 12900 2635 12952 2644
rect 12900 2601 12909 2635
rect 12909 2601 12943 2635
rect 12943 2601 12952 2635
rect 12900 2592 12952 2601
rect 14372 2592 14424 2644
rect 15660 2592 15712 2644
rect 16948 2635 17000 2644
rect 16948 2601 16957 2635
rect 16957 2601 16991 2635
rect 16991 2601 17000 2635
rect 16948 2592 17000 2601
rect 17684 2635 17736 2644
rect 17684 2601 17693 2635
rect 17693 2601 17727 2635
rect 17727 2601 17736 2635
rect 17684 2592 17736 2601
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 18972 2592 19024 2644
rect 22652 2635 22704 2644
rect 22652 2601 22661 2635
rect 22661 2601 22695 2635
rect 22695 2601 22704 2635
rect 22652 2592 22704 2601
rect 24768 2635 24820 2644
rect 24768 2601 24777 2635
rect 24777 2601 24811 2635
rect 24811 2601 24820 2635
rect 24768 2592 24820 2601
rect 1676 2524 1728 2576
rect 4528 2524 4580 2576
rect 1492 2499 1544 2508
rect 1492 2465 1501 2499
rect 1501 2465 1535 2499
rect 1535 2465 1544 2499
rect 4068 2499 4120 2508
rect 1492 2456 1544 2465
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 6644 2499 6696 2508
rect 6644 2465 6653 2499
rect 6653 2465 6687 2499
rect 6687 2465 6696 2499
rect 9680 2524 9732 2576
rect 6644 2456 6696 2465
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 8668 2431 8720 2440
rect 7472 2388 7524 2397
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 12072 2456 12124 2508
rect 12716 2499 12768 2508
rect 12716 2465 12725 2499
rect 12725 2465 12759 2499
rect 12759 2465 12768 2499
rect 12716 2456 12768 2465
rect 9864 2388 9916 2440
rect 10692 2388 10744 2440
rect 10784 2388 10836 2440
rect 10968 2320 11020 2372
rect 13544 2320 13596 2372
rect 15292 2524 15344 2576
rect 14648 2388 14700 2440
rect 13820 2363 13872 2372
rect 13820 2329 13829 2363
rect 13829 2329 13863 2363
rect 13863 2329 13872 2363
rect 13820 2320 13872 2329
rect 3516 2295 3568 2304
rect 3516 2261 3525 2295
rect 3525 2261 3559 2295
rect 3559 2261 3568 2295
rect 3516 2252 3568 2261
rect 14556 2252 14608 2304
rect 21640 2524 21692 2576
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 19616 2499 19668 2508
rect 19616 2465 19625 2499
rect 19625 2465 19659 2499
rect 19659 2465 19668 2499
rect 19616 2456 19668 2465
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 22468 2499 22520 2508
rect 22468 2465 22477 2499
rect 22477 2465 22511 2499
rect 22511 2465 22520 2499
rect 22468 2456 22520 2465
rect 24124 2456 24176 2508
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 19800 2431 19852 2440
rect 19800 2397 19809 2431
rect 19809 2397 19843 2431
rect 19843 2397 19852 2431
rect 19800 2388 19852 2397
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 16580 2252 16632 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 8668 1368 8720 1420
rect 9588 1368 9640 1420
rect 11796 552 11848 604
rect 13084 552 13136 604
<< metal2 >>
rect 2778 27704 2834 27713
rect 2778 27639 2834 27648
rect 2686 26072 2742 26081
rect 2686 26007 2742 26016
rect 1582 25528 1638 25537
rect 1582 25463 1638 25472
rect 1490 24984 1546 24993
rect 1596 24954 1624 25463
rect 1490 24919 1546 24928
rect 1584 24948 1636 24954
rect 1504 24410 1532 24919
rect 1584 24890 1636 24896
rect 2136 24608 2188 24614
rect 2136 24550 2188 24556
rect 1492 24404 1544 24410
rect 1492 24346 1544 24352
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 1412 23526 1440 24210
rect 2042 24168 2098 24177
rect 2042 24103 2044 24112
rect 2096 24103 2098 24112
rect 2044 24074 2096 24080
rect 2056 23746 2084 24074
rect 1964 23718 2084 23746
rect 1964 23662 1992 23718
rect 1952 23656 2004 23662
rect 1952 23598 2004 23604
rect 1400 23520 1452 23526
rect 1400 23462 1452 23468
rect 1952 23520 2004 23526
rect 1952 23462 2004 23468
rect 1490 23216 1546 23225
rect 1490 23151 1546 23160
rect 1676 23180 1728 23186
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 1412 21350 1440 22034
rect 1504 21690 1532 23151
rect 1676 23122 1728 23128
rect 1688 22574 1716 23122
rect 1964 22642 1992 23462
rect 2148 23254 2176 24550
rect 2700 24410 2728 26007
rect 2792 25498 2820 27639
rect 3330 27160 3386 27169
rect 3330 27095 3386 27104
rect 3344 26722 3372 27095
rect 3332 26716 3384 26722
rect 3332 26658 3384 26664
rect 5448 26716 5500 26722
rect 5448 26658 5500 26664
rect 3238 26616 3294 26625
rect 3238 26551 3294 26560
rect 2780 25492 2832 25498
rect 2780 25434 2832 25440
rect 2962 24440 3018 24449
rect 2688 24404 2740 24410
rect 2962 24375 3018 24384
rect 2688 24346 2740 24352
rect 2504 24268 2556 24274
rect 2504 24210 2556 24216
rect 2516 23866 2544 24210
rect 2686 23896 2742 23905
rect 2504 23860 2556 23866
rect 2686 23831 2742 23840
rect 2504 23802 2556 23808
rect 2136 23248 2188 23254
rect 2136 23190 2188 23196
rect 1952 22636 2004 22642
rect 1952 22578 2004 22584
rect 1676 22568 1728 22574
rect 1674 22536 1676 22545
rect 1728 22536 1730 22545
rect 1674 22471 1730 22480
rect 2596 22432 2648 22438
rect 2594 22400 2596 22409
rect 2648 22400 2650 22409
rect 2594 22335 2650 22344
rect 2412 22092 2464 22098
rect 2412 22034 2464 22040
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 1492 21684 1544 21690
rect 1492 21626 1544 21632
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1596 21049 1624 21830
rect 1676 21480 1728 21486
rect 1676 21422 1728 21428
rect 2044 21480 2096 21486
rect 2424 21457 2452 22034
rect 2700 21962 2728 23831
rect 2976 22778 3004 24375
rect 3252 23866 3280 26551
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3698 23760 3754 23769
rect 3698 23695 3700 23704
rect 3752 23695 3754 23704
rect 3700 23666 3752 23672
rect 2964 22772 3016 22778
rect 2964 22714 3016 22720
rect 3422 22672 3478 22681
rect 3422 22607 3478 22616
rect 3436 22001 3464 22607
rect 3700 22432 3752 22438
rect 3700 22374 3752 22380
rect 4434 22400 4490 22409
rect 3422 21992 3478 22001
rect 2688 21956 2740 21962
rect 3422 21927 3478 21936
rect 2688 21898 2740 21904
rect 2688 21616 2740 21622
rect 2686 21584 2688 21593
rect 2740 21584 2742 21593
rect 2686 21519 2742 21528
rect 2044 21422 2096 21428
rect 2410 21448 2466 21457
rect 1582 21040 1638 21049
rect 1582 20975 1638 20984
rect 1688 20942 1716 21422
rect 1768 21004 1820 21010
rect 1768 20946 1820 20952
rect 1676 20936 1728 20942
rect 1674 20904 1676 20913
rect 1728 20904 1730 20913
rect 1674 20839 1730 20848
rect 1780 20262 1808 20946
rect 2056 20466 2084 21422
rect 2410 21383 2412 21392
rect 2464 21383 2466 21392
rect 2412 21354 2464 21360
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1688 19174 1716 19858
rect 1780 19825 1808 20198
rect 1766 19816 1822 19825
rect 1766 19751 1822 19760
rect 2516 19378 2544 21286
rect 2688 20936 2740 20942
rect 2688 20878 2740 20884
rect 2594 20632 2650 20641
rect 2594 20567 2596 20576
rect 2648 20567 2650 20576
rect 2596 20538 2648 20544
rect 2608 20398 2636 20538
rect 2700 20505 2728 20878
rect 2686 20496 2742 20505
rect 2686 20431 2742 20440
rect 2596 20392 2648 20398
rect 2780 20392 2832 20398
rect 2596 20334 2648 20340
rect 2700 20340 2780 20346
rect 2700 20334 2832 20340
rect 2700 20318 2820 20334
rect 2504 19372 2556 19378
rect 2504 19314 2556 19320
rect 2700 19310 2728 20318
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 3252 19961 3280 20198
rect 3712 20097 3740 22374
rect 4434 22335 4490 22344
rect 4066 22128 4122 22137
rect 4066 22063 4122 22072
rect 4080 20618 4108 22063
rect 4080 20602 4200 20618
rect 4080 20596 4212 20602
rect 4080 20590 4160 20596
rect 4160 20538 4212 20544
rect 4158 20496 4214 20505
rect 4158 20431 4214 20440
rect 4172 20398 4200 20431
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 4250 20224 4306 20233
rect 4250 20159 4306 20168
rect 3698 20088 3754 20097
rect 4264 20058 4292 20159
rect 3698 20023 3754 20032
rect 4252 20052 4304 20058
rect 4252 19994 4304 20000
rect 3238 19952 3294 19961
rect 2964 19916 3016 19922
rect 3238 19887 3294 19896
rect 4068 19916 4120 19922
rect 2964 19858 3016 19864
rect 4068 19858 4120 19864
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 1676 19168 1728 19174
rect 1674 19136 1676 19145
rect 2688 19168 2740 19174
rect 1728 19136 1730 19145
rect 2688 19110 2740 19116
rect 1674 19071 1730 19080
rect 2700 19009 2728 19110
rect 2686 19000 2742 19009
rect 1492 18964 1544 18970
rect 2686 18935 2742 18944
rect 1492 18906 1544 18912
rect 1504 18222 1532 18906
rect 2596 18828 2648 18834
rect 2596 18770 2648 18776
rect 1768 18692 1820 18698
rect 1768 18634 1820 18640
rect 1780 18290 1808 18634
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1492 18216 1544 18222
rect 1492 18158 1544 18164
rect 2332 17882 2360 18566
rect 2608 18290 2636 18770
rect 2596 18284 2648 18290
rect 2596 18226 2648 18232
rect 1860 17876 1912 17882
rect 1860 17818 1912 17824
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1596 16046 1624 16623
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1398 15872 1454 15881
rect 1398 15807 1454 15816
rect 1412 15706 1440 15807
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 14618 1440 14894
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1412 11354 1440 14214
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1504 12782 1532 13262
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1504 12238 1532 12718
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1504 8906 1532 11494
rect 1596 9178 1624 15982
rect 1688 14482 1716 16934
rect 1780 16794 1808 16934
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1872 14074 1900 17818
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 14550 1992 17478
rect 2148 17202 2176 17614
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2148 17082 2176 17138
rect 2056 17054 2176 17082
rect 2056 16794 2084 17054
rect 2516 16998 2544 17682
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 1952 14544 2004 14550
rect 1952 14486 2004 14492
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 2056 13462 2084 16730
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 1858 13152 1914 13161
rect 1858 13087 1914 13096
rect 1872 12986 1900 13087
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 2056 12442 2084 13398
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1780 10606 1808 12038
rect 2148 11880 2176 16934
rect 2332 16674 2360 16934
rect 2608 16810 2636 18226
rect 2884 18193 2912 19654
rect 2976 18698 3004 19858
rect 4080 19514 4108 19858
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 2964 18692 3016 18698
rect 2964 18634 3016 18640
rect 3056 18624 3108 18630
rect 3056 18566 3108 18572
rect 2870 18184 2926 18193
rect 2870 18119 2926 18128
rect 2688 18080 2740 18086
rect 2688 18022 2740 18028
rect 2700 17626 2728 18022
rect 3068 17649 3096 18566
rect 3054 17640 3110 17649
rect 2700 17598 2820 17626
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2056 11852 2176 11880
rect 2240 16646 2360 16674
rect 2516 16782 2636 16810
rect 2412 16652 2464 16658
rect 1950 11792 2006 11801
rect 1950 11727 2006 11736
rect 1964 11694 1992 11727
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 2056 11506 2084 11852
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 1964 11478 2084 11506
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1766 10160 1822 10169
rect 1676 10124 1728 10130
rect 1766 10095 1822 10104
rect 1676 10066 1728 10072
rect 1688 9722 1716 10066
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1492 8900 1544 8906
rect 1492 8842 1544 8848
rect 1504 8430 1532 8842
rect 1780 8498 1808 10095
rect 1964 8514 1992 11478
rect 2148 11354 2176 11698
rect 2240 11354 2268 16646
rect 2412 16594 2464 16600
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 2332 15706 2360 16526
rect 2424 16250 2452 16594
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2412 15972 2464 15978
rect 2412 15914 2464 15920
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2318 15056 2374 15065
rect 2318 14991 2374 15000
rect 2332 14550 2360 14991
rect 2320 14544 2372 14550
rect 2424 14521 2452 15914
rect 2516 15162 2544 16782
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2608 15706 2636 16662
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2608 14906 2636 15302
rect 2700 15026 2728 17478
rect 2792 16794 2820 17598
rect 3054 17575 3110 17584
rect 3160 17542 3188 18770
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 3160 16590 3188 16934
rect 3148 16584 3200 16590
rect 3252 16561 3280 19110
rect 4066 19000 4122 19009
rect 4066 18935 4122 18944
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3712 18426 3740 18702
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3896 18222 3924 18566
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3332 17264 3384 17270
rect 3332 17206 3384 17212
rect 3148 16526 3200 16532
rect 3238 16552 3294 16561
rect 3056 15972 3108 15978
rect 3056 15914 3108 15920
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2792 15065 2820 15506
rect 3068 15502 3096 15914
rect 3160 15910 3188 16526
rect 3238 16487 3294 16496
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2778 15056 2834 15065
rect 2688 15020 2740 15026
rect 2778 14991 2834 15000
rect 2688 14962 2740 14968
rect 2608 14890 2820 14906
rect 2608 14884 2832 14890
rect 2608 14878 2780 14884
rect 2780 14826 2832 14832
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2516 14657 2544 14758
rect 2884 14657 2912 15438
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2502 14648 2558 14657
rect 2502 14583 2558 14592
rect 2870 14648 2926 14657
rect 2870 14583 2926 14592
rect 2320 14486 2372 14492
rect 2410 14512 2466 14521
rect 2410 14447 2466 14456
rect 2412 14340 2464 14346
rect 2412 14282 2464 14288
rect 2318 13968 2374 13977
rect 2318 13903 2320 13912
rect 2372 13903 2374 13912
rect 2320 13874 2372 13880
rect 2424 13462 2452 14282
rect 2976 14278 3004 14758
rect 3068 14550 3096 15438
rect 3056 14544 3108 14550
rect 3056 14486 3108 14492
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 3252 14074 3280 14350
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2412 13456 2464 13462
rect 2412 13398 2464 13404
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2516 12850 2544 13330
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2700 12322 2728 13874
rect 3252 13530 3280 14010
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3252 12986 3280 13466
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 2962 12744 3018 12753
rect 2962 12679 2964 12688
rect 3016 12679 3018 12688
rect 2964 12650 3016 12656
rect 2608 12306 2728 12322
rect 2596 12300 2728 12306
rect 2648 12294 2728 12300
rect 2596 12242 2648 12248
rect 2608 11898 2636 12242
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11354 2544 11494
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 2056 10538 2084 10950
rect 2044 10532 2096 10538
rect 2044 10474 2096 10480
rect 2056 10266 2084 10474
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2056 8974 2084 10202
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2148 8634 2176 11290
rect 2976 11150 3004 11834
rect 3238 11520 3294 11529
rect 3238 11455 3294 11464
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2688 10804 2740 10810
rect 2884 10792 2912 11086
rect 2976 10810 3004 11086
rect 2740 10764 2912 10792
rect 2688 10746 2740 10752
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2332 9926 2360 10542
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2332 9625 2360 9862
rect 2596 9648 2648 9654
rect 2318 9616 2374 9625
rect 2596 9590 2648 9596
rect 2318 9551 2374 9560
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2332 9110 2360 9318
rect 2320 9104 2372 9110
rect 2226 9072 2282 9081
rect 2320 9046 2372 9052
rect 2226 9007 2228 9016
rect 2280 9007 2282 9016
rect 2228 8978 2280 8984
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 1768 8492 1820 8498
rect 1964 8486 2176 8514
rect 1768 8434 1820 8440
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 2044 8288 2096 8294
rect 1398 8256 1454 8265
rect 2044 8230 2096 8236
rect 1398 8191 1454 8200
rect 1412 8090 1440 8191
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1780 7274 1808 7754
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1768 7268 1820 7274
rect 1768 7210 1820 7216
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1596 5574 1624 6258
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1504 4622 1532 5102
rect 1596 4690 1624 5510
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 296 4004 348 4010
rect 296 3946 348 3952
rect 308 480 336 3946
rect 846 2000 902 2009
rect 846 1935 902 1944
rect 860 480 888 1935
rect 1412 480 1440 4014
rect 1504 3534 1532 4558
rect 1688 4282 1716 6054
rect 1780 5234 1808 7210
rect 1872 7206 1900 7686
rect 2056 7410 2084 8230
rect 2148 7993 2176 8486
rect 2608 8090 2636 9590
rect 2700 9518 2728 9930
rect 2884 9761 2912 10764
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 3054 9888 3110 9897
rect 3054 9823 3110 9832
rect 2870 9752 2926 9761
rect 2870 9687 2926 9696
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2700 9042 2728 9318
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2134 7984 2190 7993
rect 2134 7919 2190 7928
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1872 5953 1900 7142
rect 1950 6352 2006 6361
rect 2056 6322 2084 7346
rect 1950 6287 2006 6296
rect 2044 6316 2096 6322
rect 1964 6254 1992 6287
rect 2044 6258 2096 6264
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1858 5944 1914 5953
rect 1964 5914 1992 6190
rect 1858 5879 1914 5888
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 2148 3641 2176 7919
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2516 7206 2544 7822
rect 2792 7426 2820 8366
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2700 7398 2820 7426
rect 2700 7342 2728 7398
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2504 7200 2556 7206
rect 2502 7168 2504 7177
rect 2556 7168 2558 7177
rect 2502 7103 2558 7112
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2608 5930 2636 6802
rect 2700 6662 2728 7278
rect 2884 6730 2912 8298
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2976 7478 3004 8026
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2870 6624 2926 6633
rect 2792 6254 2820 6598
rect 2870 6559 2926 6568
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2608 5902 2728 5930
rect 2700 5846 2728 5902
rect 2596 5840 2648 5846
rect 2596 5782 2648 5788
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2228 5636 2280 5642
rect 2228 5578 2280 5584
rect 2240 4146 2268 5578
rect 2424 5030 2452 5646
rect 2608 5030 2636 5782
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2240 3670 2268 4082
rect 2228 3664 2280 3670
rect 2134 3632 2190 3641
rect 2228 3606 2280 3612
rect 2134 3567 2190 3576
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1504 2514 1532 3470
rect 2240 3194 2268 3606
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 1674 3088 1730 3097
rect 1674 3023 1730 3032
rect 1688 2922 1716 3023
rect 1950 2952 2006 2961
rect 1676 2916 1728 2922
rect 1950 2887 2006 2896
rect 1676 2858 1728 2864
rect 1688 2582 1716 2858
rect 1676 2576 1728 2582
rect 1676 2518 1728 2524
rect 1492 2508 1544 2514
rect 1492 2450 1544 2456
rect 1964 480 1992 2887
rect 2424 1578 2452 4966
rect 2608 4865 2636 4966
rect 2594 4856 2650 4865
rect 2594 4791 2650 4800
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2608 3738 2636 4626
rect 2884 4128 2912 6559
rect 2792 4100 2912 4128
rect 2686 3904 2742 3913
rect 2686 3839 2742 3848
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2700 3194 2728 3839
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2792 2145 2820 4100
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2884 3738 2912 3946
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 2884 2650 2912 3062
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 2502 1592 2558 1601
rect 2424 1550 2502 1578
rect 2502 1527 2558 1536
rect 2516 480 2544 1527
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 2976 377 3004 7414
rect 3068 6905 3096 9823
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3160 7886 3188 8230
rect 3252 7886 3280 11455
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3160 7274 3188 7822
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7546 3280 7686
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3160 7002 3188 7210
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3054 6896 3110 6905
rect 3054 6831 3110 6840
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3068 4185 3096 6666
rect 3160 6458 3188 6938
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3160 5914 3188 6258
rect 3252 6254 3280 7482
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3238 5944 3294 5953
rect 3148 5908 3200 5914
rect 3238 5879 3294 5888
rect 3148 5850 3200 5856
rect 3160 5166 3188 5850
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3160 4826 3188 5102
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3054 4176 3110 4185
rect 3054 4111 3110 4120
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3068 2990 3096 3470
rect 3160 3058 3188 3674
rect 3252 3233 3280 5879
rect 3344 4146 3372 17206
rect 3436 17134 3464 17478
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3974 17096 4030 17105
rect 3436 16046 3464 17070
rect 3974 17031 4030 17040
rect 3792 16720 3844 16726
rect 3790 16688 3792 16697
rect 3844 16688 3846 16697
rect 3790 16623 3846 16632
rect 3698 16416 3754 16425
rect 3698 16351 3754 16360
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 3436 12481 3464 13631
rect 3606 13016 3662 13025
rect 3606 12951 3662 12960
rect 3514 12608 3570 12617
rect 3514 12543 3570 12552
rect 3422 12472 3478 12481
rect 3422 12407 3478 12416
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3436 11218 3464 11766
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3436 10810 3464 11154
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3436 8514 3464 10746
rect 3528 10577 3556 12543
rect 3514 10568 3570 10577
rect 3514 10503 3570 10512
rect 3514 9616 3570 9625
rect 3514 9551 3570 9560
rect 3528 9518 3556 9551
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3528 9194 3556 9454
rect 3620 9353 3648 12951
rect 3712 11393 3740 16351
rect 3988 16153 4016 17031
rect 4080 16794 4108 18935
rect 4172 18290 4200 19246
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 4250 18728 4306 18737
rect 4250 18663 4252 18672
rect 4304 18663 4306 18672
rect 4252 18634 4304 18640
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4264 17542 4292 18158
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 3974 16144 4030 16153
rect 3974 16079 4030 16088
rect 3790 16008 3846 16017
rect 3790 15943 3846 15952
rect 3804 12209 3832 15943
rect 4080 15706 4108 16594
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4080 15178 4108 15438
rect 4080 15150 4200 15178
rect 4264 15162 4292 15574
rect 4172 15026 4200 15150
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4356 14074 4384 18906
rect 4448 18193 4476 22335
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4618 19408 4674 19417
rect 4618 19343 4674 19352
rect 4632 19174 4660 19343
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4434 18184 4490 18193
rect 4434 18119 4490 18128
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4448 16794 4476 17478
rect 4632 16794 4660 17682
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4448 16250 4476 16594
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4528 14884 4580 14890
rect 4528 14826 4580 14832
rect 4540 14346 4568 14826
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4632 13977 4660 16730
rect 4816 16658 4844 19790
rect 5460 19700 5488 26658
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 24766 25120 24822 25129
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 24289 25052 24585 25072
rect 24766 25055 24822 25064
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 11978 24168 12034 24177
rect 11978 24103 12034 24112
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 10782 22536 10838 22545
rect 10782 22471 10838 22480
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 8574 21992 8630 22001
rect 8574 21927 8630 21936
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 8588 21690 8616 21927
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 7300 21457 7328 21490
rect 8760 21480 8812 21486
rect 7286 21448 7342 21457
rect 8760 21422 8812 21428
rect 7286 21383 7342 21392
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 7378 20088 7434 20097
rect 7378 20023 7434 20032
rect 7392 19990 7420 20023
rect 7380 19984 7432 19990
rect 7380 19926 7432 19932
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 5092 19672 5488 19700
rect 6920 19712 6972 19718
rect 4988 18148 5040 18154
rect 4988 18090 5040 18096
rect 5000 17678 5028 18090
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 5000 17338 5028 17614
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4908 14618 4936 14758
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 5092 14056 5120 19672
rect 6920 19654 6972 19660
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6932 19378 6960 19654
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 6472 19174 6500 19246
rect 6460 19168 6512 19174
rect 6828 19168 6880 19174
rect 6460 19110 6512 19116
rect 6826 19136 6828 19145
rect 6880 19136 6882 19145
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5552 18086 5580 18838
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5540 18080 5592 18086
rect 5460 18028 5540 18034
rect 5460 18022 5592 18028
rect 5460 18006 5580 18022
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5368 16998 5396 17682
rect 5356 16992 5408 16998
rect 5262 16960 5318 16969
rect 5356 16934 5408 16940
rect 5262 16895 5318 16904
rect 5276 16794 5304 16895
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5368 16697 5396 16934
rect 5354 16688 5410 16697
rect 5354 16623 5410 16632
rect 5460 16590 5488 18006
rect 6000 17604 6052 17610
rect 6000 17546 6052 17552
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6012 17202 6040 17546
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6012 16794 6040 17138
rect 6472 16794 6500 19110
rect 6826 19071 6882 19080
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6748 17814 6776 18566
rect 7392 17882 7420 19314
rect 7668 19174 7696 19858
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7668 18426 7696 19110
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7852 17882 7880 21286
rect 7932 21004 7984 21010
rect 7932 20946 7984 20952
rect 7944 20262 7972 20946
rect 8116 20936 8168 20942
rect 8114 20904 8116 20913
rect 8168 20904 8170 20913
rect 8114 20839 8170 20848
rect 8772 20466 8800 21422
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6748 17338 6776 17750
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5460 16250 5488 16526
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5552 16046 5580 16594
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6090 16416 6146 16425
rect 5622 16348 5918 16368
rect 6090 16351 6146 16360
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5092 14028 5212 14056
rect 4804 14000 4856 14006
rect 4250 13968 4306 13977
rect 4250 13903 4306 13912
rect 4618 13968 4674 13977
rect 4804 13942 4856 13948
rect 4618 13903 4674 13912
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3790 12200 3846 12209
rect 3790 12135 3846 12144
rect 3884 12096 3936 12102
rect 3790 12064 3846 12073
rect 3884 12038 3936 12044
rect 3790 11999 3846 12008
rect 3804 11642 3832 11999
rect 3896 11762 3924 12038
rect 4080 11830 4108 13806
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3976 11688 4028 11694
rect 3804 11614 3924 11642
rect 3976 11630 4028 11636
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3698 11384 3754 11393
rect 3698 11319 3754 11328
rect 3698 10432 3754 10441
rect 3698 10367 3754 10376
rect 3606 9344 3662 9353
rect 3606 9279 3662 9288
rect 3528 9166 3648 9194
rect 3436 8486 3556 8514
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3436 6730 3464 8366
rect 3528 8090 3556 8486
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3514 6896 3570 6905
rect 3514 6831 3570 6840
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3528 6390 3556 6831
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3436 4826 3464 6122
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3528 5681 3556 6054
rect 3514 5672 3570 5681
rect 3514 5607 3570 5616
rect 3514 4856 3570 4865
rect 3424 4820 3476 4826
rect 3620 4826 3648 9166
rect 3712 8650 3740 10367
rect 3804 9042 3832 11494
rect 3896 10441 3924 11614
rect 3988 11286 4016 11630
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3882 10432 3938 10441
rect 3882 10367 3938 10376
rect 4080 10266 4108 11290
rect 4172 11218 4200 12582
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4158 10568 4214 10577
rect 4158 10503 4214 10512
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3896 9178 3924 9386
rect 3974 9208 4030 9217
rect 3884 9172 3936 9178
rect 4080 9178 4108 10066
rect 3974 9143 4030 9152
rect 4068 9172 4120 9178
rect 3884 9114 3936 9120
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3712 8622 3832 8650
rect 3896 8634 3924 9114
rect 3698 8392 3754 8401
rect 3698 8327 3754 8336
rect 3514 4791 3570 4800
rect 3608 4820 3660 4826
rect 3424 4762 3476 4768
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3238 3224 3294 3233
rect 3528 3210 3556 4791
rect 3608 4762 3660 4768
rect 3606 4448 3662 4457
rect 3606 4383 3662 4392
rect 3238 3159 3294 3168
rect 3436 3182 3556 3210
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 3054 2816 3110 2825
rect 3054 2751 3110 2760
rect 3068 480 3096 2751
rect 3436 1442 3464 3182
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3528 2310 3556 2994
rect 3620 2553 3648 4383
rect 3606 2544 3662 2553
rect 3606 2479 3662 2488
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3712 1465 3740 8327
rect 3804 6610 3832 8622
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3988 8129 4016 9143
rect 4068 9114 4120 9120
rect 4172 8945 4200 10503
rect 4264 9178 4292 13903
rect 4620 13728 4672 13734
rect 4712 13728 4764 13734
rect 4620 13670 4672 13676
rect 4710 13696 4712 13705
rect 4764 13696 4766 13705
rect 4632 13190 4660 13670
rect 4710 13631 4766 13640
rect 4724 13530 4752 13631
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4620 13184 4672 13190
rect 4618 13152 4620 13161
rect 4672 13152 4674 13161
rect 4618 13087 4674 13096
rect 4620 12708 4672 12714
rect 4724 12696 4752 13262
rect 4672 12668 4752 12696
rect 4620 12650 4672 12656
rect 4632 12306 4660 12650
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 11801 4384 12038
rect 4342 11792 4398 11801
rect 4342 11727 4398 11736
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4448 10577 4476 11290
rect 4632 11150 4660 11698
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4434 10568 4490 10577
rect 4434 10503 4490 10512
rect 4448 10470 4476 10503
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4356 9382 4384 10134
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4158 8936 4214 8945
rect 4158 8871 4214 8880
rect 4264 8634 4292 9114
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4264 8401 4292 8570
rect 4250 8392 4306 8401
rect 4250 8327 4306 8336
rect 3974 8120 4030 8129
rect 3974 8055 4030 8064
rect 3882 7576 3938 7585
rect 3882 7511 3938 7520
rect 3896 6905 3924 7511
rect 4356 7478 4384 9318
rect 3976 7472 4028 7478
rect 4344 7472 4396 7478
rect 3976 7414 4028 7420
rect 4342 7440 4344 7449
rect 4396 7440 4398 7449
rect 3882 6896 3938 6905
rect 3988 6866 4016 7414
rect 4342 7375 4398 7384
rect 4448 7290 4476 10406
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4540 9722 4568 9998
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4632 9450 4660 11086
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4724 10606 4752 10950
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4632 9178 4660 9386
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4816 9042 4844 13942
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5092 13394 5120 13874
rect 5184 13546 5212 14028
rect 5276 13938 5304 14418
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5368 13870 5396 14350
rect 5356 13864 5408 13870
rect 5354 13832 5356 13841
rect 5408 13832 5410 13841
rect 5354 13767 5410 13776
rect 5184 13518 5396 13546
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 4908 12918 4936 13330
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4908 12374 4936 12854
rect 5092 12646 5120 13330
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 4908 11898 4936 12310
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 5172 11688 5224 11694
rect 5276 11676 5304 13518
rect 5368 13394 5396 13518
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5460 11694 5488 15914
rect 5552 12986 5580 15982
rect 6104 15910 6132 16351
rect 6564 15910 6592 16526
rect 6656 16425 6684 16594
rect 6748 16522 6776 17274
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6840 16794 6868 17138
rect 7392 17066 7420 17818
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6826 16552 6882 16561
rect 6736 16516 6788 16522
rect 6826 16487 6882 16496
rect 6736 16458 6788 16464
rect 6642 16416 6698 16425
rect 6642 16351 6698 16360
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5998 14920 6054 14929
rect 5998 14855 6054 14864
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5722 13968 5778 13977
rect 5722 13903 5724 13912
rect 5776 13903 5778 13912
rect 5724 13874 5776 13880
rect 6012 13433 6040 14855
rect 5998 13424 6054 13433
rect 5998 13359 6054 13368
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 12442 5580 12582
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5538 12200 5594 12209
rect 5538 12135 5594 12144
rect 5552 11898 5580 12135
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5224 11648 5304 11676
rect 5448 11688 5500 11694
rect 5172 11630 5224 11636
rect 5448 11630 5500 11636
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 4816 8022 4844 8978
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4356 7262 4476 7290
rect 4066 7032 4122 7041
rect 4066 6967 4122 6976
rect 3882 6831 3938 6840
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4080 6746 4108 6967
rect 4160 6792 4212 6798
rect 4080 6740 4160 6746
rect 4080 6734 4212 6740
rect 4080 6718 4200 6734
rect 4252 6656 4304 6662
rect 3804 6582 4016 6610
rect 4252 6598 4304 6604
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3804 4593 3832 6326
rect 3882 4720 3938 4729
rect 3882 4655 3938 4664
rect 3790 4584 3846 4593
rect 3790 4519 3846 4528
rect 3896 3618 3924 4655
rect 3804 3590 3924 3618
rect 3698 1456 3754 1465
rect 3436 1414 3648 1442
rect 3620 480 3648 1414
rect 3698 1391 3754 1400
rect 3804 921 3832 3590
rect 3882 3496 3938 3505
rect 3882 3431 3884 3440
rect 3936 3431 3938 3440
rect 3884 3402 3936 3408
rect 3988 1737 4016 6582
rect 4068 6384 4120 6390
rect 4264 6361 4292 6598
rect 4068 6326 4120 6332
rect 4250 6352 4306 6361
rect 4080 3738 4108 6326
rect 4250 6287 4306 6296
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4172 4457 4200 6190
rect 4356 5953 4384 7262
rect 4724 7177 4752 7686
rect 4526 7168 4582 7177
rect 4526 7103 4582 7112
rect 4710 7168 4766 7177
rect 4710 7103 4766 7112
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 4448 6254 4476 6938
rect 4540 6746 4568 7103
rect 4816 7002 4844 7958
rect 5000 7002 5028 11494
rect 5814 11384 5870 11393
rect 5814 11319 5816 11328
rect 5868 11319 5870 11328
rect 5816 11290 5868 11296
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 5092 10674 5120 10950
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5092 9722 5120 10610
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 10062 5212 10406
rect 5172 10056 5224 10062
rect 5170 10024 5172 10033
rect 5224 10024 5226 10033
rect 5170 9959 5226 9968
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5092 9518 5120 9658
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5276 9081 5304 10678
rect 5368 10470 5396 11154
rect 5448 11144 5500 11150
rect 5500 11092 5580 11098
rect 5448 11086 5580 11092
rect 5460 11070 5580 11086
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5460 10606 5488 10950
rect 5552 10810 5580 11070
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10305 5396 10406
rect 5354 10296 5410 10305
rect 5354 10231 5410 10240
rect 5552 10198 5580 10746
rect 5540 10192 5592 10198
rect 6012 10169 6040 11154
rect 6104 10266 6132 15846
rect 6564 15337 6592 15846
rect 6748 15706 6776 16458
rect 6840 16250 6868 16487
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6932 16114 6960 16662
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7010 16144 7066 16153
rect 6920 16108 6972 16114
rect 7484 16114 7512 16390
rect 7010 16079 7066 16088
rect 7472 16108 7524 16114
rect 6920 16050 6972 16056
rect 6932 15706 6960 16050
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6828 15360 6880 15366
rect 6550 15328 6606 15337
rect 6828 15302 6880 15308
rect 6550 15263 6606 15272
rect 6274 15192 6330 15201
rect 6274 15127 6276 15136
rect 6328 15127 6330 15136
rect 6276 15098 6328 15104
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 13734 6224 14350
rect 6288 14006 6316 15098
rect 6840 15065 6868 15302
rect 6826 15056 6882 15065
rect 6826 14991 6882 15000
rect 6840 14958 6868 14991
rect 6828 14952 6880 14958
rect 6458 14920 6514 14929
rect 6828 14894 6880 14900
rect 6458 14855 6514 14864
rect 6736 14884 6788 14890
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 13530 6224 13670
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6184 12708 6236 12714
rect 6184 12650 6236 12656
rect 6196 11830 6224 12650
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6380 11898 6408 12242
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6274 10296 6330 10305
rect 6092 10260 6144 10266
rect 6144 10240 6274 10248
rect 6144 10231 6330 10240
rect 6144 10220 6316 10231
rect 6092 10202 6144 10208
rect 5540 10134 5592 10140
rect 5630 10160 5686 10169
rect 5630 10095 5632 10104
rect 5684 10095 5686 10104
rect 5998 10160 6054 10169
rect 5998 10095 6054 10104
rect 5632 10066 5684 10072
rect 6104 10044 6132 10202
rect 6012 10016 6132 10044
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5446 9752 5502 9761
rect 5622 9744 5918 9764
rect 5502 9710 5580 9738
rect 5446 9687 5502 9696
rect 5262 9072 5318 9081
rect 5262 9007 5318 9016
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5184 8634 5212 8774
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5184 8362 5212 8570
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5276 8022 5304 9007
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5552 8514 5580 9710
rect 6012 9382 6040 10016
rect 6472 9994 6500 14855
rect 6736 14826 6788 14832
rect 6644 14816 6696 14822
rect 6642 14784 6644 14793
rect 6696 14784 6698 14793
rect 6642 14719 6698 14728
rect 6748 14618 6776 14826
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6550 14512 6606 14521
rect 6840 14482 6868 14894
rect 6550 14447 6606 14456
rect 6828 14476 6880 14482
rect 6564 14074 6592 14447
rect 6828 14418 6880 14424
rect 7024 14074 7052 16079
rect 7472 16050 7524 16056
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 7208 15881 7236 15914
rect 7194 15872 7250 15881
rect 7194 15807 7250 15816
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7392 15201 7420 15506
rect 7378 15192 7434 15201
rect 7484 15162 7512 16050
rect 7760 15502 7788 16934
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7378 15127 7434 15136
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7484 14550 7512 15098
rect 7576 14793 7604 15438
rect 7760 14890 7788 15438
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7562 14784 7618 14793
rect 7562 14719 7618 14728
rect 7838 14648 7894 14657
rect 7838 14583 7894 14592
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 7484 14074 7512 14486
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 6564 13870 6592 14010
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 7378 13832 7434 13841
rect 7378 13767 7434 13776
rect 7286 13696 7342 13705
rect 7286 13631 7342 13640
rect 7300 13530 7328 13631
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6564 12850 6592 13330
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6932 12646 6960 13126
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6736 12096 6788 12102
rect 6642 12064 6698 12073
rect 6736 12038 6788 12044
rect 6642 11999 6698 12008
rect 6656 11694 6684 11999
rect 6748 11830 6776 12038
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6550 10432 6606 10441
rect 6550 10367 6606 10376
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6472 9722 6500 9930
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5460 8090 5488 8502
rect 5552 8486 5672 8514
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5264 8016 5316 8022
rect 5644 8004 5672 8486
rect 5722 8392 5778 8401
rect 5722 8327 5724 8336
rect 5776 8327 5778 8336
rect 5724 8298 5776 8304
rect 5264 7958 5316 7964
rect 5552 7976 5672 8004
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5276 7546 5304 7822
rect 5264 7540 5316 7546
rect 5184 7500 5264 7528
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 4802 6896 4858 6905
rect 4802 6831 4858 6840
rect 4540 6718 4752 6746
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4632 6497 4660 6598
rect 4618 6488 4674 6497
rect 4618 6423 4674 6432
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4342 5944 4398 5953
rect 4342 5879 4398 5888
rect 4448 4554 4476 6054
rect 4540 5370 4568 6258
rect 4632 6254 4660 6423
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4252 4480 4304 4486
rect 4158 4448 4214 4457
rect 4252 4422 4304 4428
rect 4158 4383 4214 4392
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4172 3194 4200 4218
rect 4264 4146 4292 4422
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4448 3074 4476 4490
rect 4540 3641 4568 5306
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4526 3632 4582 3641
rect 4526 3567 4582 3576
rect 4172 3046 4476 3074
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4080 2514 4108 2926
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 3974 1728 4030 1737
rect 3974 1663 4030 1672
rect 3790 912 3846 921
rect 3790 847 3846 856
rect 4172 480 4200 3046
rect 4540 2582 4568 3567
rect 4632 3505 4660 4626
rect 4618 3496 4674 3505
rect 4618 3431 4674 3440
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 4724 480 4752 6718
rect 4816 5817 4844 6831
rect 5184 6730 5212 7500
rect 5264 7482 5316 7488
rect 5368 7274 5396 7890
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5448 6996 5500 7002
rect 5368 6934 5396 6965
rect 5448 6938 5500 6944
rect 5356 6928 5408 6934
rect 5276 6876 5356 6882
rect 5276 6870 5408 6876
rect 5276 6854 5396 6870
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5184 5914 5212 6666
rect 5276 6202 5304 6854
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5368 6458 5396 6734
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5276 6186 5396 6202
rect 5276 6180 5408 6186
rect 5276 6174 5356 6180
rect 5356 6122 5408 6128
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 4802 5808 4858 5817
rect 4802 5743 4858 5752
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4908 5166 4936 5714
rect 5368 5234 5396 6122
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4816 4282 4844 4558
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4908 3398 4936 4626
rect 5368 4486 5396 5034
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5092 3942 5120 4422
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 4988 3936 5040 3942
rect 5080 3936 5132 3942
rect 4988 3878 5040 3884
rect 5078 3904 5080 3913
rect 5132 3904 5134 3913
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4908 2689 4936 3334
rect 4894 2680 4950 2689
rect 4894 2615 4950 2624
rect 5000 2417 5028 3878
rect 5078 3839 5134 3848
rect 5184 3738 5212 4082
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5276 3670 5304 4082
rect 5264 3664 5316 3670
rect 5184 3612 5264 3618
rect 5184 3606 5316 3612
rect 5184 3590 5304 3606
rect 5368 3602 5396 4422
rect 5356 3596 5408 3602
rect 5184 3194 5212 3590
rect 5356 3538 5408 3544
rect 5460 3482 5488 6938
rect 5276 3454 5488 3482
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4986 2408 5042 2417
rect 4986 2343 5042 2352
rect 5276 480 5304 3454
rect 5552 1034 5580 7976
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5644 6866 5672 7414
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5736 7041 5764 7142
rect 5722 7032 5778 7041
rect 5722 6967 5778 6976
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 6012 6769 6040 9318
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6104 8634 6132 8978
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6092 7744 6144 7750
rect 6090 7712 6092 7721
rect 6144 7712 6146 7721
rect 6090 7647 6146 7656
rect 6196 7585 6224 7754
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6182 7576 6238 7585
rect 6182 7511 6238 7520
rect 6196 7342 6224 7511
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6092 7268 6144 7274
rect 6092 7210 6144 7216
rect 5998 6760 6054 6769
rect 5998 6695 6054 6704
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6254 6040 6598
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6104 4826 6132 7210
rect 6182 6896 6238 6905
rect 6182 6831 6238 6840
rect 6196 5166 6224 6831
rect 6288 6769 6316 7686
rect 6380 6866 6408 9046
rect 6472 9042 6500 9386
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6564 8242 6592 10367
rect 6748 10010 6776 11766
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6840 11218 6868 11630
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6932 10810 6960 12582
rect 7116 12442 7144 12650
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7024 11082 7052 12174
rect 7208 12170 7236 12786
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 7116 11286 7144 11562
rect 7104 11280 7156 11286
rect 7102 11248 7104 11257
rect 7156 11248 7158 11257
rect 7102 11183 7158 11192
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7024 10266 7052 11018
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6748 9994 7052 10010
rect 6748 9988 7064 9994
rect 6748 9982 7012 9988
rect 6642 9616 6698 9625
rect 6642 9551 6698 9560
rect 6472 8214 6592 8242
rect 6472 7970 6500 8214
rect 6550 8120 6606 8129
rect 6550 8055 6552 8064
rect 6604 8055 6606 8064
rect 6552 8026 6604 8032
rect 6472 7942 6592 7970
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6274 6760 6330 6769
rect 6274 6695 6330 6704
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6012 4214 6040 4490
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 6104 4010 6132 4626
rect 6196 4554 6224 5102
rect 6366 4992 6422 5001
rect 6366 4927 6422 4936
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 6196 4282 6224 4490
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6288 4078 6316 4558
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 6288 3777 6316 4014
rect 6274 3768 6330 3777
rect 6274 3703 6330 3712
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5552 1006 5856 1034
rect 5828 480 5856 1006
rect 6380 480 6408 4927
rect 6472 4690 6500 7482
rect 6564 6225 6592 7942
rect 6550 6216 6606 6225
rect 6550 6151 6606 6160
rect 6656 4729 6684 9551
rect 6748 9518 6776 9982
rect 7012 9930 7064 9936
rect 7116 9926 7144 10474
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7116 9722 7144 9862
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6920 9444 6972 9450
rect 7208 9432 7236 12106
rect 7288 10464 7340 10470
rect 7286 10432 7288 10441
rect 7340 10432 7342 10441
rect 7286 10367 7342 10376
rect 6972 9404 7236 9432
rect 6920 9386 6972 9392
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 7546 6776 7822
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 5914 6776 6802
rect 6828 6112 6880 6118
rect 6826 6080 6828 6089
rect 6880 6080 6882 6089
rect 6826 6015 6882 6024
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6642 4720 6698 4729
rect 6460 4684 6512 4690
rect 6642 4655 6698 4664
rect 6460 4626 6512 4632
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6748 3738 6776 4218
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6550 3632 6606 3641
rect 6550 3567 6606 3576
rect 6564 3194 6592 3567
rect 6932 3346 6960 8434
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 7024 7546 7052 7958
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 5846 7144 6598
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 7116 5710 7144 5782
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7010 5264 7066 5273
rect 7010 5199 7066 5208
rect 7024 4146 7052 5199
rect 7208 5137 7236 8298
rect 7286 7984 7342 7993
rect 7286 7919 7288 7928
rect 7340 7919 7342 7928
rect 7288 7890 7340 7896
rect 7300 7546 7328 7890
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7286 7168 7342 7177
rect 7286 7103 7342 7112
rect 7300 6322 7328 7103
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7300 5914 7328 6258
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7194 5128 7250 5137
rect 7194 5063 7250 5072
rect 7288 5092 7340 5098
rect 7208 4865 7236 5063
rect 7288 5034 7340 5040
rect 7194 4856 7250 4865
rect 7194 4791 7250 4800
rect 7300 4554 7328 5034
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7300 4146 7328 4490
rect 7012 4140 7064 4146
rect 7288 4140 7340 4146
rect 7012 4082 7064 4088
rect 7116 4100 7288 4128
rect 6932 3318 7052 3346
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6564 2854 6592 3130
rect 6932 2961 6960 3130
rect 6918 2952 6974 2961
rect 6918 2887 6974 2896
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6918 2680 6974 2689
rect 6918 2615 6920 2624
rect 6972 2615 6974 2624
rect 6920 2586 6972 2592
rect 6642 2544 6698 2553
rect 6642 2479 6644 2488
rect 6696 2479 6698 2488
rect 6644 2450 6696 2456
rect 7024 1601 7052 3318
rect 7116 3058 7144 4100
rect 7288 4082 7340 4088
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7208 3641 7236 3878
rect 7288 3664 7340 3670
rect 7194 3632 7250 3641
rect 7288 3606 7340 3612
rect 7194 3567 7250 3576
rect 7300 3194 7328 3606
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7102 2952 7158 2961
rect 7102 2887 7104 2896
rect 7156 2887 7158 2896
rect 7104 2858 7156 2864
rect 7010 1592 7066 1601
rect 7010 1527 7066 1536
rect 7392 1306 7420 13767
rect 7656 13252 7708 13258
rect 7656 13194 7708 13200
rect 7668 12646 7696 13194
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7484 11626 7512 12106
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7484 10674 7512 11562
rect 7562 10704 7618 10713
rect 7472 10668 7524 10674
rect 7562 10639 7618 10648
rect 7472 10610 7524 10616
rect 7484 9518 7512 10610
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 9353 7512 9454
rect 7470 9344 7526 9353
rect 7470 9279 7526 9288
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7484 7750 7512 8434
rect 7576 7993 7604 10639
rect 7562 7984 7618 7993
rect 7562 7919 7618 7928
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 6905 7512 7686
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7470 6896 7526 6905
rect 7470 6831 7526 6840
rect 7576 6730 7604 7278
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7472 6656 7524 6662
rect 7576 6633 7604 6666
rect 7472 6598 7524 6604
rect 7562 6624 7618 6633
rect 7484 6322 7512 6598
rect 7562 6559 7618 6568
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7484 6186 7512 6258
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7484 5846 7512 6122
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7484 5370 7512 5782
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4049 7512 4966
rect 7576 4826 7604 5034
rect 7668 5001 7696 12582
rect 7760 11257 7788 14214
rect 7852 12866 7880 14583
rect 7944 14074 7972 20198
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 8036 18222 8064 18702
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 8220 18329 8248 18566
rect 8206 18320 8262 18329
rect 8206 18255 8208 18264
rect 8260 18255 8262 18264
rect 8208 18226 8260 18232
rect 8024 18216 8076 18222
rect 8220 18195 8248 18226
rect 9324 18222 9352 18566
rect 9312 18216 9364 18222
rect 8024 18158 8076 18164
rect 9312 18158 9364 18164
rect 8116 18080 8168 18086
rect 8114 18048 8116 18057
rect 8168 18048 8170 18057
rect 8114 17983 8170 17992
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 8036 16794 8064 17818
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8772 16998 8800 17682
rect 9324 17610 9352 18158
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9324 17202 9352 17546
rect 9312 17196 9364 17202
rect 9140 17156 9312 17184
rect 8760 16992 8812 16998
rect 8758 16960 8760 16969
rect 8812 16960 8814 16969
rect 8758 16895 8814 16904
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8114 16552 8170 16561
rect 8114 16487 8170 16496
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7944 12986 7972 13262
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7852 12838 7972 12866
rect 7838 11792 7894 11801
rect 7838 11727 7894 11736
rect 7746 11248 7802 11257
rect 7746 11183 7802 11192
rect 7852 8090 7880 11727
rect 7944 8276 7972 12838
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 11286 8064 11494
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 8036 10577 8064 11222
rect 8022 10568 8078 10577
rect 8022 10503 8024 10512
rect 8076 10503 8078 10512
rect 8024 10474 8076 10480
rect 8022 8664 8078 8673
rect 8022 8599 8078 8608
rect 8036 8401 8064 8599
rect 8022 8392 8078 8401
rect 8022 8327 8078 8336
rect 7944 8248 8064 8276
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7746 7848 7802 7857
rect 7746 7783 7748 7792
rect 7800 7783 7802 7792
rect 7932 7812 7984 7818
rect 7748 7754 7800 7760
rect 7932 7754 7984 7760
rect 7760 7342 7788 7754
rect 7944 7449 7972 7754
rect 7930 7440 7986 7449
rect 7930 7375 7986 7384
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7760 7002 7788 7278
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7944 6458 7972 7375
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 8036 5114 8064 8248
rect 7760 5086 8064 5114
rect 7654 4992 7710 5001
rect 7654 4927 7710 4936
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7470 4040 7526 4049
rect 7470 3975 7526 3984
rect 7472 3528 7524 3534
rect 7760 3482 7788 5086
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7838 4720 7894 4729
rect 7838 4655 7840 4664
rect 7892 4655 7894 4664
rect 7840 4626 7892 4632
rect 7472 3470 7524 3476
rect 7484 2854 7512 3470
rect 7576 3454 7788 3482
rect 7838 3496 7894 3505
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7484 2446 7512 2790
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 6932 1278 7420 1306
rect 6932 480 6960 1278
rect 7576 480 7604 3454
rect 7838 3431 7840 3440
rect 7892 3431 7894 3440
rect 7840 3402 7892 3408
rect 7944 2938 7972 4966
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 8036 4214 8064 4558
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7852 2910 7972 2938
rect 7852 1737 7880 2910
rect 7930 2816 7986 2825
rect 8036 2802 8064 3470
rect 7986 2774 8064 2802
rect 7930 2751 7986 2760
rect 7944 2650 7972 2751
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 7838 1728 7894 1737
rect 7838 1663 7894 1672
rect 8128 480 8156 16487
rect 8312 16250 8340 16662
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8404 15348 8432 16526
rect 8496 15706 8524 16594
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8680 16250 8708 16526
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 9140 16114 9168 17156
rect 9312 17138 9364 17144
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8944 15428 8996 15434
rect 8944 15370 8996 15376
rect 8484 15360 8536 15366
rect 8404 15320 8484 15348
rect 8484 15302 8536 15308
rect 8496 15065 8524 15302
rect 8482 15056 8538 15065
rect 8482 14991 8538 15000
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 8404 13938 8432 14826
rect 8496 14618 8524 14991
rect 8850 14920 8906 14929
rect 8850 14855 8906 14864
rect 8864 14822 8892 14855
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8956 14550 8984 15370
rect 9140 15366 9168 16050
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9140 14958 9168 15302
rect 9218 15056 9274 15065
rect 9218 14991 9220 15000
rect 9272 14991 9274 15000
rect 9220 14962 9272 14968
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 8956 14346 8984 14486
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 9048 14074 9076 14418
rect 9140 14414 9168 14894
rect 9218 14784 9274 14793
rect 9218 14719 9274 14728
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 8942 13968 8998 13977
rect 8392 13932 8444 13938
rect 8942 13903 8944 13912
rect 8392 13874 8444 13880
rect 8996 13903 8998 13912
rect 8944 13874 8996 13880
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8220 12617 8248 13330
rect 8312 13297 8340 13670
rect 8404 13530 8432 13874
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8298 13288 8354 13297
rect 8298 13223 8354 13232
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8588 12646 8616 13126
rect 8392 12640 8444 12646
rect 8206 12608 8262 12617
rect 8392 12582 8444 12588
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8206 12543 8262 12552
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8220 12186 8248 12242
rect 8220 12158 8340 12186
rect 8208 10192 8260 10198
rect 8206 10160 8208 10169
rect 8260 10160 8262 10169
rect 8206 10095 8262 10104
rect 8220 9110 8248 10095
rect 8312 9178 8340 12158
rect 8404 11801 8432 12582
rect 8588 12170 8616 12582
rect 9048 12306 9076 14010
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8588 11937 8616 12106
rect 8668 12096 8720 12102
rect 8666 12064 8668 12073
rect 8720 12064 8722 12073
rect 8666 11999 8722 12008
rect 8574 11928 8630 11937
rect 8574 11863 8630 11872
rect 8390 11792 8446 11801
rect 8390 11727 8446 11736
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 11218 8524 11494
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8390 10704 8446 10713
rect 8390 10639 8446 10648
rect 8404 10266 8432 10639
rect 8496 10606 8524 11154
rect 9048 11082 9076 12242
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8404 9722 8432 10202
rect 8496 9926 8524 10542
rect 8772 10538 8800 10950
rect 8760 10532 8812 10538
rect 8760 10474 8812 10480
rect 8772 10169 8800 10474
rect 8758 10160 8814 10169
rect 8758 10095 8814 10104
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8220 8430 8248 9046
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8206 8256 8262 8265
rect 8206 8191 8262 8200
rect 8220 8090 8248 8191
rect 8208 8084 8260 8090
rect 8260 8044 8340 8072
rect 8208 8026 8260 8032
rect 8312 6866 8340 8044
rect 8404 7585 8432 8502
rect 8496 8090 8524 9862
rect 8864 9178 8892 9998
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8864 8362 8892 9114
rect 9048 8634 9076 11018
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8390 7576 8446 7585
rect 8390 7511 8446 7520
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8574 6624 8630 6633
rect 8574 6559 8630 6568
rect 8588 6254 8616 6559
rect 8864 6254 8892 7142
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8298 5264 8354 5273
rect 8298 5199 8354 5208
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8220 3097 8248 5102
rect 8312 4826 8340 5199
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8392 4616 8444 4622
rect 8576 4616 8628 4622
rect 8444 4576 8524 4604
rect 8392 4558 8444 4564
rect 8300 3936 8352 3942
rect 8352 3896 8432 3924
rect 8300 3878 8352 3884
rect 8206 3088 8262 3097
rect 8206 3023 8262 3032
rect 8404 2922 8432 3896
rect 8496 3505 8524 4576
rect 8576 4558 8628 4564
rect 8588 4010 8616 4558
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 8588 3738 8616 3946
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8588 3534 8616 3674
rect 8576 3528 8628 3534
rect 8482 3496 8538 3505
rect 8576 3470 8628 3476
rect 8482 3431 8538 3440
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8404 2650 8432 2858
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8668 2440 8720 2446
rect 8666 2408 8668 2417
rect 8720 2408 8722 2417
rect 8666 2343 8722 2352
rect 8668 1420 8720 1426
rect 8668 1362 8720 1368
rect 8680 480 8708 1362
rect 9232 480 9260 14719
rect 9416 12986 9444 20198
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10600 18896 10652 18902
rect 10600 18838 10652 18844
rect 10612 18358 10640 18838
rect 10600 18352 10652 18358
rect 10598 18320 10600 18329
rect 10652 18320 10654 18329
rect 10598 18255 10654 18264
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9678 18048 9734 18057
rect 9678 17983 9734 17992
rect 9692 17882 9720 17983
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9784 17814 9812 18090
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 10140 17672 10192 17678
rect 10138 17640 10140 17649
rect 10692 17672 10744 17678
rect 10192 17640 10194 17649
rect 10692 17614 10744 17620
rect 10138 17575 10194 17584
rect 10048 17332 10100 17338
rect 10152 17320 10180 17575
rect 10704 17338 10732 17614
rect 10100 17292 10180 17320
rect 10692 17332 10744 17338
rect 10048 17274 10100 17280
rect 10692 17274 10744 17280
rect 9588 17060 9640 17066
rect 9588 17002 9640 17008
rect 9600 16454 9628 17002
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16794 10732 17274
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10612 16250 10640 16390
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 10152 15586 10180 15914
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10796 15706 10824 22471
rect 11992 19310 12020 24103
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24780 23866 24808 25055
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 12714 23760 12770 23769
rect 12714 23695 12770 23704
rect 12728 23254 12756 23695
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 12716 23248 12768 23254
rect 12716 23190 12768 23196
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12452 22438 12480 23122
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 12898 20496 12954 20505
rect 12898 20431 12954 20440
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11164 16794 11192 18022
rect 11808 17814 11836 18566
rect 12176 18426 12204 19110
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12176 18222 12204 18362
rect 12544 18290 12572 18566
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12438 18184 12494 18193
rect 12438 18119 12494 18128
rect 12452 18086 12480 18119
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12544 17882 12572 18226
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11348 17134 11376 17614
rect 11808 17338 11836 17750
rect 12544 17354 12572 17818
rect 12622 17640 12678 17649
rect 12622 17575 12678 17584
rect 12452 17338 12572 17354
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 12440 17332 12572 17338
rect 12492 17326 12572 17332
rect 12440 17274 12492 17280
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11348 16726 11376 17070
rect 11336 16720 11388 16726
rect 11336 16662 11388 16668
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11532 16425 11560 16594
rect 11808 16590 11836 17274
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11518 16416 11574 16425
rect 11518 16351 11574 16360
rect 11532 16250 11560 16351
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11520 15904 11572 15910
rect 11624 15892 11652 16526
rect 11808 16250 11836 16526
rect 12452 16454 12480 17070
rect 12544 17066 12572 17326
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12636 16946 12664 17575
rect 12544 16918 12664 16946
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11572 15864 11652 15892
rect 11980 15904 12032 15910
rect 11520 15846 11572 15852
rect 11980 15846 12032 15852
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 9956 15564 10008 15570
rect 10152 15558 10272 15586
rect 9956 15506 10008 15512
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9586 15328 9642 15337
rect 9508 14929 9536 15302
rect 9586 15263 9642 15272
rect 9494 14920 9550 14929
rect 9494 14855 9496 14864
rect 9548 14855 9550 14864
rect 9496 14826 9548 14832
rect 9508 14795 9536 14826
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9508 13530 9536 13670
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9508 12782 9536 13126
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9600 12594 9628 15263
rect 9968 14822 9996 15506
rect 10244 15502 10272 15558
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10152 15065 10180 15438
rect 10244 15162 10272 15438
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10138 15056 10194 15065
rect 10138 14991 10194 15000
rect 11150 14920 11206 14929
rect 11150 14855 11206 14864
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9784 13326 9812 14350
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9416 12566 9628 12594
rect 9416 7970 9444 12566
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9496 12096 9548 12102
rect 9494 12064 9496 12073
rect 9548 12064 9550 12073
rect 9494 11999 9550 12008
rect 9600 11694 9628 12106
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9692 11354 9720 12718
rect 9864 12640 9916 12646
rect 9770 12608 9826 12617
rect 9864 12582 9916 12588
rect 9770 12543 9826 12552
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9784 10985 9812 12543
rect 9876 12073 9904 12582
rect 9862 12064 9918 12073
rect 9862 11999 9918 12008
rect 9968 11914 9996 14758
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 11164 14618 11192 14855
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11440 14482 11468 15506
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 10060 13938 10088 14418
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13530 10732 13670
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10336 12850 10364 13330
rect 11072 13297 11100 13670
rect 11058 13288 11114 13297
rect 11058 13223 11114 13232
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10980 12594 11008 12650
rect 11336 12640 11388 12646
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10796 12374 10824 12582
rect 10980 12566 11100 12594
rect 11336 12582 11388 12588
rect 11072 12442 11100 12566
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 9876 11886 9996 11914
rect 10336 11898 10364 12174
rect 11058 11928 11114 11937
rect 10324 11892 10376 11898
rect 9770 10976 9826 10985
rect 9770 10911 9826 10920
rect 9678 10432 9734 10441
rect 9678 10367 9734 10376
rect 9692 10266 9720 10367
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9784 9518 9812 10911
rect 9876 10130 9904 11886
rect 11058 11863 11114 11872
rect 10324 11834 10376 11840
rect 9954 11656 10010 11665
rect 9954 11591 9956 11600
rect 10008 11591 10010 11600
rect 9956 11562 10008 11568
rect 9968 10810 9996 11562
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 11072 11354 11100 11863
rect 11164 11558 11192 12242
rect 11242 12064 11298 12073
rect 11242 11999 11298 12008
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10152 10810 10180 11086
rect 10796 10810 10824 11154
rect 11164 11082 11192 11494
rect 11256 11354 11284 11999
rect 11348 11898 11376 12582
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10046 10296 10102 10305
rect 10046 10231 10048 10240
rect 10100 10231 10102 10240
rect 10048 10202 10100 10208
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9678 9344 9734 9353
rect 9678 9279 9734 9288
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9600 8090 9628 8842
rect 9692 8634 9720 9279
rect 9784 9178 9812 9454
rect 10060 9178 10088 10202
rect 10152 10198 10180 10746
rect 11060 10464 11112 10470
rect 10888 10412 11060 10418
rect 10888 10406 11112 10412
rect 10888 10390 11100 10406
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10138 9752 10194 9761
rect 10244 9738 10272 9998
rect 10194 9710 10272 9738
rect 10138 9687 10194 9696
rect 10152 9586 10180 9687
rect 10520 9654 10548 10066
rect 10508 9648 10560 9654
rect 10506 9616 10508 9625
rect 10560 9616 10562 9625
rect 10140 9580 10192 9586
rect 10506 9551 10562 9560
rect 10140 9522 10192 9528
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10704 9353 10732 9386
rect 10690 9344 10746 9353
rect 10289 9276 10585 9296
rect 10690 9279 10746 9288
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10598 9072 10654 9081
rect 10598 9007 10600 9016
rect 10652 9007 10654 9016
rect 10782 9072 10838 9081
rect 10782 9007 10838 9016
rect 10600 8978 10652 8984
rect 10232 8832 10284 8838
rect 9770 8800 9826 8809
rect 10232 8774 10284 8780
rect 9770 8735 9826 8744
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9416 7942 9628 7970
rect 9494 6896 9550 6905
rect 9494 6831 9496 6840
rect 9548 6831 9550 6840
rect 9496 6802 9548 6808
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 5574 9352 6598
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5166 9352 5510
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9324 4690 9352 5102
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9416 4214 9444 5034
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9508 3194 9536 5238
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9494 3088 9550 3097
rect 9494 3023 9550 3032
rect 9508 2854 9536 3023
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9600 1426 9628 7942
rect 9692 7478 9720 8366
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9692 2582 9720 6802
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9588 1420 9640 1426
rect 9588 1362 9640 1368
rect 9784 480 9812 8735
rect 10244 8537 10272 8774
rect 10612 8566 10640 8978
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10704 8634 10732 8910
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10600 8560 10652 8566
rect 10230 8528 10286 8537
rect 10600 8502 10652 8508
rect 10230 8463 10286 8472
rect 10138 8256 10194 8265
rect 10138 8191 10194 8200
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9968 7546 9996 8026
rect 10152 8022 10180 8191
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8090 10732 8570
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10140 8016 10192 8022
rect 10796 7970 10824 9007
rect 10140 7958 10192 7964
rect 10152 7546 10180 7958
rect 10612 7942 10824 7970
rect 9956 7540 10008 7546
rect 9876 7500 9956 7528
rect 9876 6866 9904 7500
rect 9956 7482 10008 7488
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10612 7426 10640 7942
rect 10690 7576 10746 7585
rect 10690 7511 10692 7520
rect 10744 7511 10746 7520
rect 10692 7482 10744 7488
rect 10152 7398 10640 7426
rect 10046 7032 10102 7041
rect 10046 6967 10102 6976
rect 10060 6934 10088 6967
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9862 6760 9918 6769
rect 9862 6695 9864 6704
rect 9916 6695 9918 6704
rect 9956 6724 10008 6730
rect 9864 6666 9916 6672
rect 9956 6666 10008 6672
rect 9876 6390 9904 6666
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9968 6254 9996 6666
rect 10060 6458 10088 6870
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9876 5098 9904 6054
rect 9968 5914 9996 6190
rect 10046 6080 10102 6089
rect 10046 6015 10102 6024
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9956 5704 10008 5710
rect 10060 5681 10088 6015
rect 9956 5646 10008 5652
rect 10046 5672 10102 5681
rect 9968 5522 9996 5646
rect 10046 5607 10102 5616
rect 9968 5494 10088 5522
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 10060 4486 10088 5494
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 4026 10088 4422
rect 9876 3998 10088 4026
rect 9876 2446 9904 3998
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9954 3768 10010 3777
rect 10060 3738 10088 3878
rect 9954 3703 10010 3712
rect 10048 3732 10100 3738
rect 9968 3369 9996 3703
rect 10048 3674 10100 3680
rect 9954 3360 10010 3369
rect 9954 3295 10010 3304
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 10152 1442 10180 7398
rect 10704 7342 10732 7482
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10782 7304 10838 7313
rect 10782 7239 10838 7248
rect 10796 7206 10824 7239
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 6089 10824 6598
rect 10782 6080 10838 6089
rect 10289 6012 10585 6032
rect 10782 6015 10838 6024
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10690 5808 10746 5817
rect 10690 5743 10692 5752
rect 10744 5743 10746 5752
rect 10692 5714 10744 5720
rect 10782 5400 10838 5409
rect 10782 5335 10784 5344
rect 10836 5335 10838 5344
rect 10784 5306 10836 5312
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10704 5001 10732 5034
rect 10690 4992 10746 5001
rect 10289 4924 10585 4944
rect 10690 4927 10746 4936
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10796 4758 10824 5306
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 10520 4146 10548 4490
rect 10690 4312 10746 4321
rect 10796 4282 10824 4694
rect 10690 4247 10746 4256
rect 10784 4276 10836 4282
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10506 4040 10562 4049
rect 10506 3975 10508 3984
rect 10560 3975 10562 3984
rect 10508 3946 10560 3952
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10244 3126 10272 3606
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10428 3126 10456 3538
rect 10704 3534 10732 4247
rect 10784 4218 10836 4224
rect 10782 3768 10838 3777
rect 10782 3703 10838 3712
rect 10796 3670 10824 3703
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2650 10732 3470
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10796 2854 10824 3402
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10704 2446 10732 2586
rect 10796 2446 10824 2790
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10152 1414 10364 1442
rect 10336 480 10364 1414
rect 10888 480 10916 10390
rect 11164 10266 11192 11018
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11256 8514 11284 8910
rect 11348 8634 11376 9318
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11256 8486 11376 8514
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11058 8120 11114 8129
rect 11058 8055 11114 8064
rect 11072 8022 11100 8055
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10966 7712 11022 7721
rect 10966 7647 11022 7656
rect 10980 6066 11008 7647
rect 11072 7177 11100 7822
rect 11164 7342 11192 8230
rect 11348 7886 11376 8486
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 11256 7410 11284 7754
rect 11348 7478 11376 7822
rect 11336 7472 11388 7478
rect 11336 7414 11388 7420
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11058 7168 11114 7177
rect 11058 7103 11114 7112
rect 11164 6934 11192 7278
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 11336 6112 11388 6118
rect 10980 6038 11100 6066
rect 11336 6054 11388 6060
rect 10966 5944 11022 5953
rect 10966 5879 10968 5888
rect 11020 5879 11022 5888
rect 10968 5850 11020 5856
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10980 5386 11008 5714
rect 11072 5658 11100 6038
rect 11072 5630 11284 5658
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 10980 5370 11100 5386
rect 10980 5364 11112 5370
rect 10980 5358 11060 5364
rect 11060 5306 11112 5312
rect 11164 5250 11192 5510
rect 10980 5222 11192 5250
rect 10980 4758 11008 5222
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10968 4480 11020 4486
rect 11256 4457 11284 5630
rect 11348 5273 11376 6054
rect 11334 5264 11390 5273
rect 11334 5199 11390 5208
rect 10968 4422 11020 4428
rect 11242 4448 11298 4457
rect 10980 3913 11008 4422
rect 11242 4383 11298 4392
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11060 4072 11112 4078
rect 11058 4040 11060 4049
rect 11112 4040 11114 4049
rect 11058 3975 11114 3984
rect 10966 3904 11022 3913
rect 10966 3839 11022 3848
rect 11152 3732 11204 3738
rect 11256 3720 11284 4082
rect 11204 3692 11284 3720
rect 11152 3674 11204 3680
rect 11164 3058 11192 3674
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10980 2378 11008 2926
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 11440 480 11468 13942
rect 11532 7256 11560 15846
rect 11992 15706 12020 15846
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11992 15162 12020 15642
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11978 15056 12034 15065
rect 11978 14991 12034 15000
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 13025 11928 13126
rect 11886 13016 11942 13025
rect 11886 12951 11888 12960
rect 11940 12951 11942 12960
rect 11888 12922 11940 12928
rect 11886 11248 11942 11257
rect 11612 11212 11664 11218
rect 11886 11183 11942 11192
rect 11612 11154 11664 11160
rect 11624 10985 11652 11154
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11610 10976 11666 10985
rect 11610 10911 11666 10920
rect 11624 10810 11652 10911
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11612 10532 11664 10538
rect 11612 10474 11664 10480
rect 11624 10130 11652 10474
rect 11716 10470 11744 11086
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11702 10296 11758 10305
rect 11702 10231 11758 10240
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11624 9722 11652 10066
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11716 9602 11744 10231
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11624 9574 11744 9602
rect 11624 8498 11652 9574
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11716 8974 11744 9454
rect 11808 9382 11836 10134
rect 11900 10062 11928 11183
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11808 8809 11836 9318
rect 11900 9110 11928 9998
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11794 8800 11850 8809
rect 11794 8735 11850 8744
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11716 7410 11744 7890
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11532 7228 11652 7256
rect 11518 7168 11574 7177
rect 11518 7103 11574 7112
rect 11532 6905 11560 7103
rect 11518 6896 11574 6905
rect 11518 6831 11520 6840
rect 11572 6831 11574 6840
rect 11520 6802 11572 6808
rect 11532 6458 11560 6802
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11624 4570 11652 7228
rect 11808 5914 11836 8434
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11716 5370 11744 5578
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11808 5166 11836 5850
rect 11900 5710 11928 6598
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4729 11928 4966
rect 11886 4720 11942 4729
rect 11886 4655 11942 4664
rect 11624 4542 11836 4570
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11716 3670 11744 4422
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11610 3088 11666 3097
rect 11610 3023 11666 3032
rect 11624 2650 11652 3023
rect 11716 2854 11744 3606
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11716 2553 11744 2790
rect 11702 2544 11758 2553
rect 11702 2479 11758 2488
rect 11808 610 11836 4542
rect 11796 604 11848 610
rect 11796 546 11848 552
rect 11992 480 12020 14991
rect 12084 14618 12112 15438
rect 12268 14822 12296 15438
rect 12438 15192 12494 15201
rect 12438 15127 12494 15136
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12084 14074 12112 14554
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12268 14006 12296 14758
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12452 13802 12480 15127
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 12452 13530 12480 13738
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12176 11898 12204 12242
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12254 10568 12310 10577
rect 12452 10538 12480 11154
rect 12254 10503 12310 10512
rect 12440 10532 12492 10538
rect 12268 10062 12296 10503
rect 12440 10474 12492 10480
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12176 8673 12204 9318
rect 12268 9178 12296 9998
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12360 9450 12388 9862
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12360 9178 12388 9386
rect 12452 9382 12480 10066
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12162 8664 12218 8673
rect 12162 8599 12218 8608
rect 12360 8498 12388 9114
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12452 8401 12480 8502
rect 12438 8392 12494 8401
rect 12438 8327 12494 8336
rect 12348 7200 12400 7206
rect 12400 7160 12480 7188
rect 12348 7142 12400 7148
rect 12452 6730 12480 7160
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12084 3602 12112 3878
rect 12176 3641 12204 6054
rect 12360 5522 12388 6598
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 12452 5817 12480 6326
rect 12438 5808 12494 5817
rect 12438 5743 12494 5752
rect 12360 5494 12480 5522
rect 12452 5166 12480 5494
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12162 3632 12218 3641
rect 12072 3596 12124 3602
rect 12162 3567 12218 3576
rect 12072 3538 12124 3544
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12360 3058 12388 3334
rect 12452 3194 12480 3878
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12070 2680 12126 2689
rect 12070 2615 12126 2624
rect 12438 2680 12494 2689
rect 12438 2615 12494 2624
rect 12084 2514 12112 2615
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 12452 2281 12480 2615
rect 12438 2272 12494 2281
rect 12438 2207 12494 2216
rect 12544 480 12572 16918
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12636 15366 12664 16390
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 14890 12664 15302
rect 12728 14958 12756 15642
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12636 14618 12664 14826
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12728 13938 12756 14894
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12820 14550 12848 14758
rect 12808 14544 12860 14550
rect 12808 14486 12860 14492
rect 12912 14362 12940 20431
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12820 14334 12940 14362
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12728 13530 12756 13874
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12820 13410 12848 14334
rect 12636 13382 12848 13410
rect 12900 13388 12952 13394
rect 12636 10266 12664 13382
rect 12900 13330 12952 13336
rect 12912 12986 12940 13330
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12728 12374 12756 12718
rect 13004 12442 13032 19246
rect 13372 13530 13400 22374
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 15382 19816 15438 19825
rect 15382 19751 15438 19760
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13728 15700 13780 15706
rect 13832 15688 13860 16934
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 13780 15660 13860 15688
rect 13728 15642 13780 15648
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13464 14074 13492 14418
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13266 13288 13322 13297
rect 13266 13223 13322 13232
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13188 12782 13216 13126
rect 13280 12986 13308 13223
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 12728 11694 12756 12310
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12820 11354 12848 12174
rect 13372 11898 13400 12174
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13266 11520 13322 11529
rect 13266 11455 13322 11464
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 13280 10266 13308 11455
rect 13372 11286 13400 11834
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13372 10470 13400 11086
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13096 9722 13124 10066
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12898 8528 12954 8537
rect 13004 8498 13032 9114
rect 12898 8463 12954 8472
rect 12992 8492 13044 8498
rect 12912 8430 12940 8463
rect 12992 8434 13044 8440
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12622 7984 12678 7993
rect 12622 7919 12678 7928
rect 12636 4826 12664 7919
rect 12806 7848 12862 7857
rect 12806 7783 12808 7792
rect 12860 7783 12862 7792
rect 12808 7754 12860 7760
rect 12912 7546 12940 8366
rect 13372 8265 13400 10406
rect 13358 8256 13414 8265
rect 13358 8191 13414 8200
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 13358 7440 13414 7449
rect 13358 7375 13414 7384
rect 13372 7342 13400 7375
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12636 4078 12664 4762
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12622 3632 12678 3641
rect 12622 3567 12678 3576
rect 12636 3398 12664 3567
rect 12624 3392 12676 3398
rect 12912 3369 12940 7142
rect 13372 7002 13400 7278
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 13004 5409 13032 6258
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12990 5400 13046 5409
rect 12990 5335 13046 5344
rect 13096 4826 13124 6122
rect 13358 5128 13414 5137
rect 13358 5063 13414 5072
rect 13372 4865 13400 5063
rect 13358 4856 13414 4865
rect 13084 4820 13136 4826
rect 13358 4791 13414 4800
rect 13084 4762 13136 4768
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13280 4593 13308 4626
rect 13360 4616 13412 4622
rect 13266 4584 13322 4593
rect 13360 4558 13412 4564
rect 13266 4519 13322 4528
rect 13280 4214 13308 4519
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13372 3942 13400 4558
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13372 3777 13400 3878
rect 13358 3768 13414 3777
rect 13358 3703 13414 3712
rect 13464 3618 13492 13806
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13740 13394 13768 13670
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13648 12306 13676 12650
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13832 12238 13860 13262
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13924 11778 13952 14214
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14004 13320 14056 13326
rect 14002 13288 14004 13297
rect 15292 13320 15344 13326
rect 14056 13288 14058 13297
rect 15292 13262 15344 13268
rect 14002 13223 14058 13232
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12986 15332 13262
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15304 12889 15332 12922
rect 14002 12880 14058 12889
rect 14002 12815 14058 12824
rect 15290 12880 15346 12889
rect 15290 12815 15346 12824
rect 13740 11750 13952 11778
rect 13740 11694 13768 11750
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 11150 13768 11630
rect 14016 11354 14044 12815
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14384 11558 14412 12242
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15396 11898 15424 19751
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24674 19544 24730 19553
rect 24674 19479 24730 19488
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 24030 15600 24086 15609
rect 24030 15535 24086 15544
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 23662 14376 23718 14385
rect 23662 14311 23718 14320
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 23386 13424 23442 13433
rect 15844 13388 15896 13394
rect 23386 13359 23388 13368
rect 15844 13330 15896 13336
rect 23440 13359 23442 13368
rect 23388 13330 23440 13336
rect 15856 12714 15884 13330
rect 16670 13288 16726 13297
rect 16670 13223 16672 13232
rect 16724 13223 16726 13232
rect 16672 13194 16724 13200
rect 23400 12986 23428 13330
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23676 12782 23704 14311
rect 24044 13870 24072 15535
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 15856 12238 15884 12650
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 22282 12336 22338 12345
rect 22282 12271 22284 12280
rect 22336 12271 22338 12280
rect 22284 12242 22336 12248
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15488 11626 15516 12174
rect 15566 11792 15622 11801
rect 15566 11727 15622 11736
rect 15752 11756 15804 11762
rect 15580 11694 15608 11727
rect 15752 11698 15804 11704
rect 15568 11688 15620 11694
rect 15764 11665 15792 11698
rect 15568 11630 15620 11636
rect 15750 11656 15806 11665
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 13924 10713 13952 11018
rect 13910 10704 13966 10713
rect 13740 10662 13910 10690
rect 13740 10606 13768 10662
rect 13910 10639 13966 10648
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13818 10160 13874 10169
rect 13740 9330 13768 10134
rect 14384 10130 14412 11494
rect 14476 11354 14504 11562
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14476 10305 14504 10406
rect 14462 10296 14518 10305
rect 14462 10231 14518 10240
rect 13818 10095 13874 10104
rect 14372 10124 14424 10130
rect 13832 10062 13860 10095
rect 14372 10066 14424 10072
rect 13820 10056 13872 10062
rect 13872 10016 13952 10044
rect 13820 9998 13872 10004
rect 13818 9752 13874 9761
rect 13818 9687 13874 9696
rect 13832 9654 13860 9687
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13740 9302 13860 9330
rect 13832 9110 13860 9302
rect 13924 9178 13952 10016
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 14016 9518 14044 9862
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14384 9382 14412 10066
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13820 9104 13872 9110
rect 13818 9072 13820 9081
rect 13872 9072 13874 9081
rect 13544 9036 13596 9042
rect 13818 9007 13874 9016
rect 13544 8978 13596 8984
rect 13556 8566 13584 8978
rect 13544 8560 13596 8566
rect 13542 8528 13544 8537
rect 13596 8528 13598 8537
rect 13542 8463 13598 8472
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13648 7410 13676 7686
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13740 7041 13768 7142
rect 13726 7032 13782 7041
rect 13726 6967 13782 6976
rect 13832 6458 13860 7346
rect 13924 7274 13952 8298
rect 14278 8256 14334 8265
rect 14278 8191 14334 8200
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 14016 6934 14044 7686
rect 14200 7002 14228 7822
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14004 6928 14056 6934
rect 14004 6870 14056 6876
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13924 5710 13952 6802
rect 14016 6633 14044 6870
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14002 6624 14058 6633
rect 14002 6559 14058 6568
rect 14200 6361 14228 6734
rect 14186 6352 14242 6361
rect 14186 6287 14242 6296
rect 13912 5704 13964 5710
rect 13910 5672 13912 5681
rect 13964 5672 13966 5681
rect 13910 5607 13966 5616
rect 14186 5672 14242 5681
rect 14186 5607 14242 5616
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13648 5137 13676 5510
rect 13634 5128 13690 5137
rect 13634 5063 13636 5072
rect 13688 5063 13690 5072
rect 13728 5092 13780 5098
rect 13636 5034 13688 5040
rect 13728 5034 13780 5040
rect 13634 4992 13690 5001
rect 13634 4927 13690 4936
rect 13740 4978 13768 5034
rect 13740 4950 13860 4978
rect 13648 4622 13676 4927
rect 13740 4758 13768 4950
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13648 3738 13676 4558
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13464 3590 13676 3618
rect 12624 3334 12676 3340
rect 12898 3360 12954 3369
rect 12636 2922 12664 3334
rect 12898 3295 12954 3304
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 12898 2816 12954 2825
rect 12898 2751 12954 2760
rect 12714 2680 12770 2689
rect 12912 2650 12940 2751
rect 12714 2615 12770 2624
rect 12900 2644 12952 2650
rect 12728 2514 12756 2615
rect 12900 2586 12952 2592
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 13542 2408 13598 2417
rect 13542 2343 13544 2352
rect 13596 2343 13598 2352
rect 13544 2314 13596 2320
rect 13542 1728 13598 1737
rect 13542 1663 13598 1672
rect 13556 1465 13584 1663
rect 13542 1456 13598 1465
rect 13542 1391 13598 1400
rect 13084 604 13136 610
rect 13084 546 13136 552
rect 13096 480 13124 546
rect 13648 480 13676 3590
rect 13740 3482 13768 4218
rect 13832 3942 13860 4950
rect 14094 4720 14150 4729
rect 14094 4655 14096 4664
rect 14148 4655 14150 4664
rect 14096 4626 14148 4632
rect 14108 4078 14136 4626
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13832 3602 13860 3878
rect 14200 3670 14228 5607
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13740 3454 13860 3482
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 2281 13768 3334
rect 13832 3126 13860 3454
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13818 2408 13874 2417
rect 13818 2343 13820 2352
rect 13872 2343 13874 2352
rect 13820 2314 13872 2320
rect 13726 2272 13782 2281
rect 13726 2207 13782 2216
rect 13740 1737 13768 2207
rect 13726 1728 13782 1737
rect 13726 1663 13782 1672
rect 14292 480 14320 8191
rect 14384 8129 14412 9318
rect 14462 8936 14518 8945
rect 14462 8871 14464 8880
rect 14516 8871 14518 8880
rect 14464 8842 14516 8848
rect 14476 8430 14504 8842
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14370 8120 14426 8129
rect 14370 8055 14426 8064
rect 14476 6866 14504 8230
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6322 14412 6598
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14384 5914 14412 6258
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14476 5846 14504 6802
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14462 5536 14518 5545
rect 14462 5471 14518 5480
rect 14476 5001 14504 5471
rect 14462 4992 14518 5001
rect 14462 4927 14518 4936
rect 14568 4570 14596 11562
rect 15580 11354 15608 11630
rect 15750 11591 15806 11600
rect 15660 11552 15712 11558
rect 15658 11520 15660 11529
rect 15712 11520 15714 11529
rect 15658 11455 15714 11464
rect 15856 11354 15884 12174
rect 22296 11898 22324 12242
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 15292 10056 15344 10062
rect 15290 10024 15292 10033
rect 15344 10024 15346 10033
rect 15290 9959 15346 9968
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14660 9722 14688 9862
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 8566 14780 8774
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14752 7750 14780 8502
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14738 7032 14794 7041
rect 14738 6967 14794 6976
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14660 5370 14688 6190
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14752 4826 14780 6967
rect 14844 5914 14872 9318
rect 15396 9042 15424 9590
rect 15474 9344 15530 9353
rect 15474 9279 15530 9288
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15396 8634 15424 8978
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15108 8492 15160 8498
rect 15396 8480 15424 8570
rect 15108 8434 15160 8440
rect 15304 8452 15424 8480
rect 15120 7954 15148 8434
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15304 7886 15332 8452
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 7426 15332 7822
rect 15028 7398 15332 7426
rect 15028 7342 15056 7398
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15382 6760 15438 6769
rect 15382 6695 15384 6704
rect 15436 6695 15438 6704
rect 15384 6666 15436 6672
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15382 6080 15438 6089
rect 15382 6015 15438 6024
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 5370 15332 5850
rect 15396 5545 15424 6015
rect 15382 5536 15438 5545
rect 15382 5471 15438 5480
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14568 4542 14780 4570
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14660 4010 14688 4422
rect 14648 4004 14700 4010
rect 14648 3946 14700 3952
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14384 2650 14412 3130
rect 14660 2922 14688 3946
rect 14648 2916 14700 2922
rect 14648 2858 14700 2864
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14660 2446 14688 2858
rect 14752 2802 14780 4542
rect 14844 3738 14872 4966
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14832 3596 14884 3602
rect 14936 3584 14964 3946
rect 15304 3777 15332 4422
rect 15290 3768 15346 3777
rect 15290 3703 15346 3712
rect 14884 3556 14964 3584
rect 14832 3538 14884 3544
rect 14844 2990 14872 3538
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 14752 2774 14872 2802
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 14568 1873 14596 2246
rect 14554 1864 14610 1873
rect 14554 1799 14610 1808
rect 14844 480 14872 2774
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15304 2310 15332 2518
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15304 1601 15332 2246
rect 15290 1592 15346 1601
rect 15290 1527 15346 1536
rect 15488 626 15516 9279
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15672 8362 15700 8978
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16302 8664 16358 8673
rect 16302 8599 16358 8608
rect 16316 8498 16344 8599
rect 16776 8537 16804 8774
rect 22282 8664 22338 8673
rect 17224 8628 17276 8634
rect 22282 8599 22338 8608
rect 17224 8570 17276 8576
rect 16762 8528 16818 8537
rect 16304 8492 16356 8498
rect 16762 8463 16818 8472
rect 16304 8434 16356 8440
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15580 7721 15608 7890
rect 15566 7712 15622 7721
rect 15566 7647 15622 7656
rect 15580 7546 15608 7647
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15844 7268 15896 7274
rect 15844 7210 15896 7216
rect 15750 7032 15806 7041
rect 15750 6967 15806 6976
rect 15764 5914 15792 6967
rect 15856 6118 15884 7210
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15856 5710 15884 6054
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15948 5642 15976 8366
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16684 7750 16712 8230
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16304 7200 16356 7206
rect 16302 7168 16304 7177
rect 16356 7168 16358 7177
rect 16302 7103 16358 7112
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 6458 16068 6734
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16316 6390 16344 6938
rect 16684 6458 16712 7686
rect 17236 7546 17264 8570
rect 20904 8424 20956 8430
rect 20902 8392 20904 8401
rect 20956 8392 20958 8401
rect 20902 8327 20958 8336
rect 22008 8356 22060 8362
rect 22008 8298 22060 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19154 7712 19210 7721
rect 19154 7647 19210 7656
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16868 6662 16896 7142
rect 17236 7002 17264 7482
rect 18052 7336 18104 7342
rect 18050 7304 18052 7313
rect 18104 7304 18106 7313
rect 18050 7239 18106 7248
rect 18328 7268 18380 7274
rect 18328 7210 18380 7216
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16304 6384 16356 6390
rect 16304 6326 16356 6332
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16302 5944 16358 5953
rect 16302 5879 16304 5888
rect 16356 5879 16358 5888
rect 16304 5850 16356 5856
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 15658 5264 15714 5273
rect 15658 5199 15660 5208
rect 15712 5199 15714 5208
rect 15660 5170 15712 5176
rect 16316 5166 16344 5850
rect 16488 5704 16540 5710
rect 16868 5681 16896 6190
rect 16488 5646 16540 5652
rect 16854 5672 16910 5681
rect 16500 5370 16528 5646
rect 16854 5607 16856 5616
rect 16908 5607 16910 5616
rect 16856 5578 16908 5584
rect 17236 5574 17264 6598
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 17776 6248 17828 6254
rect 17774 6216 17776 6225
rect 17828 6216 17830 6225
rect 17774 6151 17830 6160
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17500 5840 17552 5846
rect 17500 5782 17552 5788
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 16304 5160 16356 5166
rect 16408 5137 16436 5170
rect 16304 5102 16356 5108
rect 16394 5128 16450 5137
rect 16394 5063 16450 5072
rect 15750 4856 15806 4865
rect 16408 4826 16436 5063
rect 15750 4791 15752 4800
rect 15804 4791 15806 4800
rect 16396 4820 16448 4826
rect 15752 4762 15804 4768
rect 16396 4762 16448 4768
rect 15658 4720 15714 4729
rect 15658 4655 15660 4664
rect 15712 4655 15714 4664
rect 15660 4626 15712 4632
rect 15672 4282 15700 4626
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 15764 3738 15792 4762
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15856 3942 15884 4558
rect 17144 3942 17172 4626
rect 17236 4486 17264 5510
rect 17512 5370 17540 5782
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 18064 5098 18092 6054
rect 18052 5092 18104 5098
rect 18052 5034 18104 5040
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15856 3670 15884 3878
rect 16868 3670 16896 3878
rect 16960 3738 16988 3878
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 16856 3664 16908 3670
rect 16856 3606 16908 3612
rect 16868 3194 16896 3606
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 15658 3088 15714 3097
rect 15658 3023 15714 3032
rect 15672 2650 15700 3023
rect 15934 2816 15990 2825
rect 15934 2751 15990 2760
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15396 598 15516 626
rect 15396 480 15424 598
rect 15948 480 15976 2751
rect 16960 2650 16988 3538
rect 17144 3398 17172 3878
rect 17696 3670 17724 4422
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17776 3936 17828 3942
rect 17972 3913 18000 3946
rect 17776 3878 17828 3884
rect 17958 3904 18014 3913
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 17788 3505 17816 3878
rect 17958 3839 18014 3848
rect 17972 3670 18000 3839
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 18050 3632 18106 3641
rect 18050 3567 18106 3576
rect 17774 3496 17830 3505
rect 17774 3431 17830 3440
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17038 3224 17094 3233
rect 17144 3194 17172 3334
rect 17038 3159 17094 3168
rect 17132 3188 17184 3194
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 16026 2544 16082 2553
rect 16026 2479 16082 2488
rect 16040 2446 16068 2479
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16580 2304 16632 2310
rect 16580 2246 16632 2252
rect 16592 1442 16620 2246
rect 16500 1414 16620 1442
rect 16500 480 16528 1414
rect 17052 480 17080 3159
rect 17132 3130 17184 3136
rect 17774 2952 17830 2961
rect 17774 2887 17776 2896
rect 17828 2887 17830 2896
rect 17776 2858 17828 2864
rect 18064 2854 18092 3567
rect 18052 2848 18104 2854
rect 17590 2816 17646 2825
rect 18052 2790 18104 2796
rect 17590 2751 17646 2760
rect 17604 480 17632 2751
rect 17682 2680 17738 2689
rect 18064 2650 18092 2790
rect 17682 2615 17684 2624
rect 17736 2615 17738 2624
rect 18052 2644 18104 2650
rect 17684 2586 17736 2592
rect 18052 2586 18104 2592
rect 18156 480 18184 6326
rect 18340 4049 18368 7210
rect 19168 7002 19196 7647
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 19076 6458 19104 6802
rect 20916 6769 20944 6802
rect 21180 6792 21232 6798
rect 20902 6760 20958 6769
rect 21180 6734 21232 6740
rect 20902 6695 20958 6704
rect 20916 6458 20944 6695
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18708 5846 18736 6258
rect 19076 5914 19104 6394
rect 20534 6352 20590 6361
rect 20534 6287 20590 6296
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18524 4282 18552 4966
rect 18708 4826 18736 5782
rect 19076 5234 19104 5850
rect 19522 5808 19578 5817
rect 19522 5743 19578 5752
rect 19064 5228 19116 5234
rect 19064 5170 19116 5176
rect 19338 4992 19394 5001
rect 19338 4927 19394 4936
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 18708 4282 18736 4762
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18696 4276 18748 4282
rect 18696 4218 18748 4224
rect 18326 4040 18382 4049
rect 18326 3975 18382 3984
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18524 3641 18552 3946
rect 18694 3768 18750 3777
rect 19260 3738 19288 4422
rect 18694 3703 18750 3712
rect 19064 3732 19116 3738
rect 18708 3670 18736 3703
rect 19064 3674 19116 3680
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 18696 3664 18748 3670
rect 18510 3632 18566 3641
rect 18696 3606 18748 3612
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 18510 3567 18566 3576
rect 18788 3528 18840 3534
rect 18694 3496 18750 3505
rect 18788 3470 18840 3476
rect 18694 3431 18750 3440
rect 18510 3088 18566 3097
rect 18510 3023 18566 3032
rect 18604 3052 18656 3058
rect 18524 2990 18552 3023
rect 18604 2994 18656 3000
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18616 2854 18644 2994
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 18340 1873 18368 2450
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18326 1864 18382 1873
rect 18326 1799 18382 1808
rect 18524 1737 18552 2382
rect 18510 1728 18566 1737
rect 18510 1663 18566 1672
rect 18708 480 18736 3431
rect 18800 3194 18828 3470
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18984 2650 19012 3606
rect 19076 3194 19104 3674
rect 19246 3360 19302 3369
rect 19246 3295 19302 3304
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 19260 480 19288 3295
rect 19352 3058 19380 4927
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19444 3942 19472 4626
rect 19536 4078 19564 5743
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19444 3126 19472 3878
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20074 3768 20130 3777
rect 20074 3703 20076 3712
rect 20128 3703 20130 3712
rect 20076 3674 20128 3680
rect 19982 3224 20038 3233
rect 19982 3159 20038 3168
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19340 2916 19392 2922
rect 19340 2858 19392 2864
rect 19352 2689 19380 2858
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19338 2680 19394 2689
rect 19622 2672 19918 2692
rect 19338 2615 19394 2624
rect 19798 2544 19854 2553
rect 19616 2508 19668 2514
rect 19798 2479 19854 2488
rect 19616 2450 19668 2456
rect 19628 1465 19656 2450
rect 19812 2446 19840 2479
rect 19800 2440 19852 2446
rect 19800 2382 19852 2388
rect 19614 1456 19670 1465
rect 19614 1391 19670 1400
rect 19996 762 20024 3159
rect 19812 734 20024 762
rect 19812 480 19840 734
rect 20364 480 20392 4422
rect 20548 2553 20576 6287
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20810 5536 20866 5545
rect 20810 5471 20866 5480
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20640 4026 20668 4558
rect 20640 4010 20760 4026
rect 20640 4004 20772 4010
rect 20640 3998 20720 4004
rect 20720 3946 20772 3952
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 20732 3194 20760 3402
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 20824 2990 20852 5471
rect 20916 5370 20944 5714
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20916 4282 20944 4626
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20904 4072 20956 4078
rect 20902 4040 20904 4049
rect 21100 4049 21128 5510
rect 21192 4690 21220 6734
rect 21548 5024 21600 5030
rect 21548 4966 21600 4972
rect 21640 5024 21692 5030
rect 21640 4966 21692 4972
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 20956 4040 20958 4049
rect 20902 3975 20958 3984
rect 21086 4040 21142 4049
rect 21086 3975 21142 3984
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20534 2544 20590 2553
rect 20534 2479 20590 2488
rect 20916 480 20944 3674
rect 21100 3369 21128 3878
rect 21180 3528 21232 3534
rect 21180 3470 21232 3476
rect 21086 3360 21142 3369
rect 21086 3295 21142 3304
rect 21192 3097 21220 3470
rect 21178 3088 21234 3097
rect 21178 3023 21234 3032
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21192 2417 21220 2450
rect 21178 2408 21234 2417
rect 21178 2343 21234 2352
rect 21560 480 21588 4966
rect 21652 2582 21680 4966
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 21836 4282 21864 4626
rect 22020 4298 22048 8298
rect 21824 4276 21876 4282
rect 22020 4270 22140 4298
rect 21824 4218 21876 4224
rect 22112 3670 22140 4270
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22204 3738 22232 3878
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22100 3664 22152 3670
rect 22100 3606 22152 3612
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22204 3194 22232 3538
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22296 2990 22324 8599
rect 22480 5681 22508 12038
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 22834 10704 22890 10713
rect 22834 10639 22890 10648
rect 22466 5672 22522 5681
rect 22466 5607 22522 5616
rect 22558 4040 22614 4049
rect 22558 3975 22614 3984
rect 22466 3496 22522 3505
rect 22466 3431 22522 3440
rect 22376 3392 22428 3398
rect 22376 3334 22428 3340
rect 22388 3233 22416 3334
rect 22374 3224 22430 3233
rect 22480 3194 22508 3431
rect 22374 3159 22430 3168
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 22284 2984 22336 2990
rect 22284 2926 22336 2932
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 21640 2576 21692 2582
rect 21640 2518 21692 2524
rect 22112 480 22140 2858
rect 22466 2544 22522 2553
rect 22572 2530 22600 3975
rect 22650 2952 22706 2961
rect 22650 2887 22706 2896
rect 22664 2650 22692 2887
rect 22848 2825 22876 10639
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24214 8392 24270 8401
rect 24214 8327 24270 8336
rect 24124 6928 24176 6934
rect 24124 6870 24176 6876
rect 24030 5672 24086 5681
rect 24030 5607 24086 5616
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 22834 2816 22890 2825
rect 22834 2751 22890 2760
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 22572 2502 22692 2530
rect 22466 2479 22468 2488
rect 22520 2479 22522 2488
rect 22468 2450 22520 2456
rect 22664 480 22692 2502
rect 23216 480 23244 4422
rect 23952 4214 23980 4558
rect 23940 4208 23992 4214
rect 23940 4150 23992 4156
rect 23952 3777 23980 4150
rect 23938 3768 23994 3777
rect 23938 3703 23994 3712
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 23308 3194 23336 3538
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23662 3088 23718 3097
rect 23662 3023 23718 3032
rect 23676 2990 23704 3023
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 23768 480 23796 3334
rect 24044 1986 24072 5607
rect 24136 2514 24164 6870
rect 24228 4758 24256 8327
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 6934 24716 19479
rect 24860 14000 24912 14006
rect 24766 13968 24822 13977
rect 24860 13942 24912 13948
rect 24766 13903 24822 13912
rect 24780 13297 24808 13903
rect 24766 13288 24822 13297
rect 24766 13223 24822 13232
rect 24676 6928 24728 6934
rect 24676 6870 24728 6876
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24216 4752 24268 4758
rect 24216 4694 24268 4700
rect 24228 4282 24256 4694
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24216 4276 24268 4282
rect 24216 4218 24268 4224
rect 24674 4176 24730 4185
rect 24674 4111 24730 4120
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 2990 24716 4111
rect 24872 3670 24900 13942
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24860 3664 24912 3670
rect 24860 3606 24912 3612
rect 24964 3602 24992 13126
rect 25044 12912 25096 12918
rect 25044 12854 25096 12860
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 25056 3482 25084 12854
rect 25318 4584 25374 4593
rect 25318 4519 25320 4528
rect 25372 4519 25374 4528
rect 25320 4490 25372 4496
rect 25964 3664 26016 3670
rect 25964 3606 26016 3612
rect 25412 3596 25464 3602
rect 25412 3538 25464 3544
rect 24872 3454 25084 3482
rect 24766 3088 24822 3097
rect 24766 3023 24822 3032
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 24780 2650 24808 3023
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24044 1958 24348 1986
rect 24320 480 24348 1958
rect 24872 480 24900 3454
rect 25424 480 25452 3538
rect 25976 480 26004 3606
rect 26516 3120 26568 3126
rect 26516 3062 26568 3068
rect 27618 3088 27674 3097
rect 26528 480 26556 3062
rect 27618 3023 27674 3032
rect 27066 2952 27122 2961
rect 27066 2887 27122 2896
rect 27080 480 27108 2887
rect 27632 480 27660 3023
rect 2962 368 3018 377
rect 2962 303 3018 312
rect 3054 0 3110 480
rect 3606 0 3662 480
rect 4158 0 4214 480
rect 4710 0 4766 480
rect 5262 0 5318 480
rect 5814 0 5870 480
rect 6366 0 6422 480
rect 6918 0 6974 480
rect 7562 0 7618 480
rect 8114 0 8170 480
rect 8666 0 8722 480
rect 9218 0 9274 480
rect 9770 0 9826 480
rect 10322 0 10378 480
rect 10874 0 10930 480
rect 11426 0 11482 480
rect 11978 0 12034 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14278 0 14334 480
rect 14830 0 14886 480
rect 15382 0 15438 480
rect 15934 0 15990 480
rect 16486 0 16542 480
rect 17038 0 17094 480
rect 17590 0 17646 480
rect 18142 0 18198 480
rect 18694 0 18750 480
rect 19246 0 19302 480
rect 19798 0 19854 480
rect 20350 0 20406 480
rect 20902 0 20958 480
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22650 0 22706 480
rect 23202 0 23258 480
rect 23754 0 23810 480
rect 24306 0 24362 480
rect 24858 0 24914 480
rect 25410 0 25466 480
rect 25962 0 26018 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 2778 27648 2834 27704
rect 2686 26016 2742 26072
rect 1582 25472 1638 25528
rect 1490 24928 1546 24984
rect 2042 24132 2098 24168
rect 2042 24112 2044 24132
rect 2044 24112 2096 24132
rect 2096 24112 2098 24132
rect 1490 23160 1546 23216
rect 3330 27104 3386 27160
rect 3238 26560 3294 26616
rect 2962 24384 3018 24440
rect 2686 23840 2742 23896
rect 1674 22516 1676 22536
rect 1676 22516 1728 22536
rect 1728 22516 1730 22536
rect 1674 22480 1730 22516
rect 2594 22380 2596 22400
rect 2596 22380 2648 22400
rect 2648 22380 2650 22400
rect 2594 22344 2650 22380
rect 3698 23724 3754 23760
rect 3698 23704 3700 23724
rect 3700 23704 3752 23724
rect 3752 23704 3754 23724
rect 3422 22616 3478 22672
rect 3422 21936 3478 21992
rect 2686 21564 2688 21584
rect 2688 21564 2740 21584
rect 2740 21564 2742 21584
rect 2686 21528 2742 21564
rect 1582 20984 1638 21040
rect 1674 20884 1676 20904
rect 1676 20884 1728 20904
rect 1728 20884 1730 20904
rect 1674 20848 1730 20884
rect 2410 21412 2466 21448
rect 2410 21392 2412 21412
rect 2412 21392 2464 21412
rect 2464 21392 2466 21412
rect 1766 19760 1822 19816
rect 2594 20596 2650 20632
rect 2594 20576 2596 20596
rect 2596 20576 2648 20596
rect 2648 20576 2650 20596
rect 2686 20440 2742 20496
rect 4434 22344 4490 22400
rect 4066 22072 4122 22128
rect 4158 20440 4214 20496
rect 4250 20168 4306 20224
rect 3698 20032 3754 20088
rect 3238 19896 3294 19952
rect 1674 19116 1676 19136
rect 1676 19116 1728 19136
rect 1728 19116 1730 19136
rect 1674 19080 1730 19116
rect 2686 18944 2742 19000
rect 1582 16632 1638 16688
rect 1398 15816 1454 15872
rect 1858 13096 1914 13152
rect 2870 18128 2926 18184
rect 1950 11736 2006 11792
rect 1766 10104 1822 10160
rect 2318 15000 2374 15056
rect 3054 17584 3110 17640
rect 4066 18944 4122 19000
rect 3238 16496 3294 16552
rect 2778 15000 2834 15056
rect 2502 14592 2558 14648
rect 2870 14592 2926 14648
rect 2410 14456 2466 14512
rect 2318 13932 2374 13968
rect 2318 13912 2320 13932
rect 2320 13912 2372 13932
rect 2372 13912 2374 13932
rect 2962 12708 3018 12744
rect 2962 12688 2964 12708
rect 2964 12688 3016 12708
rect 3016 12688 3018 12708
rect 3238 11464 3294 11520
rect 2318 9560 2374 9616
rect 2226 9036 2282 9072
rect 2226 9016 2228 9036
rect 2228 9016 2280 9036
rect 2280 9016 2282 9036
rect 1398 8200 1454 8256
rect 846 1944 902 2000
rect 3054 9832 3110 9888
rect 2870 9696 2926 9752
rect 2134 7928 2190 7984
rect 1950 6296 2006 6352
rect 1858 5888 1914 5944
rect 2502 7148 2504 7168
rect 2504 7148 2556 7168
rect 2556 7148 2558 7168
rect 2502 7112 2558 7148
rect 2870 6568 2926 6624
rect 2134 3576 2190 3632
rect 1674 3032 1730 3088
rect 1950 2896 2006 2952
rect 2594 4800 2650 4856
rect 2686 3848 2742 3904
rect 2778 2080 2834 2136
rect 2502 1536 2558 1592
rect 3054 6840 3110 6896
rect 3238 5888 3294 5944
rect 3054 4120 3110 4176
rect 3974 17040 4030 17096
rect 3790 16668 3792 16688
rect 3792 16668 3844 16688
rect 3844 16668 3846 16688
rect 3790 16632 3846 16668
rect 3698 16360 3754 16416
rect 3422 13640 3478 13696
rect 3606 12960 3662 13016
rect 3514 12552 3570 12608
rect 3422 12416 3478 12472
rect 3514 10512 3570 10568
rect 3514 9560 3570 9616
rect 4250 18692 4306 18728
rect 4250 18672 4252 18692
rect 4252 18672 4304 18692
rect 4304 18672 4306 18692
rect 3974 16088 4030 16144
rect 3790 15952 3846 16008
rect 4618 19352 4674 19408
rect 4434 18128 4490 18184
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 24766 25064 24822 25120
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 11978 24112 12034 24168
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 10782 22480 10838 22536
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 8574 21936 8630 21992
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 7286 21392 7342 21448
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 7378 20032 7434 20088
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 6826 19116 6828 19136
rect 6828 19116 6880 19136
rect 6880 19116 6882 19136
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5262 16904 5318 16960
rect 5354 16632 5410 16688
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 6826 19080 6882 19116
rect 8114 20884 8116 20904
rect 8116 20884 8168 20904
rect 8168 20884 8170 20904
rect 8114 20848 8170 20884
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 6090 16360 6146 16416
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 4250 13912 4306 13968
rect 4618 13912 4674 13968
rect 3790 12144 3846 12200
rect 3790 12008 3846 12064
rect 3698 11328 3754 11384
rect 3698 10376 3754 10432
rect 3606 9288 3662 9344
rect 3514 6840 3570 6896
rect 3514 5616 3570 5672
rect 3514 4800 3570 4856
rect 3882 10376 3938 10432
rect 4158 10512 4214 10568
rect 3974 9152 4030 9208
rect 3698 8336 3754 8392
rect 3238 3168 3294 3224
rect 3606 4392 3662 4448
rect 3054 2760 3110 2816
rect 3606 2488 3662 2544
rect 4710 13676 4712 13696
rect 4712 13676 4764 13696
rect 4764 13676 4766 13696
rect 4710 13640 4766 13676
rect 4618 13132 4620 13152
rect 4620 13132 4672 13152
rect 4672 13132 4674 13152
rect 4618 13096 4674 13132
rect 4342 11736 4398 11792
rect 4434 10512 4490 10568
rect 4158 8880 4214 8936
rect 4250 8336 4306 8392
rect 3974 8064 4030 8120
rect 3882 7520 3938 7576
rect 4342 7420 4344 7440
rect 4344 7420 4396 7440
rect 4396 7420 4398 7440
rect 3882 6840 3938 6896
rect 4342 7384 4398 7420
rect 5354 13812 5356 13832
rect 5356 13812 5408 13832
rect 5408 13812 5410 13832
rect 5354 13776 5410 13812
rect 6826 16496 6882 16552
rect 6642 16360 6698 16416
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5998 14864 6054 14920
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5722 13932 5778 13968
rect 5722 13912 5724 13932
rect 5724 13912 5776 13932
rect 5776 13912 5778 13932
rect 5998 13368 6054 13424
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5538 12144 5594 12200
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 4066 6976 4122 7032
rect 3882 4664 3938 4720
rect 3790 4528 3846 4584
rect 3698 1400 3754 1456
rect 3882 3460 3938 3496
rect 3882 3440 3884 3460
rect 3884 3440 3936 3460
rect 3936 3440 3938 3460
rect 4250 6296 4306 6352
rect 4526 7112 4582 7168
rect 4710 7112 4766 7168
rect 5814 11348 5870 11384
rect 5814 11328 5816 11348
rect 5816 11328 5868 11348
rect 5868 11328 5870 11348
rect 5170 10004 5172 10024
rect 5172 10004 5224 10024
rect 5224 10004 5226 10024
rect 5170 9968 5226 10004
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5354 10240 5410 10296
rect 7010 16088 7066 16144
rect 6550 15272 6606 15328
rect 6274 15156 6330 15192
rect 6274 15136 6276 15156
rect 6276 15136 6328 15156
rect 6328 15136 6330 15156
rect 6826 15000 6882 15056
rect 6458 14864 6514 14920
rect 6274 10240 6330 10296
rect 5630 10124 5686 10160
rect 5630 10104 5632 10124
rect 5632 10104 5684 10124
rect 5684 10104 5686 10124
rect 5998 10104 6054 10160
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5446 9696 5502 9752
rect 5262 9016 5318 9072
rect 6642 14764 6644 14784
rect 6644 14764 6696 14784
rect 6696 14764 6698 14784
rect 6642 14728 6698 14764
rect 6550 14456 6606 14512
rect 7194 15816 7250 15872
rect 7378 15136 7434 15192
rect 7562 14728 7618 14784
rect 7838 14592 7894 14648
rect 7378 13776 7434 13832
rect 7286 13640 7342 13696
rect 6642 12008 6698 12064
rect 6550 10376 6606 10432
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5722 8356 5778 8392
rect 5722 8336 5724 8356
rect 5724 8336 5776 8356
rect 5776 8336 5778 8356
rect 4802 6840 4858 6896
rect 4618 6432 4674 6488
rect 4342 5888 4398 5944
rect 4158 4392 4214 4448
rect 4526 3576 4582 3632
rect 3974 1672 4030 1728
rect 3790 856 3846 912
rect 4618 3440 4674 3496
rect 4802 5752 4858 5808
rect 5078 3884 5080 3904
rect 5080 3884 5132 3904
rect 5132 3884 5134 3904
rect 4894 2624 4950 2680
rect 5078 3848 5134 3884
rect 4986 2352 5042 2408
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5722 6976 5778 7032
rect 6090 7692 6092 7712
rect 6092 7692 6144 7712
rect 6144 7692 6146 7712
rect 6090 7656 6146 7692
rect 6182 7520 6238 7576
rect 5998 6704 6054 6760
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 6182 6840 6238 6896
rect 7102 11228 7104 11248
rect 7104 11228 7156 11248
rect 7156 11228 7158 11248
rect 7102 11192 7158 11228
rect 6642 9560 6698 9616
rect 6550 8084 6606 8120
rect 6550 8064 6552 8084
rect 6552 8064 6604 8084
rect 6604 8064 6606 8084
rect 6274 6704 6330 6760
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 6366 4936 6422 4992
rect 6274 3712 6330 3768
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6550 6160 6606 6216
rect 7286 10412 7288 10432
rect 7288 10412 7340 10432
rect 7340 10412 7342 10432
rect 7286 10376 7342 10412
rect 6826 6060 6828 6080
rect 6828 6060 6880 6080
rect 6880 6060 6882 6080
rect 6826 6024 6882 6060
rect 6642 4664 6698 4720
rect 6550 3576 6606 3632
rect 7010 5208 7066 5264
rect 7286 7948 7342 7984
rect 7286 7928 7288 7948
rect 7288 7928 7340 7948
rect 7340 7928 7342 7948
rect 7286 7112 7342 7168
rect 7194 5072 7250 5128
rect 7194 4800 7250 4856
rect 6918 2896 6974 2952
rect 6918 2644 6974 2680
rect 6918 2624 6920 2644
rect 6920 2624 6972 2644
rect 6972 2624 6974 2644
rect 6642 2508 6698 2544
rect 6642 2488 6644 2508
rect 6644 2488 6696 2508
rect 6696 2488 6698 2508
rect 7194 3576 7250 3632
rect 7102 2916 7158 2952
rect 7102 2896 7104 2916
rect 7104 2896 7156 2916
rect 7156 2896 7158 2916
rect 7010 1536 7066 1592
rect 7562 10648 7618 10704
rect 7470 9288 7526 9344
rect 7562 7928 7618 7984
rect 7470 6840 7526 6896
rect 7562 6568 7618 6624
rect 8206 18284 8262 18320
rect 8206 18264 8208 18284
rect 8208 18264 8260 18284
rect 8260 18264 8262 18284
rect 8114 18028 8116 18048
rect 8116 18028 8168 18048
rect 8168 18028 8170 18048
rect 8114 17992 8170 18028
rect 8758 16940 8760 16960
rect 8760 16940 8812 16960
rect 8812 16940 8814 16960
rect 8758 16904 8814 16940
rect 8114 16496 8170 16552
rect 7838 11736 7894 11792
rect 7746 11192 7802 11248
rect 8022 10532 8078 10568
rect 8022 10512 8024 10532
rect 8024 10512 8076 10532
rect 8076 10512 8078 10532
rect 8022 8608 8078 8664
rect 8022 8336 8078 8392
rect 7746 7812 7802 7848
rect 7746 7792 7748 7812
rect 7748 7792 7800 7812
rect 7800 7792 7802 7812
rect 7930 7384 7986 7440
rect 7654 4936 7710 4992
rect 7470 3984 7526 4040
rect 7838 4684 7894 4720
rect 7838 4664 7840 4684
rect 7840 4664 7892 4684
rect 7892 4664 7894 4684
rect 7838 3460 7894 3496
rect 7838 3440 7840 3460
rect 7840 3440 7892 3460
rect 7892 3440 7894 3460
rect 7930 2760 7986 2816
rect 7838 1672 7894 1728
rect 8482 15000 8538 15056
rect 8850 14864 8906 14920
rect 9218 15020 9274 15056
rect 9218 15000 9220 15020
rect 9220 15000 9272 15020
rect 9272 15000 9274 15020
rect 9218 14728 9274 14784
rect 8942 13932 8998 13968
rect 8942 13912 8944 13932
rect 8944 13912 8996 13932
rect 8996 13912 8998 13932
rect 8298 13232 8354 13288
rect 8206 12552 8262 12608
rect 8206 10140 8208 10160
rect 8208 10140 8260 10160
rect 8260 10140 8262 10160
rect 8206 10104 8262 10140
rect 8666 12044 8668 12064
rect 8668 12044 8720 12064
rect 8720 12044 8722 12064
rect 8666 12008 8722 12044
rect 8574 11872 8630 11928
rect 8390 11736 8446 11792
rect 8390 10648 8446 10704
rect 8758 10104 8814 10160
rect 8206 8200 8262 8256
rect 8390 7520 8446 7576
rect 8574 6568 8630 6624
rect 8298 5208 8354 5264
rect 8206 3032 8262 3088
rect 8482 3440 8538 3496
rect 8666 2388 8668 2408
rect 8668 2388 8720 2408
rect 8720 2388 8722 2408
rect 8666 2352 8722 2388
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10598 18300 10600 18320
rect 10600 18300 10652 18320
rect 10652 18300 10654 18320
rect 10598 18264 10654 18300
rect 9678 17992 9734 18048
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10138 17620 10140 17640
rect 10140 17620 10192 17640
rect 10192 17620 10194 17640
rect 10138 17584 10194 17620
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 12714 23704 12770 23760
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 12898 20440 12954 20496
rect 12438 18128 12494 18184
rect 12622 17584 12678 17640
rect 11518 16360 11574 16416
rect 9586 15272 9642 15328
rect 9494 14884 9550 14920
rect 9494 14864 9496 14884
rect 9496 14864 9548 14884
rect 9548 14864 9550 14884
rect 10138 15000 10194 15056
rect 11150 14864 11206 14920
rect 9494 12044 9496 12064
rect 9496 12044 9548 12064
rect 9548 12044 9550 12064
rect 9494 12008 9550 12044
rect 9770 12552 9826 12608
rect 9862 12008 9918 12064
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 11058 13232 11114 13288
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 9770 10920 9826 10976
rect 9678 10376 9734 10432
rect 11058 11872 11114 11928
rect 9954 11620 10010 11656
rect 9954 11600 9956 11620
rect 9956 11600 10008 11620
rect 10008 11600 10010 11620
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 11242 12008 11298 12064
rect 10046 10260 10102 10296
rect 10046 10240 10048 10260
rect 10048 10240 10100 10260
rect 10100 10240 10102 10260
rect 9678 9288 9734 9344
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10138 9696 10194 9752
rect 10506 9596 10508 9616
rect 10508 9596 10560 9616
rect 10560 9596 10562 9616
rect 10506 9560 10562 9596
rect 10690 9288 10746 9344
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10598 9036 10654 9072
rect 10598 9016 10600 9036
rect 10600 9016 10652 9036
rect 10652 9016 10654 9036
rect 10782 9016 10838 9072
rect 9770 8744 9826 8800
rect 9494 6860 9550 6896
rect 9494 6840 9496 6860
rect 9496 6840 9548 6860
rect 9548 6840 9550 6860
rect 9494 3032 9550 3088
rect 10230 8472 10286 8528
rect 10138 8200 10194 8256
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10690 7540 10746 7576
rect 10690 7520 10692 7540
rect 10692 7520 10744 7540
rect 10744 7520 10746 7540
rect 10046 6976 10102 7032
rect 9862 6724 9918 6760
rect 9862 6704 9864 6724
rect 9864 6704 9916 6724
rect 9916 6704 9918 6724
rect 10046 6024 10102 6080
rect 10046 5616 10102 5672
rect 9954 3712 10010 3768
rect 9954 3304 10010 3360
rect 10782 7248 10838 7304
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10782 6024 10838 6080
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10690 5772 10746 5808
rect 10690 5752 10692 5772
rect 10692 5752 10744 5772
rect 10744 5752 10746 5772
rect 10782 5364 10838 5400
rect 10782 5344 10784 5364
rect 10784 5344 10836 5364
rect 10836 5344 10838 5364
rect 10690 4936 10746 4992
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10690 4256 10746 4312
rect 10506 4004 10562 4040
rect 10506 3984 10508 4004
rect 10508 3984 10560 4004
rect 10560 3984 10562 4004
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10782 3712 10838 3768
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11058 8064 11114 8120
rect 10966 7656 11022 7712
rect 11058 7112 11114 7168
rect 10966 5908 11022 5944
rect 10966 5888 10968 5908
rect 10968 5888 11020 5908
rect 11020 5888 11022 5908
rect 11334 5208 11390 5264
rect 11242 4392 11298 4448
rect 11058 4020 11060 4040
rect 11060 4020 11112 4040
rect 11112 4020 11114 4040
rect 11058 3984 11114 4020
rect 10966 3848 11022 3904
rect 11978 15000 12034 15056
rect 11886 12980 11942 13016
rect 11886 12960 11888 12980
rect 11888 12960 11940 12980
rect 11940 12960 11942 12980
rect 11886 11192 11942 11248
rect 11610 10920 11666 10976
rect 11702 10240 11758 10296
rect 11794 8744 11850 8800
rect 11518 7112 11574 7168
rect 11518 6860 11574 6896
rect 11518 6840 11520 6860
rect 11520 6840 11572 6860
rect 11572 6840 11574 6860
rect 11886 4664 11942 4720
rect 11610 3032 11666 3088
rect 11702 2488 11758 2544
rect 12438 15136 12494 15192
rect 12254 10512 12310 10568
rect 12162 8608 12218 8664
rect 12438 8336 12494 8392
rect 12438 5752 12494 5808
rect 12162 3576 12218 3632
rect 12070 2624 12126 2680
rect 12438 2624 12494 2680
rect 12438 2216 12494 2272
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 15382 19760 15438 19816
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 13266 13232 13322 13288
rect 13266 11464 13322 11520
rect 12898 8472 12954 8528
rect 12622 7928 12678 7984
rect 12806 7812 12862 7848
rect 12806 7792 12808 7812
rect 12808 7792 12860 7812
rect 12860 7792 12862 7812
rect 13358 8200 13414 8256
rect 13358 7384 13414 7440
rect 12622 3576 12678 3632
rect 12990 5344 13046 5400
rect 13358 5072 13414 5128
rect 13358 4800 13414 4856
rect 13266 4528 13322 4584
rect 13358 3712 13414 3768
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14002 13268 14004 13288
rect 14004 13268 14056 13288
rect 14056 13268 14058 13288
rect 14002 13232 14058 13268
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14002 12824 14058 12880
rect 15290 12824 15346 12880
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24674 19488 24730 19544
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 24030 15544 24086 15600
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 23662 14320 23718 14376
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 23386 13388 23442 13424
rect 23386 13368 23388 13388
rect 23388 13368 23440 13388
rect 23440 13368 23442 13388
rect 16670 13252 16726 13288
rect 16670 13232 16672 13252
rect 16672 13232 16724 13252
rect 16724 13232 16726 13252
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 22282 12300 22338 12336
rect 22282 12280 22284 12300
rect 22284 12280 22336 12300
rect 22336 12280 22338 12300
rect 15566 11736 15622 11792
rect 13910 10648 13966 10704
rect 13818 10104 13874 10160
rect 14462 10240 14518 10296
rect 13818 9696 13874 9752
rect 13818 9052 13820 9072
rect 13820 9052 13872 9072
rect 13872 9052 13874 9072
rect 13818 9016 13874 9052
rect 13542 8508 13544 8528
rect 13544 8508 13596 8528
rect 13596 8508 13598 8528
rect 13542 8472 13598 8508
rect 13726 6976 13782 7032
rect 14278 8200 14334 8256
rect 14002 6568 14058 6624
rect 14186 6296 14242 6352
rect 13910 5652 13912 5672
rect 13912 5652 13964 5672
rect 13964 5652 13966 5672
rect 13910 5616 13966 5652
rect 14186 5616 14242 5672
rect 13634 5092 13690 5128
rect 13634 5072 13636 5092
rect 13636 5072 13688 5092
rect 13688 5072 13690 5092
rect 13634 4936 13690 4992
rect 12898 3304 12954 3360
rect 12898 2760 12954 2816
rect 12714 2624 12770 2680
rect 13542 2372 13598 2408
rect 13542 2352 13544 2372
rect 13544 2352 13596 2372
rect 13596 2352 13598 2372
rect 13542 1672 13598 1728
rect 13542 1400 13598 1456
rect 14094 4684 14150 4720
rect 14094 4664 14096 4684
rect 14096 4664 14148 4684
rect 14148 4664 14150 4684
rect 13818 2372 13874 2408
rect 13818 2352 13820 2372
rect 13820 2352 13872 2372
rect 13872 2352 13874 2372
rect 13726 2216 13782 2272
rect 13726 1672 13782 1728
rect 14462 8900 14518 8936
rect 14462 8880 14464 8900
rect 14464 8880 14516 8900
rect 14516 8880 14518 8900
rect 14370 8064 14426 8120
rect 14462 5480 14518 5536
rect 14462 4936 14518 4992
rect 15750 11600 15806 11656
rect 15658 11500 15660 11520
rect 15660 11500 15712 11520
rect 15712 11500 15714 11520
rect 15658 11464 15714 11500
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 15290 10004 15292 10024
rect 15292 10004 15344 10024
rect 15344 10004 15346 10024
rect 15290 9968 15346 10004
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14738 6976 14794 7032
rect 15474 9288 15530 9344
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15382 6724 15438 6760
rect 15382 6704 15384 6724
rect 15384 6704 15436 6724
rect 15436 6704 15438 6724
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15382 6024 15438 6080
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15382 5480 15438 5536
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15290 3712 15346 3768
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14554 1808 14610 1864
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15290 1536 15346 1592
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 16302 8608 16358 8664
rect 22282 8608 22338 8664
rect 16762 8472 16818 8528
rect 15566 7656 15622 7712
rect 15750 6976 15806 7032
rect 16302 7148 16304 7168
rect 16304 7148 16356 7168
rect 16356 7148 16358 7168
rect 16302 7112 16358 7148
rect 20902 8372 20904 8392
rect 20904 8372 20956 8392
rect 20956 8372 20958 8392
rect 20902 8336 20958 8372
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19154 7656 19210 7712
rect 18050 7284 18052 7304
rect 18052 7284 18104 7304
rect 18104 7284 18106 7304
rect 18050 7248 18106 7284
rect 16302 5908 16358 5944
rect 16302 5888 16304 5908
rect 16304 5888 16356 5908
rect 16356 5888 16358 5908
rect 15658 5228 15714 5264
rect 15658 5208 15660 5228
rect 15660 5208 15712 5228
rect 15712 5208 15714 5228
rect 16854 5636 16910 5672
rect 16854 5616 16856 5636
rect 16856 5616 16908 5636
rect 16908 5616 16910 5636
rect 17774 6196 17776 6216
rect 17776 6196 17828 6216
rect 17828 6196 17830 6216
rect 17774 6160 17830 6196
rect 16394 5072 16450 5128
rect 15750 4820 15806 4856
rect 15750 4800 15752 4820
rect 15752 4800 15804 4820
rect 15804 4800 15806 4820
rect 15658 4684 15714 4720
rect 15658 4664 15660 4684
rect 15660 4664 15712 4684
rect 15712 4664 15714 4684
rect 15658 3032 15714 3088
rect 15934 2760 15990 2816
rect 17958 3848 18014 3904
rect 18050 3576 18106 3632
rect 17774 3440 17830 3496
rect 17038 3168 17094 3224
rect 16026 2488 16082 2544
rect 17774 2916 17830 2952
rect 17774 2896 17776 2916
rect 17776 2896 17828 2916
rect 17828 2896 17830 2916
rect 17590 2760 17646 2816
rect 17682 2644 17738 2680
rect 17682 2624 17684 2644
rect 17684 2624 17736 2644
rect 17736 2624 17738 2644
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 20902 6704 20958 6760
rect 20534 6296 20590 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19522 5752 19578 5808
rect 19338 4936 19394 4992
rect 18326 3984 18382 4040
rect 18694 3712 18750 3768
rect 18510 3576 18566 3632
rect 18694 3440 18750 3496
rect 18510 3032 18566 3088
rect 18326 1808 18382 1864
rect 18510 1672 18566 1728
rect 19246 3304 19302 3360
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20074 3732 20130 3768
rect 20074 3712 20076 3732
rect 20076 3712 20128 3732
rect 20128 3712 20130 3732
rect 19982 3168 20038 3224
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19338 2624 19394 2680
rect 19798 2488 19854 2544
rect 19614 1400 19670 1456
rect 20810 5480 20866 5536
rect 20902 4020 20904 4040
rect 20904 4020 20956 4040
rect 20956 4020 20958 4040
rect 20902 3984 20958 4020
rect 21086 3984 21142 4040
rect 20534 2488 20590 2544
rect 21086 3304 21142 3360
rect 21178 3032 21234 3088
rect 21178 2352 21234 2408
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 22834 10648 22890 10704
rect 22466 5616 22522 5672
rect 22558 3984 22614 4040
rect 22466 3440 22522 3496
rect 22374 3168 22430 3224
rect 22466 2508 22522 2544
rect 22466 2488 22468 2508
rect 22468 2488 22520 2508
rect 22520 2488 22522 2508
rect 22650 2896 22706 2952
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24214 8336 24270 8392
rect 24030 5616 24086 5672
rect 22834 2760 22890 2816
rect 23938 3712 23994 3768
rect 23662 3032 23718 3088
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24766 13912 24822 13968
rect 24766 13232 24822 13288
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24674 4120 24730 4176
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 25318 4548 25374 4584
rect 25318 4528 25320 4548
rect 25320 4528 25372 4548
rect 25372 4528 25374 4548
rect 24766 3032 24822 3088
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 27618 3032 27674 3088
rect 27066 2896 27122 2952
rect 2962 312 3018 368
<< metal3 >>
rect 0 27706 480 27736
rect 2773 27706 2839 27709
rect 0 27704 2839 27706
rect 0 27648 2778 27704
rect 2834 27648 2839 27704
rect 0 27646 2839 27648
rect 0 27616 480 27646
rect 2773 27643 2839 27646
rect 0 27162 480 27192
rect 3325 27162 3391 27165
rect 0 27160 3391 27162
rect 0 27104 3330 27160
rect 3386 27104 3391 27160
rect 0 27102 3391 27104
rect 0 27072 480 27102
rect 3325 27099 3391 27102
rect 0 26618 480 26648
rect 3233 26618 3299 26621
rect 0 26616 3299 26618
rect 0 26560 3238 26616
rect 3294 26560 3299 26616
rect 0 26558 3299 26560
rect 0 26528 480 26558
rect 3233 26555 3299 26558
rect 0 26074 480 26104
rect 2681 26074 2747 26077
rect 0 26072 2747 26074
rect 0 26016 2686 26072
rect 2742 26016 2747 26072
rect 0 26014 2747 26016
rect 0 25984 480 26014
rect 2681 26011 2747 26014
rect 10277 25600 10597 25601
rect 0 25530 480 25560
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 1577 25530 1643 25533
rect 0 25528 1643 25530
rect 0 25472 1582 25528
rect 1638 25472 1643 25528
rect 0 25470 1643 25472
rect 0 25440 480 25470
rect 1577 25467 1643 25470
rect 24761 25122 24827 25125
rect 27520 25122 28000 25152
rect 24761 25120 28000 25122
rect 24761 25064 24766 25120
rect 24822 25064 28000 25120
rect 24761 25062 28000 25064
rect 24761 25059 24827 25062
rect 5610 25056 5930 25057
rect 0 24986 480 25016
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 27520 25032 28000 25062
rect 24277 24991 24597 24992
rect 1485 24986 1551 24989
rect 0 24984 1551 24986
rect 0 24928 1490 24984
rect 1546 24928 1551 24984
rect 0 24926 1551 24928
rect 0 24896 480 24926
rect 1485 24923 1551 24926
rect 10277 24512 10597 24513
rect 0 24442 480 24472
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 2957 24442 3023 24445
rect 0 24440 3023 24442
rect 0 24384 2962 24440
rect 3018 24384 3023 24440
rect 0 24382 3023 24384
rect 0 24352 480 24382
rect 2957 24379 3023 24382
rect 2037 24170 2103 24173
rect 11973 24170 12039 24173
rect 2037 24168 12039 24170
rect 2037 24112 2042 24168
rect 2098 24112 11978 24168
rect 12034 24112 12039 24168
rect 2037 24110 12039 24112
rect 2037 24107 2103 24110
rect 11973 24107 12039 24110
rect 5610 23968 5930 23969
rect 0 23898 480 23928
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 2681 23898 2747 23901
rect 0 23896 2747 23898
rect 0 23840 2686 23896
rect 2742 23840 2747 23896
rect 0 23838 2747 23840
rect 0 23808 480 23838
rect 2681 23835 2747 23838
rect 3693 23762 3759 23765
rect 12709 23762 12775 23765
rect 3693 23760 12775 23762
rect 3693 23704 3698 23760
rect 3754 23704 12714 23760
rect 12770 23704 12775 23760
rect 3693 23702 12775 23704
rect 3693 23699 3759 23702
rect 12709 23699 12775 23702
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23218 480 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 480 23158
rect 1485 23155 1551 23158
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 0 22674 480 22704
rect 3417 22674 3483 22677
rect 0 22672 3483 22674
rect 0 22616 3422 22672
rect 3478 22616 3483 22672
rect 0 22614 3483 22616
rect 0 22584 480 22614
rect 3417 22611 3483 22614
rect 1669 22538 1735 22541
rect 10777 22538 10843 22541
rect 1669 22536 10843 22538
rect 1669 22480 1674 22536
rect 1730 22480 10782 22536
rect 10838 22480 10843 22536
rect 1669 22478 10843 22480
rect 1669 22475 1735 22478
rect 10777 22475 10843 22478
rect 2589 22402 2655 22405
rect 4429 22402 4495 22405
rect 2589 22400 4495 22402
rect 2589 22344 2594 22400
rect 2650 22344 4434 22400
rect 4490 22344 4495 22400
rect 2589 22342 4495 22344
rect 2589 22339 2655 22342
rect 4429 22339 4495 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 0 22130 480 22160
rect 4061 22130 4127 22133
rect 0 22128 4127 22130
rect 0 22072 4066 22128
rect 4122 22072 4127 22128
rect 0 22070 4127 22072
rect 0 22040 480 22070
rect 4061 22067 4127 22070
rect 3417 21994 3483 21997
rect 8569 21994 8635 21997
rect 3417 21992 8635 21994
rect 3417 21936 3422 21992
rect 3478 21936 8574 21992
rect 8630 21936 8635 21992
rect 3417 21934 8635 21936
rect 3417 21931 3483 21934
rect 8569 21931 8635 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21586 480 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 480 21526
rect 2681 21523 2747 21526
rect 2405 21450 2471 21453
rect 7281 21450 7347 21453
rect 2405 21448 7347 21450
rect 2405 21392 2410 21448
rect 2466 21392 7286 21448
rect 7342 21392 7347 21448
rect 2405 21390 7347 21392
rect 2405 21387 2471 21390
rect 7281 21387 7347 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 0 21042 480 21072
rect 1577 21042 1643 21045
rect 0 21040 1643 21042
rect 0 20984 1582 21040
rect 1638 20984 1643 21040
rect 0 20982 1643 20984
rect 0 20952 480 20982
rect 1577 20979 1643 20982
rect 1669 20906 1735 20909
rect 8109 20906 8175 20909
rect 1669 20904 8175 20906
rect 1669 20848 1674 20904
rect 1730 20848 8114 20904
rect 8170 20848 8175 20904
rect 1669 20846 8175 20848
rect 1669 20843 1735 20846
rect 8109 20843 8175 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 2589 20634 2655 20637
rect 2589 20632 4354 20634
rect 2589 20576 2594 20632
rect 2650 20576 4354 20632
rect 2589 20574 4354 20576
rect 2589 20571 2655 20574
rect 0 20498 480 20528
rect 2681 20498 2747 20501
rect 4153 20498 4219 20501
rect 0 20438 2514 20498
rect 0 20408 480 20438
rect 2454 20226 2514 20438
rect 2681 20496 4219 20498
rect 2681 20440 2686 20496
rect 2742 20440 4158 20496
rect 4214 20440 4219 20496
rect 2681 20438 4219 20440
rect 4294 20498 4354 20574
rect 12893 20498 12959 20501
rect 4294 20496 12959 20498
rect 4294 20440 12898 20496
rect 12954 20440 12959 20496
rect 4294 20438 12959 20440
rect 2681 20435 2747 20438
rect 4153 20435 4219 20438
rect 12893 20435 12959 20438
rect 4245 20226 4311 20229
rect 2454 20224 4311 20226
rect 2454 20168 4250 20224
rect 4306 20168 4311 20224
rect 2454 20166 4311 20168
rect 4245 20163 4311 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 3693 20090 3759 20093
rect 7373 20090 7439 20093
rect 3693 20088 7439 20090
rect 3693 20032 3698 20088
rect 3754 20032 7378 20088
rect 7434 20032 7439 20088
rect 3693 20030 7439 20032
rect 3693 20027 3759 20030
rect 7373 20027 7439 20030
rect 0 19954 480 19984
rect 3233 19954 3299 19957
rect 0 19952 3299 19954
rect 0 19896 3238 19952
rect 3294 19896 3299 19952
rect 0 19894 3299 19896
rect 0 19864 480 19894
rect 3233 19891 3299 19894
rect 1761 19818 1827 19821
rect 15377 19818 15443 19821
rect 1761 19816 15443 19818
rect 1761 19760 1766 19816
rect 1822 19760 15382 19816
rect 15438 19760 15443 19816
rect 1761 19758 15443 19760
rect 1761 19755 1827 19758
rect 15377 19755 15443 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 24669 19546 24735 19549
rect 27520 19546 28000 19576
rect 24669 19544 28000 19546
rect 24669 19488 24674 19544
rect 24730 19488 28000 19544
rect 24669 19486 28000 19488
rect 24669 19483 24735 19486
rect 27520 19456 28000 19486
rect 0 19410 480 19440
rect 4613 19410 4679 19413
rect 0 19408 4679 19410
rect 0 19352 4618 19408
rect 4674 19352 4679 19408
rect 0 19350 4679 19352
rect 0 19320 480 19350
rect 4613 19347 4679 19350
rect 1669 19138 1735 19141
rect 6821 19138 6887 19141
rect 1669 19136 6887 19138
rect 1669 19080 1674 19136
rect 1730 19080 6826 19136
rect 6882 19080 6887 19136
rect 1669 19078 6887 19080
rect 1669 19075 1735 19078
rect 6821 19075 6887 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 2681 19002 2747 19005
rect 4061 19002 4127 19005
rect 2681 19000 4127 19002
rect 2681 18944 2686 19000
rect 2742 18944 4066 19000
rect 4122 18944 4127 19000
rect 2681 18942 4127 18944
rect 2681 18939 2747 18942
rect 4061 18939 4127 18942
rect 0 18730 480 18760
rect 4245 18730 4311 18733
rect 0 18728 4311 18730
rect 0 18672 4250 18728
rect 4306 18672 4311 18728
rect 0 18670 4311 18672
rect 0 18640 480 18670
rect 4245 18667 4311 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 8201 18322 8267 18325
rect 10593 18322 10659 18325
rect 8201 18320 10659 18322
rect 8201 18264 8206 18320
rect 8262 18264 10598 18320
rect 10654 18264 10659 18320
rect 8201 18262 10659 18264
rect 8201 18259 8267 18262
rect 10593 18259 10659 18262
rect 0 18186 480 18216
rect 2865 18186 2931 18189
rect 0 18184 2931 18186
rect 0 18128 2870 18184
rect 2926 18128 2931 18184
rect 0 18126 2931 18128
rect 0 18096 480 18126
rect 2865 18123 2931 18126
rect 4429 18186 4495 18189
rect 12433 18186 12499 18189
rect 4429 18184 12499 18186
rect 4429 18128 4434 18184
rect 4490 18128 12438 18184
rect 12494 18128 12499 18184
rect 4429 18126 12499 18128
rect 4429 18123 4495 18126
rect 12433 18123 12499 18126
rect 8109 18050 8175 18053
rect 9673 18050 9739 18053
rect 8109 18048 9739 18050
rect 8109 17992 8114 18048
rect 8170 17992 9678 18048
rect 9734 17992 9739 18048
rect 8109 17990 9739 17992
rect 8109 17987 8175 17990
rect 9673 17987 9739 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 0 17642 480 17672
rect 3049 17642 3115 17645
rect 0 17640 3115 17642
rect 0 17584 3054 17640
rect 3110 17584 3115 17640
rect 0 17582 3115 17584
rect 0 17552 480 17582
rect 3049 17579 3115 17582
rect 10133 17642 10199 17645
rect 12617 17642 12683 17645
rect 10133 17640 12683 17642
rect 10133 17584 10138 17640
rect 10194 17584 12622 17640
rect 12678 17584 12683 17640
rect 10133 17582 12683 17584
rect 10133 17579 10199 17582
rect 12617 17579 12683 17582
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 0 17098 480 17128
rect 3969 17098 4035 17101
rect 0 17096 4035 17098
rect 0 17040 3974 17096
rect 4030 17040 4035 17096
rect 0 17038 4035 17040
rect 0 17008 480 17038
rect 3969 17035 4035 17038
rect 5257 16962 5323 16965
rect 8753 16962 8819 16965
rect 5257 16960 8819 16962
rect 5257 16904 5262 16960
rect 5318 16904 8758 16960
rect 8814 16904 8819 16960
rect 5257 16902 8819 16904
rect 5257 16899 5323 16902
rect 8753 16899 8819 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 1577 16690 1643 16693
rect 3785 16690 3851 16693
rect 1577 16688 3851 16690
rect 1577 16632 1582 16688
rect 1638 16632 3790 16688
rect 3846 16632 3851 16688
rect 1577 16630 3851 16632
rect 1577 16627 1643 16630
rect 3785 16627 3851 16630
rect 5349 16690 5415 16693
rect 5349 16688 7114 16690
rect 5349 16632 5354 16688
rect 5410 16632 7114 16688
rect 5349 16630 7114 16632
rect 5349 16627 5415 16630
rect 0 16554 480 16584
rect 3233 16554 3299 16557
rect 6821 16554 6887 16557
rect 0 16494 3112 16554
rect 0 16464 480 16494
rect 3052 16418 3112 16494
rect 3233 16552 6887 16554
rect 3233 16496 3238 16552
rect 3294 16496 6826 16552
rect 6882 16496 6887 16552
rect 3233 16494 6887 16496
rect 7054 16554 7114 16630
rect 8109 16554 8175 16557
rect 7054 16552 8175 16554
rect 7054 16496 8114 16552
rect 8170 16496 8175 16552
rect 7054 16494 8175 16496
rect 3233 16491 3299 16494
rect 6821 16491 6887 16494
rect 8109 16491 8175 16494
rect 3693 16418 3759 16421
rect 3052 16416 3759 16418
rect 3052 16360 3698 16416
rect 3754 16360 3759 16416
rect 3052 16358 3759 16360
rect 3693 16355 3759 16358
rect 6085 16418 6151 16421
rect 6637 16418 6703 16421
rect 11513 16418 11579 16421
rect 6085 16416 11579 16418
rect 6085 16360 6090 16416
rect 6146 16360 6642 16416
rect 6698 16360 11518 16416
rect 11574 16360 11579 16416
rect 6085 16358 11579 16360
rect 6085 16355 6151 16358
rect 6637 16355 6703 16358
rect 11513 16355 11579 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 3969 16146 4035 16149
rect 7005 16146 7071 16149
rect 3969 16144 7071 16146
rect 3969 16088 3974 16144
rect 4030 16088 7010 16144
rect 7066 16088 7071 16144
rect 3969 16086 7071 16088
rect 3969 16083 4035 16086
rect 7005 16083 7071 16086
rect 0 16010 480 16040
rect 3785 16010 3851 16013
rect 0 16008 3851 16010
rect 0 15952 3790 16008
rect 3846 15952 3851 16008
rect 0 15950 3851 15952
rect 0 15920 480 15950
rect 3785 15947 3851 15950
rect 1393 15874 1459 15877
rect 7189 15874 7255 15877
rect 1393 15872 7255 15874
rect 1393 15816 1398 15872
rect 1454 15816 7194 15872
rect 7250 15816 7255 15872
rect 1393 15814 7255 15816
rect 1393 15811 1459 15814
rect 7189 15811 7255 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 24025 15602 24091 15605
rect 3512 15600 24091 15602
rect 3512 15544 24030 15600
rect 24086 15544 24091 15600
rect 3512 15542 24091 15544
rect 0 15466 480 15496
rect 3512 15466 3572 15542
rect 24025 15539 24091 15542
rect 0 15406 3572 15466
rect 0 15376 480 15406
rect 6545 15330 6611 15333
rect 9581 15330 9647 15333
rect 6545 15328 9647 15330
rect 6545 15272 6550 15328
rect 6606 15272 9586 15328
rect 9642 15272 9647 15328
rect 6545 15270 9647 15272
rect 6545 15267 6611 15270
rect 9581 15267 9647 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 6269 15194 6335 15197
rect 7373 15194 7439 15197
rect 12433 15194 12499 15197
rect 6269 15192 12499 15194
rect 6269 15136 6274 15192
rect 6330 15136 7378 15192
rect 7434 15136 12438 15192
rect 12494 15136 12499 15192
rect 6269 15134 12499 15136
rect 6269 15131 6335 15134
rect 7373 15131 7439 15134
rect 12433 15131 12499 15134
rect 2313 15058 2379 15061
rect 2773 15058 2839 15061
rect 6821 15058 6887 15061
rect 8477 15058 8543 15061
rect 2313 15056 6194 15058
rect 2313 15000 2318 15056
rect 2374 15000 2778 15056
rect 2834 15000 6194 15056
rect 2313 14998 6194 15000
rect 2313 14995 2379 14998
rect 2773 14995 2839 14998
rect 0 14922 480 14952
rect 5993 14922 6059 14925
rect 0 14920 6059 14922
rect 0 14864 5998 14920
rect 6054 14864 6059 14920
rect 0 14862 6059 14864
rect 6134 14922 6194 14998
rect 6821 15056 8543 15058
rect 6821 15000 6826 15056
rect 6882 15000 8482 15056
rect 8538 15000 8543 15056
rect 6821 14998 8543 15000
rect 6821 14995 6887 14998
rect 8477 14995 8543 14998
rect 9213 15058 9279 15061
rect 10133 15058 10199 15061
rect 11973 15058 12039 15061
rect 9213 15056 12039 15058
rect 9213 15000 9218 15056
rect 9274 15000 10138 15056
rect 10194 15000 11978 15056
rect 12034 15000 12039 15056
rect 9213 14998 12039 15000
rect 9213 14995 9279 14998
rect 10133 14995 10199 14998
rect 11973 14995 12039 14998
rect 6453 14922 6519 14925
rect 8845 14922 8911 14925
rect 6134 14920 8911 14922
rect 6134 14864 6458 14920
rect 6514 14864 8850 14920
rect 8906 14864 8911 14920
rect 6134 14862 8911 14864
rect 0 14832 480 14862
rect 5993 14859 6059 14862
rect 6453 14859 6519 14862
rect 8845 14859 8911 14862
rect 9489 14922 9555 14925
rect 11145 14922 11211 14925
rect 9489 14920 11211 14922
rect 9489 14864 9494 14920
rect 9550 14864 11150 14920
rect 11206 14864 11211 14920
rect 9489 14862 11211 14864
rect 9489 14859 9555 14862
rect 11145 14859 11211 14862
rect 6637 14786 6703 14789
rect 7557 14786 7623 14789
rect 9213 14786 9279 14789
rect 6637 14784 9279 14786
rect 6637 14728 6642 14784
rect 6698 14728 7562 14784
rect 7618 14728 9218 14784
rect 9274 14728 9279 14784
rect 6637 14726 9279 14728
rect 6637 14723 6703 14726
rect 7557 14723 7623 14726
rect 9213 14723 9279 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 2497 14650 2563 14653
rect 2865 14650 2931 14653
rect 7833 14650 7899 14653
rect 2497 14648 7899 14650
rect 2497 14592 2502 14648
rect 2558 14592 2870 14648
rect 2926 14592 7838 14648
rect 7894 14592 7899 14648
rect 2497 14590 7899 14592
rect 2497 14587 2563 14590
rect 2865 14587 2931 14590
rect 7833 14587 7899 14590
rect 2405 14514 2471 14517
rect 6545 14514 6611 14517
rect 2405 14512 6611 14514
rect 2405 14456 2410 14512
rect 2466 14456 6550 14512
rect 6606 14456 6611 14512
rect 2405 14454 6611 14456
rect 2405 14451 2471 14454
rect 6545 14451 6611 14454
rect 0 14378 480 14408
rect 23657 14378 23723 14381
rect 0 14376 23723 14378
rect 0 14320 23662 14376
rect 23718 14320 23723 14376
rect 0 14318 23723 14320
rect 0 14288 480 14318
rect 23657 14315 23723 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 2313 13970 2379 13973
rect 4245 13970 4311 13973
rect 4613 13970 4679 13973
rect 2313 13968 4679 13970
rect 2313 13912 2318 13968
rect 2374 13912 4250 13968
rect 4306 13912 4618 13968
rect 4674 13912 4679 13968
rect 2313 13910 4679 13912
rect 2313 13907 2379 13910
rect 4245 13907 4311 13910
rect 4613 13907 4679 13910
rect 5717 13970 5783 13973
rect 8937 13970 9003 13973
rect 5717 13968 9003 13970
rect 5717 13912 5722 13968
rect 5778 13912 8942 13968
rect 8998 13912 9003 13968
rect 5717 13910 9003 13912
rect 5717 13907 5783 13910
rect 8937 13907 9003 13910
rect 24761 13970 24827 13973
rect 27520 13970 28000 14000
rect 24761 13968 28000 13970
rect 24761 13912 24766 13968
rect 24822 13912 28000 13968
rect 24761 13910 28000 13912
rect 24761 13907 24827 13910
rect 27520 13880 28000 13910
rect 5349 13834 5415 13837
rect 7373 13834 7439 13837
rect 5349 13832 7439 13834
rect 5349 13776 5354 13832
rect 5410 13776 7378 13832
rect 7434 13776 7439 13832
rect 5349 13774 7439 13776
rect 5349 13771 5415 13774
rect 7373 13771 7439 13774
rect 0 13698 480 13728
rect 3417 13698 3483 13701
rect 0 13696 3483 13698
rect 0 13640 3422 13696
rect 3478 13640 3483 13696
rect 0 13638 3483 13640
rect 0 13608 480 13638
rect 3417 13635 3483 13638
rect 4705 13698 4771 13701
rect 7281 13698 7347 13701
rect 4705 13696 7347 13698
rect 4705 13640 4710 13696
rect 4766 13640 7286 13696
rect 7342 13640 7347 13696
rect 4705 13638 7347 13640
rect 4705 13635 4771 13638
rect 7281 13635 7347 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 5993 13426 6059 13429
rect 23381 13426 23447 13429
rect 5993 13424 23447 13426
rect 5993 13368 5998 13424
rect 6054 13368 23386 13424
rect 23442 13368 23447 13424
rect 5993 13366 23447 13368
rect 5993 13363 6059 13366
rect 23381 13363 23447 13366
rect 8293 13290 8359 13293
rect 11053 13290 11119 13293
rect 8293 13288 11119 13290
rect 8293 13232 8298 13288
rect 8354 13232 11058 13288
rect 11114 13232 11119 13288
rect 8293 13230 11119 13232
rect 8293 13227 8359 13230
rect 11053 13227 11119 13230
rect 13261 13290 13327 13293
rect 13997 13290 14063 13293
rect 16665 13290 16731 13293
rect 24761 13290 24827 13293
rect 13261 13288 24827 13290
rect 13261 13232 13266 13288
rect 13322 13232 14002 13288
rect 14058 13232 16670 13288
rect 16726 13232 24766 13288
rect 24822 13232 24827 13288
rect 13261 13230 24827 13232
rect 13261 13227 13327 13230
rect 13997 13227 14063 13230
rect 16665 13227 16731 13230
rect 24761 13227 24827 13230
rect 0 13154 480 13184
rect 1853 13154 1919 13157
rect 4613 13154 4679 13157
rect 0 13094 1778 13154
rect 0 13064 480 13094
rect 1718 13018 1778 13094
rect 1853 13152 4679 13154
rect 1853 13096 1858 13152
rect 1914 13096 4618 13152
rect 4674 13096 4679 13152
rect 1853 13094 4679 13096
rect 1853 13091 1919 13094
rect 4613 13091 4679 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 3601 13018 3667 13021
rect 1718 13016 3667 13018
rect 1718 12960 3606 13016
rect 3662 12960 3667 13016
rect 1718 12958 3667 12960
rect 3601 12955 3667 12958
rect 11881 13018 11947 13021
rect 11881 13016 14842 13018
rect 11881 12960 11886 13016
rect 11942 12960 14842 13016
rect 11881 12958 14842 12960
rect 11881 12955 11947 12958
rect 13997 12882 14063 12885
rect 9860 12880 14063 12882
rect 9860 12824 14002 12880
rect 14058 12824 14063 12880
rect 9860 12822 14063 12824
rect 14782 12882 14842 12958
rect 15285 12882 15351 12885
rect 14782 12880 15351 12882
rect 14782 12824 15290 12880
rect 15346 12824 15351 12880
rect 14782 12822 15351 12824
rect 2957 12746 3023 12749
rect 9860 12746 9920 12822
rect 13997 12819 14063 12822
rect 15285 12819 15351 12822
rect 2957 12744 9920 12746
rect 2957 12688 2962 12744
rect 3018 12688 9920 12744
rect 2957 12686 9920 12688
rect 9998 12686 12450 12746
rect 2957 12683 3023 12686
rect 0 12610 480 12640
rect 3509 12610 3575 12613
rect 0 12608 3575 12610
rect 0 12552 3514 12608
rect 3570 12552 3575 12608
rect 0 12550 3575 12552
rect 0 12520 480 12550
rect 3509 12547 3575 12550
rect 8201 12610 8267 12613
rect 9765 12610 9831 12613
rect 8201 12608 9831 12610
rect 8201 12552 8206 12608
rect 8262 12552 9770 12608
rect 9826 12552 9831 12608
rect 8201 12550 9831 12552
rect 8201 12547 8267 12550
rect 9765 12547 9831 12550
rect 3417 12474 3483 12477
rect 9998 12474 10058 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 3417 12472 10058 12474
rect 3417 12416 3422 12472
rect 3478 12416 10058 12472
rect 3417 12414 10058 12416
rect 3417 12411 3483 12414
rect 12390 12338 12450 12686
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 22277 12338 22343 12341
rect 12390 12336 22343 12338
rect 12390 12280 22282 12336
rect 22338 12280 22343 12336
rect 12390 12278 22343 12280
rect 22277 12275 22343 12278
rect 3785 12202 3851 12205
rect 5533 12202 5599 12205
rect 3785 12200 5599 12202
rect 3785 12144 3790 12200
rect 3846 12144 5538 12200
rect 5594 12144 5599 12200
rect 3785 12142 5599 12144
rect 3785 12139 3851 12142
rect 5533 12139 5599 12142
rect 0 12066 480 12096
rect 3785 12066 3851 12069
rect 0 12064 3851 12066
rect 0 12008 3790 12064
rect 3846 12008 3851 12064
rect 0 12006 3851 12008
rect 0 11976 480 12006
rect 3785 12003 3851 12006
rect 6637 12066 6703 12069
rect 8661 12066 8727 12069
rect 6637 12064 8727 12066
rect 6637 12008 6642 12064
rect 6698 12008 8666 12064
rect 8722 12008 8727 12064
rect 6637 12006 8727 12008
rect 6637 12003 6703 12006
rect 8661 12003 8727 12006
rect 9489 12066 9555 12069
rect 9857 12066 9923 12069
rect 11237 12066 11303 12069
rect 9489 12064 11303 12066
rect 9489 12008 9494 12064
rect 9550 12008 9862 12064
rect 9918 12008 11242 12064
rect 11298 12008 11303 12064
rect 9489 12006 11303 12008
rect 9489 12003 9555 12006
rect 9857 12003 9923 12006
rect 11237 12003 11303 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 8569 11930 8635 11933
rect 11053 11930 11119 11933
rect 8569 11928 11119 11930
rect 8569 11872 8574 11928
rect 8630 11872 11058 11928
rect 11114 11872 11119 11928
rect 8569 11870 11119 11872
rect 8569 11867 8635 11870
rect 11053 11867 11119 11870
rect 1945 11794 2011 11797
rect 4337 11794 4403 11797
rect 7833 11794 7899 11797
rect 1945 11792 7899 11794
rect 1945 11736 1950 11792
rect 2006 11736 4342 11792
rect 4398 11736 7838 11792
rect 7894 11736 7899 11792
rect 1945 11734 7899 11736
rect 1945 11731 2011 11734
rect 4337 11731 4403 11734
rect 7833 11731 7899 11734
rect 8385 11794 8451 11797
rect 15561 11794 15627 11797
rect 8385 11792 15627 11794
rect 8385 11736 8390 11792
rect 8446 11736 15566 11792
rect 15622 11736 15627 11792
rect 8385 11734 15627 11736
rect 8385 11731 8451 11734
rect 15561 11731 15627 11734
rect 9949 11658 10015 11661
rect 15745 11658 15811 11661
rect 9949 11656 15811 11658
rect 9949 11600 9954 11656
rect 10010 11600 15750 11656
rect 15806 11600 15811 11656
rect 9949 11598 15811 11600
rect 9949 11595 10015 11598
rect 15745 11595 15811 11598
rect 0 11522 480 11552
rect 3233 11522 3299 11525
rect 0 11520 3299 11522
rect 0 11464 3238 11520
rect 3294 11464 3299 11520
rect 0 11462 3299 11464
rect 0 11432 480 11462
rect 3233 11459 3299 11462
rect 13261 11522 13327 11525
rect 15653 11522 15719 11525
rect 13261 11520 15719 11522
rect 13261 11464 13266 11520
rect 13322 11464 15658 11520
rect 15714 11464 15719 11520
rect 13261 11462 15719 11464
rect 13261 11459 13327 11462
rect 15653 11459 15719 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3693 11386 3759 11389
rect 5809 11386 5875 11389
rect 3693 11384 5875 11386
rect 3693 11328 3698 11384
rect 3754 11328 5814 11384
rect 5870 11328 5875 11384
rect 3693 11326 5875 11328
rect 3693 11323 3759 11326
rect 5809 11323 5875 11326
rect 7097 11250 7163 11253
rect 7741 11250 7807 11253
rect 11881 11250 11947 11253
rect 7097 11248 11947 11250
rect 7097 11192 7102 11248
rect 7158 11192 7746 11248
rect 7802 11192 11886 11248
rect 11942 11192 11947 11248
rect 7097 11190 11947 11192
rect 7097 11187 7163 11190
rect 7741 11187 7807 11190
rect 11881 11187 11947 11190
rect 0 10978 480 11008
rect 9765 10978 9831 10981
rect 11605 10978 11671 10981
rect 0 10918 3572 10978
rect 0 10888 480 10918
rect 3512 10706 3572 10918
rect 9765 10976 11671 10978
rect 9765 10920 9770 10976
rect 9826 10920 11610 10976
rect 11666 10920 11671 10976
rect 9765 10918 11671 10920
rect 9765 10915 9831 10918
rect 11605 10915 11671 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 7557 10706 7623 10709
rect 8385 10706 8451 10709
rect 3512 10704 7623 10706
rect 3512 10648 7562 10704
rect 7618 10648 7623 10704
rect 3512 10646 7623 10648
rect 7557 10643 7623 10646
rect 7790 10704 8451 10706
rect 7790 10648 8390 10704
rect 8446 10648 8451 10704
rect 7790 10646 8451 10648
rect 3509 10570 3575 10573
rect 4153 10570 4219 10573
rect 3509 10568 4219 10570
rect 3509 10512 3514 10568
rect 3570 10512 4158 10568
rect 4214 10512 4219 10568
rect 3509 10510 4219 10512
rect 3509 10507 3575 10510
rect 4153 10507 4219 10510
rect 4429 10570 4495 10573
rect 7790 10570 7850 10646
rect 8385 10643 8451 10646
rect 13905 10706 13971 10709
rect 22829 10706 22895 10709
rect 13905 10704 22895 10706
rect 13905 10648 13910 10704
rect 13966 10648 22834 10704
rect 22890 10648 22895 10704
rect 13905 10646 22895 10648
rect 13905 10643 13971 10646
rect 22829 10643 22895 10646
rect 4429 10568 7850 10570
rect 4429 10512 4434 10568
rect 4490 10512 7850 10568
rect 4429 10510 7850 10512
rect 8017 10570 8083 10573
rect 12249 10570 12315 10573
rect 8017 10568 12315 10570
rect 8017 10512 8022 10568
rect 8078 10512 12254 10568
rect 12310 10512 12315 10568
rect 8017 10510 12315 10512
rect 4429 10507 4495 10510
rect 8017 10507 8083 10510
rect 12249 10507 12315 10510
rect 0 10434 480 10464
rect 3693 10434 3759 10437
rect 0 10432 3759 10434
rect 0 10376 3698 10432
rect 3754 10376 3759 10432
rect 0 10374 3759 10376
rect 0 10344 480 10374
rect 3693 10371 3759 10374
rect 3877 10434 3943 10437
rect 6545 10434 6611 10437
rect 3877 10432 6611 10434
rect 3877 10376 3882 10432
rect 3938 10376 6550 10432
rect 6606 10376 6611 10432
rect 3877 10374 6611 10376
rect 3877 10371 3943 10374
rect 6545 10371 6611 10374
rect 7281 10434 7347 10437
rect 9673 10434 9739 10437
rect 7281 10432 9739 10434
rect 7281 10376 7286 10432
rect 7342 10376 9678 10432
rect 9734 10376 9739 10432
rect 7281 10374 9739 10376
rect 7281 10371 7347 10374
rect 9673 10371 9739 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 5349 10298 5415 10301
rect 6269 10298 6335 10301
rect 10041 10298 10107 10301
rect 5349 10296 6194 10298
rect 5349 10240 5354 10296
rect 5410 10240 6194 10296
rect 5349 10238 6194 10240
rect 5349 10235 5415 10238
rect 1761 10162 1827 10165
rect 5625 10162 5691 10165
rect 5993 10162 6059 10165
rect 1761 10160 6059 10162
rect 1761 10104 1766 10160
rect 1822 10104 5630 10160
rect 5686 10104 5998 10160
rect 6054 10104 6059 10160
rect 1761 10102 6059 10104
rect 6134 10162 6194 10238
rect 6269 10296 10107 10298
rect 6269 10240 6274 10296
rect 6330 10240 10046 10296
rect 10102 10240 10107 10296
rect 6269 10238 10107 10240
rect 6269 10235 6335 10238
rect 10041 10235 10107 10238
rect 11697 10298 11763 10301
rect 14457 10298 14523 10301
rect 11697 10296 14523 10298
rect 11697 10240 11702 10296
rect 11758 10240 14462 10296
rect 14518 10240 14523 10296
rect 11697 10238 14523 10240
rect 11697 10235 11763 10238
rect 14457 10235 14523 10238
rect 8201 10162 8267 10165
rect 6134 10160 8267 10162
rect 6134 10104 8206 10160
rect 8262 10104 8267 10160
rect 6134 10102 8267 10104
rect 1761 10099 1827 10102
rect 5625 10099 5691 10102
rect 5993 10099 6059 10102
rect 8201 10099 8267 10102
rect 8753 10162 8819 10165
rect 13813 10162 13879 10165
rect 8753 10160 13879 10162
rect 8753 10104 8758 10160
rect 8814 10104 13818 10160
rect 13874 10104 13879 10160
rect 8753 10102 13879 10104
rect 8753 10099 8819 10102
rect 13813 10099 13879 10102
rect 5165 10026 5231 10029
rect 15285 10026 15351 10029
rect 5165 10024 15351 10026
rect 5165 9968 5170 10024
rect 5226 9968 15290 10024
rect 15346 9968 15351 10024
rect 5165 9966 15351 9968
rect 5165 9963 5231 9966
rect 15285 9963 15351 9966
rect 0 9890 480 9920
rect 3049 9890 3115 9893
rect 0 9888 3115 9890
rect 0 9832 3054 9888
rect 3110 9832 3115 9888
rect 0 9830 3115 9832
rect 0 9800 480 9830
rect 3049 9827 3115 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 2865 9754 2931 9757
rect 5441 9754 5507 9757
rect 2865 9752 5507 9754
rect 2865 9696 2870 9752
rect 2926 9696 5446 9752
rect 5502 9696 5507 9752
rect 2865 9694 5507 9696
rect 2865 9691 2931 9694
rect 5441 9691 5507 9694
rect 10133 9754 10199 9757
rect 13813 9754 13879 9757
rect 10133 9752 13879 9754
rect 10133 9696 10138 9752
rect 10194 9696 13818 9752
rect 13874 9696 13879 9752
rect 10133 9694 13879 9696
rect 10133 9691 10199 9694
rect 13813 9691 13879 9694
rect 2313 9618 2379 9621
rect 3509 9618 3575 9621
rect 2313 9616 3575 9618
rect 2313 9560 2318 9616
rect 2374 9560 3514 9616
rect 3570 9560 3575 9616
rect 2313 9558 3575 9560
rect 2313 9555 2379 9558
rect 3509 9555 3575 9558
rect 6637 9618 6703 9621
rect 10501 9618 10567 9621
rect 6637 9616 10567 9618
rect 6637 9560 6642 9616
rect 6698 9560 10506 9616
rect 10562 9560 10567 9616
rect 6637 9558 10567 9560
rect 6637 9555 6703 9558
rect 10501 9555 10567 9558
rect 3601 9346 3667 9349
rect 7465 9346 7531 9349
rect 9673 9346 9739 9349
rect 3601 9344 5458 9346
rect 3601 9288 3606 9344
rect 3662 9288 5458 9344
rect 3601 9286 5458 9288
rect 3601 9283 3667 9286
rect 0 9210 480 9240
rect 3969 9210 4035 9213
rect 0 9208 4035 9210
rect 0 9152 3974 9208
rect 4030 9152 4035 9208
rect 0 9150 4035 9152
rect 0 9120 480 9150
rect 3969 9147 4035 9150
rect 2221 9074 2287 9077
rect 5257 9074 5323 9077
rect 2221 9072 5323 9074
rect 2221 9016 2226 9072
rect 2282 9016 5262 9072
rect 5318 9016 5323 9072
rect 2221 9014 5323 9016
rect 5398 9074 5458 9286
rect 7465 9344 9739 9346
rect 7465 9288 7470 9344
rect 7526 9288 9678 9344
rect 9734 9288 9739 9344
rect 7465 9286 9739 9288
rect 7465 9283 7531 9286
rect 9673 9283 9739 9286
rect 10685 9346 10751 9349
rect 15469 9346 15535 9349
rect 10685 9344 15535 9346
rect 10685 9288 10690 9344
rect 10746 9288 15474 9344
rect 15530 9288 15535 9344
rect 10685 9286 15535 9288
rect 10685 9283 10751 9286
rect 15469 9283 15535 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 10593 9074 10659 9077
rect 5398 9072 10659 9074
rect 5398 9016 10598 9072
rect 10654 9016 10659 9072
rect 5398 9014 10659 9016
rect 2221 9011 2287 9014
rect 5257 9011 5323 9014
rect 10593 9011 10659 9014
rect 10777 9074 10843 9077
rect 13813 9074 13879 9077
rect 10777 9072 13879 9074
rect 10777 9016 10782 9072
rect 10838 9016 13818 9072
rect 13874 9016 13879 9072
rect 10777 9014 13879 9016
rect 10777 9011 10843 9014
rect 13813 9011 13879 9014
rect 4153 8938 4219 8941
rect 14457 8938 14523 8941
rect 4153 8936 14523 8938
rect 4153 8880 4158 8936
rect 4214 8880 14462 8936
rect 14518 8880 14523 8936
rect 4153 8878 14523 8880
rect 4153 8875 4219 8878
rect 14457 8875 14523 8878
rect 9765 8802 9831 8805
rect 11789 8802 11855 8805
rect 9765 8800 11855 8802
rect 9765 8744 9770 8800
rect 9826 8744 11794 8800
rect 11850 8744 11855 8800
rect 9765 8742 11855 8744
rect 9765 8739 9831 8742
rect 11789 8739 11855 8742
rect 5610 8736 5930 8737
rect 0 8666 480 8696
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 8017 8666 8083 8669
rect 12157 8666 12223 8669
rect 0 8606 3572 8666
rect 0 8576 480 8606
rect 3512 8530 3572 8606
rect 8017 8664 12223 8666
rect 8017 8608 8022 8664
rect 8078 8608 12162 8664
rect 12218 8608 12223 8664
rect 8017 8606 12223 8608
rect 8017 8603 8083 8606
rect 12157 8603 12223 8606
rect 16297 8666 16363 8669
rect 22277 8666 22343 8669
rect 16297 8664 22343 8666
rect 16297 8608 16302 8664
rect 16358 8608 22282 8664
rect 22338 8608 22343 8664
rect 16297 8606 22343 8608
rect 16297 8603 16363 8606
rect 22277 8603 22343 8606
rect 10225 8530 10291 8533
rect 12893 8530 12959 8533
rect 3512 8470 8218 8530
rect 3693 8394 3759 8397
rect 4245 8394 4311 8397
rect 3693 8392 4311 8394
rect 3693 8336 3698 8392
rect 3754 8336 4250 8392
rect 4306 8336 4311 8392
rect 3693 8334 4311 8336
rect 3693 8331 3759 8334
rect 4245 8331 4311 8334
rect 5717 8394 5783 8397
rect 8017 8394 8083 8397
rect 5717 8392 8083 8394
rect 5717 8336 5722 8392
rect 5778 8336 8022 8392
rect 8078 8336 8083 8392
rect 5717 8334 8083 8336
rect 8158 8394 8218 8470
rect 10225 8528 12959 8530
rect 10225 8472 10230 8528
rect 10286 8472 12898 8528
rect 12954 8472 12959 8528
rect 10225 8470 12959 8472
rect 10225 8467 10291 8470
rect 12893 8467 12959 8470
rect 13537 8530 13603 8533
rect 16757 8530 16823 8533
rect 13537 8528 16823 8530
rect 13537 8472 13542 8528
rect 13598 8472 16762 8528
rect 16818 8472 16823 8528
rect 13537 8470 16823 8472
rect 13537 8467 13603 8470
rect 16757 8467 16823 8470
rect 12433 8394 12499 8397
rect 20897 8394 20963 8397
rect 8158 8334 8402 8394
rect 5717 8331 5783 8334
rect 8017 8331 8083 8334
rect 1393 8258 1459 8261
rect 8201 8258 8267 8261
rect 1393 8256 8267 8258
rect 1393 8200 1398 8256
rect 1454 8200 8206 8256
rect 8262 8200 8267 8256
rect 1393 8198 8267 8200
rect 8342 8258 8402 8334
rect 12433 8392 20963 8394
rect 12433 8336 12438 8392
rect 12494 8336 20902 8392
rect 20958 8336 20963 8392
rect 12433 8334 20963 8336
rect 12433 8331 12499 8334
rect 20897 8331 20963 8334
rect 24209 8394 24275 8397
rect 27520 8394 28000 8424
rect 24209 8392 28000 8394
rect 24209 8336 24214 8392
rect 24270 8336 28000 8392
rect 24209 8334 28000 8336
rect 24209 8331 24275 8334
rect 27520 8304 28000 8334
rect 10133 8258 10199 8261
rect 8342 8256 10199 8258
rect 8342 8200 10138 8256
rect 10194 8200 10199 8256
rect 8342 8198 10199 8200
rect 1393 8195 1459 8198
rect 8201 8195 8267 8198
rect 10133 8195 10199 8198
rect 13353 8258 13419 8261
rect 14273 8258 14339 8261
rect 13353 8256 14339 8258
rect 13353 8200 13358 8256
rect 13414 8200 14278 8256
rect 14334 8200 14339 8256
rect 13353 8198 14339 8200
rect 13353 8195 13419 8198
rect 14273 8195 14339 8198
rect 10277 8192 10597 8193
rect 0 8122 480 8152
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 3969 8122 4035 8125
rect 6545 8122 6611 8125
rect 0 8062 1226 8122
rect 0 8032 480 8062
rect 1166 7714 1226 8062
rect 3969 8120 6611 8122
rect 3969 8064 3974 8120
rect 4030 8064 6550 8120
rect 6606 8064 6611 8120
rect 3969 8062 6611 8064
rect 3969 8059 4035 8062
rect 6545 8059 6611 8062
rect 11053 8122 11119 8125
rect 14365 8122 14431 8125
rect 11053 8120 14431 8122
rect 11053 8064 11058 8120
rect 11114 8064 14370 8120
rect 14426 8064 14431 8120
rect 11053 8062 14431 8064
rect 11053 8059 11119 8062
rect 14365 8059 14431 8062
rect 2129 7986 2195 7989
rect 7281 7986 7347 7989
rect 2129 7984 7347 7986
rect 2129 7928 2134 7984
rect 2190 7928 7286 7984
rect 7342 7928 7347 7984
rect 2129 7926 7347 7928
rect 2129 7923 2195 7926
rect 7281 7923 7347 7926
rect 7557 7986 7623 7989
rect 12617 7986 12683 7989
rect 7557 7984 12683 7986
rect 7557 7928 7562 7984
rect 7618 7928 12622 7984
rect 12678 7928 12683 7984
rect 7557 7926 12683 7928
rect 7557 7923 7623 7926
rect 12617 7923 12683 7926
rect 7741 7850 7807 7853
rect 12801 7850 12867 7853
rect 7741 7848 12867 7850
rect 7741 7792 7746 7848
rect 7802 7792 12806 7848
rect 12862 7792 12867 7848
rect 7741 7790 12867 7792
rect 7741 7787 7807 7790
rect 12801 7787 12867 7790
rect 6085 7714 6151 7717
rect 10961 7714 11027 7717
rect 1166 7654 4170 7714
rect 0 7578 480 7608
rect 3877 7578 3943 7581
rect 0 7576 3943 7578
rect 0 7520 3882 7576
rect 3938 7520 3943 7576
rect 0 7518 3943 7520
rect 0 7488 480 7518
rect 3877 7515 3943 7518
rect 4110 7306 4170 7654
rect 6085 7712 11027 7714
rect 6085 7656 6090 7712
rect 6146 7656 10966 7712
rect 11022 7656 11027 7712
rect 6085 7654 11027 7656
rect 6085 7651 6151 7654
rect 10961 7651 11027 7654
rect 15561 7714 15627 7717
rect 19149 7714 19215 7717
rect 15561 7712 19215 7714
rect 15561 7656 15566 7712
rect 15622 7656 19154 7712
rect 19210 7656 19215 7712
rect 15561 7654 19215 7656
rect 15561 7651 15627 7654
rect 19149 7651 19215 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 6177 7578 6243 7581
rect 8385 7578 8451 7581
rect 10685 7578 10751 7581
rect 6177 7576 10751 7578
rect 6177 7520 6182 7576
rect 6238 7520 8390 7576
rect 8446 7520 10690 7576
rect 10746 7520 10751 7576
rect 6177 7518 10751 7520
rect 6177 7515 6243 7518
rect 8385 7515 8451 7518
rect 10685 7515 10751 7518
rect 4337 7442 4403 7445
rect 7925 7442 7991 7445
rect 13353 7442 13419 7445
rect 4337 7440 7991 7442
rect 4337 7384 4342 7440
rect 4398 7384 7930 7440
rect 7986 7384 7991 7440
rect 4337 7382 7991 7384
rect 4337 7379 4403 7382
rect 7925 7379 7991 7382
rect 10550 7440 13419 7442
rect 10550 7384 13358 7440
rect 13414 7384 13419 7440
rect 10550 7382 13419 7384
rect 10550 7306 10610 7382
rect 13353 7379 13419 7382
rect 4110 7246 10610 7306
rect 10777 7306 10843 7309
rect 18045 7306 18111 7309
rect 10777 7304 18111 7306
rect 10777 7248 10782 7304
rect 10838 7248 18050 7304
rect 18106 7248 18111 7304
rect 10777 7246 18111 7248
rect 10777 7243 10843 7246
rect 18045 7243 18111 7246
rect 2497 7170 2563 7173
rect 4521 7170 4587 7173
rect 2497 7168 4587 7170
rect 2497 7112 2502 7168
rect 2558 7112 4526 7168
rect 4582 7112 4587 7168
rect 2497 7110 4587 7112
rect 2497 7107 2563 7110
rect 4521 7107 4587 7110
rect 4705 7170 4771 7173
rect 7281 7170 7347 7173
rect 4705 7168 7347 7170
rect 4705 7112 4710 7168
rect 4766 7112 7286 7168
rect 7342 7112 7347 7168
rect 4705 7110 7347 7112
rect 4705 7107 4771 7110
rect 7281 7107 7347 7110
rect 11053 7170 11119 7173
rect 11513 7170 11579 7173
rect 16297 7170 16363 7173
rect 11053 7168 16363 7170
rect 11053 7112 11058 7168
rect 11114 7112 11518 7168
rect 11574 7112 16302 7168
rect 16358 7112 16363 7168
rect 11053 7110 16363 7112
rect 11053 7107 11119 7110
rect 11513 7107 11579 7110
rect 16297 7107 16363 7110
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 4061 7034 4127 7037
rect 0 7032 4127 7034
rect 0 6976 4066 7032
rect 4122 6976 4127 7032
rect 0 6974 4127 6976
rect 0 6944 480 6974
rect 4061 6971 4127 6974
rect 5717 7034 5783 7037
rect 10041 7034 10107 7037
rect 5717 7032 10107 7034
rect 5717 6976 5722 7032
rect 5778 6976 10046 7032
rect 10102 6976 10107 7032
rect 5717 6974 10107 6976
rect 5717 6971 5783 6974
rect 10041 6971 10107 6974
rect 13721 7034 13787 7037
rect 14733 7034 14799 7037
rect 15745 7034 15811 7037
rect 13721 7032 15811 7034
rect 13721 6976 13726 7032
rect 13782 6976 14738 7032
rect 14794 6976 15750 7032
rect 15806 6976 15811 7032
rect 13721 6974 15811 6976
rect 13721 6971 13787 6974
rect 14733 6971 14799 6974
rect 15745 6971 15811 6974
rect 3049 6898 3115 6901
rect 3509 6898 3575 6901
rect 3049 6896 3575 6898
rect 3049 6840 3054 6896
rect 3110 6840 3514 6896
rect 3570 6840 3575 6896
rect 3049 6838 3575 6840
rect 3049 6835 3115 6838
rect 3509 6835 3575 6838
rect 3877 6898 3943 6901
rect 4797 6898 4863 6901
rect 3877 6896 4863 6898
rect 3877 6840 3882 6896
rect 3938 6840 4802 6896
rect 4858 6840 4863 6896
rect 3877 6838 4863 6840
rect 3877 6835 3943 6838
rect 4797 6835 4863 6838
rect 6177 6898 6243 6901
rect 7465 6898 7531 6901
rect 6177 6896 7531 6898
rect 6177 6840 6182 6896
rect 6238 6840 7470 6896
rect 7526 6840 7531 6896
rect 6177 6838 7531 6840
rect 6177 6835 6243 6838
rect 7465 6835 7531 6838
rect 9489 6898 9555 6901
rect 11513 6898 11579 6901
rect 9489 6896 11579 6898
rect 9489 6840 9494 6896
rect 9550 6840 11518 6896
rect 11574 6840 11579 6896
rect 9489 6838 11579 6840
rect 9489 6835 9555 6838
rect 11513 6835 11579 6838
rect 5993 6762 6059 6765
rect 3926 6760 6059 6762
rect 3926 6704 5998 6760
rect 6054 6704 6059 6760
rect 3926 6702 6059 6704
rect 2865 6626 2931 6629
rect 3926 6626 3986 6702
rect 5993 6699 6059 6702
rect 6269 6762 6335 6765
rect 9857 6762 9923 6765
rect 6269 6760 9923 6762
rect 6269 6704 6274 6760
rect 6330 6704 9862 6760
rect 9918 6704 9923 6760
rect 6269 6702 9923 6704
rect 6269 6699 6335 6702
rect 9857 6699 9923 6702
rect 15377 6762 15443 6765
rect 20897 6762 20963 6765
rect 15377 6760 20963 6762
rect 15377 6704 15382 6760
rect 15438 6704 20902 6760
rect 20958 6704 20963 6760
rect 15377 6702 20963 6704
rect 15377 6699 15443 6702
rect 20897 6699 20963 6702
rect 2865 6624 3986 6626
rect 2865 6568 2870 6624
rect 2926 6568 3986 6624
rect 2865 6566 3986 6568
rect 7557 6626 7623 6629
rect 8569 6626 8635 6629
rect 13997 6626 14063 6629
rect 7557 6624 14063 6626
rect 7557 6568 7562 6624
rect 7618 6568 8574 6624
rect 8630 6568 14002 6624
rect 14058 6568 14063 6624
rect 7557 6566 14063 6568
rect 2865 6563 2931 6566
rect 7557 6563 7623 6566
rect 8569 6563 8635 6566
rect 13997 6563 14063 6566
rect 5610 6560 5930 6561
rect 0 6490 480 6520
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 4613 6490 4679 6493
rect 0 6488 4679 6490
rect 0 6432 4618 6488
rect 4674 6432 4679 6488
rect 0 6430 4679 6432
rect 0 6400 480 6430
rect 4613 6427 4679 6430
rect 1945 6354 2011 6357
rect 4245 6354 4311 6357
rect 1945 6352 4311 6354
rect 1945 6296 1950 6352
rect 2006 6296 4250 6352
rect 4306 6296 4311 6352
rect 1945 6294 4311 6296
rect 1945 6291 2011 6294
rect 4245 6291 4311 6294
rect 14181 6354 14247 6357
rect 20529 6354 20595 6357
rect 14181 6352 20595 6354
rect 14181 6296 14186 6352
rect 14242 6296 20534 6352
rect 20590 6296 20595 6352
rect 14181 6294 20595 6296
rect 14181 6291 14247 6294
rect 20529 6291 20595 6294
rect 6545 6218 6611 6221
rect 17769 6218 17835 6221
rect 6545 6216 17835 6218
rect 6545 6160 6550 6216
rect 6606 6160 17774 6216
rect 17830 6160 17835 6216
rect 6545 6158 17835 6160
rect 6545 6155 6611 6158
rect 17769 6155 17835 6158
rect 6821 6082 6887 6085
rect 10041 6082 10107 6085
rect 6821 6080 10107 6082
rect 6821 6024 6826 6080
rect 6882 6024 10046 6080
rect 10102 6024 10107 6080
rect 6821 6022 10107 6024
rect 6821 6019 6887 6022
rect 10041 6019 10107 6022
rect 10777 6082 10843 6085
rect 15377 6082 15443 6085
rect 10777 6080 15443 6082
rect 10777 6024 10782 6080
rect 10838 6024 15382 6080
rect 15438 6024 15443 6080
rect 10777 6022 15443 6024
rect 10777 6019 10843 6022
rect 15377 6019 15443 6022
rect 10277 6016 10597 6017
rect 0 5946 480 5976
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 1853 5946 1919 5949
rect 0 5944 1919 5946
rect 0 5888 1858 5944
rect 1914 5888 1919 5944
rect 0 5886 1919 5888
rect 0 5856 480 5886
rect 1853 5883 1919 5886
rect 3233 5946 3299 5949
rect 4337 5946 4403 5949
rect 3233 5944 4403 5946
rect 3233 5888 3238 5944
rect 3294 5888 4342 5944
rect 4398 5888 4403 5944
rect 3233 5886 4403 5888
rect 3233 5883 3299 5886
rect 4337 5883 4403 5886
rect 10961 5946 11027 5949
rect 16297 5946 16363 5949
rect 10961 5944 16363 5946
rect 10961 5888 10966 5944
rect 11022 5888 16302 5944
rect 16358 5888 16363 5944
rect 10961 5886 16363 5888
rect 10961 5883 11027 5886
rect 16297 5883 16363 5886
rect 4797 5810 4863 5813
rect 10685 5810 10751 5813
rect 4797 5808 10751 5810
rect 4797 5752 4802 5808
rect 4858 5752 10690 5808
rect 10746 5752 10751 5808
rect 4797 5750 10751 5752
rect 4797 5747 4863 5750
rect 10685 5747 10751 5750
rect 12433 5810 12499 5813
rect 19517 5810 19583 5813
rect 12433 5808 19583 5810
rect 12433 5752 12438 5808
rect 12494 5752 19522 5808
rect 19578 5752 19583 5808
rect 12433 5750 19583 5752
rect 12433 5747 12499 5750
rect 19517 5747 19583 5750
rect 3509 5674 3575 5677
rect 10041 5674 10107 5677
rect 13905 5674 13971 5677
rect 3509 5672 9506 5674
rect 3509 5616 3514 5672
rect 3570 5616 9506 5672
rect 3509 5614 9506 5616
rect 3509 5611 3575 5614
rect 9446 5538 9506 5614
rect 10041 5672 13971 5674
rect 10041 5616 10046 5672
rect 10102 5616 13910 5672
rect 13966 5616 13971 5672
rect 10041 5614 13971 5616
rect 10041 5611 10107 5614
rect 13905 5611 13971 5614
rect 14181 5674 14247 5677
rect 16849 5674 16915 5677
rect 14181 5672 16915 5674
rect 14181 5616 14186 5672
rect 14242 5616 16854 5672
rect 16910 5616 16915 5672
rect 14181 5614 16915 5616
rect 14181 5611 14247 5614
rect 16849 5611 16915 5614
rect 22461 5674 22527 5677
rect 24025 5674 24091 5677
rect 22461 5672 24091 5674
rect 22461 5616 22466 5672
rect 22522 5616 24030 5672
rect 24086 5616 24091 5672
rect 22461 5614 24091 5616
rect 22461 5611 22527 5614
rect 24025 5611 24091 5614
rect 14457 5538 14523 5541
rect 9446 5536 14523 5538
rect 9446 5480 14462 5536
rect 14518 5480 14523 5536
rect 9446 5478 14523 5480
rect 14457 5475 14523 5478
rect 15377 5538 15443 5541
rect 20805 5538 20871 5541
rect 15377 5536 20871 5538
rect 15377 5480 15382 5536
rect 15438 5480 20810 5536
rect 20866 5480 20871 5536
rect 15377 5478 20871 5480
rect 15377 5475 15443 5478
rect 20805 5475 20871 5478
rect 5610 5472 5930 5473
rect 0 5402 480 5432
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 10777 5402 10843 5405
rect 12985 5402 13051 5405
rect 0 5342 3066 5402
rect 0 5312 480 5342
rect 3006 5266 3066 5342
rect 10777 5400 13051 5402
rect 10777 5344 10782 5400
rect 10838 5344 12990 5400
rect 13046 5344 13051 5400
rect 10777 5342 13051 5344
rect 10777 5339 10843 5342
rect 12985 5339 13051 5342
rect 7005 5266 7071 5269
rect 8293 5266 8359 5269
rect 3006 5264 8359 5266
rect 3006 5208 7010 5264
rect 7066 5208 8298 5264
rect 8354 5208 8359 5264
rect 3006 5206 8359 5208
rect 7005 5203 7071 5206
rect 8293 5203 8359 5206
rect 11329 5266 11395 5269
rect 15653 5266 15719 5269
rect 11329 5264 15719 5266
rect 11329 5208 11334 5264
rect 11390 5208 15658 5264
rect 15714 5208 15719 5264
rect 11329 5206 15719 5208
rect 11329 5203 11395 5206
rect 15653 5203 15719 5206
rect 7189 5130 7255 5133
rect 13353 5130 13419 5133
rect 7189 5128 13419 5130
rect 7189 5072 7194 5128
rect 7250 5072 13358 5128
rect 13414 5072 13419 5128
rect 7189 5070 13419 5072
rect 7189 5067 7255 5070
rect 13353 5067 13419 5070
rect 13629 5130 13695 5133
rect 16389 5130 16455 5133
rect 13629 5128 16455 5130
rect 13629 5072 13634 5128
rect 13690 5072 16394 5128
rect 16450 5072 16455 5128
rect 13629 5070 16455 5072
rect 13629 5067 13695 5070
rect 16389 5067 16455 5070
rect 6361 4994 6427 4997
rect 7649 4994 7715 4997
rect 6361 4992 7715 4994
rect 6361 4936 6366 4992
rect 6422 4936 7654 4992
rect 7710 4936 7715 4992
rect 6361 4934 7715 4936
rect 6361 4931 6427 4934
rect 7649 4931 7715 4934
rect 10685 4994 10751 4997
rect 13629 4994 13695 4997
rect 10685 4992 13695 4994
rect 10685 4936 10690 4992
rect 10746 4936 13634 4992
rect 13690 4936 13695 4992
rect 10685 4934 13695 4936
rect 10685 4931 10751 4934
rect 13629 4931 13695 4934
rect 14457 4994 14523 4997
rect 19333 4994 19399 4997
rect 14457 4992 19399 4994
rect 14457 4936 14462 4992
rect 14518 4936 19338 4992
rect 19394 4936 19399 4992
rect 14457 4934 19399 4936
rect 14457 4931 14523 4934
rect 19333 4931 19399 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 2589 4858 2655 4861
rect 3509 4858 3575 4861
rect 7189 4858 7255 4861
rect 2589 4856 7255 4858
rect 2589 4800 2594 4856
rect 2650 4800 3514 4856
rect 3570 4800 7194 4856
rect 7250 4800 7255 4856
rect 2589 4798 7255 4800
rect 2589 4795 2655 4798
rect 3509 4795 3575 4798
rect 7189 4795 7255 4798
rect 13353 4858 13419 4861
rect 15745 4858 15811 4861
rect 13353 4856 15811 4858
rect 13353 4800 13358 4856
rect 13414 4800 15750 4856
rect 15806 4800 15811 4856
rect 13353 4798 15811 4800
rect 13353 4795 13419 4798
rect 15745 4795 15811 4798
rect 0 4722 480 4752
rect 3877 4722 3943 4725
rect 6637 4722 6703 4725
rect 0 4662 3434 4722
rect 0 4632 480 4662
rect 0 4178 480 4208
rect 3049 4178 3115 4181
rect 0 4176 3115 4178
rect 0 4120 3054 4176
rect 3110 4120 3115 4176
rect 0 4118 3115 4120
rect 3374 4178 3434 4662
rect 3877 4720 6703 4722
rect 3877 4664 3882 4720
rect 3938 4664 6642 4720
rect 6698 4664 6703 4720
rect 3877 4662 6703 4664
rect 3877 4659 3943 4662
rect 6637 4659 6703 4662
rect 7833 4722 7899 4725
rect 11881 4722 11947 4725
rect 14089 4722 14155 4725
rect 15653 4722 15719 4725
rect 7833 4720 14155 4722
rect 7833 4664 7838 4720
rect 7894 4664 11886 4720
rect 11942 4664 14094 4720
rect 14150 4664 14155 4720
rect 7833 4662 14155 4664
rect 7833 4659 7899 4662
rect 11881 4659 11947 4662
rect 14089 4659 14155 4662
rect 14598 4720 15719 4722
rect 14598 4664 15658 4720
rect 15714 4664 15719 4720
rect 14598 4662 15719 4664
rect 3785 4586 3851 4589
rect 13261 4586 13327 4589
rect 3785 4584 13327 4586
rect 3785 4528 3790 4584
rect 3846 4528 13266 4584
rect 13322 4528 13327 4584
rect 3785 4526 13327 4528
rect 3785 4523 3851 4526
rect 13261 4523 13327 4526
rect 3601 4450 3667 4453
rect 4153 4450 4219 4453
rect 3601 4448 4219 4450
rect 3601 4392 3606 4448
rect 3662 4392 4158 4448
rect 4214 4392 4219 4448
rect 3601 4390 4219 4392
rect 3601 4387 3667 4390
rect 4153 4387 4219 4390
rect 11237 4450 11303 4453
rect 14598 4450 14658 4662
rect 15653 4659 15719 4662
rect 25313 4586 25379 4589
rect 11237 4448 14658 4450
rect 11237 4392 11242 4448
rect 11298 4392 14658 4448
rect 11237 4390 14658 4392
rect 14782 4584 25379 4586
rect 14782 4528 25318 4584
rect 25374 4528 25379 4584
rect 14782 4526 25379 4528
rect 11237 4387 11303 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 10685 4314 10751 4317
rect 14782 4314 14842 4526
rect 25313 4523 25379 4526
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10685 4312 14842 4314
rect 10685 4256 10690 4312
rect 10746 4256 14842 4312
rect 10685 4254 14842 4256
rect 10685 4251 10751 4254
rect 24669 4178 24735 4181
rect 3374 4176 24735 4178
rect 3374 4120 24674 4176
rect 24730 4120 24735 4176
rect 3374 4118 24735 4120
rect 0 4088 480 4118
rect 3049 4115 3115 4118
rect 24669 4115 24735 4118
rect 7465 4042 7531 4045
rect 10501 4042 10567 4045
rect 11053 4042 11119 4045
rect 7465 4040 11119 4042
rect 7465 3984 7470 4040
rect 7526 3984 10506 4040
rect 10562 3984 11058 4040
rect 11114 3984 11119 4040
rect 7465 3982 11119 3984
rect 7465 3979 7531 3982
rect 10501 3979 10567 3982
rect 11053 3979 11119 3982
rect 18321 4042 18387 4045
rect 20897 4042 20963 4045
rect 18321 4040 20963 4042
rect 18321 3984 18326 4040
rect 18382 3984 20902 4040
rect 20958 3984 20963 4040
rect 18321 3982 20963 3984
rect 18321 3979 18387 3982
rect 20897 3979 20963 3982
rect 21081 4042 21147 4045
rect 22553 4042 22619 4045
rect 21081 4040 22619 4042
rect 21081 3984 21086 4040
rect 21142 3984 22558 4040
rect 22614 3984 22619 4040
rect 21081 3982 22619 3984
rect 21081 3979 21147 3982
rect 22553 3979 22619 3982
rect 2681 3906 2747 3909
rect 5073 3906 5139 3909
rect 2681 3904 5139 3906
rect 2681 3848 2686 3904
rect 2742 3848 5078 3904
rect 5134 3848 5139 3904
rect 2681 3846 5139 3848
rect 2681 3843 2747 3846
rect 5073 3843 5139 3846
rect 10961 3906 11027 3909
rect 17953 3906 18019 3909
rect 10961 3904 18019 3906
rect 10961 3848 10966 3904
rect 11022 3848 17958 3904
rect 18014 3848 18019 3904
rect 10961 3846 18019 3848
rect 10961 3843 11027 3846
rect 17953 3843 18019 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 6269 3770 6335 3773
rect 9949 3770 10015 3773
rect 6269 3768 10015 3770
rect 6269 3712 6274 3768
rect 6330 3712 9954 3768
rect 10010 3712 10015 3768
rect 6269 3710 10015 3712
rect 6269 3707 6335 3710
rect 9949 3707 10015 3710
rect 10777 3770 10843 3773
rect 13353 3770 13419 3773
rect 10777 3768 13419 3770
rect 10777 3712 10782 3768
rect 10838 3712 13358 3768
rect 13414 3712 13419 3768
rect 10777 3710 13419 3712
rect 10777 3707 10843 3710
rect 13353 3707 13419 3710
rect 15285 3770 15351 3773
rect 18689 3770 18755 3773
rect 15285 3768 18755 3770
rect 15285 3712 15290 3768
rect 15346 3712 18694 3768
rect 18750 3712 18755 3768
rect 15285 3710 18755 3712
rect 15285 3707 15351 3710
rect 18689 3707 18755 3710
rect 20069 3770 20135 3773
rect 23933 3770 23999 3773
rect 20069 3768 23999 3770
rect 20069 3712 20074 3768
rect 20130 3712 23938 3768
rect 23994 3712 23999 3768
rect 20069 3710 23999 3712
rect 20069 3707 20135 3710
rect 23933 3707 23999 3710
rect 0 3634 480 3664
rect 2129 3634 2195 3637
rect 0 3632 2195 3634
rect 0 3576 2134 3632
rect 2190 3576 2195 3632
rect 0 3574 2195 3576
rect 0 3544 480 3574
rect 2129 3571 2195 3574
rect 4521 3634 4587 3637
rect 6545 3634 6611 3637
rect 4521 3632 6611 3634
rect 4521 3576 4526 3632
rect 4582 3576 6550 3632
rect 6606 3576 6611 3632
rect 4521 3574 6611 3576
rect 4521 3571 4587 3574
rect 6545 3571 6611 3574
rect 7189 3634 7255 3637
rect 12157 3634 12223 3637
rect 7189 3632 12223 3634
rect 7189 3576 7194 3632
rect 7250 3576 12162 3632
rect 12218 3576 12223 3632
rect 7189 3574 12223 3576
rect 7189 3571 7255 3574
rect 12157 3571 12223 3574
rect 12617 3634 12683 3637
rect 18045 3634 18111 3637
rect 12617 3632 18111 3634
rect 12617 3576 12622 3632
rect 12678 3576 18050 3632
rect 18106 3576 18111 3632
rect 12617 3574 18111 3576
rect 12617 3571 12683 3574
rect 18045 3571 18111 3574
rect 18505 3634 18571 3637
rect 18505 3632 23858 3634
rect 18505 3576 18510 3632
rect 18566 3576 23858 3632
rect 18505 3574 23858 3576
rect 18505 3571 18571 3574
rect 3877 3498 3943 3501
rect 4613 3498 4679 3501
rect 7833 3498 7899 3501
rect 3877 3496 7899 3498
rect 3877 3440 3882 3496
rect 3938 3440 4618 3496
rect 4674 3440 7838 3496
rect 7894 3440 7899 3496
rect 3877 3438 7899 3440
rect 3877 3435 3943 3438
rect 4613 3435 4679 3438
rect 7833 3435 7899 3438
rect 8477 3498 8543 3501
rect 17769 3498 17835 3501
rect 8477 3496 17835 3498
rect 8477 3440 8482 3496
rect 8538 3440 17774 3496
rect 17830 3440 17835 3496
rect 8477 3438 17835 3440
rect 8477 3435 8543 3438
rect 17769 3435 17835 3438
rect 18689 3498 18755 3501
rect 22461 3498 22527 3501
rect 18689 3496 22527 3498
rect 18689 3440 18694 3496
rect 18750 3440 22466 3496
rect 22522 3440 22527 3496
rect 18689 3438 22527 3440
rect 18689 3435 18755 3438
rect 22461 3435 22527 3438
rect 9949 3362 10015 3365
rect 12893 3362 12959 3365
rect 9949 3360 12959 3362
rect 9949 3304 9954 3360
rect 10010 3304 12898 3360
rect 12954 3304 12959 3360
rect 9949 3302 12959 3304
rect 9949 3299 10015 3302
rect 12893 3299 12959 3302
rect 19241 3362 19307 3365
rect 21081 3362 21147 3365
rect 19241 3360 21147 3362
rect 19241 3304 19246 3360
rect 19302 3304 21086 3360
rect 21142 3304 21147 3360
rect 19241 3302 21147 3304
rect 19241 3299 19307 3302
rect 21081 3299 21147 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 3233 3226 3299 3229
rect 17033 3226 17099 3229
rect 1350 3224 3299 3226
rect 1350 3168 3238 3224
rect 3294 3168 3299 3224
rect 1350 3166 3299 3168
rect 0 3090 480 3120
rect 1350 3090 1410 3166
rect 3233 3163 3299 3166
rect 15334 3224 17099 3226
rect 15334 3168 17038 3224
rect 17094 3168 17099 3224
rect 15334 3166 17099 3168
rect 0 3030 1410 3090
rect 1669 3090 1735 3093
rect 8201 3090 8267 3093
rect 9489 3090 9555 3093
rect 1669 3088 9555 3090
rect 1669 3032 1674 3088
rect 1730 3032 8206 3088
rect 8262 3032 9494 3088
rect 9550 3032 9555 3088
rect 1669 3030 9555 3032
rect 0 3000 480 3030
rect 1669 3027 1735 3030
rect 8201 3027 8267 3030
rect 9489 3027 9555 3030
rect 11605 3090 11671 3093
rect 15334 3090 15394 3166
rect 17033 3163 17099 3166
rect 19977 3226 20043 3229
rect 22369 3226 22435 3229
rect 19977 3224 22435 3226
rect 19977 3168 19982 3224
rect 20038 3168 22374 3224
rect 22430 3168 22435 3224
rect 19977 3166 22435 3168
rect 19977 3163 20043 3166
rect 22369 3163 22435 3166
rect 11605 3088 15394 3090
rect 11605 3032 11610 3088
rect 11666 3032 15394 3088
rect 11605 3030 15394 3032
rect 15653 3090 15719 3093
rect 18505 3090 18571 3093
rect 15653 3088 18571 3090
rect 15653 3032 15658 3088
rect 15714 3032 18510 3088
rect 18566 3032 18571 3088
rect 15653 3030 18571 3032
rect 11605 3027 11671 3030
rect 15653 3027 15719 3030
rect 18505 3027 18571 3030
rect 21173 3090 21239 3093
rect 23657 3090 23723 3093
rect 21173 3088 23723 3090
rect 21173 3032 21178 3088
rect 21234 3032 23662 3088
rect 23718 3032 23723 3088
rect 21173 3030 23723 3032
rect 21173 3027 21239 3030
rect 23657 3027 23723 3030
rect 1945 2954 2011 2957
rect 6913 2954 6979 2957
rect 1945 2952 6979 2954
rect 1945 2896 1950 2952
rect 2006 2896 6918 2952
rect 6974 2896 6979 2952
rect 1945 2894 6979 2896
rect 1945 2891 2011 2894
rect 6913 2891 6979 2894
rect 7097 2954 7163 2957
rect 17769 2954 17835 2957
rect 22645 2954 22711 2957
rect 7097 2952 17835 2954
rect 7097 2896 7102 2952
rect 7158 2896 17774 2952
rect 17830 2896 17835 2952
rect 7097 2894 17835 2896
rect 7097 2891 7163 2894
rect 17769 2891 17835 2894
rect 17910 2952 22711 2954
rect 17910 2896 22650 2952
rect 22706 2896 22711 2952
rect 17910 2894 22711 2896
rect 23798 2954 23858 3574
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 24761 3090 24827 3093
rect 27613 3090 27679 3093
rect 24761 3088 27679 3090
rect 24761 3032 24766 3088
rect 24822 3032 27618 3088
rect 27674 3032 27679 3088
rect 24761 3030 27679 3032
rect 24761 3027 24827 3030
rect 27613 3027 27679 3030
rect 27061 2954 27127 2957
rect 23798 2952 27127 2954
rect 23798 2896 27066 2952
rect 27122 2896 27127 2952
rect 23798 2894 27127 2896
rect 3049 2818 3115 2821
rect 7925 2818 7991 2821
rect 3049 2816 7991 2818
rect 3049 2760 3054 2816
rect 3110 2760 7930 2816
rect 7986 2760 7991 2816
rect 3049 2758 7991 2760
rect 3049 2755 3115 2758
rect 7925 2755 7991 2758
rect 12893 2818 12959 2821
rect 15929 2818 15995 2821
rect 12893 2816 15995 2818
rect 12893 2760 12898 2816
rect 12954 2760 15934 2816
rect 15990 2760 15995 2816
rect 12893 2758 15995 2760
rect 12893 2755 12959 2758
rect 15929 2755 15995 2758
rect 17585 2818 17651 2821
rect 17910 2818 17970 2894
rect 22645 2891 22711 2894
rect 27061 2891 27127 2894
rect 17585 2816 17970 2818
rect 17585 2760 17590 2816
rect 17646 2760 17970 2816
rect 17585 2758 17970 2760
rect 22829 2818 22895 2821
rect 27520 2818 28000 2848
rect 22829 2816 28000 2818
rect 22829 2760 22834 2816
rect 22890 2760 28000 2816
rect 22829 2758 28000 2760
rect 17585 2755 17651 2758
rect 22829 2755 22895 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 27520 2728 28000 2758
rect 19610 2687 19930 2688
rect 4889 2682 4955 2685
rect 6913 2682 6979 2685
rect 4889 2680 6979 2682
rect 4889 2624 4894 2680
rect 4950 2624 6918 2680
rect 6974 2624 6979 2680
rect 4889 2622 6979 2624
rect 4889 2619 4955 2622
rect 6913 2619 6979 2622
rect 12065 2682 12131 2685
rect 12433 2682 12499 2685
rect 12065 2680 12499 2682
rect 12065 2624 12070 2680
rect 12126 2624 12438 2680
rect 12494 2624 12499 2680
rect 12065 2622 12499 2624
rect 12065 2619 12131 2622
rect 12433 2619 12499 2622
rect 12709 2682 12775 2685
rect 17677 2682 17743 2685
rect 19333 2682 19399 2685
rect 12709 2680 16314 2682
rect 12709 2624 12714 2680
rect 12770 2624 16314 2680
rect 12709 2622 16314 2624
rect 12709 2619 12775 2622
rect 0 2546 480 2576
rect 3601 2546 3667 2549
rect 6637 2546 6703 2549
rect 0 2544 3667 2546
rect 0 2488 3606 2544
rect 3662 2488 3667 2544
rect 0 2486 3667 2488
rect 0 2456 480 2486
rect 3601 2483 3667 2486
rect 4846 2544 6703 2546
rect 4846 2488 6642 2544
rect 6698 2488 6703 2544
rect 4846 2486 6703 2488
rect 2773 2138 2839 2141
rect 614 2136 2839 2138
rect 614 2080 2778 2136
rect 2834 2080 2839 2136
rect 614 2078 2839 2080
rect 0 2002 480 2032
rect 614 2002 674 2078
rect 2773 2075 2839 2078
rect 0 1942 674 2002
rect 841 2002 907 2005
rect 4846 2002 4906 2486
rect 6637 2483 6703 2486
rect 11697 2546 11763 2549
rect 16021 2546 16087 2549
rect 11697 2544 16087 2546
rect 11697 2488 11702 2544
rect 11758 2488 16026 2544
rect 16082 2488 16087 2544
rect 11697 2486 16087 2488
rect 16254 2546 16314 2622
rect 17677 2680 19399 2682
rect 17677 2624 17682 2680
rect 17738 2624 19338 2680
rect 19394 2624 19399 2680
rect 17677 2622 19399 2624
rect 17677 2619 17743 2622
rect 19333 2619 19399 2622
rect 19793 2546 19859 2549
rect 16254 2544 19859 2546
rect 16254 2488 19798 2544
rect 19854 2488 19859 2544
rect 16254 2486 19859 2488
rect 11697 2483 11763 2486
rect 16021 2483 16087 2486
rect 19793 2483 19859 2486
rect 20529 2546 20595 2549
rect 22461 2546 22527 2549
rect 20529 2544 22527 2546
rect 20529 2488 20534 2544
rect 20590 2488 22466 2544
rect 22522 2488 22527 2544
rect 20529 2486 22527 2488
rect 20529 2483 20595 2486
rect 22461 2483 22527 2486
rect 4981 2410 5047 2413
rect 8661 2410 8727 2413
rect 13537 2410 13603 2413
rect 4981 2408 6194 2410
rect 4981 2352 4986 2408
rect 5042 2352 6194 2408
rect 4981 2350 6194 2352
rect 4981 2347 5047 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 6134 2138 6194 2350
rect 8661 2408 13603 2410
rect 8661 2352 8666 2408
rect 8722 2352 13542 2408
rect 13598 2352 13603 2408
rect 8661 2350 13603 2352
rect 8661 2347 8727 2350
rect 13537 2347 13603 2350
rect 13813 2410 13879 2413
rect 21173 2410 21239 2413
rect 13813 2408 21239 2410
rect 13813 2352 13818 2408
rect 13874 2352 21178 2408
rect 21234 2352 21239 2408
rect 13813 2350 21239 2352
rect 13813 2347 13879 2350
rect 21173 2347 21239 2350
rect 12433 2274 12499 2277
rect 13721 2274 13787 2277
rect 12433 2272 13787 2274
rect 12433 2216 12438 2272
rect 12494 2216 13726 2272
rect 13782 2216 13787 2272
rect 12433 2214 13787 2216
rect 12433 2211 12499 2214
rect 13721 2211 13787 2214
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 6134 2078 14842 2138
rect 841 2000 4906 2002
rect 841 1944 846 2000
rect 902 1944 4906 2000
rect 841 1942 4906 1944
rect 0 1912 480 1942
rect 841 1939 907 1942
rect 14549 1866 14615 1869
rect 6870 1864 14615 1866
rect 6870 1808 14554 1864
rect 14610 1808 14615 1864
rect 6870 1806 14615 1808
rect 14782 1866 14842 2078
rect 18321 1866 18387 1869
rect 14782 1864 18387 1866
rect 14782 1808 18326 1864
rect 18382 1808 18387 1864
rect 14782 1806 18387 1808
rect 3969 1730 4035 1733
rect 6870 1730 6930 1806
rect 14549 1803 14615 1806
rect 18321 1803 18387 1806
rect 3969 1728 6930 1730
rect 3969 1672 3974 1728
rect 4030 1672 6930 1728
rect 3969 1670 6930 1672
rect 7833 1730 7899 1733
rect 13537 1730 13603 1733
rect 7833 1728 13603 1730
rect 7833 1672 7838 1728
rect 7894 1672 13542 1728
rect 13598 1672 13603 1728
rect 7833 1670 13603 1672
rect 3969 1667 4035 1670
rect 7833 1667 7899 1670
rect 13537 1667 13603 1670
rect 13721 1730 13787 1733
rect 18505 1730 18571 1733
rect 13721 1728 18571 1730
rect 13721 1672 13726 1728
rect 13782 1672 18510 1728
rect 18566 1672 18571 1728
rect 13721 1670 18571 1672
rect 13721 1667 13787 1670
rect 18505 1667 18571 1670
rect 2497 1594 2563 1597
rect 7005 1594 7071 1597
rect 15285 1594 15351 1597
rect 2497 1592 15351 1594
rect 2497 1536 2502 1592
rect 2558 1536 7010 1592
rect 7066 1536 15290 1592
rect 15346 1536 15351 1592
rect 2497 1534 15351 1536
rect 2497 1531 2563 1534
rect 7005 1531 7071 1534
rect 15285 1531 15351 1534
rect 0 1458 480 1488
rect 3693 1458 3759 1461
rect 0 1456 3759 1458
rect 0 1400 3698 1456
rect 3754 1400 3759 1456
rect 0 1398 3759 1400
rect 0 1368 480 1398
rect 3693 1395 3759 1398
rect 13537 1458 13603 1461
rect 19609 1458 19675 1461
rect 13537 1456 19675 1458
rect 13537 1400 13542 1456
rect 13598 1400 19614 1456
rect 19670 1400 19675 1456
rect 13537 1398 19675 1400
rect 13537 1395 13603 1398
rect 19609 1395 19675 1398
rect 0 914 480 944
rect 3785 914 3851 917
rect 0 912 3851 914
rect 0 856 3790 912
rect 3846 856 3851 912
rect 0 854 3851 856
rect 0 824 480 854
rect 3785 851 3851 854
rect 0 370 480 400
rect 2957 370 3023 373
rect 0 368 3023 370
rect 0 312 2962 368
rect 3018 312 3023 368
rect 0 310 3023 312
rect 0 280 480 310
rect 2957 307 3023 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1472 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_30
timestamp 1604681595
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1604681595
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4232 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1604681595
transform 1 0 5796 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1604681595
transform 1 0 6164 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_72
timestamp 1604681595
transform 1 0 7728 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1604681595
transform 1 0 7360 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _062_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 1604681595
transform 1 0 8004 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1604681595
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604681595
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8096 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_99
timestamp 1604681595
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_95
timestamp 1604681595
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1604681595
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_112
timestamp 1604681595
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1604681595
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107
timestamp 1604681595
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_116
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 12696 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_130
timestamp 1604681595
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1604681595
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1604681595
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1604681595
transform 1 0 17020 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1604681595
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp 1604681595
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1604681595
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1604681595
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1604681595
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1604681595
transform 1 0 19228 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_207
timestamp 1604681595
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1604681595
transform 1 0 20148 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_211
timestamp 1604681595
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20700 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1604681595
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1604681595
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1604681595
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_224
timestamp 1604681595
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21896 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 22172 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1604681595
transform 1 0 22908 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_233
timestamp 1604681595
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_236
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 22724 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 22448 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1604681595
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_240 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 23276 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_249
timestamp 1604681595
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_253
timestamp 1604681595
transform 1 0 24380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_259
timestamp 1604681595
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_261
timestamp 1604681595
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_265 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_263
timestamp 1604681595
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_275
timestamp 1604681595
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1472 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1604681595
transform 1 0 4324 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_38
timestamp 1604681595
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5336 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_42
timestamp 1604681595
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7820 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_65
timestamp 1604681595
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_69
timestamp 1604681595
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1604681595
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_86
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1604681595
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11224 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_106
timestamp 1604681595
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_133
timestamp 1604681595
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_137
timestamp 1604681595
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15732 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1604681595
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_158
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18216 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1604681595
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_195
timestamp 1604681595
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_199
timestamp 1604681595
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 22172 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_211
timestamp 1604681595
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_221
timestamp 1604681595
transform 1 0 21436 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 23276 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_233
timestamp 1604681595
transform 1 0 22540 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_245
timestamp 1604681595
transform 1 0 23644 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_257
timestamp 1604681595
transform 1 0 24748 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_269
timestamp 1604681595
transform 1 0 25852 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1656 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_19
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1604681595
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_30
timestamp 1604681595
transform 1 0 3864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1604681595
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_48
timestamp 1604681595
transform 1 0 5520 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1604681595
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604681595
transform 1 0 7176 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8188 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1604681595
transform 1 0 7452 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_73
timestamp 1604681595
transform 1 0 7820 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_76
timestamp 1604681595
transform 1 0 8096 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_96
timestamp 1604681595
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_100
timestamp 1604681595
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1604681595
transform 1 0 11500 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14444 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13984 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_136
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp 1604681595
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_164
timestamp 1604681595
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604681595
transform 1 0 16928 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_168
timestamp 1604681595
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_207
timestamp 1604681595
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 21988 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1604681595
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_219
timestamp 1604681595
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_223
timestamp 1604681595
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23920 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_231
timestamp 1604681595
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_235
timestamp 1604681595
transform 1 0 22724 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1604681595
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_250
timestamp 1604681595
transform 1 0 24104 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24288 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_254
timestamp 1604681595
transform 1 0 24472 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_266
timestamp 1604681595
transform 1 0 25576 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_274
timestamp 1604681595
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1472 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4232 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5796 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_43
timestamp 1604681595
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_47
timestamp 1604681595
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_60
timestamp 1604681595
transform 1 0 6624 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7912 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 7636 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_64
timestamp 1604681595
transform 1 0 6992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_67
timestamp 1604681595
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_83
timestamp 1604681595
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1604681595
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 1604681595
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_98
timestamp 1604681595
transform 1 0 10120 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9936 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10304 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10580 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_122
timestamp 1604681595
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13064 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1604681595
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_139
timestamp 1604681595
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_143
timestamp 1604681595
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_147
timestamp 1604681595
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1604681595
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 17020 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_167
timestamp 1604681595
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_171
timestamp 1604681595
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_192
timestamp 1604681595
transform 1 0 18768 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_196
timestamp 1604681595
transform 1 0 19136 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_219
timestamp 1604681595
transform 1 0 21252 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23920 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_4_231
timestamp 1604681595
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_243
timestamp 1604681595
transform 1 0 23460 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_247
timestamp 1604681595
transform 1 0 23828 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_267
timestamp 1604681595
transform 1 0 25668 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1604681595
transform 1 0 1656 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_10
timestamp 1604681595
transform 1 0 2024 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_13
timestamp 1604681595
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_17
timestamp 1604681595
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_38
timestamp 1604681595
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_42
timestamp 1604681595
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_46
timestamp 1604681595
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604681595
transform 1 0 6900 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1604681595
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_70
timestamp 1604681595
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_83
timestamp 1604681595
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9476 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_87
timestamp 1604681595
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1604681595
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13340 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_127
timestamp 1604681595
transform 1 0 12788 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15824 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1604681595
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_173
timestamp 1604681595
transform 1 0 17020 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19780 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_197
timestamp 1604681595
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_201
timestamp 1604681595
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 21068 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_209
timestamp 1604681595
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_213
timestamp 1604681595
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1604681595
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1604681595
transform 1 0 21804 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_237
timestamp 1604681595
transform 1 0 22908 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_243
timestamp 1604681595
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_7
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1564 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_18
timestamp 1604681595
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_14
timestamp 1604681595
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2116 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_20
timestamp 1604681595
transform 1 0 2944 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1604681595
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_28
timestamp 1604681595
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_24
timestamp 1604681595
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3128 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3128 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4600 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_48
timestamp 1604681595
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_56
timestamp 1604681595
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_52
timestamp 1604681595
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_61
timestamp 1604681595
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_57
timestamp 1604681595
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8556 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7084 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_88
timestamp 1604681595
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_100
timestamp 1604681595
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_97
timestamp 1604681595
transform 1 0 10028 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10304 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1604681595
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_108
timestamp 1604681595
transform 1 0 11040 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_113
timestamp 1604681595
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1604681595
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1604681595
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1604681595
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_136
timestamp 1604681595
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_136
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14352 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16284 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1604681595
transform 1 0 14536 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_150
timestamp 1604681595
transform 1 0 14904 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1604681595
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_163
timestamp 1604681595
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_167
timestamp 1604681595
transform 1 0 16468 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_167
timestamp 1604681595
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_173
timestamp 1604681595
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_177
timestamp 1604681595
transform 1 0 17388 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604681595
transform 1 0 19596 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1604681595
transform 1 0 19228 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604681595
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_204
timestamp 1604681595
transform 1 0 19872 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1604681595
transform 1 0 20332 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1604681595
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_219
timestamp 1604681595
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_212
timestamp 1604681595
transform 1 0 20608 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_217
timestamp 1604681595
transform 1 0 21068 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_229
timestamp 1604681595
transform 1 0 22172 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_231
timestamp 1604681595
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_243
timestamp 1604681595
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_241
timestamp 1604681595
transform 1 0 23276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_255
timestamp 1604681595
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_267
timestamp 1604681595
transform 1 0 25668 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1472 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4876 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6440 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5888 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_50
timestamp 1604681595
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_54
timestamp 1604681595
transform 1 0 6072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_77
timestamp 1604681595
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_81
timestamp 1604681595
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1604681595
transform 1 0 8924 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp 1604681595
transform 1 0 9292 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11224 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_107
timestamp 1604681595
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15364 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_164
timestamp 1604681595
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 17756 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_168
timestamp 1604681595
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_172
timestamp 1604681595
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_176
timestamp 1604681595
transform 1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_200
timestamp 1604681595
transform 1 0 19504 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1604681595
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1604681595
transform 1 0 21436 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1604681595
transform 1 0 22540 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_245
timestamp 1604681595
transform 1 0 23644 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_257
timestamp 1604681595
transform 1 0 24748 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_269
timestamp 1604681595
transform 1 0 25852 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2944 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_12
timestamp 1604681595
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_16
timestamp 1604681595
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604681595
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 5428 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_43
timestamp 1604681595
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1604681595
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7636 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_66
timestamp 1604681595
transform 1 0 7176 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 10488 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_90
timestamp 1604681595
transform 1 0 9384 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_94
timestamp 1604681595
transform 1 0 9752 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1604681595
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_101
timestamp 1604681595
transform 1 0 10396 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13340 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_127
timestamp 1604681595
transform 1 0 12788 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_142
timestamp 1604681595
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14904 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_146
timestamp 1604681595
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1604681595
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_173
timestamp 1604681595
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_177
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_190
timestamp 1604681595
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_194
timestamp 1604681595
transform 1 0 18952 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_206
timestamp 1604681595
transform 1 0 20056 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_218
timestamp 1604681595
transform 1 0 21160 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_230
timestamp 1604681595
transform 1 0 22264 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_242
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_6
timestamp 1604681595
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_10
timestamp 1604681595
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4692 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_36
timestamp 1604681595
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_48
timestamp 1604681595
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1604681595
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7820 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1604681595
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_69
timestamp 1604681595
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1604681595
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_86
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_104
timestamp 1604681595
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11408 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11224 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_108
timestamp 1604681595
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1604681595
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_131
timestamp 1604681595
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_135
timestamp 1604681595
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_139
timestamp 1604681595
transform 1 0 13892 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1604681595
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_173
timestamp 1604681595
transform 1 0 17020 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_185
timestamp 1604681595
transform 1 0 18124 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1604681595
transform 1 0 19228 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1604681595
transform 1 0 20332 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2760 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_9
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_13
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_37
timestamp 1604681595
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1604681595
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_45
timestamp 1604681595
transform 1 0 5244 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 5704 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8648 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1604681595
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1604681595
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1604681595
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_105
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604681595
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14444 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_136
timestamp 1604681595
transform 1 0 13616 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_141
timestamp 1604681595
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16008 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1604681595
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_158
timestamp 1604681595
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_168
timestamp 1604681595
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1604681595
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_176
timestamp 1604681595
transform 1 0 17296 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1604681595
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_214
timestamp 1604681595
transform 1 0 20792 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1604681595
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1604681595
transform 1 0 21804 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_237
timestamp 1604681595
transform 1 0 22908 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1604681595
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1840 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_17
timestamp 1604681595
transform 1 0 2668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_21
timestamp 1604681595
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_25
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5796 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_45
timestamp 1604681595
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 8280 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_70
timestamp 1604681595
transform 1 0 7544 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_76
timestamp 1604681595
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_81
timestamp 1604681595
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10212 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1604681595
transform 1 0 8924 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1604681595
transform 1 0 9292 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1604681595
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11776 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_108
timestamp 1604681595
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_112
timestamp 1604681595
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_135
timestamp 1604681595
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_139
timestamp 1604681595
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_143
timestamp 1604681595
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15364 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_147
timestamp 1604681595
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_174
timestamp 1604681595
transform 1 0 17112 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_186
timestamp 1604681595
transform 1 0 18216 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_198
timestamp 1604681595
transform 1 0 19320 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1604681595
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2208 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_26
timestamp 1604681595
transform 1 0 3496 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1604681595
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_25
timestamp 1604681595
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_21
timestamp 1604681595
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 3772 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_45
timestamp 1604681595
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_52
timestamp 1604681595
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_48
timestamp 1604681595
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5612 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_62
timestamp 1604681595
transform 1 0 6808 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1604681595
transform 1 0 6440 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_69
timestamp 1604681595
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_65
timestamp 1604681595
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_73
timestamp 1604681595
transform 1 0 7820 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1604681595
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7912 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_83
timestamp 1604681595
transform 1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1604681595
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_85
timestamp 1604681595
transform 1 0 8924 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9476 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_100
timestamp 1604681595
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_104
timestamp 1604681595
transform 1 0 10672 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_106
timestamp 1604681595
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_108
timestamp 1604681595
transform 1 0 11040 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1604681595
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_119
timestamp 1604681595
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_142
timestamp 1604681595
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_153
timestamp 1604681595
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_146
timestamp 1604681595
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604681595
transform 1 0 14904 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_157
timestamp 1604681595
transform 1 0 15548 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_157
timestamp 1604681595
transform 1 0 15548 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1604681595
transform 1 0 16652 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_169
timestamp 1604681595
transform 1 0 16652 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_181
timestamp 1604681595
transform 1 0 17756 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_193
timestamp 1604681595
transform 1 0 18860 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_205
timestamp 1604681595
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4232 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_26
timestamp 1604681595
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1604681595
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_43
timestamp 1604681595
transform 1 0 5060 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_47
timestamp 1604681595
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8464 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_72
timestamp 1604681595
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_76
timestamp 1604681595
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1604681595
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_103
timestamp 1604681595
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 10948 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13156 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_129
timestamp 1604681595
transform 1 0 12972 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_151
timestamp 1604681595
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_163
timestamp 1604681595
transform 1 0 16100 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_232
timestamp 1604681595
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_6
timestamp 1604681595
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_10
timestamp 1604681595
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_45
timestamp 1604681595
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_53
timestamp 1604681595
transform 1 0 5980 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_57
timestamp 1604681595
transform 1 0 6348 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1604681595
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7084 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_16_64
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_88
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_102
timestamp 1604681595
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_106
timestamp 1604681595
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_119
timestamp 1604681595
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_123
timestamp 1604681595
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 13984 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_136
timestamp 1604681595
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1604681595
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_147
timestamp 1604681595
transform 1 0 14628 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_158
timestamp 1604681595
transform 1 0 15640 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_162
timestamp 1604681595
transform 1 0 16008 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_174
timestamp 1604681595
transform 1 0 17112 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_186
timestamp 1604681595
transform 1 0 18216 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_198
timestamp 1604681595
transform 1 0 19320 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1604681595
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1564 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_14
timestamp 1604681595
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_18
timestamp 1604681595
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3772 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_22
timestamp 1604681595
transform 1 0 3128 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_26
timestamp 1604681595
transform 1 0 3496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_38
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_50
timestamp 1604681595
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_42
timestamp 1604681595
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 5336 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1604681595
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1604681595
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9660 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 9384 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_85
timestamp 1604681595
transform 1 0 8924 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_112
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12696 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1604681595
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15180 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_149
timestamp 1604681595
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1604681595
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_170
timestamp 1604681595
transform 1 0 16744 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1604681595
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_228
timestamp 1604681595
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_232
timestamp 1604681595
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1472 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4600 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_36
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_57
timestamp 1604681595
transform 1 0 6348 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_61
timestamp 1604681595
transform 1 0 6716 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7084 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 8648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_64
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_74
timestamp 1604681595
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_78
timestamp 1604681595
transform 1 0 8280 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10304 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1604681595
transform 1 0 8924 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1604681595
transform 1 0 9292 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_97
timestamp 1604681595
transform 1 0 10028 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_119
timestamp 1604681595
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_123
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_136
timestamp 1604681595
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_140
timestamp 1604681595
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_144
timestamp 1604681595
transform 1 0 14352 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1604681595
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_175
timestamp 1604681595
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_187
timestamp 1604681595
transform 1 0 18308 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_199
timestamp 1604681595
transform 1 0 19412 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_211
timestamp 1604681595
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_227
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 22264 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_234
timestamp 1604681595
transform 1 0 22632 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_246
timestamp 1604681595
transform 1 0 23736 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_258
timestamp 1604681595
transform 1 0 24840 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_270
timestamp 1604681595
transform 1 0 25944 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1604681595
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1472 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1604681595
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_21
timestamp 1604681595
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_36
timestamp 1604681595
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3404 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_19_48
timestamp 1604681595
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_44
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_59
timestamp 1604681595
transform 1 0 6532 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_52
timestamp 1604681595
transform 1 0 5888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_64
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_76
timestamp 1604681595
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_82
timestamp 1604681595
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_75
timestamp 1604681595
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9384 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_103
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_99
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10028 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_19_107
timestamp 1604681595
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_116
timestamp 1604681595
transform 1 0 11776 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_122
timestamp 1604681595
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13340 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13340 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_129
timestamp 1604681595
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_142
timestamp 1604681595
transform 1 0 14168 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1604681595
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_156
timestamp 1604681595
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_160
timestamp 1604681595
transform 1 0 15824 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1604681595
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_172
timestamp 1604681595
transform 1 0 16928 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1604681595
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_173
timestamp 1604681595
transform 1 0 17020 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_185
timestamp 1604681595
transform 1 0 18124 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1604681595
transform 1 0 19228 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1604681595
transform 1 0 20332 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 23368 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_232
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_249
timestamp 1604681595
transform 1 0 24012 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_239
timestamp 1604681595
transform 1 0 23092 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_246
timestamp 1604681595
transform 1 0 23736 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 24196 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_253
timestamp 1604681595
transform 1 0 24380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_265
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_258
timestamp 1604681595
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_270
timestamp 1604681595
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_274
timestamp 1604681595
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 1840 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_17
timestamp 1604681595
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_21
timestamp 1604681595
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_25
timestamp 1604681595
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_29
timestamp 1604681595
transform 1 0 3772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_43
timestamp 1604681595
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_47
timestamp 1604681595
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_55
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_66
timestamp 1604681595
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_70
timestamp 1604681595
transform 1 0 7544 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9476 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_87
timestamp 1604681595
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_100
timestamp 1604681595
transform 1 0 10304 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_104
timestamp 1604681595
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 11040 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_111
timestamp 1604681595
transform 1 0 11316 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_115
timestamp 1604681595
transform 1 0 11684 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 13984 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_143
timestamp 1604681595
transform 1 0 14260 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_155
timestamp 1604681595
transform 1 0 15364 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_167
timestamp 1604681595
transform 1 0 16468 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 24012 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 24564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_253
timestamp 1604681595
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1604681595
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1472 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_13
timestamp 1604681595
transform 1 0 2300 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_17
timestamp 1604681595
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_25
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_21
timestamp 1604681595
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_40
timestamp 1604681595
transform 1 0 4784 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_36
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4876 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6716 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_50
timestamp 1604681595
transform 1 0 5704 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_54
timestamp 1604681595
transform 1 0 6072 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_57
timestamp 1604681595
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9752 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1604681595
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_113
timestamp 1604681595
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_117
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_121
timestamp 1604681595
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_142
timestamp 1604681595
transform 1 0 14168 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_150
timestamp 1604681595
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604681595
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2668 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_9
timestamp 1604681595
transform 1 0 1932 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_13
timestamp 1604681595
transform 1 0 2300 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_16
timestamp 1604681595
transform 1 0 2576 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_26
timestamp 1604681595
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_30
timestamp 1604681595
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_81
timestamp 1604681595
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9292 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_85
timestamp 1604681595
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_108
timestamp 1604681595
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_112
timestamp 1604681595
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_116
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_142
timestamp 1604681595
transform 1 0 14168 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1604681595
transform 1 0 15272 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_166
timestamp 1604681595
transform 1 0 16376 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1604681595
transform 1 0 17480 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1604681595
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_6
timestamp 1604681595
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_10
timestamp 1604681595
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6808 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_51
timestamp 1604681595
transform 1 0 5796 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_60
timestamp 1604681595
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_74
timestamp 1604681595
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_78
timestamp 1604681595
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_82
timestamp 1604681595
transform 1 0 8648 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9292 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1604681595
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1604681595
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11592 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_113
timestamp 1604681595
transform 1 0 11500 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_127
timestamp 1604681595
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_131
timestamp 1604681595
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_143
timestamp 1604681595
transform 1 0 14260 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604681595
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2668 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_9
timestamp 1604681595
transform 1 0 1932 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_13
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_16
timestamp 1604681595
transform 1 0 2576 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_36
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_50
timestamp 1604681595
transform 1 0 5704 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_56
timestamp 1604681595
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1604681595
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1604681595
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_75
timestamp 1604681595
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1604681595
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_83
timestamp 1604681595
transform 1 0 8740 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9200 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_107
timestamp 1604681595
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_111
timestamp 1604681595
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1604681595
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_119
timestamp 1604681595
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_126
timestamp 1604681595
transform 1 0 12696 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_138
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_150
timestamp 1604681595
transform 1 0 14904 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_162
timestamp 1604681595
transform 1 0 16008 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_174
timestamp 1604681595
transform 1 0 17112 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1604681595
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_6
timestamp 1604681595
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1656 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_19
timestamp 1604681595
transform 1 0 2852 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_10
timestamp 1604681595
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3312 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_45
timestamp 1604681595
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_43
timestamp 1604681595
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_49
timestamp 1604681595
transform 1 0 5612 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_47
timestamp 1604681595
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1604681595
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_53
timestamp 1604681595
transform 1 0 5980 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_67
timestamp 1604681595
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_71
timestamp 1604681595
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1604681595
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1604681595
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_88
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9292 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_104
timestamp 1604681595
transform 1 0 10672 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_100
timestamp 1604681595
transform 1 0 10304 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_96
timestamp 1604681595
transform 1 0 9936 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10120 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9292 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_108
timestamp 1604681595
transform 1 0 11040 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_108
timestamp 1604681595
transform 1 0 11040 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11132 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_117
timestamp 1604681595
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_122
timestamp 1604681595
transform 1 0 12328 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_118
timestamp 1604681595
transform 1 0 11960 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_125
timestamp 1604681595
transform 1 0 12604 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_26_137
timestamp 1604681595
transform 1 0 13708 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_142
timestamp 1604681595
transform 1 0 14168 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_154
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_166
timestamp 1604681595
transform 1 0 16376 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1604681595
transform 1 0 17480 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1604681595
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604681595
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 2852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_16
timestamp 1604681595
transform 1 0 2576 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4416 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_21
timestamp 1604681595
transform 1 0 3036 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_25
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_45
timestamp 1604681595
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_49
timestamp 1604681595
transform 1 0 5612 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_53
timestamp 1604681595
transform 1 0 5980 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_75
timestamp 1604681595
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9292 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_87
timestamp 1604681595
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1604681595
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11316 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_28_106
timestamp 1604681595
transform 1 0 10856 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_110
timestamp 1604681595
transform 1 0 11224 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_130
timestamp 1604681595
transform 1 0 13064 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_142
timestamp 1604681595
transform 1 0 14168 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_150
timestamp 1604681595
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2760 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_10
timestamp 1604681595
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_14
timestamp 1604681595
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4232 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_24
timestamp 1604681595
transform 1 0 3312 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_30
timestamp 1604681595
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_67
timestamp 1604681595
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_80
timestamp 1604681595
transform 1 0 8464 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9200 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_107
timestamp 1604681595
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_111
timestamp 1604681595
transform 1 0 11316 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_115
timestamp 1604681595
transform 1 0 11684 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_132
timestamp 1604681595
transform 1 0 13248 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_144
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_156
timestamp 1604681595
transform 1 0 15456 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_168
timestamp 1604681595
transform 1 0 16560 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1604681595
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 2852 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2300 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1604681595
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_40
timestamp 1604681595
transform 1 0 4784 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5336 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_65
timestamp 1604681595
transform 1 0 7084 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_73
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10396 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_84
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_120
timestamp 1604681595
transform 1 0 12144 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_125
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_137
timestamp 1604681595
transform 1 0 13708 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1840 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_14
timestamp 1604681595
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_18
timestamp 1604681595
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 4416 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 3128 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_28
timestamp 1604681595
transform 1 0 3680 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_34
timestamp 1604681595
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_40
timestamp 1604681595
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 5704 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_44
timestamp 1604681595
transform 1 0 5152 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_75
timestamp 1604681595
transform 1 0 8004 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_87
timestamp 1604681595
transform 1 0 9108 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_99
timestamp 1604681595
transform 1 0 10212 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 10948 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 2852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_11
timestamp 1604681595
transform 1 0 2116 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_36
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_47
timestamp 1604681595
transform 1 0 5428 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_59
timestamp 1604681595
transform 1 0 6532 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7636 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_64
timestamp 1604681595
transform 1 0 6992 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_70
timestamp 1604681595
transform 1 0 7544 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_77
timestamp 1604681595
transform 1 0 8188 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_89
timestamp 1604681595
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 1564 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_17
timestamp 1604681595
transform 1 0 2668 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 1604681595
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_13
timestamp 1604681595
transform 1 0 2300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_25
timestamp 1604681595
transform 1 0 3404 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_29
timestamp 1604681595
transform 1 0 3772 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_25
timestamp 1604681595
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 3036 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_37
timestamp 1604681595
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 4140 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_41
timestamp 1604681595
transform 1 0 4876 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_53
timestamp 1604681595
transform 1 0 5980 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7912 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_76
timestamp 1604681595
transform 1 0 8096 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_80
timestamp 1604681595
transform 1 0 8464 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_87
timestamp 1604681595
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_91
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_103
timestamp 1604681595
transform 1 0 10580 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_115
timestamp 1604681595
transform 1 0 11684 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1604681595
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_7
timestamp 1604681595
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_11
timestamp 1604681595
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_19
timestamp 1604681595
transform 1 0 2852 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 3036 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_23
timestamp 1604681595
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_35
timestamp 1604681595
transform 1 0 4324 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_47
timestamp 1604681595
transform 1 0 5428 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 8372 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7084 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_71
timestamp 1604681595
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1604681595
transform 1 0 8004 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_83
timestamp 1604681595
transform 1 0 8740 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 8924 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_87
timestamp 1604681595
transform 1 0 9108 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_99
timestamp 1604681595
transform 1 0 10212 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_111
timestamp 1604681595
transform 1 0 11316 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_119
timestamp 1604681595
transform 1 0 12052 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1604681595
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1604681595
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1604681595
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1604681595
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_7
timestamp 1604681595
transform 1 0 1748 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_19
timestamp 1604681595
transform 1 0 2852 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1604681595
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1604681595
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1604681595
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1604681595
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1604681595
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1604681595
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1604681595
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_13
timestamp 1604681595
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_17
timestamp 1604681595
transform 1 0 2668 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 3036 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_25
timestamp 1604681595
transform 1 0 3404 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_29
timestamp 1604681595
transform 1 0 3772 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_41
timestamp 1604681595
transform 1 0 4876 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_53
timestamp 1604681595
transform 1 0 5980 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604681595
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12604 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_110
timestamp 1604681595
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_127
timestamp 1604681595
transform 1 0 12788 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_139
timestamp 1604681595
transform 1 0 13892 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1604681595
transform 1 0 14996 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_163
timestamp 1604681595
transform 1 0 16100 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_175
timestamp 1604681595
transform 1 0 17204 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1604681595
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1604681595
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1604681595
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604681595
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_13
timestamp 1604681595
transform 1 0 2300 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_25
timestamp 1604681595
transform 1 0 3404 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_117
timestamp 1604681595
transform 1 0 11868 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1604681595
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1604681595
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1604681595
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1604681595
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1604681595
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1604681595
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1604681595
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1604681595
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_251
timestamp 1604681595
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1604681595
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_7
timestamp 1604681595
transform 1 0 1748 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 1564 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1604681595
transform 1 0 2116 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_17
timestamp 1604681595
transform 1 0 2668 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_13
timestamp 1604681595
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_19
timestamp 1604681595
transform 1 0 2852 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 3036 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_25
timestamp 1604681595
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_29
timestamp 1604681595
transform 1 0 3772 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_41
timestamp 1604681595
transform 1 0 4876 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_53
timestamp 1604681595
transform 1 0 5980 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604681595
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1604681595
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1604681595
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1604681595
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604681595
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_220
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1604681595
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_232
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1604681595
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_253
timestamp 1604681595
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_259
timestamp 1604681595
transform 1 0 24932 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1604681595
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1604681595
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_271
timestamp 1604681595
transform 1 0 26036 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1604681595
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_11
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_23
timestamp 1604681595
transform 1 0 3220 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_35
timestamp 1604681595
transform 1 0 4324 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_47
timestamp 1604681595
transform 1 0 5428 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1604681595
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_7
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_19
timestamp 1604681595
transform 1 0 2852 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 27520 19456 28000 19576 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 27618 0 27674 480 6 SC_IN_TOP
port 1 nsew default input
rlabel metal3 s 27520 25032 28000 25152 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal3 s 0 27616 480 27736 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_42_
port 4 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_43_
port 5 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_44_
port 6 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_45_
port 7 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_46_
port 8 nsew default input
rlabel metal2 s 3054 0 3110 480 6 bottom_left_grid_pin_47_
port 9 nsew default input
rlabel metal2 s 3606 0 3662 480 6 bottom_left_grid_pin_48_
port 10 nsew default input
rlabel metal2 s 4158 0 4214 480 6 bottom_left_grid_pin_49_
port 11 nsew default input
rlabel metal2 s 27066 0 27122 480 6 bottom_right_grid_pin_1_
port 12 nsew default input
rlabel metal3 s 27520 8304 28000 8424 6 ccff_head
port 13 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 ccff_tail
port 14 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[10]
port 16 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[11]
port 17 nsew default input
rlabel metal3 s 0 11432 480 11552 6 chanx_left_in[12]
port 18 nsew default input
rlabel metal3 s 0 11976 480 12096 6 chanx_left_in[13]
port 19 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[14]
port 20 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[15]
port 21 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[16]
port 22 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[17]
port 23 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[18]
port 24 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[19]
port 25 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[1]
port 26 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[2]
port 27 nsew default input
rlabel metal3 s 0 6400 480 6520 6 chanx_left_in[3]
port 28 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[4]
port 29 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[5]
port 30 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[6]
port 31 nsew default input
rlabel metal3 s 0 8576 480 8696 6 chanx_left_in[7]
port 32 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[8]
port 33 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_left_in[9]
port 34 nsew default input
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[0]
port 35 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[10]
port 36 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[11]
port 37 nsew default tristate
rlabel metal3 s 0 22584 480 22704 6 chanx_left_out[12]
port 38 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[13]
port 39 nsew default tristate
rlabel metal3 s 0 23808 480 23928 6 chanx_left_out[14]
port 40 nsew default tristate
rlabel metal3 s 0 24352 480 24472 6 chanx_left_out[15]
port 41 nsew default tristate
rlabel metal3 s 0 24896 480 25016 6 chanx_left_out[16]
port 42 nsew default tristate
rlabel metal3 s 0 25440 480 25560 6 chanx_left_out[17]
port 43 nsew default tristate
rlabel metal3 s 0 25984 480 26104 6 chanx_left_out[18]
port 44 nsew default tristate
rlabel metal3 s 0 26528 480 26648 6 chanx_left_out[19]
port 45 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[1]
port 46 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chanx_left_out[2]
port 47 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 chanx_left_out[3]
port 48 nsew default tristate
rlabel metal3 s 0 18096 480 18216 6 chanx_left_out[4]
port 49 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_left_out[5]
port 50 nsew default tristate
rlabel metal3 s 0 19320 480 19440 6 chanx_left_out[6]
port 51 nsew default tristate
rlabel metal3 s 0 19864 480 19984 6 chanx_left_out[7]
port 52 nsew default tristate
rlabel metal3 s 0 20408 480 20528 6 chanx_left_out[8]
port 53 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 chanx_left_out[9]
port 54 nsew default tristate
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_in[0]
port 55 nsew default input
rlabel metal2 s 10322 0 10378 480 6 chany_bottom_in[10]
port 56 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[11]
port 57 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_bottom_in[12]
port 58 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[13]
port 59 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[14]
port 60 nsew default input
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_in[15]
port 61 nsew default input
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_in[16]
port 62 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_in[17]
port 63 nsew default input
rlabel metal2 s 14830 0 14886 480 6 chany_bottom_in[18]
port 64 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[19]
port 65 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[1]
port 66 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[2]
port 67 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[3]
port 68 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[4]
port 69 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[5]
port 70 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[6]
port 71 nsew default input
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[7]
port 72 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[8]
port 73 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[9]
port 74 nsew default input
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[0]
port 75 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[10]
port 76 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[11]
port 77 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[12]
port 78 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[13]
port 79 nsew default tristate
rlabel metal2 s 23754 0 23810 480 6 chany_bottom_out[14]
port 80 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[15]
port 81 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[16]
port 82 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[17]
port 83 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[18]
port 84 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[19]
port 85 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[1]
port 86 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[2]
port 87 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 chany_bottom_out[3]
port 88 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 chany_bottom_out[4]
port 89 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_bottom_out[5]
port 90 nsew default tristate
rlabel metal2 s 19246 0 19302 480 6 chany_bottom_out[6]
port 91 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[7]
port 92 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 chany_bottom_out[8]
port 93 nsew default tristate
rlabel metal2 s 20902 0 20958 480 6 chany_bottom_out[9]
port 94 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_34_
port 95 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_35_
port 96 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_36_
port 97 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_37_
port 98 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_38_
port 99 nsew default input
rlabel metal3 s 0 3000 480 3120 6 left_bottom_grid_pin_39_
port 100 nsew default input
rlabel metal3 s 0 3544 480 3664 6 left_bottom_grid_pin_40_
port 101 nsew default input
rlabel metal3 s 0 4088 480 4208 6 left_bottom_grid_pin_41_
port 102 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_top_grid_pin_1_
port 103 nsew default input
rlabel metal3 s 27520 2728 28000 2848 6 prog_clk
port 104 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 105 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 106 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 27736
<< end >>
