VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__3_
  CLASS BLOCK ;
  FOREIGN sb_0__3_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 138.070 BY 137.320 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.760 0.000 72.040 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.900 0.000 76.180 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.580 0.000 79.860 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.720 0.000 84.000 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.860 0.000 88.140 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.540 0.000 91.820 2.400 ;
    END
  END address[5]
  PIN bottom_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.780 0.000 20.060 2.400 ;
    END
  END bottom_left_grid_pin_11_
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.920 0.000 24.200 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.600 0.000 27.880 2.400 ;
    END
  END bottom_left_grid_pin_15_
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.000 0.280 2.400 ;
    END
  END bottom_left_grid_pin_1_
  PIN bottom_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.680 0.000 3.960 2.400 ;
    END
  END bottom_left_grid_pin_3_
  PIN bottom_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.820 0.000 8.100 2.400 ;
    END
  END bottom_left_grid_pin_5_
  PIN bottom_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.960 0.000 12.240 2.400 ;
    END
  END bottom_left_grid_pin_7_
  PIN bottom_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.640 0.000 15.920 2.400 ;
    END
  END bottom_left_grid_pin_9_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.700 0.000 135.980 2.400 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 2.080 138.070 2.680 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 6.840 138.070 7.440 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 12.280 138.070 12.880 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 17.040 138.070 17.640 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 22.480 138.070 23.080 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 27.920 138.070 28.520 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 32.680 138.070 33.280 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 38.120 138.070 38.720 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 43.560 138.070 44.160 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 95.240 138.070 95.840 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 100.000 138.070 100.600 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 105.440 138.070 106.040 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 110.880 138.070 111.480 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 115.640 138.070 116.240 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 121.080 138.070 121.680 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 126.520 138.070 127.120 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 131.280 138.070 131.880 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 136.720 138.070 137.320 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.740 0.000 32.020 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.880 0.000 36.160 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.560 0.000 39.840 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.700 0.000 43.980 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.840 0.000 48.120 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.520 0.000 51.800 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.660 0.000 55.940 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.800 0.000 60.080 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.480 0.000 63.760 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.820 0.000 100.100 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.500 0.000 103.780 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.640 0.000 107.920 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.780 0.000 112.060 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.460 0.000 115.740 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.600 0.000 119.880 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.740 0.000 124.020 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.420 0.000 127.700 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.560 0.000 131.840 2.400 ;
    END
  END chany_bottom_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.680 0.000 95.960 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.620 0.000 67.900 2.400 ;
    END
  END enable
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 89.800 138.070 90.400 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 74.160 138.070 74.760 ;
    END
  END right_top_grid_pin_11_
  PIN right_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 79.600 138.070 80.200 ;
    END
  END right_top_grid_pin_13_
  PIN right_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 85.040 138.070 85.640 ;
    END
  END right_top_grid_pin_15_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 48.320 138.070 48.920 ;
    END
  END right_top_grid_pin_1_
  PIN right_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 53.760 138.070 54.360 ;
    END
  END right_top_grid_pin_3_
  PIN right_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 58.520 138.070 59.120 ;
    END
  END right_top_grid_pin_5_
  PIN right_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 63.960 138.070 64.560 ;
    END
  END right_top_grid_pin_7_
  PIN right_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 69.400 138.070 70.000 ;
    END
  END right_top_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 26.125 10.640 27.725 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 49.455 10.640 51.055 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 3.590 10.795 132.390 127.925 ;
      LAYER met1 ;
        RECT 1.360 0.040 136.460 128.080 ;
      LAYER met2 ;
        RECT 0.280 2.680 136.440 134.485 ;
        RECT 0.560 0.010 3.400 2.680 ;
        RECT 4.240 0.010 7.540 2.680 ;
        RECT 8.380 0.010 11.680 2.680 ;
        RECT 12.520 0.010 15.360 2.680 ;
        RECT 16.200 0.010 19.500 2.680 ;
        RECT 20.340 0.010 23.640 2.680 ;
        RECT 24.480 0.010 27.320 2.680 ;
        RECT 28.160 0.010 31.460 2.680 ;
        RECT 32.300 0.010 35.600 2.680 ;
        RECT 36.440 0.010 39.280 2.680 ;
        RECT 40.120 0.010 43.420 2.680 ;
        RECT 44.260 0.010 47.560 2.680 ;
        RECT 48.400 0.010 51.240 2.680 ;
        RECT 52.080 0.010 55.380 2.680 ;
        RECT 56.220 0.010 59.520 2.680 ;
        RECT 60.360 0.010 63.200 2.680 ;
        RECT 64.040 0.010 67.340 2.680 ;
        RECT 68.180 0.010 71.480 2.680 ;
        RECT 72.320 0.010 75.620 2.680 ;
        RECT 76.460 0.010 79.300 2.680 ;
        RECT 80.140 0.010 83.440 2.680 ;
        RECT 84.280 0.010 87.580 2.680 ;
        RECT 88.420 0.010 91.260 2.680 ;
        RECT 92.100 0.010 95.400 2.680 ;
        RECT 96.240 0.010 99.540 2.680 ;
        RECT 100.380 0.010 103.220 2.680 ;
        RECT 104.060 0.010 107.360 2.680 ;
        RECT 108.200 0.010 111.500 2.680 ;
        RECT 112.340 0.010 115.180 2.680 ;
        RECT 116.020 0.010 119.320 2.680 ;
        RECT 120.160 0.010 123.460 2.680 ;
        RECT 124.300 0.010 127.140 2.680 ;
        RECT 127.980 0.010 131.280 2.680 ;
        RECT 132.120 0.010 135.420 2.680 ;
        RECT 136.260 0.010 136.440 2.680 ;
      LAYER met3 ;
        RECT 10.555 136.320 135.270 136.720 ;
        RECT 10.555 132.280 136.720 136.320 ;
        RECT 10.555 130.880 135.270 132.280 ;
        RECT 10.555 127.520 136.720 130.880 ;
        RECT 10.555 126.120 135.270 127.520 ;
        RECT 10.555 122.080 136.720 126.120 ;
        RECT 10.555 120.680 135.270 122.080 ;
        RECT 10.555 116.640 136.720 120.680 ;
        RECT 10.555 115.240 135.270 116.640 ;
        RECT 10.555 111.880 136.720 115.240 ;
        RECT 10.555 110.480 135.270 111.880 ;
        RECT 10.555 106.440 136.720 110.480 ;
        RECT 10.555 105.040 135.270 106.440 ;
        RECT 10.555 101.000 136.720 105.040 ;
        RECT 10.555 99.600 135.270 101.000 ;
        RECT 10.555 96.240 136.720 99.600 ;
        RECT 10.555 94.840 135.270 96.240 ;
        RECT 10.555 90.800 136.720 94.840 ;
        RECT 10.555 89.400 135.270 90.800 ;
        RECT 10.555 86.040 136.720 89.400 ;
        RECT 10.555 84.640 135.270 86.040 ;
        RECT 10.555 80.600 136.720 84.640 ;
        RECT 10.555 79.200 135.270 80.600 ;
        RECT 10.555 75.160 136.720 79.200 ;
        RECT 10.555 73.760 135.270 75.160 ;
        RECT 10.555 70.400 136.720 73.760 ;
        RECT 10.555 69.000 135.270 70.400 ;
        RECT 10.555 64.960 136.720 69.000 ;
        RECT 10.555 63.560 135.270 64.960 ;
        RECT 10.555 59.520 136.720 63.560 ;
        RECT 10.555 58.120 135.270 59.520 ;
        RECT 10.555 54.760 136.720 58.120 ;
        RECT 10.555 53.360 135.270 54.760 ;
        RECT 10.555 49.320 136.720 53.360 ;
        RECT 10.555 47.920 135.270 49.320 ;
        RECT 10.555 44.560 136.720 47.920 ;
        RECT 10.555 43.160 135.270 44.560 ;
        RECT 10.555 39.120 136.720 43.160 ;
        RECT 10.555 37.720 135.270 39.120 ;
        RECT 10.555 33.680 136.720 37.720 ;
        RECT 10.555 32.280 135.270 33.680 ;
        RECT 10.555 28.920 136.720 32.280 ;
        RECT 10.555 27.520 135.270 28.920 ;
        RECT 10.555 23.480 136.720 27.520 ;
        RECT 10.555 22.080 135.270 23.480 ;
        RECT 10.555 18.040 136.720 22.080 ;
        RECT 10.555 16.640 135.270 18.040 ;
        RECT 10.555 13.280 136.720 16.640 ;
        RECT 10.555 11.880 135.270 13.280 ;
        RECT 10.555 7.840 136.720 11.880 ;
        RECT 10.555 6.440 135.270 7.840 ;
        RECT 10.555 3.080 136.720 6.440 ;
        RECT 10.555 1.680 135.270 3.080 ;
        RECT 10.555 0.175 136.720 1.680 ;
      LAYER met4 ;
        RECT 10.820 10.240 25.725 128.080 ;
        RECT 28.125 10.240 49.055 128.080 ;
        RECT 51.455 10.240 137.120 128.080 ;
        RECT 10.820 1.110 137.120 10.240 ;
      LAYER met5 ;
        RECT 10.610 0.900 137.330 60.300 ;
  END
END sb_0__3_
END LIBRARY

