* NGSPICE file created from sb_1__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand3_4 abstract view
.subckt scs8hd_nand3_4 A B C Y vgnd vpwr
.ends

.subckt sb_1__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] chanx_left_in[0] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_bottom_grid_pin_11_ left_bottom_grid_pin_13_ left_bottom_grid_pin_15_ left_bottom_grid_pin_1_
+ left_bottom_grid_pin_3_ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_
+ left_top_grid_pin_10_ right_bottom_grid_pin_11_ right_bottom_grid_pin_13_ right_bottom_grid_pin_15_
+ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_ right_bottom_grid_pin_7_
+ right_bottom_grid_pin_9_ right_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_
+ vpwr vgnd
XFILLER_39_233 vgnd vpwr scs8hd_decap_8
XFILLER_39_211 vgnd vpwr scs8hd_decap_12
XFILLER_22_144 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_115 vpwr vgnd scs8hd_fill_2
XFILLER_13_199 vpwr vgnd scs8hd_fill_2
XANTENNA__113__B _112_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_181 vpwr vgnd scs8hd_fill_2
XFILLER_27_258 vgnd vpwr scs8hd_decap_12
XFILLER_27_236 vpwr vgnd scs8hd_fill_2
XFILLER_27_225 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_118 vgnd vpwr scs8hd_decap_8
XFILLER_10_103 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_18_247 vgnd vpwr scs8hd_decap_3
XANTENNA__108__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_206 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__209__A _209_/A vgnd vpwr scs8hd_diode_2
X_200_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_217 vgnd vpwr scs8hd_fill_1
X_131_ _113_/A _128_/X _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XANTENNA__119__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_21_209 vpwr vgnd scs8hd_fill_2
XFILLER_12_209 vgnd vpwr scs8hd_decap_4
XFILLER_20_242 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_20 vgnd vpwr scs8hd_decap_8
XFILLER_18_64 vpwr vgnd scs8hd_fill_2
XFILLER_34_30 vgnd vpwr scs8hd_fill_1
XFILLER_11_231 vgnd vpwr scs8hd_decap_3
X_114_ _114_/A _112_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_128 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__121__B _124_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_10 vpwr vgnd scs8hd_fill_2
XFILLER_20_21 vgnd vpwr scs8hd_decap_4
XANTENNA__116__B _112_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_172 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _106_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _179_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_25_175 vgnd vpwr scs8hd_decap_6
XFILLER_25_142 vgnd vpwr scs8hd_decap_4
XFILLER_15_21 vgnd vpwr scs8hd_decap_4
XFILLER_15_32 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_fill_1
XFILLER_31_31 vpwr vgnd scs8hd_fill_2
XFILLER_31_97 vpwr vgnd scs8hd_fill_2
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XFILLER_0_274 vgnd vpwr scs8hd_decap_3
XFILLER_31_123 vgnd vpwr scs8hd_decap_8
XFILLER_31_101 vgnd vpwr scs8hd_decap_3
XANTENNA__127__A address[4] vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_223 vpwr vgnd scs8hd_fill_2
XFILLER_39_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_112 vgnd vpwr scs8hd_decap_6
XFILLER_22_189 vgnd vpwr scs8hd_decap_4
XFILLER_13_101 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_3
XFILLER_13_156 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_127 vgnd vpwr scs8hd_fill_1
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_44 vgnd vpwr scs8hd_decap_6
XFILLER_12_88 vpwr vgnd scs8hd_fill_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_3
XFILLER_18_259 vgnd vpwr scs8hd_decap_12
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XFILLER_5_174 vpwr vgnd scs8hd_fill_2
XFILLER_5_141 vpwr vgnd scs8hd_fill_2
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_7_ mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_207 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_130_ _112_/A _128_/X _130_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XANTENNA__119__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__135__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_273 vpwr vgnd scs8hd_fill_2
XFILLER_20_232 vgnd vpwr scs8hd_fill_1
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_32 vgnd vpwr scs8hd_fill_1
X_113_ _113_/A _112_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_210 vpwr vgnd scs8hd_fill_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_5_ mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_4_228 vgnd vpwr scs8hd_decap_12
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XANTENNA__132__B _128_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_151 vpwr vgnd scs8hd_fill_2
XFILLER_19_184 vpwr vgnd scs8hd_fill_2
XFILLER_19_195 vpwr vgnd scs8hd_fill_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_198 vgnd vpwr scs8hd_decap_4
XFILLER_31_65 vpwr vgnd scs8hd_fill_2
XFILLER_15_88 vpwr vgnd scs8hd_fill_2
XFILLER_31_87 vgnd vpwr scs8hd_decap_4
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__127__B _163_/B vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_187 vgnd vpwr scs8hd_decap_6
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_190 vpwr vgnd scs8hd_fill_2
XFILLER_22_168 vgnd vpwr scs8hd_decap_8
XFILLER_26_32 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _144_/Y mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_9_139 vpwr vgnd scs8hd_fill_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_161 vpwr vgnd scs8hd_fill_2
XFILLER_8_150 vgnd vpwr scs8hd_decap_3
XFILLER_8_194 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_37_31 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_41_263 vgnd vpwr scs8hd_decap_12
XANTENNA__140__B _136_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_77 vgnd vpwr scs8hd_decap_6
XFILLER_23_44 vgnd vpwr scs8hd_decap_4
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XANTENNA__119__C address[5] vgnd vpwr scs8hd_diode_2
XFILLER_14_230 vgnd vpwr scs8hd_decap_4
X_189_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__135__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__151__A _151_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _144_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_8
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _181_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_88 vgnd vpwr scs8hd_decap_4
X_112_ _112_/A _112_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_204 vgnd vpwr scs8hd_decap_12
XFILLER_15_8 vpwr vgnd scs8hd_fill_2
XANTENNA__146__A _146_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_119 vgnd vpwr scs8hd_fill_1
XFILLER_29_108 vgnd vpwr scs8hd_decap_4
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_20_56 vpwr vgnd scs8hd_fill_2
XFILLER_20_67 vpwr vgnd scs8hd_fill_2
XFILLER_29_76 vpwr vgnd scs8hd_fill_2
XFILLER_29_43 vpwr vgnd scs8hd_fill_2
XFILLER_28_152 vgnd vpwr scs8hd_fill_1
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_188 vgnd vpwr scs8hd_fill_1
XFILLER_15_45 vpwr vgnd scs8hd_fill_2
XFILLER_15_56 vgnd vpwr scs8hd_decap_3
XFILLER_15_67 vpwr vgnd scs8hd_fill_2
XFILLER_31_44 vpwr vgnd scs8hd_fill_2
XFILLER_31_22 vpwr vgnd scs8hd_fill_2
XFILLER_31_11 vgnd vpwr scs8hd_decap_4
XFILLER_16_144 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _176_/HI mem_right_track_0.LATCH_2_.latch/Q
+ mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C address[5] vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_177 vgnd vpwr scs8hd_fill_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_66 vgnd vpwr scs8hd_decap_6
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_88 vgnd vpwr scs8hd_decap_4
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_147 vpwr vgnd scs8hd_fill_2
XFILLER_13_169 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_21_191 vpwr vgnd scs8hd_fill_2
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__138__B _136_/X vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_128 vpwr vgnd scs8hd_fill_2
XFILLER_18_206 vgnd vpwr scs8hd_fill_1
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_37_43 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_275 vpwr vgnd scs8hd_fill_2
XFILLER_41_253 vpwr vgnd scs8hd_fill_2
XFILLER_5_110 vpwr vgnd scs8hd_fill_2
XFILLER_38_7 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _157_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A _149_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A left_bottom_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XFILLER_23_220 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__119__D _135_/D vgnd vpwr scs8hd_diode_2
X_188_ _188_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__135__C address[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_4
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
X_111_ _111_/A _112_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_216 vgnd vpwr scs8hd_decap_12
XFILLER_11_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _144_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__162__A _095_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_153 vgnd vpwr scs8hd_fill_1
XANTENNA__072__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_29_22 vpwr vgnd scs8hd_fill_2
XFILLER_20_46 vgnd vpwr scs8hd_decap_8
XFILLER_28_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_6 vpwr vgnd scs8hd_fill_2
XFILLER_20_7 vgnd vpwr scs8hd_fill_1
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vpwr vgnd scs8hd_fill_2
XFILLER_25_101 vpwr vgnd scs8hd_fill_2
XFILLER_25_134 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_16_167 vpwr vgnd scs8hd_fill_2
XFILLER_31_159 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__D _135_/D vgnd vpwr scs8hd_diode_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_45 vgnd vpwr scs8hd_decap_8
XFILLER_26_23 vgnd vpwr scs8hd_decap_3
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_119 vgnd vpwr scs8hd_decap_3
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XANTENNA__154__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _087_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_229 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_107 vpwr vgnd scs8hd_fill_2
XANTENNA__080__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_229 vgnd vpwr scs8hd_decap_4
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_5_133 vpwr vgnd scs8hd_fill_2
XANTENNA__149__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_17_262 vgnd vpwr scs8hd_decap_4
XFILLER_17_273 vgnd vpwr scs8hd_decap_4
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_23_265 vpwr vgnd scs8hd_fill_2
XFILLER_23_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__075__A _074_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_14_243 vpwr vgnd scs8hd_fill_2
XFILLER_14_254 vgnd vpwr scs8hd_decap_8
XFILLER_14_265 vgnd vpwr scs8hd_decap_8
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__135__D _135_/D vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_224 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_68 vgnd vpwr scs8hd_decap_4
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _110_/A _112_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_228 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_121 vgnd vpwr scs8hd_fill_1
XFILLER_37_110 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_187 vpwr vgnd scs8hd_fill_2
XFILLER_28_154 vgnd vpwr scs8hd_fill_1
XFILLER_28_121 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_220 vgnd vpwr scs8hd_decap_4
XFILLER_19_132 vgnd vpwr scs8hd_decap_4
XANTENNA__157__B _157_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_146 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XANTENNA__067__B _067_/B vgnd vpwr scs8hd_diode_2
XANTENNA__083__A _082_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_25 vgnd vpwr scs8hd_fill_1
XFILLER_31_79 vpwr vgnd scs8hd_fill_2
XFILLER_31_138 vgnd vpwr scs8hd_decap_4
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_113 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_249 vgnd vpwr scs8hd_decap_4
XANTENNA__168__A _080_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_190 vpwr vgnd scs8hd_fill_2
XFILLER_22_127 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_271 vgnd vpwr scs8hd_decap_4
XANTENNA__078__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_182 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XFILLER_12_171 vgnd vpwr scs8hd_fill_1
XANTENNA__170__B _169_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vpwr vgnd scs8hd_fill_2
XFILLER_35_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__080__B _080_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
XFILLER_26_252 vgnd vpwr scs8hd_decap_8
XFILLER_26_241 vgnd vpwr scs8hd_decap_4
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _090_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_track_8.LATCH_1_.latch data_in _145_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_178 vgnd vpwr scs8hd_decap_4
XFILLER_5_123 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__149__C address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__165__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_8
XFILLER_23_14 vpwr vgnd scs8hd_fill_2
XFILLER_23_25 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_9_16 vgnd vpwr scs8hd_decap_12
X_186_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_36_6 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_247 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A _085_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_203 vpwr vgnd scs8hd_fill_2
XFILLER_11_214 vpwr vgnd scs8hd_fill_2
XFILLER_11_236 vgnd vpwr scs8hd_decap_8
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
XANTENNA__162__C _085_/C vgnd vpwr scs8hd_diode_2
X_169_ _101_/A _169_/B _169_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_166 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_243 vgnd vpwr scs8hd_fill_1
XFILLER_19_100 vgnd vpwr scs8hd_decap_3
XFILLER_19_155 vpwr vgnd scs8hd_fill_2
XFILLER_19_199 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_158 vpwr vgnd scs8hd_fill_2
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XANTENNA__067__C _082_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_69 vpwr vgnd scs8hd_fill_2
XFILLER_31_106 vgnd vpwr scs8hd_decap_4
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vgnd vpwr scs8hd_decap_3
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _169_/B vgnd vpwr scs8hd_diode_2
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_194 vgnd vpwr scs8hd_decap_6
XFILLER_30_161 vgnd vpwr scs8hd_decap_3
XFILLER_15_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__078__B _067_/B vgnd vpwr scs8hd_diode_2
XANTENNA__094__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_13_139 vpwr vgnd scs8hd_fill_2
Xmem_top_track_14.LATCH_0_.latch data_in _148_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_161 vpwr vgnd scs8hd_fill_2
XFILLER_12_150 vgnd vpwr scs8hd_decap_3
XFILLER_8_165 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _143_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_275 vpwr vgnd scs8hd_fill_2
XFILLER_35_253 vpwr vgnd scs8hd_fill_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XANTENNA__089__A _088_/X vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _169_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_5_ mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_209 vgnd vpwr scs8hd_decap_3
XFILLER_41_245 vgnd vpwr scs8hd_decap_8
XFILLER_5_157 vpwr vgnd scs8hd_fill_2
XFILLER_5_146 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XFILLER_17_220 vgnd vpwr scs8hd_decap_3
XANTENNA__165__C _074_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_48 vgnd vpwr scs8hd_fill_1
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XANTENNA__091__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_185_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_9_28 vgnd vpwr scs8hd_decap_12
XFILLER_13_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_259 vgnd vpwr scs8hd_decap_12
XFILLER_24_91 vgnd vpwr scs8hd_fill_1
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
X_168_ _080_/B _169_/B _168_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_3 vpwr vgnd scs8hd_fill_2
X_099_ _080_/B _112_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_156 vgnd vpwr scs8hd_decap_12
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XANTENNA__187__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
XFILLER_29_47 vgnd vpwr scs8hd_decap_3
XANTENNA__097__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_93 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_33_170 vgnd vpwr scs8hd_decap_12
XFILLER_15_49 vgnd vpwr scs8hd_decap_4
XFILLER_31_48 vgnd vpwr scs8hd_decap_12
XFILLER_31_26 vgnd vpwr scs8hd_decap_3
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
XFILLER_16_148 vpwr vgnd scs8hd_fill_2
XFILLER_31_118 vgnd vpwr scs8hd_decap_4
XFILLER_24_170 vgnd vpwr scs8hd_decap_12
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_92 vpwr vgnd scs8hd_fill_2
XFILLER_39_229 vpwr vgnd scs8hd_fill_2
XFILLER_39_207 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_30_173 vgnd vpwr scs8hd_decap_8
XANTENNA__078__C _085_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_195 vgnd vpwr scs8hd_fill_1
XFILLER_8_177 vpwr vgnd scs8hd_fill_2
XFILLER_12_140 vgnd vpwr scs8hd_decap_4
XANTENNA__195__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XFILLER_12_17 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_213 vgnd vpwr scs8hd_decap_4
XFILLER_23_235 vpwr vgnd scs8hd_fill_2
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XANTENNA__091__C _085_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_9_ mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_15_ mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_184_ _184_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _179_/HI mem_top_track_0.LATCH_5_.latch/Q
+ mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_227 vpwr vgnd scs8hd_fill_2
XFILLER_11_249 vgnd vpwr scs8hd_decap_12
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_098_ _111_/A _106_/B _098_/Y vgnd vpwr scs8hd_nor2_4
X_167_ _152_/A _169_/B _167_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_168 vgnd vpwr scs8hd_decap_12
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_26 vpwr vgnd scs8hd_fill_2
XFILLER_28_146 vgnd vpwr scs8hd_decap_6
XFILLER_28_102 vgnd vpwr scs8hd_decap_3
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_92 vpwr vgnd scs8hd_fill_2
XFILLER_19_168 vgnd vpwr scs8hd_decap_4
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XANTENNA__198__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_33_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_138 vpwr vgnd scs8hd_fill_2
XFILLER_15_28 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_116 vgnd vpwr scs8hd_decap_6
XFILLER_24_193 vpwr vgnd scs8hd_fill_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_71 vpwr vgnd scs8hd_fill_2
XFILLER_11_7 vgnd vpwr scs8hd_fill_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_22_108 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_141 vgnd vpwr scs8hd_decap_4
XFILLER_21_174 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _174_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_263 vgnd vpwr scs8hd_decap_12
XFILLER_29_241 vgnd vpwr scs8hd_decap_3
XFILLER_29_230 vgnd vpwr scs8hd_decap_8
XFILLER_16_93 vgnd vpwr scs8hd_decap_4
XFILLER_8_145 vgnd vpwr scs8hd_decap_3
XFILLER_12_163 vpwr vgnd scs8hd_fill_2
XFILLER_12_174 vpwr vgnd scs8hd_fill_2
XFILLER_12_185 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_12_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_137 vpwr vgnd scs8hd_fill_2
XFILLER_27_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _192_/A vgnd vpwr scs8hd_inv_1
XFILLER_4_170 vpwr vgnd scs8hd_fill_2
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_23_258 vgnd vpwr scs8hd_decap_4
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _209_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_247 vgnd vpwr scs8hd_decap_4
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_206 vgnd vpwr scs8hd_decap_6
XFILLER_20_228 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _175_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_250 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_097_ _096_/X _106_/B vgnd vpwr scs8hd_buf_1
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_166_ _165_/X _169_/B vgnd vpwr scs8hd_buf_1
XFILLER_37_147 vgnd vpwr scs8hd_decap_6
XFILLER_1_31 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XFILLER_28_125 vpwr vgnd scs8hd_fill_2
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_3_224 vgnd vpwr scs8hd_fill_1
XFILLER_10_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_71 vgnd vpwr scs8hd_decap_4
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_27_191 vgnd vpwr scs8hd_decap_4
X_149_ _149_/A address[6] address[5] _150_/C vgnd vpwr scs8hd_or3_4
XFILLER_18_180 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_161 vpwr vgnd scs8hd_fill_2
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_38_253 vpwr vgnd scs8hd_fill_2
XFILLER_26_28 vgnd vpwr scs8hd_decap_3
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_275 vpwr vgnd scs8hd_fill_2
XFILLER_29_253 vpwr vgnd scs8hd_fill_2
XFILLER_8_102 vgnd vpwr scs8hd_decap_3
XFILLER_8_157 vpwr vgnd scs8hd_fill_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_204 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vpwr vgnd scs8hd_fill_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_29 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_226 vpwr vgnd scs8hd_fill_2
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_62 vgnd vpwr scs8hd_decap_4
XFILLER_13_73 vpwr vgnd scs8hd_fill_2
XFILLER_13_95 vgnd vpwr scs8hd_decap_4
XFILLER_29_9 vpwr vgnd scs8hd_fill_2
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_7 vgnd vpwr scs8hd_decap_12
X_165_ address[4] address[3] _074_/B _165_/X vgnd vpwr scs8hd_or3_4
XFILLER_10_262 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_7 vgnd vpwr scs8hd_decap_8
X_096_ _074_/B _095_/X _096_/X vgnd vpwr scs8hd_or2_4
XFILLER_37_115 vgnd vpwr scs8hd_decap_6
XFILLER_1_43 vgnd vpwr scs8hd_decap_12
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _156_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_39 vpwr vgnd scs8hd_fill_2
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_10_74 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_148_ _148_/A _148_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_3 vgnd vpwr scs8hd_decap_4
X_079_ _078_/X _080_/B vgnd vpwr scs8hd_buf_1
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_18 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _138_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_151 vpwr vgnd scs8hd_fill_2
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_154 vgnd vpwr scs8hd_decap_4
XPHY_4 vgnd vpwr scs8hd_decap_3
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 left_bottom_grid_pin_1_ mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_184 vgnd vpwr scs8hd_decap_4
XFILLER_7_97 vpwr vgnd scs8hd_fill_2
XFILLER_7_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_132 vgnd vpwr scs8hd_decap_3
XFILLER_21_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _144_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_121 vgnd vpwr scs8hd_decap_4
XFILLER_16_84 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A _087_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_224 vgnd vpwr scs8hd_decap_6
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_40_271 vgnd vpwr scs8hd_decap_4
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XANTENNA__100__B _106_/B vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_18 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_190 vgnd vpwr scs8hd_fill_1
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_62 vpwr vgnd scs8hd_fill_2
XFILLER_10_274 vgnd vpwr scs8hd_fill_1
X_164_ _163_/A _163_/B _159_/B _085_/C _164_/Y vgnd vpwr scs8hd_nor4_4
X_095_ _163_/A address[3] _095_/X vgnd vpwr scs8hd_or2_4
XFILLER_27_7 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_55 vgnd vpwr scs8hd_decap_6
XFILLER_28_138 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_171 vgnd vpwr scs8hd_decap_4
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XFILLER_27_182 vgnd vpwr scs8hd_fill_1
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_078_ address[1] _067_/B _085_/C _078_/X vgnd vpwr scs8hd_or3_4
X_147_ _147_/A _147_/Y vgnd vpwr scs8hd_inv_8
XFILLER_18_3 vpwr vgnd scs8hd_fill_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_96 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_122 vgnd vpwr scs8hd_fill_1
XFILLER_26_19 vpwr vgnd scs8hd_fill_2
XFILLER_21_100 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_200 vgnd vpwr scs8hd_decap_3
XFILLER_32_62 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_247 vpwr vgnd scs8hd_fill_2
XANTENNA__204__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_5_118 vgnd vpwr scs8hd_decap_4
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_73 vpwr vgnd scs8hd_fill_2
XFILLER_17_236 vgnd vpwr scs8hd_decap_6
XFILLER_17_258 vpwr vgnd scs8hd_fill_2
XFILLER_17_269 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_162 vgnd vpwr scs8hd_decap_3
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_239 vgnd vpwr scs8hd_decap_3
XFILLER_23_217 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_206 vgnd vpwr scs8hd_decap_6
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
X_180_ _180_/HI _180_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XFILLER_9_210 vgnd vpwr scs8hd_decap_4
XANTENNA__109__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_85 vgnd vpwr scs8hd_decap_6
XFILLER_24_41 vpwr vgnd scs8hd_fill_2
X_094_ address[4] _163_/A vgnd vpwr scs8hd_inv_8
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
X_163_ _163_/A _163_/B _159_/B _082_/C _163_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__111__B _112_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _087_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_227 vgnd vpwr scs8hd_decap_12
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_19_41 vpwr vgnd scs8hd_fill_2
XFILLER_19_96 vpwr vgnd scs8hd_fill_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XANTENNA__106__B _106_/B vgnd vpwr scs8hd_diode_2
X_077_ address[0] _085_/C vgnd vpwr scs8hd_buf_1
X_146_ _146_/A _146_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__122__A _112_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_16_109 vgnd vpwr scs8hd_decap_4
XANTENNA__207__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_24_197 vpwr vgnd scs8hd_fill_2
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_101 vgnd vpwr scs8hd_decap_12
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_175 vgnd vpwr scs8hd_decap_3
XFILLER_30_145 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A enable vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vpwr vgnd scs8hd_fill_2
X_129_ _111_/A _128_/X _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_21_145 vgnd vpwr scs8hd_fill_1
XFILLER_21_178 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_8
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_101 vgnd vpwr scs8hd_decap_3
XFILLER_16_53 vgnd vpwr scs8hd_fill_1
XFILLER_32_96 vgnd vpwr scs8hd_decap_8
XFILLER_8_127 vgnd vpwr scs8hd_decap_3
XFILLER_12_167 vgnd vpwr scs8hd_decap_4
XFILLER_12_189 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _178_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_193 vgnd vpwr scs8hd_decap_8
XFILLER_37_19 vgnd vpwr scs8hd_decap_12
XFILLER_27_52 vpwr vgnd scs8hd_fill_2
XFILLER_27_30 vpwr vgnd scs8hd_fill_2
XFILLER_17_204 vgnd vpwr scs8hd_decap_6
XFILLER_17_215 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_96 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B _112_/B vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_174 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_270 vgnd vpwr scs8hd_decap_4
XFILLER_13_10 vpwr vgnd scs8hd_fill_2
XFILLER_13_21 vpwr vgnd scs8hd_fill_2
XFILLER_13_32 vpwr vgnd scs8hd_fill_2
XFILLER_13_43 vgnd vpwr scs8hd_decap_4
XFILLER_22_273 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_3 vpwr vgnd scs8hd_fill_2
XFILLER_9_233 vgnd vpwr scs8hd_decap_8
Xmem_top_track_14.LATCH_1_.latch data_in _147_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__109__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_181 vpwr vgnd scs8hd_fill_2
XFILLER_39_170 vpwr vgnd scs8hd_fill_2
XFILLER_24_75 vpwr vgnd scs8hd_fill_2
X_162_ _095_/X _159_/B _085_/C _162_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ _090_/A _107_/A _093_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _168_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_107 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_239 vgnd vpwr scs8hd_decap_4
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_77 vgnd vpwr scs8hd_decap_4
XFILLER_10_88 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_145_ _145_/A _145_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_7 vgnd vpwr scs8hd_decap_8
XANTENNA__122__B _124_/B vgnd vpwr scs8hd_diode_2
X_076_ _111_/A _090_/A _076_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vpwr vgnd scs8hd_fill_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_21 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_165 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
X_128_ _127_/X _128_/X vgnd vpwr scs8hd_buf_1
XANTENNA__133__A _106_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_213 vgnd vpwr scs8hd_fill_1
XFILLER_21_157 vpwr vgnd scs8hd_fill_2
XFILLER_29_213 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XFILLER_16_65 vgnd vpwr scs8hd_decap_8
XFILLER_12_146 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__128__A _127_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_172 vgnd vpwr scs8hd_decap_4
Xmux_top_track_2.INVTX1_2_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_208 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__130__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_186 vgnd vpwr scs8hd_decap_12
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_252 vgnd vpwr scs8hd_decap_4
XFILLER_13_88 vgnd vpwr scs8hd_decap_4
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XANTENNA__125__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__109__C _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_252 vpwr vgnd scs8hd_fill_2
XANTENNA__141__A _106_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_161_ _095_/X _159_/B _082_/C _161_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
X_092_ _091_/X _107_/A vgnd vpwr scs8hd_buf_1
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _102_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__136__A _135_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XFILLER_19_21 vgnd vpwr scs8hd_decap_4
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_152 vpwr vgnd scs8hd_fill_2
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_075_ _074_/X _090_/A vgnd vpwr scs8hd_buf_1
X_144_ _144_/A _144_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_33_111 vgnd vpwr scs8hd_decap_8
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_158 vgnd vpwr scs8hd_fill_1
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_111 vpwr vgnd scs8hd_fill_2
XFILLER_15_144 vpwr vgnd scs8hd_fill_2
X_127_ address[4] _163_/B address[5] _135_/D _127_/X vgnd vpwr scs8hd_or4_4
XANTENNA__133__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_4
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_107 vgnd vpwr scs8hd_decap_3
XFILLER_12_125 vgnd vpwr scs8hd_fill_1
XFILLER_12_136 vpwr vgnd scs8hd_fill_2
XFILLER_16_99 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_206 vgnd vpwr scs8hd_decap_6
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _147_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_198 vgnd vpwr scs8hd_decap_12
XFILLER_4_154 vgnd vpwr scs8hd_decap_8
XFILLER_31_253 vpwr vgnd scs8hd_fill_2
XFILLER_31_242 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_209 vpwr vgnd scs8hd_fill_2
XFILLER_31_275 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XFILLER_13_264 vgnd vpwr scs8hd_decap_12
XANTENNA__141__B _136_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_22 vgnd vpwr scs8hd_decap_6
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
X_091_ address[1] address[2] _085_/C _091_/X vgnd vpwr scs8hd_or3_4
X_160_ _074_/A _159_/B _085_/C _160_/Y vgnd vpwr scs8hd_nor3_4
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_1_ mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _152_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_68 vgnd vpwr scs8hd_decap_6
XFILLER_19_77 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_27_175 vgnd vpwr scs8hd_fill_1
X_074_ _074_/A _074_/B _074_/X vgnd vpwr scs8hd_or2_4
X_143_ _143_/A _143_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_7 vpwr vgnd scs8hd_fill_2
XANTENNA__147__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_123 vpwr vgnd scs8hd_fill_2
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_34 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_126_ _108_/A _124_/B _126_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_259 vgnd vpwr scs8hd_decap_12
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_21_137 vpwr vgnd scs8hd_fill_2
XFILLER_29_259 vpwr vgnd scs8hd_fill_2
XFILLER_29_226 vpwr vgnd scs8hd_fill_2
XFILLER_8_119 vgnd vpwr scs8hd_decap_8
XFILLER_16_45 vgnd vpwr scs8hd_decap_8
XFILLER_32_77 vgnd vpwr scs8hd_decap_12
XFILLER_32_66 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_130 vgnd vpwr scs8hd_decap_4
X_109_ _163_/A _163_/B _074_/B _110_/A vgnd vpwr scs8hd_or3_4
XANTENNA__160__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_11 vpwr vgnd scs8hd_fill_2
XANTENNA__070__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_27_77 vpwr vgnd scs8hd_fill_2
XFILLER_27_22 vpwr vgnd scs8hd_fill_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_210 vgnd vpwr scs8hd_decap_12
XANTENNA__139__B _136_/X vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__065__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_22_232 vgnd vpwr scs8hd_fill_1
XFILLER_22_265 vgnd vpwr scs8hd_decap_8
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_214 vgnd vpwr scs8hd_fill_1
XFILLER_13_243 vgnd vpwr scs8hd_fill_1
XFILLER_13_276 vgnd vpwr scs8hd_fill_1
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_39_195 vpwr vgnd scs8hd_fill_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_6
XFILLER_24_45 vpwr vgnd scs8hd_fill_2
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
X_090_ _090_/A _090_/B _090_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__152__B _157_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_22 vgnd vpwr scs8hd_decap_12
XFILLER_35_11 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_45 vgnd vpwr scs8hd_decap_3
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_27_187 vpwr vgnd scs8hd_fill_2
X_142_ _108_/A _136_/X _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_073_ enable _073_/B address[5] _074_/B vgnd vpwr scs8hd_nand3_4
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XFILLER_18_110 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__A enable vgnd vpwr scs8hd_diode_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_21_79 vpwr vgnd scs8hd_fill_2
XFILLER_15_135 vpwr vgnd scs8hd_fill_2
XFILLER_30_149 vgnd vpwr scs8hd_decap_4
XFILLER_30_116 vgnd vpwr scs8hd_decap_6
XFILLER_23_190 vpwr vgnd scs8hd_fill_2
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
X_125_ _106_/A _124_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_7 vgnd vpwr scs8hd_decap_6
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_38_205 vgnd vpwr scs8hd_decap_8
XFILLER_23_6 vpwr vgnd scs8hd_fill_2
XANTENNA__158__A _150_/C vgnd vpwr scs8hd_diode_2
XFILLER_29_205 vgnd vpwr scs8hd_fill_1
XFILLER_29_238 vgnd vpwr scs8hd_fill_1
XANTENNA__068__A _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_89 vgnd vpwr scs8hd_decap_3
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _155_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_171 vgnd vpwr scs8hd_decap_8
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XFILLER_28_271 vgnd vpwr scs8hd_decap_4
X_108_ _108_/A _106_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_153 vpwr vgnd scs8hd_fill_2
XANTENNA__160__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_3
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_80 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _206_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_45 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _137_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_263 vpwr vgnd scs8hd_fill_2
XFILLER_25_252 vpwr vgnd scs8hd_fill_2
XFILLER_25_241 vgnd vpwr scs8hd_decap_3
XFILLER_4_101 vgnd vpwr scs8hd_decap_3
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_222 vgnd vpwr scs8hd_decap_12
XFILLER_16_252 vgnd vpwr scs8hd_decap_3
XFILLER_16_274 vgnd vpwr scs8hd_fill_1
XANTENNA__155__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _090_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_47 vgnd vpwr scs8hd_fill_1
XFILLER_13_69 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_7 vgnd vpwr scs8hd_decap_12
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XANTENNA__081__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_222 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_174 vgnd vpwr scs8hd_decap_4
XFILLER_39_130 vgnd vpwr scs8hd_decap_8
XFILLER_24_79 vgnd vpwr scs8hd_decap_4
XANTENNA__076__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_35_34 vgnd vpwr scs8hd_decap_12
XFILLER_27_100 vgnd vpwr scs8hd_decap_3
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
X_210_ _210_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_141_ _106_/A _136_/X _141_/Y vgnd vpwr scs8hd_nor2_4
X_072_ address[6] _073_/B vgnd vpwr scs8hd_inv_8
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _145_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_133 vgnd vpwr scs8hd_fill_1
XFILLER_33_158 vgnd vpwr scs8hd_decap_12
XFILLER_33_147 vgnd vpwr scs8hd_decap_4
XFILLER_18_188 vgnd vpwr scs8hd_decap_3
XANTENNA__163__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XFILLER_24_158 vgnd vpwr scs8hd_fill_1
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_128 vgnd vpwr scs8hd_decap_8
XFILLER_15_169 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
X_124_ _114_/A _124_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_91 vpwr vgnd scs8hd_fill_2
XFILLER_38_239 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_46 vgnd vpwr scs8hd_decap_12
XFILLER_32_35 vpwr vgnd scs8hd_fill_2
XFILLER_12_128 vgnd vpwr scs8hd_fill_1
XANTENNA__084__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_150 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_176 vgnd vpwr scs8hd_fill_1
XFILLER_11_161 vpwr vgnd scs8hd_fill_2
X_107_ _107_/A _108_/A vgnd vpwr scs8hd_buf_1
XANTENNA__160__C _085_/C vgnd vpwr scs8hd_diode_2
XANTENNA__169__A _101_/A vgnd vpwr scs8hd_diode_2
XANTENNA__079__A _078_/X vgnd vpwr scs8hd_diode_2
XFILLER_25_275 vpwr vgnd scs8hd_fill_2
XFILLER_4_113 vgnd vpwr scs8hd_decap_12
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_8
XFILLER_31_234 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _146_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__171__B _169_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_58 vpwr vgnd scs8hd_fill_2
XFILLER_10_204 vpwr vgnd scs8hd_fill_2
XFILLER_10_226 vgnd vpwr scs8hd_decap_12
XANTENNA__076__B _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_25 vgnd vpwr scs8hd_fill_1
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_35_46 vgnd vpwr scs8hd_decap_12
XFILLER_27_178 vpwr vgnd scs8hd_fill_2
XFILLER_27_167 vpwr vgnd scs8hd_fill_2
XFILLER_27_145 vgnd vpwr scs8hd_decap_4
XFILLER_27_134 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _090_/A vgnd vpwr scs8hd_diode_2
X_140_ _114_/A _136_/X _140_/Y vgnd vpwr scs8hd_nor2_4
X_071_ address[4] _163_/B _074_/A vgnd vpwr scs8hd_or2_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_145 vpwr vgnd scs8hd_fill_2
XFILLER_18_167 vgnd vpwr scs8hd_decap_4
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__C _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_24_137 vgnd vpwr scs8hd_decap_12
XANTENNA__073__C address[5] vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_115 vgnd vpwr scs8hd_decap_4
XFILLER_15_148 vpwr vgnd scs8hd_fill_2
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
X_123_ _113_/A _124_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_7 vgnd vpwr scs8hd_fill_1
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA__190__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_240 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _084_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_58 vgnd vpwr scs8hd_decap_4
XANTENNA__084__B _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
X_106_ _106_/A _106_/B _106_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_195 vpwr vgnd scs8hd_fill_2
XANTENNA__169__B _169_/B vgnd vpwr scs8hd_diode_2
XANTENNA__185__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_213 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_17_91 vpwr vgnd scs8hd_fill_2
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_202 vpwr vgnd scs8hd_fill_2
XFILLER_22_224 vgnd vpwr scs8hd_decap_8
XFILLER_22_235 vpwr vgnd scs8hd_fill_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_9_217 vgnd vpwr scs8hd_decap_3
XFILLER_13_235 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_250 vgnd vpwr scs8hd_decap_12
XFILLER_39_143 vpwr vgnd scs8hd_fill_2
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_5_94 vgnd vpwr scs8hd_fill_1
XFILLER_39_165 vgnd vpwr scs8hd_fill_1
XFILLER_10_238 vgnd vpwr scs8hd_decap_12
XFILLER_1_19 vgnd vpwr scs8hd_decap_12
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_10_17 vgnd vpwr scs8hd_decap_12
XFILLER_19_37 vpwr vgnd scs8hd_fill_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_35_58 vgnd vpwr scs8hd_decap_3
XANTENNA__087__B _087_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_070_ address[3] _163_/B vgnd vpwr scs8hd_inv_8
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_top_in[6] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _148_/A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__163__D _082_/C vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_127 vgnd vpwr scs8hd_fill_1
XFILLER_32_193 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_38 vgnd vpwr scs8hd_decap_4
XANTENNA__098__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_127 vgnd vpwr scs8hd_fill_1
X_122_ _112_/A _124_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_171 vgnd vpwr scs8hd_fill_1
XFILLER_14_193 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _167_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_263 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_163 vpwr vgnd scs8hd_fill_2
XFILLER_28_241 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_101 vpwr vgnd scs8hd_fill_2
XFILLER_11_130 vpwr vgnd scs8hd_fill_2
XFILLER_11_174 vpwr vgnd scs8hd_fill_2
X_105_ _090_/B _106_/A vgnd vpwr scs8hd_buf_1
XFILLER_27_26 vpwr vgnd scs8hd_fill_2
XFILLER_25_233 vpwr vgnd scs8hd_fill_2
XFILLER_25_222 vpwr vgnd scs8hd_fill_2
XFILLER_40_247 vgnd vpwr scs8hd_decap_8
XANTENNA__095__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_137 vgnd vpwr scs8hd_decap_12
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_181 vpwr vgnd scs8hd_fill_2
XANTENNA__196__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_13_ mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_17 vpwr vgnd scs8hd_fill_2
XFILLER_13_28 vpwr vgnd scs8hd_fill_2
XFILLER_13_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_203 vpwr vgnd scs8hd_fill_2
XFILLER_9_229 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_8_262 vgnd vpwr scs8hd_decap_12
XFILLER_39_199 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_81 vpwr vgnd scs8hd_fill_2
XFILLER_30_70 vgnd vpwr scs8hd_decap_8
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_10_29 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XFILLER_18_125 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_92 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
XFILLER_32_183 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_17 vpwr vgnd scs8hd_fill_2
XANTENNA__098__B _106_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_139 vgnd vpwr scs8hd_decap_3
XFILLER_23_194 vpwr vgnd scs8hd_fill_2
XFILLER_23_150 vpwr vgnd scs8hd_fill_2
X_121_ _111_/A _124_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_50 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_14_183 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__199__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_29_209 vpwr vgnd scs8hd_fill_2
XFILLER_37_275 vpwr vgnd scs8hd_fill_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _100_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_7_168 vpwr vgnd scs8hd_fill_2
XFILLER_11_142 vgnd vpwr scs8hd_decap_4
Xmem_top_track_2.LATCH_0_.latch data_in _144_/A _160_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_104_ _114_/A _106_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_82 vgnd vpwr scs8hd_decap_3
XFILLER_14_6 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_27_49 vgnd vpwr scs8hd_fill_1
XFILLER_25_267 vgnd vpwr scs8hd_decap_8
XFILLER_40_259 vgnd vpwr scs8hd_decap_12
XFILLER_4_149 vgnd vpwr scs8hd_decap_4
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_259 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _175_/HI mem_left_track_9.LATCH_2_.latch/Q
+ mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_248 vpwr vgnd scs8hd_fill_2
XFILLER_13_248 vpwr vgnd scs8hd_fill_2
XFILLER_13_259 vgnd vpwr scs8hd_decap_3
Xmux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ _144_/A mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_8_274 vgnd vpwr scs8hd_fill_1
XFILLER_39_178 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_28 vgnd vpwr scs8hd_fill_1
XFILLER_14_61 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_9_ mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 left_bottom_grid_pin_3_ mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_17 vpwr vgnd scs8hd_fill_2
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _180_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_71 vgnd vpwr scs8hd_decap_4
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
X_197_ _197_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_107 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _202_/A vgnd vpwr scs8hd_inv_1
XFILLER_23_184 vgnd vpwr scs8hd_decap_3
XFILLER_23_173 vpwr vgnd scs8hd_fill_2
X_120_ _119_/X _124_/B vgnd vpwr scs8hd_buf_1
XFILLER_11_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _145_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _180_/HI _147_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_243 vgnd vpwr scs8hd_fill_1
XFILLER_37_232 vgnd vpwr scs8hd_decap_8
XFILLER_32_39 vgnd vpwr scs8hd_decap_4
XFILLER_20_121 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
X_103_ _087_/B _114_/A vgnd vpwr scs8hd_buf_1
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_19_254 vpwr vgnd scs8hd_fill_2
XFILLER_19_265 vgnd vpwr scs8hd_decap_12
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_202 vgnd vpwr scs8hd_fill_1
XFILLER_16_224 vpwr vgnd scs8hd_fill_2
XFILLER_17_72 vpwr vgnd scs8hd_fill_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _146_/A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_260 vgnd vpwr scs8hd_decap_12
XFILLER_5_97 vpwr vgnd scs8hd_fill_2
XFILLER_5_86 vgnd vpwr scs8hd_decap_8
XFILLER_24_18 vpwr vgnd scs8hd_fill_2
XFILLER_10_208 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _197_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_73 vpwr vgnd scs8hd_fill_2
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_27_149 vgnd vpwr scs8hd_fill_1
XFILLER_27_138 vpwr vgnd scs8hd_fill_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_149 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XFILLER_33_119 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_182 vgnd vpwr scs8hd_fill_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_119 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_119 vgnd vpwr scs8hd_fill_1
XFILLER_11_74 vpwr vgnd scs8hd_fill_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_163 vpwr vgnd scs8hd_fill_2
XFILLER_14_196 vgnd vpwr scs8hd_fill_1
X_179_ _179_/HI _179_/LO vgnd vpwr scs8hd_conb_1
XFILLER_16_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_126 vpwr vgnd scs8hd_fill_2
XFILLER_11_199 vpwr vgnd scs8hd_fill_2
X_102_ _113_/A _106_/B _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_51 vgnd vpwr scs8hd_decap_3
XFILLER_19_222 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_4
XFILLER_16_236 vpwr vgnd scs8hd_fill_2
XFILLER_16_247 vgnd vpwr scs8hd_decap_3
XFILLER_16_258 vgnd vpwr scs8hd_decap_12
XFILLER_17_62 vgnd vpwr scs8hd_decap_3
XFILLER_17_95 vgnd vpwr scs8hd_decap_4
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _076_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__104__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_206 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_239 vpwr vgnd scs8hd_fill_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _154_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_12_272 vgnd vpwr scs8hd_decap_3
XFILLER_39_147 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_96 vpwr vgnd scs8hd_fill_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_106 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_194 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_37_7 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_131 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _172_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_14_142 vgnd vpwr scs8hd_decap_4
XANTENNA__107__A _107_/A vgnd vpwr scs8hd_diode_2
X_178_ _178_/HI _178_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_28_3 vgnd vpwr scs8hd_decap_4
XFILLER_32_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_145 vgnd vpwr scs8hd_decap_3
XFILLER_20_167 vpwr vgnd scs8hd_fill_2
XFILLER_20_189 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_112 vpwr vgnd scs8hd_fill_2
XFILLER_11_134 vpwr vgnd scs8hd_fill_2
XFILLER_11_178 vgnd vpwr scs8hd_decap_3
X_101_ _101_/A _113_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_149 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XFILLER_25_248 vpwr vgnd scs8hd_fill_2
XFILLER_25_237 vpwr vgnd scs8hd_fill_2
XFILLER_25_226 vpwr vgnd scs8hd_fill_2
XFILLER_40_207 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_259 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__210__A _210_/A vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_30 vpwr vgnd scs8hd_fill_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_95 vpwr vgnd scs8hd_fill_2
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _119_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _111_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_21_240 vpwr vgnd scs8hd_fill_2
XANTENNA__205__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_28_84 vgnd vpwr scs8hd_decap_8
XFILLER_28_73 vpwr vgnd scs8hd_fill_2
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XANTENNA__115__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_222 vpwr vgnd scs8hd_fill_2
XFILLER_39_159 vgnd vpwr scs8hd_decap_6
XFILLER_39_126 vpwr vgnd scs8hd_fill_2
XFILLER_40_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_181 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_41 vgnd vpwr scs8hd_decap_8
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _183_/HI _145_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_30_96 vgnd vpwr scs8hd_decap_3
XFILLER_30_85 vgnd vpwr scs8hd_decap_6
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XFILLER_29_170 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _146_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_52 vpwr vgnd scs8hd_fill_2
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA__112__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_165 vgnd vpwr scs8hd_decap_12
XFILLER_17_151 vpwr vgnd scs8hd_fill_2
XFILLER_17_184 vgnd vpwr scs8hd_decap_3
XFILLER_23_154 vpwr vgnd scs8hd_fill_2
XFILLER_11_65 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_13_ mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_121 vgnd vpwr scs8hd_decap_4
X_177_ _177_/HI _177_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_187 vgnd vpwr scs8hd_decap_6
XANTENNA__123__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_102 vgnd vpwr scs8hd_decap_3
XFILLER_20_135 vgnd vpwr scs8hd_fill_1
XFILLER_20_179 vgnd vpwr scs8hd_fill_1
XFILLER_28_224 vpwr vgnd scs8hd_fill_2
XANTENNA__208__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_100_ _112_/A _106_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_157 vpwr vgnd scs8hd_fill_2
XFILLER_19_235 vpwr vgnd scs8hd_fill_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _149_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_88 vpwr vgnd scs8hd_fill_2
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _148_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_11_ mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_274 vgnd vpwr scs8hd_fill_1
XFILLER_38_19 vgnd vpwr scs8hd_decap_12
XFILLER_21_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _080_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_230 vgnd vpwr scs8hd_decap_4
XANTENNA__115__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_138 vpwr vgnd scs8hd_fill_2
XANTENNA__131__A _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_193 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_21 vgnd vpwr scs8hd_decap_8
XFILLER_14_32 vgnd vpwr scs8hd_decap_3
XFILLER_14_65 vgnd vpwr scs8hd_decap_8
XFILLER_30_53 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _181_/HI mem_top_track_16.LATCH_5_.latch/Q
+ mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XANTENNA__126__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_174 vgnd vpwr scs8hd_decap_8
XFILLER_26_163 vpwr vgnd scs8hd_fill_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
X_193_ _193_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_97 vpwr vgnd scs8hd_fill_2
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_177 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_177 vgnd vpwr scs8hd_decap_4
XFILLER_2_6 vgnd vpwr scs8hd_decap_12
XFILLER_11_11 vpwr vgnd scs8hd_fill_2
XFILLER_11_22 vpwr vgnd scs8hd_fill_2
XFILLER_14_100 vpwr vgnd scs8hd_fill_2
X_176_ _176_/HI _176_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__123__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_22_21 vgnd vpwr scs8hd_decap_4
XFILLER_22_32 vgnd vpwr scs8hd_fill_1
XFILLER_22_65 vpwr vgnd scs8hd_fill_2
XFILLER_22_87 vgnd vpwr scs8hd_decap_3
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_203 vpwr vgnd scs8hd_fill_2
XFILLER_19_258 vgnd vpwr scs8hd_decap_4
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_162 vpwr vgnd scs8hd_fill_2
X_159_ _074_/A _159_/B _082_/C _159_/Y vgnd vpwr scs8hd_nor3_4
Xmux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__134__A _108_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _174_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vgnd vpwr scs8hd_decap_6
XFILLER_16_228 vgnd vpwr scs8hd_decap_8
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_6
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_250 vgnd vpwr scs8hd_decap_4
XFILLER_17_87 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_242 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_53 vgnd vpwr scs8hd_fill_1
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XANTENNA__131__B _128_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_44 vgnd vpwr scs8hd_decap_8
XFILLER_14_88 vpwr vgnd scs8hd_fill_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _148_/Y mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _108_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_131 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_17_164 vpwr vgnd scs8hd_fill_2
XFILLER_32_145 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_123 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _178_/HI mem_right_track_8.LATCH_2_.latch/Q
+ mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_78 vpwr vgnd scs8hd_fill_2
XFILLER_14_167 vgnd vpwr scs8hd_decap_4
X_175_ _175_/HI _175_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_7 vpwr vgnd scs8hd_fill_2
XFILLER_37_259 vpwr vgnd scs8hd_fill_2
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
XFILLER_28_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_44 vgnd vpwr scs8hd_decap_4
XFILLER_27_270 vgnd vpwr scs8hd_decap_6
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
X_089_ _088_/X _090_/B vgnd vpwr scs8hd_buf_1
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
X_158_ _150_/C _159_/B vgnd vpwr scs8hd_buf_1
XANTENNA__134__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_4
XANTENNA__150__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_22 vpwr vgnd scs8hd_fill_2
XFILLER_17_55 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XFILLER_30_254 vgnd vpwr scs8hd_decap_12
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_254 vpwr vgnd scs8hd_fill_2
XFILLER_21_265 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_65 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _098_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _143_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_6 vgnd vpwr scs8hd_decap_8
Xmem_top_track_2.LATCH_1_.latch data_in _143_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_140 vgnd vpwr scs8hd_decap_12
XFILLER_30_22 vgnd vpwr scs8hd_decap_8
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_3
XFILLER_29_151 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _177_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__B _136_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_272 vgnd vpwr scs8hd_decap_3
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_25_77 vgnd vpwr scs8hd_decap_4
XFILLER_25_22 vpwr vgnd scs8hd_fill_2
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XFILLER_32_157 vgnd vpwr scs8hd_decap_6
XANTENNA__137__B _136_/X vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_146 vpwr vgnd scs8hd_fill_2
XFILLER_23_135 vpwr vgnd scs8hd_fill_2
XFILLER_23_113 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vgnd vpwr scs8hd_decap_4
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_146 vgnd vpwr scs8hd_fill_1
X_174_ _174_/HI _174_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__148__A _148_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_161 vpwr vgnd scs8hd_fill_2
XFILLER_11_116 vgnd vpwr scs8hd_decap_4
XFILLER_11_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _108_/A _157_/B _157_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_142 vpwr vgnd scs8hd_fill_2
XFILLER_10_193 vpwr vgnd scs8hd_fill_2
XANTENNA__150__B address[3] vgnd vpwr scs8hd_diode_2
X_088_ address[1] address[2] _082_/C _088_/X vgnd vpwr scs8hd_or3_4
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_263 vgnd vpwr scs8hd_decap_12
XFILLER_18_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_45 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_99 vgnd vpwr scs8hd_decap_12
XFILLER_33_33 vgnd vpwr scs8hd_decap_12
XFILLER_33_22 vpwr vgnd scs8hd_fill_2
XFILLER_33_11 vpwr vgnd scs8hd_fill_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_274 vgnd vpwr scs8hd_fill_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _182_/HI _144_/Y mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_200 vgnd vpwr scs8hd_fill_1
X_209_ _209_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_30_266 vgnd vpwr scs8hd_decap_8
XANTENNA__161__A _095_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _145_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_222 vpwr vgnd scs8hd_fill_2
XANTENNA__071__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_28_22 vgnd vpwr scs8hd_decap_6
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_4
XFILLER_8_226 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__156__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_152 vgnd vpwr scs8hd_fill_1
XANTENNA__066__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_29_196 vpwr vgnd scs8hd_fill_2
XFILLER_29_174 vgnd vpwr scs8hd_decap_3
XFILLER_4_240 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_80 vgnd vpwr scs8hd_decap_8
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
X_190_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_199 vpwr vgnd scs8hd_fill_2
XFILLER_25_56 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XANTENNA__153__B _157_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 chany_top_in[6] mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_169 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _147_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_69 vgnd vpwr scs8hd_decap_3
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_125 vgnd vpwr scs8hd_fill_1
X_173_ _173_/HI _173_/LO vgnd vpwr scs8hd_conb_1
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__164__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_228 vgnd vpwr scs8hd_decap_4
XFILLER_28_206 vgnd vpwr scs8hd_decap_8
XANTENNA__074__A _074_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_239 vgnd vpwr scs8hd_decap_3
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_6_154 vpwr vgnd scs8hd_fill_2
XFILLER_10_150 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_087_ _090_/A _087_/B _087_/Y vgnd vpwr scs8hd_nor2_4
X_156_ _106_/A _157_/B _156_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_7 vgnd vpwr scs8hd_decap_12
XANTENNA__150__C _150_/C vgnd vpwr scs8hd_diode_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XFILLER_25_209 vpwr vgnd scs8hd_fill_2
XANTENNA__159__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_275 vpwr vgnd scs8hd_fill_2
XFILLER_33_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _152_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_68 vpwr vgnd scs8hd_fill_2
XFILLER_33_45 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _146_/Y mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_231 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_208_ chanx_right_in[4] chany_top_out[2] vgnd vpwr scs8hd_buf_2
X_139_ _113_/A _136_/X _139_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XFILLER_9_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _173_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XANTENNA__071__B _163_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_45 vgnd vpwr scs8hd_decap_8
XFILLER_8_205 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XFILLER_8_238 vgnd vpwr scs8hd_decap_12
XANTENNA__172__A _107_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _182_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__156__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_57 vpwr vgnd scs8hd_fill_2
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_11 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_252 vgnd vpwr scs8hd_decap_12
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__167__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_167 vpwr vgnd scs8hd_fill_2
XFILLER_26_145 vgnd vpwr scs8hd_decap_8
XFILLER_26_112 vgnd vpwr scs8hd_decap_4
XFILLER_25_35 vpwr vgnd scs8hd_fill_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A address[0] vgnd vpwr scs8hd_diode_2
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_17_101 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vpwr vgnd scs8hd_fill_2
XFILLER_17_189 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_11_ mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _153_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_15 vgnd vpwr scs8hd_decap_4
XFILLER_11_26 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
X_172_ _107_/A _169_/B _172_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__164__B _163_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_107 vgnd vpwr scs8hd_decap_3
XFILLER_20_129 vgnd vpwr scs8hd_decap_6
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XANTENNA__074__B _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_69 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A _090_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
XFILLER_19_218 vpwr vgnd scs8hd_fill_2
XFILLER_6_166 vpwr vgnd scs8hd_fill_2
X_086_ _085_/X _087_/B vgnd vpwr scs8hd_buf_1
X_155_ _114_/A _157_/B _155_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_240 vgnd vpwr scs8hd_decap_4
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_57 vgnd vpwr scs8hd_decap_4
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_254 vgnd vpwr scs8hd_fill_1
XFILLER_24_232 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_169 vgnd vpwr scs8hd_decap_12
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _171_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_207_ chanx_right_in[5] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_30_224 vgnd vpwr scs8hd_decap_12
XFILLER_15_254 vpwr vgnd scs8hd_fill_2
XFILLER_15_265 vpwr vgnd scs8hd_fill_2
X_138_ _112_/A _136_/X _138_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__C _082_/C vgnd vpwr scs8hd_diode_2
X_069_ _152_/A _111_/A vgnd vpwr scs8hd_buf_1
XFILLER_24_3 vgnd vpwr scs8hd_decap_4
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XFILLER_12_202 vgnd vpwr scs8hd_decap_4
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__172__B _169_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__082__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_29_132 vgnd vpwr scs8hd_decap_4
XFILLER_4_264 vgnd vpwr scs8hd_decap_8
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__167__B _169_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _210_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_135 vgnd vpwr scs8hd_fill_1
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_2_18 vgnd vpwr scs8hd_decap_12
XFILLER_32_149 vgnd vpwr scs8hd_decap_4
XFILLER_17_168 vpwr vgnd scs8hd_fill_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_31_193 vpwr vgnd scs8hd_fill_2
XFILLER_11_38 vgnd vpwr scs8hd_decap_12
XANTENNA__088__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_149 vpwr vgnd scs8hd_fill_2
X_171_ _090_/B _169_/B _171_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XANTENNA__164__C _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_193 vgnd vpwr scs8hd_decap_4
XFILLER_9_197 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_15_ mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_11_108 vpwr vgnd scs8hd_fill_2
XFILLER_22_48 vgnd vpwr scs8hd_fill_1
XANTENNA__090__B _090_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_101 vgnd vpwr scs8hd_decap_3
X_154_ _113_/A _157_/B _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_163 vpwr vgnd scs8hd_fill_2
XFILLER_10_174 vpwr vgnd scs8hd_fill_2
X_085_ _085_/A address[2] _085_/C _085_/X vgnd vpwr scs8hd_or3_4
XFILLER_26_7 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__159__C _082_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__191__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_26 vpwr vgnd scs8hd_fill_2
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__085__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_159 vgnd vpwr scs8hd_decap_8
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _108_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_206_ _206_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_30_236 vgnd vpwr scs8hd_decap_3
X_137_ _111_/A _136_/X _137_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_068_ _067_/X _152_/A vgnd vpwr scs8hd_buf_1
XFILLER_17_3 vgnd vpwr scs8hd_decap_4
XANTENNA__186__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_60 vgnd vpwr scs8hd_fill_1
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
XFILLER_21_258 vpwr vgnd scs8hd_fill_2
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _184_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XFILLER_28_69 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _074_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_240 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__082__C _082_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_210 vgnd vpwr scs8hd_decap_4
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _148_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _188_/A vgnd vpwr scs8hd_inv_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _107_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_147 vpwr vgnd scs8hd_fill_2
XFILLER_40_183 vgnd vpwr scs8hd_decap_12
XFILLER_32_139 vgnd vpwr scs8hd_decap_3
XFILLER_15_92 vpwr vgnd scs8hd_fill_2
XFILLER_31_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__194__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_23_139 vgnd vpwr scs8hd_decap_4
XFILLER_23_117 vgnd vpwr scs8hd_decap_3
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _076_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_172 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__088__B address[2] vgnd vpwr scs8hd_diode_2
X_170_ _087_/B _169_/B _170_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_128 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_143 vgnd vpwr scs8hd_decap_3
XFILLER_9_165 vgnd vpwr scs8hd_fill_1
XANTENNA__164__D _085_/C vgnd vpwr scs8hd_diode_2
XANTENNA__189__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A _080_/B vgnd vpwr scs8hd_diode_2
X_153_ _112_/A _157_/B _153_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_120 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _144_/A mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_6_179 vgnd vpwr scs8hd_decap_6
XFILLER_6_146 vgnd vpwr scs8hd_decap_6
XFILLER_10_197 vgnd vpwr scs8hd_decap_4
XFILLER_12_60 vgnd vpwr scs8hd_decap_12
X_084_ _090_/A _101_/A _084_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_245 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_201 vpwr vgnd scs8hd_fill_2
XFILLER_17_49 vgnd vpwr scs8hd_decap_4
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _177_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__085__C _085_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_205_ chanx_left_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
X_136_ _135_/X _136_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_067_ address[1] _067_/B _082_/C _067_/X vgnd vpwr scs8hd_or3_4
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_83 vpwr vgnd scs8hd_fill_2
XFILLER_9_94 vpwr vgnd scs8hd_fill_2
XFILLER_21_226 vpwr vgnd scs8hd_fill_2
XANTENNA__096__B _095_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_226 vpwr vgnd scs8hd_fill_2
XFILLER_8_219 vgnd vpwr scs8hd_fill_1
XFILLER_12_237 vgnd vpwr scs8hd_decap_8
XFILLER_12_248 vgnd vpwr scs8hd_decap_12
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
X_119_ address[4] address[3] address[5] _135_/D _119_/X vgnd vpwr scs8hd_or4_4
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_30_49 vgnd vpwr scs8hd_fill_1
XFILLER_29_112 vgnd vpwr scs8hd_fill_1
XFILLER_20_71 vpwr vgnd scs8hd_fill_2
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XFILLER_29_91 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XFILLER_9_6 vpwr vgnd scs8hd_fill_2
XFILLER_32_107 vgnd vpwr scs8hd_decap_12
XFILLER_40_195 vgnd vpwr scs8hd_decap_12
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XANTENNA__088__C _082_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _176_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _144_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_111 vpwr vgnd scs8hd_fill_2
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_17 vpwr vgnd scs8hd_fill_2
XFILLER_27_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_254 vpwr vgnd scs8hd_fill_2
XFILLER_8_19 vgnd vpwr scs8hd_decap_12
XFILLER_6_158 vgnd vpwr scs8hd_fill_1
XFILLER_10_132 vgnd vpwr scs8hd_decap_4
XFILLER_12_50 vgnd vpwr scs8hd_fill_1
XFILLER_12_72 vgnd vpwr scs8hd_fill_1
X_083_ _082_/X _101_/A vgnd vpwr scs8hd_buf_1
X_152_ _152_/A _157_/B _152_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_246 vpwr vgnd scs8hd_fill_2
XFILLER_24_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_106 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_204_ chanx_left_in[4] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_15_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_066_ address[0] _082_/C vgnd vpwr scs8hd_inv_8
X_135_ _163_/A address[3] address[5] _135_/D _135_/X vgnd vpwr scs8hd_or4_4
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_9_40 vgnd vpwr scs8hd_decap_12
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_21_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_271 vgnd vpwr scs8hd_decap_4
XFILLER_18_93 vgnd vpwr scs8hd_decap_4
X_118_ _149_/A _073_/B _135_/D vgnd vpwr scs8hd_or2_4
XFILLER_38_157 vgnd vpwr scs8hd_decap_12
XFILLER_22_3 vgnd vpwr scs8hd_decap_3
XFILLER_14_29 vpwr vgnd scs8hd_fill_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_7_ mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_223 vpwr vgnd scs8hd_fill_2
XFILLER_26_127 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_39 vpwr vgnd scs8hd_fill_2
XPHY_39 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_119 vgnd vpwr scs8hd_decap_12
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_31_60 vgnd vpwr scs8hd_fill_1
XFILLER_16_171 vgnd vpwr scs8hd_decap_6
XFILLER_39_241 vgnd vpwr scs8hd_decap_3
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
XFILLER_22_185 vpwr vgnd scs8hd_fill_2
XFILLER_26_93 vgnd vpwr scs8hd_decap_6
XFILLER_9_123 vgnd vpwr scs8hd_decap_4
XFILLER_13_152 vpwr vgnd scs8hd_fill_2
XFILLER_13_174 vgnd vpwr scs8hd_decap_3
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
XFILLER_6_126 vgnd vpwr scs8hd_decap_3
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
X_151_ _151_/A _157_/B vgnd vpwr scs8hd_buf_1
X_082_ _085_/A address[2] _082_/C _082_/X vgnd vpwr scs8hd_or3_4
XFILLER_18_244 vgnd vpwr scs8hd_fill_1
XFILLER_17_18 vpwr vgnd scs8hd_fill_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_258 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _173_/HI mem_left_track_1.LATCH_2_.latch/Q
+ mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_118 vgnd vpwr scs8hd_decap_4
XFILLER_15_203 vpwr vgnd scs8hd_fill_2
X_203_ _203_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_30_206 vgnd vpwr scs8hd_decap_8
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
XFILLER_15_258 vgnd vpwr scs8hd_decap_4
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _143_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_065_ address[2] _067_/B vgnd vpwr scs8hd_inv_8
X_134_ _108_/A _128_/X _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_52 vgnd vpwr scs8hd_decap_8
XFILLER_9_74 vgnd vpwr scs8hd_decap_6
XFILLER_28_28 vgnd vpwr scs8hd_fill_1
XFILLER_12_206 vgnd vpwr scs8hd_fill_1
XFILLER_18_72 vgnd vpwr scs8hd_fill_1
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_117_ enable _149_/A vgnd vpwr scs8hd_inv_8
XFILLER_11_261 vgnd vpwr scs8hd_decap_12
XFILLER_38_169 vgnd vpwr scs8hd_decap_12
XFILLER_15_3 vgnd vpwr scs8hd_decap_3
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _126_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_37_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_71 vgnd vpwr scs8hd_decap_3
XFILLER_28_191 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_18 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XFILLER_15_84 vpwr vgnd scs8hd_fill_2
XFILLER_17_128 vpwr vgnd scs8hd_fill_2
XFILLER_31_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_197 vpwr vgnd scs8hd_fill_2
XFILLER_31_131 vgnd vpwr scs8hd_fill_1
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_36_17 vgnd vpwr scs8hd_decap_12
XFILLER_22_131 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_3_ mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_72 vgnd vpwr scs8hd_fill_1
XFILLER_9_157 vpwr vgnd scs8hd_fill_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_98 vgnd vpwr scs8hd_decap_6
XFILLER_27_212 vpwr vgnd scs8hd_fill_2
X_150_ address[4] address[3] _150_/C _151_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_138 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vgnd vpwr scs8hd_decap_3
XFILLER_10_167 vpwr vgnd scs8hd_fill_2
XFILLER_10_178 vgnd vpwr scs8hd_decap_4
XFILLER_12_96 vgnd vpwr scs8hd_decap_3
X_081_ address[1] _085_/A vgnd vpwr scs8hd_inv_8
XFILLER_33_259 vpwr vgnd scs8hd_fill_2
XFILLER_5_182 vgnd vpwr scs8hd_fill_1
XFILLER_33_29 vpwr vgnd scs8hd_fill_2
XFILLER_33_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__200__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
X_202_ _202_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_23_73 vpwr vgnd scs8hd_fill_2
X_133_ _106_/A _128_/X _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_51 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _147_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_18 vpwr vgnd scs8hd_fill_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
X_116_ _108_/A _112_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_273 vgnd vpwr scs8hd_decap_4
XANTENNA__105__A _090_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XFILLER_29_115 vgnd vpwr scs8hd_decap_4
XFILLER_20_41 vgnd vpwr scs8hd_decap_3
XFILLER_28_170 vgnd vpwr scs8hd_decap_6
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_0_.latch data_in _146_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_184 vpwr vgnd scs8hd_fill_2
XFILLER_25_162 vpwr vgnd scs8hd_fill_2
XFILLER_15_96 vpwr vgnd scs8hd_fill_2
XFILLER_31_73 vgnd vpwr scs8hd_decap_3
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__102__B _106_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_110 vgnd vpwr scs8hd_fill_1
XFILLER_31_176 vgnd vpwr scs8hd_fill_1
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_29 vpwr vgnd scs8hd_fill_2
XFILLER_22_154 vgnd vpwr scs8hd_decap_3
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vpwr vgnd scs8hd_fill_2
XFILLER_26_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_13_143 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_10_124 vpwr vgnd scs8hd_fill_2
X_080_ _090_/A _080_/B _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _201_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_202 vgnd vpwr scs8hd_decap_4
XFILLER_18_235 vpwr vgnd scs8hd_fill_2
XANTENNA__108__A _108_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_161 vpwr vgnd scs8hd_fill_2
XFILLER_5_150 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_227 vpwr vgnd scs8hd_fill_2
X_201_ _201_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _152_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_96 vpwr vgnd scs8hd_fill_2
X_132_ _114_/A _128_/X _132_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _193_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_9_10 vgnd vpwr scs8hd_decap_4
XFILLER_9_87 vpwr vgnd scs8hd_fill_2
XFILLER_9_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_30 vgnd vpwr scs8hd_fill_1
XFILLER_18_52 vgnd vpwr scs8hd_fill_1
X_115_ _106_/A _112_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XFILLER_7_201 vgnd vpwr scs8hd_fill_1
XFILLER_38_116 vgnd vpwr scs8hd_decap_12
XFILLER_38_105 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A left_bottom_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__121__A _111_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _143_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_95 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_26_108 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _170_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_3 vgnd vpwr scs8hd_decap_4
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_53 vgnd vpwr scs8hd_fill_1
XFILLER_0_262 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_130 vgnd vpwr scs8hd_decap_3
XFILLER_16_152 vgnd vpwr scs8hd_fill_1
XFILLER_16_163 vpwr vgnd scs8hd_fill_2
XFILLER_31_155 vpwr vgnd scs8hd_fill_2
XFILLER_31_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

