magic
tech sky130A
magscale 1 2
timestamp 1609017204
<< locali >>
rect 12357 20247 12391 20349
rect 13737 20247 13771 20349
rect 14381 20315 14415 20553
rect 15301 20247 15335 20417
rect 16497 20247 16531 20417
rect 17601 20247 17635 20349
rect 20729 19873 20821 19907
rect 9873 19703 9907 19805
rect 20729 19703 20763 19873
rect 8493 19159 8527 19329
rect 18061 18683 18095 18921
rect 12265 18275 12299 18377
rect 14197 18071 14231 18377
rect 12173 16983 12207 17085
rect 16129 16439 16163 16609
rect 19993 14943 20027 15113
rect 19717 14263 19751 14569
rect 17785 11611 17819 11713
rect 8769 9367 8803 9605
rect 12817 8891 12851 8993
rect 16129 8823 16163 8993
rect 9505 7939 9539 8041
rect 9413 7735 9447 7837
rect 8217 7191 8251 7497
rect 12173 6103 12207 6341
rect 16129 6171 16163 6409
rect 17233 5559 17267 5661
rect 19533 5015 19567 5185
rect 9873 3383 9907 3485
rect 12265 2907 12299 3077
rect 15669 1887 15703 2057
<< viali >>
rect 11161 20553 11195 20587
rect 13001 20553 13035 20587
rect 14381 20553 14415 20587
rect 14657 20553 14691 20587
rect 17877 20553 17911 20587
rect 19349 20553 19383 20587
rect 19901 20553 19935 20587
rect 11713 20485 11747 20519
rect 14105 20485 14139 20519
rect 10333 20417 10367 20451
rect 10977 20349 11011 20383
rect 11529 20349 11563 20383
rect 12357 20349 12391 20383
rect 13369 20349 13403 20383
rect 13737 20349 13771 20383
rect 13921 20349 13955 20383
rect 9965 20281 9999 20315
rect 16773 20485 16807 20519
rect 17325 20485 17359 20519
rect 21189 20485 21223 20519
rect 15301 20417 15335 20451
rect 14473 20349 14507 20383
rect 14381 20281 14415 20315
rect 15025 20281 15059 20315
rect 9321 20213 9355 20247
rect 10701 20213 10735 20247
rect 12173 20213 12207 20247
rect 12357 20213 12391 20247
rect 12725 20213 12759 20247
rect 13553 20213 13587 20247
rect 13737 20213 13771 20247
rect 16497 20417 16531 20451
rect 15485 20349 15519 20383
rect 16037 20349 16071 20383
rect 16589 20349 16623 20383
rect 17141 20349 17175 20383
rect 17601 20349 17635 20383
rect 17693 20349 17727 20383
rect 18613 20349 18647 20383
rect 19165 20349 19199 20383
rect 19717 20349 19751 20383
rect 20545 20349 20579 20383
rect 15301 20213 15335 20247
rect 15669 20213 15703 20247
rect 16221 20213 16255 20247
rect 16497 20213 16531 20247
rect 17601 20213 17635 20247
rect 18797 20213 18831 20247
rect 20729 20213 20763 20247
rect 8953 20009 8987 20043
rect 13461 20009 13495 20043
rect 14289 20009 14323 20043
rect 14841 20009 14875 20043
rect 16497 20009 16531 20043
rect 17049 20009 17083 20043
rect 18061 20009 18095 20043
rect 18981 20009 19015 20043
rect 21189 19941 21223 19975
rect 10425 19873 10459 19907
rect 11161 19873 11195 19907
rect 11428 19873 11462 19907
rect 14105 19873 14139 19907
rect 14657 19873 14691 19907
rect 15669 19873 15703 19907
rect 16313 19873 16347 19907
rect 16865 19873 16899 19907
rect 17877 19873 17911 19907
rect 18429 19873 18463 19907
rect 18797 19873 18831 19907
rect 19717 19873 19751 19907
rect 20269 19873 20303 19907
rect 20821 19873 20855 19907
rect 20913 19873 20947 19907
rect 9873 19805 9907 19839
rect 10517 19805 10551 19839
rect 10609 19805 10643 19839
rect 13553 19805 13587 19839
rect 13737 19805 13771 19839
rect 15761 19805 15795 19839
rect 15853 19805 15887 19839
rect 17417 19805 17451 19839
rect 20453 19737 20487 19771
rect 9229 19669 9263 19703
rect 9781 19669 9815 19703
rect 9873 19669 9907 19703
rect 10057 19669 10091 19703
rect 12541 19669 12575 19703
rect 13093 19669 13127 19703
rect 15301 19669 15335 19703
rect 19349 19669 19383 19703
rect 19901 19669 19935 19703
rect 20729 19669 20763 19703
rect 11621 19465 11655 19499
rect 13829 19465 13863 19499
rect 15761 19465 15795 19499
rect 15485 19397 15519 19431
rect 8493 19329 8527 19363
rect 9321 19329 9355 19363
rect 11897 19329 11931 19363
rect 16313 19329 16347 19363
rect 17233 19329 17267 19363
rect 18337 19329 18371 19363
rect 20269 19329 20303 19363
rect 8309 19193 8343 19227
rect 9689 19261 9723 19295
rect 10241 19261 10275 19295
rect 12449 19261 12483 19295
rect 12705 19261 12739 19295
rect 14105 19261 14139 19295
rect 14361 19261 14395 19295
rect 16129 19261 16163 19295
rect 16957 19261 16991 19295
rect 18061 19261 18095 19295
rect 18889 19261 18923 19295
rect 19165 19261 19199 19295
rect 19901 19261 19935 19295
rect 10508 19193 10542 19227
rect 16221 19193 16255 19227
rect 8493 19125 8527 19159
rect 8677 19125 8711 19159
rect 9045 19125 9079 19159
rect 21281 19125 21315 19159
rect 11069 18921 11103 18955
rect 11805 18921 11839 18955
rect 12725 18921 12759 18955
rect 13553 18921 13587 18955
rect 14657 18921 14691 18955
rect 17325 18921 17359 18955
rect 17877 18921 17911 18955
rect 18061 18921 18095 18955
rect 15752 18853 15786 18887
rect 8861 18785 8895 18819
rect 9689 18785 9723 18819
rect 9956 18785 9990 18819
rect 11713 18785 11747 18819
rect 13369 18785 13403 18819
rect 14565 18785 14599 18819
rect 17141 18785 17175 18819
rect 17693 18785 17727 18819
rect 11897 18717 11931 18751
rect 12817 18717 12851 18751
rect 12909 18717 12943 18751
rect 14841 18717 14875 18751
rect 15485 18717 15519 18751
rect 19165 18853 19199 18887
rect 18245 18785 18279 18819
rect 20269 18785 20303 18819
rect 20913 18785 20947 18819
rect 19257 18717 19291 18751
rect 19441 18717 19475 18751
rect 11345 18649 11379 18683
rect 14197 18649 14231 18683
rect 18061 18649 18095 18683
rect 19809 18649 19843 18683
rect 8217 18581 8251 18615
rect 8493 18581 8527 18615
rect 9321 18581 9355 18615
rect 12357 18581 12391 18615
rect 16865 18581 16899 18615
rect 18429 18581 18463 18615
rect 18797 18581 18831 18615
rect 20453 18581 20487 18615
rect 21097 18581 21131 18615
rect 7113 18377 7147 18411
rect 12081 18377 12115 18411
rect 12265 18377 12299 18411
rect 7481 18309 7515 18343
rect 10057 18309 10091 18343
rect 14197 18377 14231 18411
rect 15669 18377 15703 18411
rect 16221 18377 16255 18411
rect 13921 18309 13955 18343
rect 8125 18241 8159 18275
rect 12265 18241 12299 18275
rect 13001 18241 13035 18275
rect 7849 18173 7883 18207
rect 8677 18173 8711 18207
rect 11253 18173 11287 18207
rect 12817 18173 12851 18207
rect 12909 18173 12943 18207
rect 13737 18173 13771 18207
rect 7941 18105 7975 18139
rect 8944 18105 8978 18139
rect 11529 18105 11563 18139
rect 16589 18309 16623 18343
rect 19717 18309 19751 18343
rect 17233 18241 17267 18275
rect 20269 18241 20303 18275
rect 14289 18173 14323 18207
rect 16037 18173 16071 18207
rect 16957 18173 16991 18207
rect 18061 18173 18095 18207
rect 20085 18173 20119 18207
rect 20821 18173 20855 18207
rect 14556 18105 14590 18139
rect 17601 18105 17635 18139
rect 18328 18105 18362 18139
rect 10333 18037 10367 18071
rect 10885 18037 10919 18071
rect 12449 18037 12483 18071
rect 14197 18037 14231 18071
rect 17049 18037 17083 18071
rect 19441 18037 19475 18071
rect 20177 18037 20211 18071
rect 21005 18037 21039 18071
rect 7113 17833 7147 17867
rect 9045 17833 9079 17867
rect 9689 17833 9723 17867
rect 11161 17833 11195 17867
rect 13829 17833 13863 17867
rect 17417 17833 17451 17867
rect 19349 17833 19383 17867
rect 20361 17833 20395 17867
rect 10149 17765 10183 17799
rect 13737 17765 13771 17799
rect 16304 17765 16338 17799
rect 17938 17765 17972 17799
rect 21189 17765 21223 17799
rect 7932 17697 7966 17731
rect 10057 17697 10091 17731
rect 11069 17697 11103 17731
rect 12173 17697 12207 17731
rect 14657 17697 14691 17731
rect 15301 17697 15335 17731
rect 16037 17697 16071 17731
rect 19717 17697 19751 17731
rect 20913 17697 20947 17731
rect 7665 17629 7699 17663
rect 10241 17629 10275 17663
rect 11253 17629 11287 17663
rect 12449 17629 12483 17663
rect 14013 17629 14047 17663
rect 15577 17629 15611 17663
rect 17693 17629 17727 17663
rect 19809 17629 19843 17663
rect 19901 17629 19935 17663
rect 19073 17561 19107 17595
rect 6745 17493 6779 17527
rect 10701 17493 10735 17527
rect 11805 17493 11839 17527
rect 13093 17493 13127 17527
rect 13369 17493 13403 17527
rect 14841 17493 14875 17527
rect 8401 17289 8435 17323
rect 9137 17289 9171 17323
rect 9505 17289 9539 17323
rect 11345 17289 11379 17323
rect 12449 17289 12483 17323
rect 16589 17289 16623 17323
rect 14289 17221 14323 17255
rect 14565 17221 14599 17255
rect 7021 17153 7055 17187
rect 10057 17153 10091 17187
rect 11805 17153 11839 17187
rect 11989 17153 12023 17187
rect 12909 17153 12943 17187
rect 15209 17153 15243 17187
rect 16129 17153 16163 17187
rect 17141 17153 17175 17187
rect 18337 17153 18371 17187
rect 20269 17153 20303 17187
rect 21097 17153 21131 17187
rect 9873 17085 9907 17119
rect 10517 17085 10551 17119
rect 11713 17085 11747 17119
rect 12173 17085 12207 17119
rect 12633 17085 12667 17119
rect 13176 17085 13210 17119
rect 18604 17085 18638 17119
rect 20085 17085 20119 17119
rect 20821 17085 20855 17119
rect 7288 17017 7322 17051
rect 9965 17017 9999 17051
rect 10793 17017 10827 17051
rect 15025 17017 15059 17051
rect 6469 16949 6503 16983
rect 8861 16949 8895 16983
rect 12173 16949 12207 16983
rect 14933 16949 14967 16983
rect 15577 16949 15611 16983
rect 15945 16949 15979 16983
rect 16037 16949 16071 16983
rect 16957 16949 16991 16983
rect 17049 16949 17083 16983
rect 17601 16949 17635 16983
rect 19717 16949 19751 16983
rect 5917 16745 5951 16779
rect 7021 16745 7055 16779
rect 10333 16745 10367 16779
rect 12173 16745 12207 16779
rect 13829 16745 13863 16779
rect 14105 16745 14139 16779
rect 14473 16745 14507 16779
rect 14565 16745 14599 16779
rect 15301 16745 15335 16779
rect 17141 16745 17175 16779
rect 18153 16745 18187 16779
rect 18521 16745 18555 16779
rect 21097 16745 21131 16779
rect 6653 16677 6687 16711
rect 12694 16677 12728 16711
rect 15669 16677 15703 16711
rect 20269 16677 20303 16711
rect 7297 16609 7331 16643
rect 7564 16609 7598 16643
rect 10517 16609 10551 16643
rect 10793 16609 10827 16643
rect 11060 16609 11094 16643
rect 16129 16609 16163 16643
rect 17049 16609 17083 16643
rect 17969 16609 18003 16643
rect 18889 16609 18923 16643
rect 19993 16609 20027 16643
rect 20913 16609 20947 16643
rect 12449 16541 12483 16575
rect 14749 16541 14783 16575
rect 15761 16541 15795 16575
rect 15853 16541 15887 16575
rect 17233 16541 17267 16575
rect 18981 16541 19015 16575
rect 19073 16541 19107 16575
rect 19533 16541 19567 16575
rect 6285 16405 6319 16439
rect 8677 16405 8711 16439
rect 9321 16405 9355 16439
rect 9965 16405 9999 16439
rect 16129 16405 16163 16439
rect 16313 16405 16347 16439
rect 16681 16405 16715 16439
rect 8217 16201 8251 16235
rect 9873 16201 9907 16235
rect 12449 16201 12483 16235
rect 15117 16201 15151 16235
rect 18705 16201 18739 16235
rect 19901 16201 19935 16235
rect 11529 16133 11563 16167
rect 16129 16133 16163 16167
rect 8493 16065 8527 16099
rect 12081 16065 12115 16099
rect 13093 16065 13127 16099
rect 13461 16065 13495 16099
rect 15761 16065 15795 16099
rect 16589 16065 16623 16099
rect 16681 16065 16715 16099
rect 19165 16065 19199 16099
rect 19349 16065 19383 16099
rect 20453 16065 20487 16099
rect 6837 15997 6871 16031
rect 8760 15997 8794 16031
rect 10149 15997 10183 16031
rect 13728 15997 13762 16031
rect 16497 15997 16531 16031
rect 17141 15997 17175 16031
rect 18153 15997 18187 16031
rect 19073 15997 19107 16031
rect 20913 15997 20947 16031
rect 7104 15929 7138 15963
rect 10416 15929 10450 15963
rect 12909 15929 12943 15963
rect 17417 15929 17451 15963
rect 6469 15861 6503 15895
rect 12817 15861 12851 15895
rect 14841 15861 14875 15895
rect 15485 15861 15519 15895
rect 15577 15861 15611 15895
rect 18337 15861 18371 15895
rect 20269 15861 20303 15895
rect 20361 15861 20395 15895
rect 21097 15861 21131 15895
rect 6193 15657 6227 15691
rect 6561 15657 6595 15691
rect 6929 15657 6963 15691
rect 7297 15657 7331 15691
rect 8861 15657 8895 15691
rect 10241 15657 10275 15691
rect 11253 15657 11287 15691
rect 12265 15657 12299 15691
rect 15393 15657 15427 15691
rect 16405 15657 16439 15691
rect 16957 15657 16991 15691
rect 19165 15657 19199 15691
rect 19625 15657 19659 15691
rect 7757 15589 7791 15623
rect 10609 15589 10643 15623
rect 13645 15589 13679 15623
rect 16313 15589 16347 15623
rect 17776 15589 17810 15623
rect 7665 15521 7699 15555
rect 8769 15521 8803 15555
rect 11621 15521 11655 15555
rect 12633 15521 12667 15555
rect 14289 15521 14323 15555
rect 19533 15521 19567 15555
rect 20269 15521 20303 15555
rect 20913 15521 20947 15555
rect 7941 15453 7975 15487
rect 8953 15453 8987 15487
rect 9689 15453 9723 15487
rect 10701 15453 10735 15487
rect 10793 15453 10827 15487
rect 11713 15453 11747 15487
rect 11805 15453 11839 15487
rect 12725 15453 12759 15487
rect 12909 15453 12943 15487
rect 13737 15453 13771 15487
rect 13829 15453 13863 15487
rect 14749 15453 14783 15487
rect 16497 15453 16531 15487
rect 17509 15453 17543 15487
rect 19717 15453 19751 15487
rect 13277 15385 13311 15419
rect 15945 15385 15979 15419
rect 18889 15385 18923 15419
rect 5917 15317 5951 15351
rect 8401 15317 8435 15351
rect 20453 15317 20487 15351
rect 21097 15317 21131 15351
rect 6469 15113 6503 15147
rect 6929 15113 6963 15147
rect 7849 15113 7883 15147
rect 19993 15113 20027 15147
rect 20177 15113 20211 15147
rect 11437 15045 11471 15079
rect 13369 15045 13403 15079
rect 16037 15045 16071 15079
rect 17325 15045 17359 15079
rect 7481 14977 7515 15011
rect 9045 14977 9079 15011
rect 9781 14977 9815 15011
rect 13921 14977 13955 15011
rect 14657 14977 14691 15011
rect 16865 14977 16899 15011
rect 20729 14977 20763 15011
rect 9505 14909 9539 14943
rect 10333 14909 10367 14943
rect 10701 14909 10735 14943
rect 11621 14909 11655 14943
rect 12081 14909 12115 14943
rect 12449 14909 12483 14943
rect 17509 14909 17543 14943
rect 18245 14909 18279 14943
rect 18521 14909 18555 14943
rect 18788 14909 18822 14943
rect 19993 14909 20027 14943
rect 20637 14909 20671 14943
rect 8217 14841 8251 14875
rect 8861 14841 8895 14875
rect 12725 14841 12759 14875
rect 14902 14841 14936 14875
rect 16681 14841 16715 14875
rect 20545 14841 20579 14875
rect 8493 14773 8527 14807
rect 8953 14773 8987 14807
rect 11161 14773 11195 14807
rect 11897 14773 11931 14807
rect 13737 14773 13771 14807
rect 13829 14773 13863 14807
rect 16313 14773 16347 14807
rect 16773 14773 16807 14807
rect 18061 14773 18095 14807
rect 19901 14773 19935 14807
rect 21189 14773 21223 14807
rect 6837 14569 6871 14603
rect 7297 14569 7331 14603
rect 7941 14569 7975 14603
rect 8309 14569 8343 14603
rect 8677 14569 8711 14603
rect 8769 14569 8803 14603
rect 11805 14569 11839 14603
rect 12541 14569 12575 14603
rect 19717 14569 19751 14603
rect 19809 14569 19843 14603
rect 20177 14569 20211 14603
rect 9956 14501 9990 14535
rect 9689 14433 9723 14467
rect 11713 14433 11747 14467
rect 12909 14433 12943 14467
rect 13820 14433 13854 14467
rect 15669 14433 15703 14467
rect 16764 14433 16798 14467
rect 18409 14433 18443 14467
rect 8953 14365 8987 14399
rect 11897 14365 11931 14399
rect 13001 14365 13035 14399
rect 13185 14365 13219 14399
rect 13553 14365 13587 14399
rect 15761 14365 15795 14399
rect 15853 14365 15887 14399
rect 16497 14365 16531 14399
rect 18153 14365 18187 14399
rect 11069 14297 11103 14331
rect 20269 14501 20303 14535
rect 20913 14433 20947 14467
rect 20361 14365 20395 14399
rect 7665 14229 7699 14263
rect 11345 14229 11379 14263
rect 14933 14229 14967 14263
rect 15301 14229 15335 14263
rect 17877 14229 17911 14263
rect 19533 14229 19567 14263
rect 19717 14229 19751 14263
rect 21097 14229 21131 14263
rect 6469 14025 6503 14059
rect 7297 14025 7331 14059
rect 8033 14025 8067 14059
rect 8401 14025 8435 14059
rect 9781 14025 9815 14059
rect 14105 14025 14139 14059
rect 15209 14025 15243 14059
rect 17693 14025 17727 14059
rect 6929 13957 6963 13991
rect 8769 13957 8803 13991
rect 13829 13957 13863 13991
rect 16589 13957 16623 13991
rect 20637 13957 20671 13991
rect 10241 13889 10275 13923
rect 14565 13889 14599 13923
rect 14749 13889 14783 13923
rect 15853 13889 15887 13923
rect 17049 13889 17083 13923
rect 17233 13889 17267 13923
rect 18705 13889 18739 13923
rect 21189 13889 21223 13923
rect 7573 13821 7607 13855
rect 9045 13821 9079 13855
rect 9505 13821 9539 13855
rect 9965 13821 9999 13855
rect 10508 13821 10542 13855
rect 12449 13821 12483 13855
rect 12716 13821 12750 13855
rect 15669 13821 15703 13855
rect 16221 13821 16255 13855
rect 18521 13821 18555 13855
rect 19257 13821 19291 13855
rect 19524 13821 19558 13855
rect 20913 13821 20947 13855
rect 16957 13753 16991 13787
rect 11621 13685 11655 13719
rect 11897 13685 11931 13719
rect 14473 13685 14507 13719
rect 15577 13685 15611 13719
rect 18061 13685 18095 13719
rect 18429 13685 18463 13719
rect 8125 13481 8159 13515
rect 11437 13481 11471 13515
rect 11897 13481 11931 13515
rect 12909 13481 12943 13515
rect 14565 13481 14599 13515
rect 15393 13481 15427 13515
rect 15761 13481 15795 13515
rect 17785 13481 17819 13515
rect 7481 13413 7515 13447
rect 7757 13413 7791 13447
rect 9137 13413 9171 13447
rect 10048 13413 10082 13447
rect 14657 13413 14691 13447
rect 21189 13413 21223 13447
rect 8861 13345 8895 13379
rect 9781 13345 9815 13379
rect 11805 13345 11839 13379
rect 12817 13345 12851 13379
rect 13461 13345 13495 13379
rect 16405 13345 16439 13379
rect 16672 13345 16706 13379
rect 18429 13345 18463 13379
rect 19421 13345 19455 13379
rect 20913 13345 20947 13379
rect 7113 13277 7147 13311
rect 11989 13277 12023 13311
rect 13001 13277 13035 13311
rect 13645 13277 13679 13311
rect 14749 13277 14783 13311
rect 15853 13277 15887 13311
rect 16037 13277 16071 13311
rect 18521 13277 18555 13311
rect 18705 13277 18739 13311
rect 19165 13277 19199 13311
rect 12449 13209 12483 13243
rect 14197 13209 14231 13243
rect 8585 13141 8619 13175
rect 11161 13141 11195 13175
rect 18061 13141 18095 13175
rect 20545 13141 20579 13175
rect 7849 12937 7883 12971
rect 11069 12937 11103 12971
rect 13185 12937 13219 12971
rect 16957 12937 16991 12971
rect 20085 12937 20119 12971
rect 10057 12869 10091 12903
rect 20453 12869 20487 12903
rect 7389 12801 7423 12835
rect 10517 12801 10551 12835
rect 10701 12801 10735 12835
rect 11621 12801 11655 12835
rect 12725 12801 12759 12835
rect 13829 12801 13863 12835
rect 14749 12801 14783 12835
rect 16589 12801 16623 12835
rect 17601 12801 17635 12835
rect 18705 12801 18739 12835
rect 21005 12801 21039 12835
rect 8125 12733 8159 12767
rect 8392 12733 8426 12767
rect 11437 12733 11471 12767
rect 12449 12733 12483 12767
rect 15209 12733 15243 12767
rect 16313 12733 16347 12767
rect 17417 12733 17451 12767
rect 18972 12733 19006 12767
rect 20821 12733 20855 12767
rect 10425 12665 10459 12699
rect 13553 12665 13587 12699
rect 13645 12665 13679 12699
rect 14565 12665 14599 12699
rect 15485 12665 15519 12699
rect 17325 12665 17359 12699
rect 20913 12665 20947 12699
rect 9505 12597 9539 12631
rect 11529 12597 11563 12631
rect 14197 12597 14231 12631
rect 14657 12597 14691 12631
rect 15945 12597 15979 12631
rect 16405 12597 16439 12631
rect 18061 12597 18095 12631
rect 8125 12393 8159 12427
rect 10149 12393 10183 12427
rect 14565 12393 14599 12427
rect 16957 12393 16991 12427
rect 17417 12393 17451 12427
rect 18429 12393 18463 12427
rect 20545 12393 20579 12427
rect 21097 12393 21131 12427
rect 8493 12325 8527 12359
rect 11060 12325 11094 12359
rect 13737 12325 13771 12359
rect 17325 12325 17359 12359
rect 18521 12325 18555 12359
rect 10057 12257 10091 12291
rect 12817 12257 12851 12291
rect 13461 12257 13495 12291
rect 15301 12257 15335 12291
rect 15568 12257 15602 12291
rect 19165 12257 19199 12291
rect 19432 12257 19466 12291
rect 20913 12257 20947 12291
rect 9137 12189 9171 12223
rect 10241 12189 10275 12223
rect 10793 12189 10827 12223
rect 12909 12189 12943 12223
rect 13001 12189 13035 12223
rect 14657 12189 14691 12223
rect 14841 12189 14875 12223
rect 17601 12189 17635 12223
rect 18705 12189 18739 12223
rect 8861 12053 8895 12087
rect 9689 12053 9723 12087
rect 12173 12053 12207 12087
rect 12449 12053 12483 12087
rect 14197 12053 14231 12087
rect 16681 12053 16715 12087
rect 18061 12053 18095 12087
rect 11621 11849 11655 11883
rect 20177 11849 20211 11883
rect 20545 11849 20579 11883
rect 14381 11781 14415 11815
rect 16957 11781 16991 11815
rect 12449 11713 12483 11747
rect 13001 11713 13035 11747
rect 17601 11713 17635 11747
rect 17785 11713 17819 11747
rect 18245 11713 18279 11747
rect 21097 11713 21131 11747
rect 8585 11645 8619 11679
rect 8852 11645 8886 11679
rect 10241 11645 10275 11679
rect 14657 11645 14691 11679
rect 14913 11645 14947 11679
rect 16313 11645 16347 11679
rect 17325 11645 17359 11679
rect 18061 11645 18095 11679
rect 18797 11645 18831 11679
rect 10486 11577 10520 11611
rect 13268 11577 13302 11611
rect 17785 11577 17819 11611
rect 19042 11577 19076 11611
rect 21005 11577 21039 11611
rect 9965 11509 9999 11543
rect 11989 11509 12023 11543
rect 16037 11509 16071 11543
rect 17417 11509 17451 11543
rect 20913 11509 20947 11543
rect 8861 11305 8895 11339
rect 9689 11305 9723 11339
rect 10149 11305 10183 11339
rect 11253 11305 11287 11339
rect 14473 11305 14507 11339
rect 15301 11305 15335 11339
rect 18981 11305 19015 11339
rect 19257 11305 19291 11339
rect 19625 11305 19659 11339
rect 20913 11305 20947 11339
rect 10057 11237 10091 11271
rect 16190 11237 16224 11271
rect 11529 11169 11563 11203
rect 11796 11169 11830 11203
rect 13185 11169 13219 11203
rect 17868 11169 17902 11203
rect 10333 11101 10367 11135
rect 15945 11101 15979 11135
rect 17601 11101 17635 11135
rect 19717 11101 19751 11135
rect 19901 11101 19935 11135
rect 10701 11033 10735 11067
rect 12909 11033 12943 11067
rect 20545 11033 20579 11067
rect 9229 10965 9263 10999
rect 17325 10965 17359 10999
rect 8769 10761 8803 10795
rect 10793 10761 10827 10795
rect 14749 10761 14783 10795
rect 20729 10761 20763 10795
rect 9781 10693 9815 10727
rect 15761 10693 15795 10727
rect 10425 10625 10459 10659
rect 11345 10625 11379 10659
rect 13185 10625 13219 10659
rect 13369 10625 13403 10659
rect 14289 10625 14323 10659
rect 15301 10625 15335 10659
rect 16313 10625 16347 10659
rect 17601 10625 17635 10659
rect 18705 10625 18739 10659
rect 19349 10625 19383 10659
rect 9045 10557 9079 10591
rect 13093 10557 13127 10591
rect 14197 10557 14231 10591
rect 9321 10489 9355 10523
rect 10149 10489 10183 10523
rect 11253 10489 11287 10523
rect 12081 10489 12115 10523
rect 15209 10489 15243 10523
rect 16221 10489 16255 10523
rect 17325 10489 17359 10523
rect 19616 10489 19650 10523
rect 10241 10421 10275 10455
rect 11161 10421 11195 10455
rect 12725 10421 12759 10455
rect 13737 10421 13771 10455
rect 14105 10421 14139 10455
rect 15117 10421 15151 10455
rect 16129 10421 16163 10455
rect 16957 10421 16991 10455
rect 17417 10421 17451 10455
rect 18061 10421 18095 10455
rect 18429 10421 18463 10455
rect 18521 10421 18555 10455
rect 21281 10421 21315 10455
rect 8585 10217 8619 10251
rect 8861 10217 8895 10251
rect 13369 10217 13403 10251
rect 13645 10217 13679 10251
rect 14013 10217 14047 10251
rect 15669 10217 15703 10251
rect 17141 10217 17175 10251
rect 18521 10217 18555 10251
rect 19165 10217 19199 10251
rect 19717 10217 19751 10251
rect 10578 10149 10612 10183
rect 17509 10149 17543 10183
rect 17601 10149 17635 10183
rect 20177 10149 20211 10183
rect 11989 10081 12023 10115
rect 12256 10081 12290 10115
rect 15761 10081 15795 10115
rect 16313 10081 16347 10115
rect 16589 10081 16623 10115
rect 20085 10081 20119 10115
rect 10333 10013 10367 10047
rect 14105 10013 14139 10047
rect 14289 10013 14323 10047
rect 14749 10013 14783 10047
rect 15853 10013 15887 10047
rect 17785 10013 17819 10047
rect 18613 10013 18647 10047
rect 18705 10013 18739 10047
rect 20269 10013 20303 10047
rect 9229 9945 9263 9979
rect 11713 9945 11747 9979
rect 18153 9945 18187 9979
rect 21373 9945 21407 9979
rect 10057 9877 10091 9911
rect 15301 9877 15335 9911
rect 21005 9877 21039 9911
rect 8585 9673 8619 9707
rect 10609 9673 10643 9707
rect 10885 9673 10919 9707
rect 11897 9673 11931 9707
rect 19717 9673 19751 9707
rect 8769 9605 8803 9639
rect 12449 9605 12483 9639
rect 13277 9605 13311 9639
rect 14289 9605 14323 9639
rect 17693 9605 17727 9639
rect 11345 9537 11379 9571
rect 11437 9537 11471 9571
rect 13829 9537 13863 9571
rect 15209 9537 15243 9571
rect 16313 9537 16347 9571
rect 20913 9537 20947 9571
rect 9229 9469 9263 9503
rect 9496 9469 9530 9503
rect 12081 9469 12115 9503
rect 13001 9469 13035 9503
rect 16580 9469 16614 9503
rect 18337 9469 18371 9503
rect 20821 9469 20855 9503
rect 11253 9401 11287 9435
rect 13737 9401 13771 9435
rect 15025 9401 15059 9435
rect 15669 9401 15703 9435
rect 18582 9401 18616 9435
rect 8769 9333 8803 9367
rect 8861 9333 8895 9367
rect 12817 9333 12851 9367
rect 13645 9333 13679 9367
rect 14657 9333 14691 9367
rect 15117 9333 15151 9367
rect 19993 9333 20027 9367
rect 20361 9333 20395 9367
rect 20729 9333 20763 9367
rect 9965 9129 9999 9163
rect 10425 9129 10459 9163
rect 11897 9129 11931 9163
rect 13369 9129 13403 9163
rect 13921 9129 13955 9163
rect 14289 9129 14323 9163
rect 15301 9129 15335 9163
rect 16681 9129 16715 9163
rect 18521 9129 18555 9163
rect 18797 9129 18831 9163
rect 19165 9129 19199 9163
rect 20913 9129 20947 9163
rect 9321 9061 9355 9095
rect 11805 9061 11839 9095
rect 13277 9061 13311 9095
rect 17408 9061 17442 9095
rect 20177 9061 20211 9095
rect 8953 8993 8987 9027
rect 10793 8993 10827 9027
rect 10885 8993 10919 9027
rect 12633 8993 12667 9027
rect 12817 8993 12851 9027
rect 15669 8993 15703 9027
rect 16129 8993 16163 9027
rect 16873 8993 16907 9027
rect 17141 8993 17175 9027
rect 10977 8925 11011 8959
rect 11989 8925 12023 8959
rect 13553 8925 13587 8959
rect 14381 8925 14415 8959
rect 14473 8925 14507 8959
rect 15761 8925 15795 8959
rect 15945 8925 15979 8959
rect 11437 8857 11471 8891
rect 12817 8857 12851 8891
rect 19257 8925 19291 8959
rect 19349 8925 19383 8959
rect 20269 8925 20303 8959
rect 20453 8925 20487 8959
rect 12449 8789 12483 8823
rect 12909 8789 12943 8823
rect 16129 8789 16163 8823
rect 16405 8789 16439 8823
rect 19809 8789 19843 8823
rect 8401 8585 8435 8619
rect 10793 8585 10827 8619
rect 16037 8585 16071 8619
rect 17049 8585 17083 8619
rect 21097 8585 21131 8619
rect 13829 8517 13863 8551
rect 15761 8517 15795 8551
rect 17509 8517 17543 8551
rect 18705 8517 18739 8551
rect 9413 8449 9447 8483
rect 11713 8449 11747 8483
rect 12449 8449 12483 8483
rect 16497 8449 16531 8483
rect 16681 8449 16715 8483
rect 18061 8449 18095 8483
rect 19257 8449 19291 8483
rect 19717 8449 19751 8483
rect 8769 8381 8803 8415
rect 9680 8381 9714 8415
rect 11529 8381 11563 8415
rect 14381 8381 14415 8415
rect 14648 8381 14682 8415
rect 17233 8381 17267 8415
rect 19165 8381 19199 8415
rect 19984 8381 20018 8415
rect 9045 8313 9079 8347
rect 11437 8313 11471 8347
rect 12716 8313 12750 8347
rect 16405 8313 16439 8347
rect 19073 8313 19107 8347
rect 11069 8245 11103 8279
rect 9505 8041 9539 8075
rect 9689 8041 9723 8075
rect 11069 8041 11103 8075
rect 14197 8041 14231 8075
rect 14565 8041 14599 8075
rect 14657 8041 14691 8075
rect 16681 8041 16715 8075
rect 17601 8041 17635 8075
rect 18245 8041 18279 8075
rect 20545 8041 20579 8075
rect 8585 7973 8619 8007
rect 10793 7973 10827 8007
rect 11529 7973 11563 8007
rect 12532 7973 12566 8007
rect 18337 7973 18371 8007
rect 8861 7905 8895 7939
rect 9505 7905 9539 7939
rect 10057 7905 10091 7939
rect 11437 7905 11471 7939
rect 12265 7905 12299 7939
rect 15568 7905 15602 7939
rect 17141 7905 17175 7939
rect 19432 7905 19466 7939
rect 9137 7837 9171 7871
rect 9413 7837 9447 7871
rect 10149 7837 10183 7871
rect 10333 7837 10367 7871
rect 11621 7837 11655 7871
rect 14841 7837 14875 7871
rect 15301 7837 15335 7871
rect 18429 7837 18463 7871
rect 19165 7837 19199 7871
rect 20913 7837 20947 7871
rect 17877 7769 17911 7803
rect 8125 7701 8159 7735
rect 9413 7701 9447 7735
rect 13645 7701 13679 7735
rect 16957 7701 16991 7735
rect 7665 7497 7699 7531
rect 8217 7497 8251 7531
rect 11437 7497 11471 7531
rect 11989 7497 12023 7531
rect 14473 7497 14507 7531
rect 16313 7497 16347 7531
rect 8125 7429 8159 7463
rect 14013 7361 14047 7395
rect 17601 7361 17635 7395
rect 18613 7361 18647 7395
rect 20085 7361 20119 7395
rect 21097 7361 21131 7395
rect 8401 7293 8435 7327
rect 10057 7293 10091 7327
rect 10324 7293 10358 7327
rect 13829 7293 13863 7327
rect 14933 7293 14967 7327
rect 17417 7293 17451 7327
rect 18521 7293 18555 7327
rect 19165 7293 19199 7327
rect 19901 7293 19935 7327
rect 8668 7225 8702 7259
rect 13185 7225 13219 7259
rect 15200 7225 15234 7259
rect 16681 7225 16715 7259
rect 17325 7225 17359 7259
rect 18429 7225 18463 7259
rect 21005 7225 21039 7259
rect 8217 7157 8251 7191
rect 9781 7157 9815 7191
rect 12541 7157 12575 7191
rect 13461 7157 13495 7191
rect 13921 7157 13955 7191
rect 16957 7157 16991 7191
rect 18061 7157 18095 7191
rect 19533 7157 19567 7191
rect 19993 7157 20027 7191
rect 20545 7157 20579 7191
rect 20913 7157 20947 7191
rect 7573 6953 7607 6987
rect 8953 6953 8987 6987
rect 9689 6953 9723 6987
rect 10149 6953 10183 6987
rect 10701 6953 10735 6987
rect 11069 6953 11103 6987
rect 16497 6953 16531 6987
rect 16589 6953 16623 6987
rect 18889 6953 18923 6987
rect 20545 6953 20579 6987
rect 7941 6885 7975 6919
rect 11161 6885 11195 6919
rect 12716 6885 12750 6919
rect 17408 6885 17442 6919
rect 19432 6885 19466 6919
rect 9045 6817 9079 6851
rect 10057 6817 10091 6851
rect 11897 6817 11931 6851
rect 14473 6817 14507 6851
rect 15761 6817 15795 6851
rect 17141 6817 17175 6851
rect 19165 6817 19199 6851
rect 20913 6817 20947 6851
rect 8033 6749 8067 6783
rect 8217 6749 8251 6783
rect 9137 6749 9171 6783
rect 10241 6749 10275 6783
rect 11253 6749 11287 6783
rect 12449 6749 12483 6783
rect 14565 6749 14599 6783
rect 14657 6749 14691 6783
rect 16681 6749 16715 6783
rect 6929 6681 6963 6715
rect 8585 6681 8619 6715
rect 15301 6681 15335 6715
rect 7205 6613 7239 6647
rect 11713 6613 11747 6647
rect 13829 6613 13863 6647
rect 14105 6613 14139 6647
rect 16129 6613 16163 6647
rect 18521 6613 18555 6647
rect 7205 6409 7239 6443
rect 9321 6409 9355 6443
rect 10333 6409 10367 6443
rect 14381 6409 14415 6443
rect 16129 6409 16163 6443
rect 16313 6409 16347 6443
rect 18429 6409 18463 6443
rect 11345 6341 11379 6375
rect 12173 6341 12207 6375
rect 15301 6341 15335 6375
rect 9597 6273 9631 6307
rect 10885 6273 10919 6307
rect 11989 6273 12023 6307
rect 7941 6205 7975 6239
rect 8208 6205 8242 6239
rect 10793 6137 10827 6171
rect 11805 6137 11839 6171
rect 13921 6273 13955 6307
rect 15761 6273 15795 6307
rect 15945 6273 15979 6307
rect 12541 6205 12575 6239
rect 13829 6205 13863 6239
rect 18061 6341 18095 6375
rect 16773 6273 16807 6307
rect 16865 6273 16899 6307
rect 20913 6273 20947 6307
rect 21097 6273 21131 6307
rect 18797 6205 18831 6239
rect 19064 6205 19098 6239
rect 13737 6137 13771 6171
rect 15669 6137 15703 6171
rect 16129 6137 16163 6171
rect 16681 6137 16715 6171
rect 17325 6137 17359 6171
rect 20821 6137 20855 6171
rect 7665 6069 7699 6103
rect 10701 6069 10735 6103
rect 11713 6069 11747 6103
rect 12173 6069 12207 6103
rect 12909 6069 12943 6103
rect 13369 6069 13403 6103
rect 14749 6069 14783 6103
rect 20177 6069 20211 6103
rect 20453 6069 20487 6103
rect 8217 5865 8251 5899
rect 8585 5865 8619 5899
rect 9229 5865 9263 5899
rect 10057 5865 10091 5899
rect 14105 5865 14139 5899
rect 14565 5865 14599 5899
rect 15301 5865 15335 5899
rect 16773 5865 16807 5899
rect 18705 5865 18739 5899
rect 19533 5865 19567 5899
rect 20269 5865 20303 5899
rect 8861 5797 8895 5831
rect 10600 5797 10634 5831
rect 14473 5797 14507 5831
rect 15669 5797 15703 5831
rect 17570 5797 17604 5831
rect 20177 5797 20211 5831
rect 6469 5729 6503 5763
rect 7093 5729 7127 5763
rect 10333 5729 10367 5763
rect 12081 5729 12115 5763
rect 12449 5729 12483 5763
rect 12716 5729 12750 5763
rect 16681 5729 16715 5763
rect 20913 5729 20947 5763
rect 6837 5661 6871 5695
rect 14657 5661 14691 5695
rect 15761 5661 15795 5695
rect 15853 5661 15887 5695
rect 16865 5661 16899 5695
rect 17233 5661 17267 5695
rect 17325 5661 17359 5695
rect 18981 5661 19015 5695
rect 20361 5661 20395 5695
rect 11713 5525 11747 5559
rect 13829 5525 13863 5559
rect 16313 5525 16347 5559
rect 17233 5525 17267 5559
rect 19809 5525 19843 5559
rect 21097 5525 21131 5559
rect 8401 5321 8435 5355
rect 9137 5321 9171 5355
rect 9597 5321 9631 5355
rect 9965 5321 9999 5355
rect 12449 5321 12483 5355
rect 13001 5321 13035 5355
rect 15853 5321 15887 5355
rect 19441 5321 19475 5355
rect 8861 5253 8895 5287
rect 10241 5253 10275 5287
rect 10885 5185 10919 5219
rect 11805 5185 11839 5219
rect 13461 5185 13495 5219
rect 13645 5185 13679 5219
rect 19533 5185 19567 5219
rect 19717 5185 19751 5219
rect 11621 5117 11655 5151
rect 14473 5117 14507 5151
rect 16129 5117 16163 5151
rect 16396 5117 16430 5151
rect 18061 5117 18095 5151
rect 10609 5049 10643 5083
rect 10701 5049 10735 5083
rect 11713 5049 11747 5083
rect 13369 5049 13403 5083
rect 14740 5049 14774 5083
rect 18328 5049 18362 5083
rect 19984 5049 20018 5083
rect 11253 4981 11287 5015
rect 14105 4981 14139 5015
rect 17509 4981 17543 5015
rect 19533 4981 19567 5015
rect 21097 4981 21131 5015
rect 18245 4777 18279 4811
rect 18981 4777 19015 4811
rect 20085 4777 20119 4811
rect 9956 4709 9990 4743
rect 14749 4709 14783 4743
rect 16681 4709 16715 4743
rect 16773 4709 16807 4743
rect 19993 4709 20027 4743
rect 9689 4641 9723 4675
rect 11713 4641 11747 4675
rect 13165 4641 13199 4675
rect 15669 4641 15703 4675
rect 15761 4641 15795 4675
rect 18061 4641 18095 4675
rect 19073 4641 19107 4675
rect 20913 4641 20947 4675
rect 8953 4573 8987 4607
rect 9321 4573 9355 4607
rect 11805 4573 11839 4607
rect 11897 4573 11931 4607
rect 12357 4573 12391 4607
rect 12909 4573 12943 4607
rect 15853 4573 15887 4607
rect 16865 4573 16899 4607
rect 17325 4573 17359 4607
rect 19257 4573 19291 4607
rect 20269 4573 20303 4607
rect 14289 4505 14323 4539
rect 8585 4437 8619 4471
rect 11069 4437 11103 4471
rect 11345 4437 11379 4471
rect 15301 4437 15335 4471
rect 16313 4437 16347 4471
rect 18613 4437 18647 4471
rect 19625 4437 19659 4471
rect 21097 4437 21131 4471
rect 8861 4233 8895 4267
rect 9321 4233 9355 4267
rect 11989 4233 12023 4267
rect 20269 4233 20303 4267
rect 19993 4165 20027 4199
rect 10241 4097 10275 4131
rect 16037 4097 16071 4131
rect 16221 4097 16255 4131
rect 20821 4097 20855 4131
rect 10609 4029 10643 4063
rect 12541 4029 12575 4063
rect 13277 4029 13311 4063
rect 14933 4029 14967 4063
rect 15945 4029 15979 4063
rect 16589 4029 16623 4063
rect 17141 4029 17175 4063
rect 18061 4029 18095 4063
rect 18613 4029 18647 4063
rect 21281 4029 21315 4063
rect 8585 3961 8619 3995
rect 10876 3961 10910 3995
rect 13522 3961 13556 3995
rect 18880 3961 18914 3995
rect 9597 3893 9631 3927
rect 9965 3893 9999 3927
rect 10057 3893 10091 3927
rect 12725 3893 12759 3927
rect 14657 3893 14691 3927
rect 15117 3893 15151 3927
rect 15577 3893 15611 3927
rect 16773 3893 16807 3927
rect 17325 3893 17359 3927
rect 18245 3893 18279 3927
rect 20637 3893 20671 3927
rect 20729 3893 20763 3927
rect 9321 3689 9355 3723
rect 10057 3689 10091 3723
rect 10793 3689 10827 3723
rect 14197 3689 14231 3723
rect 18061 3689 18095 3723
rect 19717 3689 19751 3723
rect 12326 3621 12360 3655
rect 13921 3621 13955 3655
rect 16037 3621 16071 3655
rect 18582 3621 18616 3655
rect 11161 3553 11195 3587
rect 11253 3553 11287 3587
rect 12081 3553 12115 3587
rect 14565 3553 14599 3587
rect 15301 3553 15335 3587
rect 15761 3553 15795 3587
rect 16948 3553 16982 3587
rect 19993 3553 20027 3587
rect 20913 3553 20947 3587
rect 9781 3485 9815 3519
rect 9873 3485 9907 3519
rect 11345 3485 11379 3519
rect 14657 3485 14691 3519
rect 14749 3485 14783 3519
rect 16681 3485 16715 3519
rect 18337 3485 18371 3519
rect 20177 3485 20211 3519
rect 9873 3349 9907 3383
rect 10517 3349 10551 3383
rect 13461 3349 13495 3383
rect 21097 3349 21131 3383
rect 9229 3145 9263 3179
rect 10793 3145 10827 3179
rect 13461 3145 13495 3179
rect 17509 3145 17543 3179
rect 19073 3145 19107 3179
rect 10425 3077 10459 3111
rect 12265 3077 12299 3111
rect 9965 3009 9999 3043
rect 11345 3009 11379 3043
rect 10241 2941 10275 2975
rect 11805 2941 11839 2975
rect 12725 3009 12759 3043
rect 14013 3009 14047 3043
rect 18613 3009 18647 3043
rect 19717 3009 19751 3043
rect 20453 3009 20487 3043
rect 12541 2941 12575 2975
rect 14473 2941 14507 2975
rect 14740 2941 14774 2975
rect 16129 2941 16163 2975
rect 18429 2941 18463 2975
rect 19441 2941 19475 2975
rect 20177 2941 20211 2975
rect 20913 2941 20947 2975
rect 8861 2873 8895 2907
rect 12265 2873 12299 2907
rect 13829 2873 13863 2907
rect 16374 2873 16408 2907
rect 19533 2873 19567 2907
rect 9505 2805 9539 2839
rect 11161 2805 11195 2839
rect 11253 2805 11287 2839
rect 11989 2805 12023 2839
rect 13921 2805 13955 2839
rect 15853 2805 15887 2839
rect 18061 2805 18095 2839
rect 18521 2805 18555 2839
rect 21097 2805 21131 2839
rect 8953 2601 8987 2635
rect 10517 2601 10551 2635
rect 16313 2601 16347 2635
rect 16957 2601 16991 2635
rect 17325 2601 17359 2635
rect 21281 2601 21315 2635
rect 10885 2533 10919 2567
rect 11437 2533 11471 2567
rect 13645 2533 13679 2567
rect 15669 2533 15703 2567
rect 16405 2533 16439 2567
rect 11161 2465 11195 2499
rect 11989 2465 12023 2499
rect 12633 2465 12667 2499
rect 13369 2465 13403 2499
rect 14105 2465 14139 2499
rect 14657 2465 14691 2499
rect 17417 2465 17451 2499
rect 18337 2465 18371 2499
rect 18889 2465 18923 2499
rect 19441 2465 19475 2499
rect 19993 2465 20027 2499
rect 20545 2465 20579 2499
rect 10149 2397 10183 2431
rect 12817 2397 12851 2431
rect 16497 2397 16531 2431
rect 17509 2397 17543 2431
rect 15945 2329 15979 2363
rect 19073 2329 19107 2363
rect 20177 2329 20211 2363
rect 8309 2261 8343 2295
rect 8677 2261 8711 2295
rect 9413 2261 9447 2295
rect 12173 2261 12207 2295
rect 14289 2261 14323 2295
rect 14841 2261 14875 2295
rect 18521 2261 18555 2295
rect 19625 2261 19659 2295
rect 20729 2261 20763 2295
rect 15669 2057 15703 2091
rect 15669 1853 15703 1887
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 11149 20587 11207 20593
rect 11149 20553 11161 20587
rect 11195 20584 11207 20587
rect 12066 20584 12072 20596
rect 11195 20556 12072 20584
rect 11195 20553 11207 20556
rect 11149 20547 11207 20553
rect 12066 20544 12072 20556
rect 12124 20544 12130 20596
rect 12342 20544 12348 20596
rect 12400 20584 12406 20596
rect 12989 20587 13047 20593
rect 12989 20584 13001 20587
rect 12400 20556 13001 20584
rect 12400 20544 12406 20556
rect 12989 20553 13001 20556
rect 13035 20584 13047 20587
rect 14369 20587 14427 20593
rect 14369 20584 14381 20587
rect 13035 20556 14381 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 14369 20553 14381 20556
rect 14415 20553 14427 20587
rect 14369 20547 14427 20553
rect 14645 20587 14703 20593
rect 14645 20553 14657 20587
rect 14691 20584 14703 20587
rect 14826 20584 14832 20596
rect 14691 20556 14832 20584
rect 14691 20553 14703 20556
rect 14645 20547 14703 20553
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 16298 20544 16304 20596
rect 16356 20584 16362 20596
rect 17770 20584 17776 20596
rect 16356 20556 17776 20584
rect 16356 20544 16362 20556
rect 17770 20544 17776 20556
rect 17828 20544 17834 20596
rect 17865 20587 17923 20593
rect 17865 20553 17877 20587
rect 17911 20584 17923 20587
rect 18138 20584 18144 20596
rect 17911 20556 18144 20584
rect 17911 20553 17923 20556
rect 17865 20547 17923 20553
rect 18138 20544 18144 20556
rect 18196 20544 18202 20596
rect 18598 20544 18604 20596
rect 18656 20584 18662 20596
rect 19334 20584 19340 20596
rect 18656 20556 18920 20584
rect 19295 20556 19340 20584
rect 18656 20544 18662 20556
rect 11701 20519 11759 20525
rect 11701 20485 11713 20519
rect 11747 20516 11759 20519
rect 12618 20516 12624 20528
rect 11747 20488 12624 20516
rect 11747 20485 11759 20488
rect 11701 20479 11759 20485
rect 12618 20476 12624 20488
rect 12676 20476 12682 20528
rect 14093 20519 14151 20525
rect 14093 20485 14105 20519
rect 14139 20516 14151 20519
rect 15378 20516 15384 20528
rect 14139 20488 15384 20516
rect 14139 20485 14151 20488
rect 14093 20479 14151 20485
rect 15378 20476 15384 20488
rect 15436 20476 15442 20528
rect 16761 20519 16819 20525
rect 16761 20485 16773 20519
rect 16807 20485 16819 20519
rect 16761 20479 16819 20485
rect 17313 20519 17371 20525
rect 17313 20485 17325 20519
rect 17359 20516 17371 20519
rect 18782 20516 18788 20528
rect 17359 20488 18788 20516
rect 17359 20485 17371 20488
rect 17313 20479 17371 20485
rect 10321 20451 10379 20457
rect 10321 20417 10333 20451
rect 10367 20448 10379 20451
rect 10686 20448 10692 20460
rect 10367 20420 10692 20448
rect 10367 20417 10379 20420
rect 10321 20411 10379 20417
rect 10686 20408 10692 20420
rect 10744 20448 10750 20460
rect 15289 20451 15347 20457
rect 10744 20420 14504 20448
rect 10744 20408 10750 20420
rect 10962 20380 10968 20392
rect 10923 20352 10968 20380
rect 10962 20340 10968 20352
rect 11020 20340 11026 20392
rect 11517 20383 11575 20389
rect 11517 20349 11529 20383
rect 11563 20380 11575 20383
rect 12066 20380 12072 20392
rect 11563 20352 12072 20380
rect 11563 20349 11575 20352
rect 11517 20343 11575 20349
rect 12066 20340 12072 20352
rect 12124 20340 12130 20392
rect 12345 20383 12403 20389
rect 12345 20349 12357 20383
rect 12391 20380 12403 20383
rect 13357 20383 13415 20389
rect 13357 20380 13369 20383
rect 12391 20352 13369 20380
rect 12391 20349 12403 20352
rect 12345 20343 12403 20349
rect 13357 20349 13369 20352
rect 13403 20349 13415 20383
rect 13357 20343 13415 20349
rect 13446 20340 13452 20392
rect 13504 20380 13510 20392
rect 14476 20389 14504 20420
rect 15289 20417 15301 20451
rect 15335 20448 15347 20451
rect 16485 20451 16543 20457
rect 16485 20448 16497 20451
rect 15335 20420 16497 20448
rect 15335 20417 15347 20420
rect 15289 20411 15347 20417
rect 13725 20383 13783 20389
rect 13725 20380 13737 20383
rect 13504 20352 13737 20380
rect 13504 20340 13510 20352
rect 13725 20349 13737 20352
rect 13771 20349 13783 20383
rect 13725 20343 13783 20349
rect 13909 20383 13967 20389
rect 13909 20349 13921 20383
rect 13955 20349 13967 20383
rect 13909 20343 13967 20349
rect 14461 20383 14519 20389
rect 14461 20349 14473 20383
rect 14507 20349 14519 20383
rect 14461 20343 14519 20349
rect 15473 20383 15531 20389
rect 15473 20349 15485 20383
rect 15519 20380 15531 20383
rect 15838 20380 15844 20392
rect 15519 20352 15844 20380
rect 15519 20349 15531 20352
rect 15473 20343 15531 20349
rect 9953 20315 10011 20321
rect 9953 20281 9965 20315
rect 9999 20312 10011 20315
rect 12250 20312 12256 20324
rect 9999 20284 12256 20312
rect 9999 20281 10011 20284
rect 9953 20275 10011 20281
rect 12250 20272 12256 20284
rect 12308 20312 12314 20324
rect 13924 20312 13952 20343
rect 15838 20340 15844 20352
rect 15896 20340 15902 20392
rect 16040 20389 16068 20420
rect 16485 20417 16497 20420
rect 16531 20417 16543 20451
rect 16776 20448 16804 20479
rect 18782 20476 18788 20488
rect 18840 20476 18846 20528
rect 18892 20516 18920 20556
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 19886 20584 19892 20596
rect 19847 20556 19892 20584
rect 19886 20544 19892 20556
rect 19944 20544 19950 20596
rect 21177 20519 21235 20525
rect 21177 20516 21189 20519
rect 18892 20488 21189 20516
rect 21177 20485 21189 20488
rect 21223 20485 21235 20519
rect 21177 20479 21235 20485
rect 19426 20448 19432 20460
rect 16776 20420 19432 20448
rect 16485 20411 16543 20417
rect 19426 20408 19432 20420
rect 19484 20408 19490 20460
rect 16025 20383 16083 20389
rect 16025 20349 16037 20383
rect 16071 20349 16083 20383
rect 16577 20383 16635 20389
rect 16577 20380 16589 20383
rect 16025 20343 16083 20349
rect 16132 20352 16589 20380
rect 12308 20284 13952 20312
rect 14369 20315 14427 20321
rect 12308 20272 12314 20284
rect 14369 20281 14381 20315
rect 14415 20312 14427 20315
rect 15013 20315 15071 20321
rect 15013 20312 15025 20315
rect 14415 20284 15025 20312
rect 14415 20281 14427 20284
rect 14369 20275 14427 20281
rect 15013 20281 15025 20284
rect 15059 20312 15071 20315
rect 16132 20312 16160 20352
rect 16577 20349 16589 20352
rect 16623 20349 16635 20383
rect 16577 20343 16635 20349
rect 17129 20383 17187 20389
rect 17129 20349 17141 20383
rect 17175 20380 17187 20383
rect 17589 20383 17647 20389
rect 17589 20380 17601 20383
rect 17175 20352 17601 20380
rect 17175 20349 17187 20352
rect 17129 20343 17187 20349
rect 17589 20349 17601 20352
rect 17635 20349 17647 20383
rect 17589 20343 17647 20349
rect 17681 20383 17739 20389
rect 17681 20349 17693 20383
rect 17727 20380 17739 20383
rect 17770 20380 17776 20392
rect 17727 20352 17776 20380
rect 17727 20349 17739 20352
rect 17681 20343 17739 20349
rect 17770 20340 17776 20352
rect 17828 20380 17834 20392
rect 18414 20380 18420 20392
rect 17828 20352 18420 20380
rect 17828 20340 17834 20352
rect 18414 20340 18420 20352
rect 18472 20340 18478 20392
rect 18598 20380 18604 20392
rect 18559 20352 18604 20380
rect 18598 20340 18604 20352
rect 18656 20340 18662 20392
rect 19150 20380 19156 20392
rect 19111 20352 19156 20380
rect 19150 20340 19156 20352
rect 19208 20340 19214 20392
rect 19518 20340 19524 20392
rect 19576 20380 19582 20392
rect 19705 20383 19763 20389
rect 19705 20380 19717 20383
rect 19576 20352 19717 20380
rect 19576 20340 19582 20352
rect 19705 20349 19717 20352
rect 19751 20349 19763 20383
rect 20530 20380 20536 20392
rect 20491 20352 20536 20380
rect 19705 20343 19763 20349
rect 20530 20340 20536 20352
rect 20588 20340 20594 20392
rect 19794 20312 19800 20324
rect 15059 20284 16160 20312
rect 16224 20284 19800 20312
rect 15059 20281 15071 20284
rect 15013 20275 15071 20281
rect 16040 20256 16068 20284
rect 7742 20204 7748 20256
rect 7800 20244 7806 20256
rect 9309 20247 9367 20253
rect 9309 20244 9321 20247
rect 7800 20216 9321 20244
rect 7800 20204 7806 20216
rect 9309 20213 9321 20216
rect 9355 20213 9367 20247
rect 9309 20207 9367 20213
rect 10410 20204 10416 20256
rect 10468 20244 10474 20256
rect 10689 20247 10747 20253
rect 10689 20244 10701 20247
rect 10468 20216 10701 20244
rect 10468 20204 10474 20216
rect 10689 20213 10701 20216
rect 10735 20244 10747 20247
rect 10778 20244 10784 20256
rect 10735 20216 10784 20244
rect 10735 20213 10747 20216
rect 10689 20207 10747 20213
rect 10778 20204 10784 20216
rect 10836 20204 10842 20256
rect 11974 20204 11980 20256
rect 12032 20244 12038 20256
rect 12161 20247 12219 20253
rect 12161 20244 12173 20247
rect 12032 20216 12173 20244
rect 12032 20204 12038 20216
rect 12161 20213 12173 20216
rect 12207 20244 12219 20247
rect 12345 20247 12403 20253
rect 12345 20244 12357 20247
rect 12207 20216 12357 20244
rect 12207 20213 12219 20216
rect 12161 20207 12219 20213
rect 12345 20213 12357 20216
rect 12391 20213 12403 20247
rect 12345 20207 12403 20213
rect 12713 20247 12771 20253
rect 12713 20213 12725 20247
rect 12759 20244 12771 20247
rect 12986 20244 12992 20256
rect 12759 20216 12992 20244
rect 12759 20213 12771 20216
rect 12713 20207 12771 20213
rect 12986 20204 12992 20216
rect 13044 20244 13050 20256
rect 13446 20244 13452 20256
rect 13044 20216 13452 20244
rect 13044 20204 13050 20216
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 13538 20204 13544 20256
rect 13596 20244 13602 20256
rect 13725 20247 13783 20253
rect 13596 20216 13641 20244
rect 13596 20204 13602 20216
rect 13725 20213 13737 20247
rect 13771 20244 13783 20247
rect 15289 20247 15347 20253
rect 15289 20244 15301 20247
rect 13771 20216 15301 20244
rect 13771 20213 13783 20216
rect 13725 20207 13783 20213
rect 15289 20213 15301 20216
rect 15335 20213 15347 20247
rect 15289 20207 15347 20213
rect 15657 20247 15715 20253
rect 15657 20213 15669 20247
rect 15703 20244 15715 20247
rect 15746 20244 15752 20256
rect 15703 20216 15752 20244
rect 15703 20213 15715 20216
rect 15657 20207 15715 20213
rect 15746 20204 15752 20216
rect 15804 20204 15810 20256
rect 16022 20204 16028 20256
rect 16080 20204 16086 20256
rect 16224 20253 16252 20284
rect 19794 20272 19800 20284
rect 19852 20272 19858 20324
rect 16209 20247 16267 20253
rect 16209 20213 16221 20247
rect 16255 20213 16267 20247
rect 16209 20207 16267 20213
rect 16485 20247 16543 20253
rect 16485 20213 16497 20247
rect 16531 20244 16543 20247
rect 17126 20244 17132 20256
rect 16531 20216 17132 20244
rect 16531 20213 16543 20216
rect 16485 20207 16543 20213
rect 17126 20204 17132 20216
rect 17184 20204 17190 20256
rect 17589 20247 17647 20253
rect 17589 20213 17601 20247
rect 17635 20244 17647 20247
rect 17954 20244 17960 20256
rect 17635 20216 17960 20244
rect 17635 20213 17647 20216
rect 17589 20207 17647 20213
rect 17954 20204 17960 20216
rect 18012 20204 18018 20256
rect 18785 20247 18843 20253
rect 18785 20213 18797 20247
rect 18831 20244 18843 20247
rect 18874 20244 18880 20256
rect 18831 20216 18880 20244
rect 18831 20213 18843 20216
rect 18785 20207 18843 20213
rect 18874 20204 18880 20216
rect 18932 20204 18938 20256
rect 20622 20204 20628 20256
rect 20680 20244 20686 20256
rect 20717 20247 20775 20253
rect 20717 20244 20729 20247
rect 20680 20216 20729 20244
rect 20680 20204 20686 20216
rect 20717 20213 20729 20216
rect 20763 20213 20775 20247
rect 20717 20207 20775 20213
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 8941 20043 8999 20049
rect 8941 20009 8953 20043
rect 8987 20040 8999 20043
rect 11238 20040 11244 20052
rect 8987 20012 11244 20040
rect 8987 20009 8999 20012
rect 8941 20003 8999 20009
rect 11238 20000 11244 20012
rect 11296 20040 11302 20052
rect 13449 20043 13507 20049
rect 13449 20040 13461 20043
rect 11296 20012 13461 20040
rect 11296 20000 11302 20012
rect 13449 20009 13461 20012
rect 13495 20009 13507 20043
rect 13449 20003 13507 20009
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 13872 20012 14289 20040
rect 13872 20000 13878 20012
rect 14277 20009 14289 20012
rect 14323 20009 14335 20043
rect 14277 20003 14335 20009
rect 14366 20000 14372 20052
rect 14424 20040 14430 20052
rect 14829 20043 14887 20049
rect 14829 20040 14841 20043
rect 14424 20012 14841 20040
rect 14424 20000 14430 20012
rect 14829 20009 14841 20012
rect 14875 20009 14887 20043
rect 14829 20003 14887 20009
rect 15930 20000 15936 20052
rect 15988 20040 15994 20052
rect 16485 20043 16543 20049
rect 16485 20040 16497 20043
rect 15988 20012 16497 20040
rect 15988 20000 15994 20012
rect 16485 20009 16497 20012
rect 16531 20009 16543 20043
rect 16485 20003 16543 20009
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 17037 20043 17095 20049
rect 17037 20040 17049 20043
rect 16632 20012 17049 20040
rect 16632 20000 16638 20012
rect 17037 20009 17049 20012
rect 17083 20009 17095 20043
rect 17037 20003 17095 20009
rect 18049 20043 18107 20049
rect 18049 20009 18061 20043
rect 18095 20040 18107 20043
rect 18690 20040 18696 20052
rect 18095 20012 18696 20040
rect 18095 20009 18107 20012
rect 18049 20003 18107 20009
rect 18690 20000 18696 20012
rect 18748 20000 18754 20052
rect 18966 20040 18972 20052
rect 18927 20012 18972 20040
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 20990 20040 20996 20052
rect 19076 20012 20996 20040
rect 9122 19932 9128 19984
rect 9180 19972 9186 19984
rect 11882 19972 11888 19984
rect 9180 19944 11888 19972
rect 9180 19932 9186 19944
rect 11882 19932 11888 19944
rect 11940 19932 11946 19984
rect 13722 19932 13728 19984
rect 13780 19972 13786 19984
rect 14458 19972 14464 19984
rect 13780 19944 13952 19972
rect 13780 19932 13786 19944
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 10413 19907 10471 19913
rect 10413 19904 10425 19907
rect 9732 19876 10425 19904
rect 9732 19864 9738 19876
rect 10413 19873 10425 19876
rect 10459 19873 10471 19907
rect 10413 19867 10471 19873
rect 11149 19907 11207 19913
rect 11149 19873 11161 19907
rect 11195 19904 11207 19907
rect 11238 19904 11244 19916
rect 11195 19876 11244 19904
rect 11195 19873 11207 19876
rect 11149 19867 11207 19873
rect 11238 19864 11244 19876
rect 11296 19864 11302 19916
rect 11416 19907 11474 19913
rect 11416 19873 11428 19907
rect 11462 19904 11474 19907
rect 11698 19904 11704 19916
rect 11462 19876 11704 19904
rect 11462 19873 11474 19876
rect 11416 19867 11474 19873
rect 11698 19864 11704 19876
rect 11756 19864 11762 19916
rect 9861 19839 9919 19845
rect 9861 19805 9873 19839
rect 9907 19836 9919 19839
rect 10505 19839 10563 19845
rect 10505 19836 10517 19839
rect 9907 19808 10517 19836
rect 9907 19805 9919 19808
rect 9861 19799 9919 19805
rect 10505 19805 10517 19808
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 10594 19796 10600 19848
rect 10652 19836 10658 19848
rect 10652 19808 10697 19836
rect 10652 19796 10658 19808
rect 12158 19796 12164 19848
rect 12216 19836 12222 19848
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 12216 19808 13553 19836
rect 12216 19796 12222 19808
rect 13541 19805 13553 19808
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19836 13783 19839
rect 13814 19836 13820 19848
rect 13771 19808 13820 19836
rect 13771 19805 13783 19808
rect 13725 19799 13783 19805
rect 13814 19796 13820 19808
rect 13872 19796 13878 19848
rect 13924 19836 13952 19944
rect 14200 19944 14464 19972
rect 14093 19907 14151 19913
rect 14093 19873 14105 19907
rect 14139 19904 14151 19907
rect 14200 19904 14228 19944
rect 14458 19932 14464 19944
rect 14516 19932 14522 19984
rect 15746 19932 15752 19984
rect 15804 19972 15810 19984
rect 19076 19972 19104 20012
rect 20990 20000 20996 20012
rect 21048 20000 21054 20052
rect 15804 19944 19104 19972
rect 15804 19932 15810 19944
rect 19150 19932 19156 19984
rect 19208 19972 19214 19984
rect 21177 19975 21235 19981
rect 21177 19972 21189 19975
rect 19208 19944 21189 19972
rect 19208 19932 19214 19944
rect 21177 19941 21189 19944
rect 21223 19941 21235 19975
rect 21177 19935 21235 19941
rect 14139 19876 14228 19904
rect 14645 19907 14703 19913
rect 14139 19873 14151 19876
rect 14093 19867 14151 19873
rect 14645 19873 14657 19907
rect 14691 19873 14703 19907
rect 15654 19904 15660 19916
rect 15615 19876 15660 19904
rect 14645 19867 14703 19873
rect 14660 19836 14688 19867
rect 15654 19864 15660 19876
rect 15712 19864 15718 19916
rect 16301 19907 16359 19913
rect 16301 19873 16313 19907
rect 16347 19904 16359 19907
rect 16390 19904 16396 19916
rect 16347 19876 16396 19904
rect 16347 19873 16359 19876
rect 16301 19867 16359 19873
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 16853 19907 16911 19913
rect 16853 19873 16865 19907
rect 16899 19904 16911 19907
rect 17310 19904 17316 19916
rect 16899 19876 17316 19904
rect 16899 19873 16911 19876
rect 16853 19867 16911 19873
rect 17310 19864 17316 19876
rect 17368 19864 17374 19916
rect 17862 19904 17868 19916
rect 17823 19876 17868 19904
rect 17862 19864 17868 19876
rect 17920 19864 17926 19916
rect 18414 19904 18420 19916
rect 18375 19876 18420 19904
rect 18414 19864 18420 19876
rect 18472 19864 18478 19916
rect 18782 19904 18788 19916
rect 18743 19876 18788 19904
rect 18782 19864 18788 19876
rect 18840 19864 18846 19916
rect 19705 19907 19763 19913
rect 19705 19904 19717 19907
rect 18892 19876 19717 19904
rect 13924 19808 14688 19836
rect 15378 19796 15384 19848
rect 15436 19836 15442 19848
rect 15749 19839 15807 19845
rect 15749 19836 15761 19839
rect 15436 19808 15761 19836
rect 15436 19796 15442 19808
rect 15749 19805 15761 19808
rect 15795 19805 15807 19839
rect 15749 19799 15807 19805
rect 15838 19796 15844 19848
rect 15896 19836 15902 19848
rect 15896 19808 15941 19836
rect 15896 19796 15902 19808
rect 16574 19796 16580 19848
rect 16632 19836 16638 19848
rect 17405 19839 17463 19845
rect 17405 19836 17417 19839
rect 16632 19808 17417 19836
rect 16632 19796 16638 19808
rect 17405 19805 17417 19808
rect 17451 19805 17463 19839
rect 17405 19799 17463 19805
rect 11146 19768 11152 19780
rect 9232 19740 11152 19768
rect 7558 19660 7564 19712
rect 7616 19700 7622 19712
rect 8386 19700 8392 19712
rect 7616 19672 8392 19700
rect 7616 19660 7622 19672
rect 8386 19660 8392 19672
rect 8444 19700 8450 19712
rect 9232 19709 9260 19740
rect 11146 19728 11152 19740
rect 11204 19728 11210 19780
rect 12084 19740 15424 19768
rect 9217 19703 9275 19709
rect 9217 19700 9229 19703
rect 8444 19672 9229 19700
rect 8444 19660 8450 19672
rect 9217 19669 9229 19672
rect 9263 19669 9275 19703
rect 9217 19663 9275 19669
rect 9769 19703 9827 19709
rect 9769 19669 9781 19703
rect 9815 19700 9827 19703
rect 9858 19700 9864 19712
rect 9815 19672 9864 19700
rect 9815 19669 9827 19672
rect 9769 19663 9827 19669
rect 9858 19660 9864 19672
rect 9916 19660 9922 19712
rect 10045 19703 10103 19709
rect 10045 19669 10057 19703
rect 10091 19700 10103 19703
rect 11790 19700 11796 19712
rect 10091 19672 11796 19700
rect 10091 19669 10103 19672
rect 10045 19663 10103 19669
rect 11790 19660 11796 19672
rect 11848 19660 11854 19712
rect 11882 19660 11888 19712
rect 11940 19700 11946 19712
rect 12084 19700 12112 19740
rect 12526 19700 12532 19712
rect 11940 19672 12112 19700
rect 12487 19672 12532 19700
rect 11940 19660 11946 19672
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 13081 19703 13139 19709
rect 13081 19669 13093 19703
rect 13127 19700 13139 19703
rect 14642 19700 14648 19712
rect 13127 19672 14648 19700
rect 13127 19669 13139 19672
rect 13081 19663 13139 19669
rect 14642 19660 14648 19672
rect 14700 19660 14706 19712
rect 15286 19700 15292 19712
rect 15247 19672 15292 19700
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 15396 19700 15424 19740
rect 18892 19700 18920 19876
rect 19705 19873 19717 19876
rect 19751 19873 19763 19907
rect 19705 19867 19763 19873
rect 20257 19907 20315 19913
rect 20257 19873 20269 19907
rect 20303 19904 20315 19907
rect 20714 19904 20720 19916
rect 20303 19876 20720 19904
rect 20303 19873 20315 19876
rect 20257 19867 20315 19873
rect 20714 19864 20720 19876
rect 20772 19864 20778 19916
rect 20809 19907 20867 19913
rect 20809 19873 20821 19907
rect 20855 19904 20867 19907
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20855 19876 20913 19904
rect 20855 19873 20867 19876
rect 20809 19867 20867 19873
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 18966 19796 18972 19848
rect 19024 19836 19030 19848
rect 21542 19836 21548 19848
rect 19024 19808 21548 19836
rect 19024 19796 19030 19808
rect 21542 19796 21548 19808
rect 21600 19796 21606 19848
rect 19242 19728 19248 19780
rect 19300 19768 19306 19780
rect 20441 19771 20499 19777
rect 20441 19768 20453 19771
rect 19300 19740 20453 19768
rect 19300 19728 19306 19740
rect 20441 19737 20453 19740
rect 20487 19737 20499 19771
rect 20441 19731 20499 19737
rect 15396 19672 18920 19700
rect 19150 19660 19156 19712
rect 19208 19700 19214 19712
rect 19337 19703 19395 19709
rect 19337 19700 19349 19703
rect 19208 19672 19349 19700
rect 19208 19660 19214 19672
rect 19337 19669 19349 19672
rect 19383 19669 19395 19703
rect 19886 19700 19892 19712
rect 19847 19672 19892 19700
rect 19337 19663 19395 19669
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 19978 19660 19984 19712
rect 20036 19700 20042 19712
rect 20717 19703 20775 19709
rect 20717 19700 20729 19703
rect 20036 19672 20729 19700
rect 20036 19660 20042 19672
rect 20717 19669 20729 19672
rect 20763 19669 20775 19703
rect 20717 19663 20775 19669
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 9490 19456 9496 19508
rect 9548 19496 9554 19508
rect 11609 19499 11667 19505
rect 9548 19468 11192 19496
rect 9548 19456 9554 19468
rect 11164 19428 11192 19468
rect 11609 19465 11621 19499
rect 11655 19496 11667 19499
rect 11698 19496 11704 19508
rect 11655 19468 11704 19496
rect 11655 19465 11667 19468
rect 11609 19459 11667 19465
rect 11698 19456 11704 19468
rect 11756 19456 11762 19508
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 13814 19496 13820 19508
rect 12492 19468 13676 19496
rect 13775 19468 13820 19496
rect 12492 19456 12498 19468
rect 12342 19428 12348 19440
rect 11164 19400 12348 19428
rect 12342 19388 12348 19400
rect 12400 19388 12406 19440
rect 13648 19428 13676 19468
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 14108 19468 15608 19496
rect 14108 19428 14136 19468
rect 13648 19400 14136 19428
rect 15473 19431 15531 19437
rect 15473 19397 15485 19431
rect 15519 19397 15531 19431
rect 15580 19428 15608 19468
rect 15654 19456 15660 19508
rect 15712 19496 15718 19508
rect 15749 19499 15807 19505
rect 15749 19496 15761 19499
rect 15712 19468 15761 19496
rect 15712 19456 15718 19468
rect 15749 19465 15761 19468
rect 15795 19465 15807 19499
rect 15749 19459 15807 19465
rect 15930 19456 15936 19508
rect 15988 19496 15994 19508
rect 21542 19496 21548 19508
rect 15988 19468 21548 19496
rect 15988 19456 15994 19468
rect 21542 19456 21548 19468
rect 21600 19456 21606 19508
rect 19150 19428 19156 19440
rect 15580 19400 19156 19428
rect 15473 19391 15531 19397
rect 8481 19363 8539 19369
rect 8481 19329 8493 19363
rect 8527 19360 8539 19363
rect 9309 19363 9367 19369
rect 9309 19360 9321 19363
rect 8527 19332 9321 19360
rect 8527 19329 8539 19332
rect 8481 19323 8539 19329
rect 9309 19329 9321 19332
rect 9355 19360 9367 19363
rect 9582 19360 9588 19372
rect 9355 19332 9588 19360
rect 9355 19329 9367 19332
rect 9309 19323 9367 19329
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 11882 19360 11888 19372
rect 11843 19332 11888 19360
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 13872 19332 14228 19360
rect 13872 19320 13878 19332
rect 290 19252 296 19304
rect 348 19292 354 19304
rect 8570 19292 8576 19304
rect 348 19264 8576 19292
rect 348 19252 354 19264
rect 8570 19252 8576 19264
rect 8628 19252 8634 19304
rect 9214 19252 9220 19304
rect 9272 19292 9278 19304
rect 9674 19292 9680 19304
rect 9272 19264 9680 19292
rect 9272 19252 9278 19264
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 9766 19252 9772 19304
rect 9824 19292 9830 19304
rect 10229 19295 10287 19301
rect 10229 19292 10241 19295
rect 9824 19264 10241 19292
rect 9824 19252 9830 19264
rect 10229 19261 10241 19264
rect 10275 19292 10287 19295
rect 11238 19292 11244 19304
rect 10275 19264 11244 19292
rect 10275 19261 10287 19264
rect 10229 19255 10287 19261
rect 11238 19252 11244 19264
rect 11296 19292 11302 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 11296 19264 12449 19292
rect 11296 19252 11302 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 12526 19252 12532 19304
rect 12584 19292 12590 19304
rect 12693 19295 12751 19301
rect 12693 19292 12705 19295
rect 12584 19264 12705 19292
rect 12584 19252 12590 19264
rect 12693 19261 12705 19264
rect 12739 19261 12751 19295
rect 14090 19292 14096 19304
rect 14051 19264 14096 19292
rect 12693 19255 12751 19261
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 14200 19292 14228 19332
rect 15194 19320 15200 19372
rect 15252 19360 15258 19372
rect 15488 19360 15516 19391
rect 19150 19388 19156 19400
rect 19208 19388 19214 19440
rect 16301 19363 16359 19369
rect 16301 19360 16313 19363
rect 15252 19332 16313 19360
rect 15252 19320 15258 19332
rect 16301 19329 16313 19332
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19360 17279 19363
rect 17862 19360 17868 19372
rect 17267 19332 17868 19360
rect 17267 19329 17279 19332
rect 17221 19323 17279 19329
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19360 18383 19363
rect 18782 19360 18788 19372
rect 18371 19332 18788 19360
rect 18371 19329 18383 19332
rect 18325 19323 18383 19329
rect 18782 19320 18788 19332
rect 18840 19320 18846 19372
rect 20257 19363 20315 19369
rect 20257 19329 20269 19363
rect 20303 19329 20315 19363
rect 20257 19323 20315 19329
rect 14349 19295 14407 19301
rect 14349 19292 14361 19295
rect 14200 19264 14361 19292
rect 14349 19261 14361 19264
rect 14395 19261 14407 19295
rect 14349 19255 14407 19261
rect 16117 19295 16175 19301
rect 16117 19261 16129 19295
rect 16163 19292 16175 19295
rect 16574 19292 16580 19304
rect 16163 19264 16580 19292
rect 16163 19261 16175 19264
rect 16117 19255 16175 19261
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 16850 19252 16856 19304
rect 16908 19292 16914 19304
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 16908 19264 16957 19292
rect 16908 19252 16914 19264
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 18046 19292 18052 19304
rect 18007 19264 18052 19292
rect 16945 19255 17003 19261
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 18877 19295 18935 19301
rect 18877 19292 18889 19295
rect 18800 19264 18889 19292
rect 18800 19236 18828 19264
rect 18877 19261 18889 19264
rect 18923 19261 18935 19295
rect 18877 19255 18935 19261
rect 19153 19295 19211 19301
rect 19153 19261 19165 19295
rect 19199 19292 19211 19295
rect 19518 19292 19524 19304
rect 19199 19264 19524 19292
rect 19199 19261 19211 19264
rect 19153 19255 19211 19261
rect 19518 19252 19524 19264
rect 19576 19252 19582 19304
rect 19889 19295 19947 19301
rect 19889 19292 19901 19295
rect 19628 19264 19901 19292
rect 8297 19227 8355 19233
rect 8297 19193 8309 19227
rect 8343 19224 8355 19227
rect 10134 19224 10140 19236
rect 8343 19196 10140 19224
rect 8343 19193 8355 19196
rect 8297 19187 8355 19193
rect 10134 19184 10140 19196
rect 10192 19184 10198 19236
rect 10502 19233 10508 19236
rect 10496 19224 10508 19233
rect 10463 19196 10508 19224
rect 10496 19187 10508 19196
rect 10502 19184 10508 19187
rect 10560 19184 10566 19236
rect 13906 19184 13912 19236
rect 13964 19224 13970 19236
rect 13964 19196 14872 19224
rect 13964 19184 13970 19196
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 8481 19159 8539 19165
rect 8481 19156 8493 19159
rect 4212 19128 8493 19156
rect 4212 19116 4218 19128
rect 8481 19125 8493 19128
rect 8527 19125 8539 19159
rect 8481 19119 8539 19125
rect 8665 19159 8723 19165
rect 8665 19125 8677 19159
rect 8711 19156 8723 19159
rect 8938 19156 8944 19168
rect 8711 19128 8944 19156
rect 8711 19125 8723 19128
rect 8665 19119 8723 19125
rect 8938 19116 8944 19128
rect 8996 19116 9002 19168
rect 9030 19116 9036 19168
rect 9088 19156 9094 19168
rect 9088 19128 9133 19156
rect 9088 19116 9094 19128
rect 10778 19116 10784 19168
rect 10836 19156 10842 19168
rect 14734 19156 14740 19168
rect 10836 19128 14740 19156
rect 10836 19116 10842 19128
rect 14734 19116 14740 19128
rect 14792 19116 14798 19168
rect 14844 19156 14872 19196
rect 16022 19184 16028 19236
rect 16080 19224 16086 19236
rect 16209 19227 16267 19233
rect 16209 19224 16221 19227
rect 16080 19196 16221 19224
rect 16080 19184 16086 19196
rect 16209 19193 16221 19196
rect 16255 19193 16267 19227
rect 16209 19187 16267 19193
rect 18782 19184 18788 19236
rect 18840 19184 18846 19236
rect 18966 19184 18972 19236
rect 19024 19224 19030 19236
rect 19628 19224 19656 19264
rect 19889 19261 19901 19264
rect 19935 19261 19947 19295
rect 19889 19255 19947 19261
rect 19024 19196 19656 19224
rect 19024 19184 19030 19196
rect 19794 19184 19800 19236
rect 19852 19224 19858 19236
rect 20272 19224 20300 19323
rect 22646 19224 22652 19236
rect 19852 19196 20300 19224
rect 20364 19196 22652 19224
rect 19852 19184 19858 19196
rect 20364 19156 20392 19196
rect 22646 19184 22652 19196
rect 22704 19184 22710 19236
rect 14844 19128 20392 19156
rect 21269 19159 21327 19165
rect 21269 19125 21281 19159
rect 21315 19156 21327 19159
rect 21450 19156 21456 19168
rect 21315 19128 21456 19156
rect 21315 19125 21327 19128
rect 21269 19119 21327 19125
rect 21450 19116 21456 19128
rect 21508 19116 21514 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 842 18912 848 18964
rect 900 18952 906 18964
rect 6362 18952 6368 18964
rect 900 18924 6368 18952
rect 900 18912 906 18924
rect 6362 18912 6368 18924
rect 6420 18912 6426 18964
rect 6454 18912 6460 18964
rect 6512 18952 6518 18964
rect 9858 18952 9864 18964
rect 6512 18924 9864 18952
rect 6512 18912 6518 18924
rect 9858 18912 9864 18924
rect 9916 18952 9922 18964
rect 10042 18952 10048 18964
rect 9916 18924 10048 18952
rect 9916 18912 9922 18924
rect 10042 18912 10048 18924
rect 10100 18912 10106 18964
rect 10502 18912 10508 18964
rect 10560 18952 10566 18964
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 10560 18924 11069 18952
rect 10560 18912 10566 18924
rect 11057 18921 11069 18924
rect 11103 18921 11115 18955
rect 11790 18952 11796 18964
rect 11751 18924 11796 18952
rect 11057 18915 11115 18921
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 11882 18912 11888 18964
rect 11940 18952 11946 18964
rect 12713 18955 12771 18961
rect 12713 18952 12725 18955
rect 11940 18924 12725 18952
rect 11940 18912 11946 18924
rect 12713 18921 12725 18924
rect 12759 18921 12771 18955
rect 12713 18915 12771 18921
rect 13170 18912 13176 18964
rect 13228 18952 13234 18964
rect 13541 18955 13599 18961
rect 13541 18952 13553 18955
rect 13228 18924 13553 18952
rect 13228 18912 13234 18924
rect 13541 18921 13553 18924
rect 13587 18921 13599 18955
rect 14642 18952 14648 18964
rect 14603 18924 14648 18952
rect 13541 18915 13599 18921
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 15672 18924 16988 18952
rect 1394 18844 1400 18896
rect 1452 18884 1458 18896
rect 6822 18884 6828 18896
rect 1452 18856 6828 18884
rect 1452 18844 1458 18856
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 9030 18844 9036 18896
rect 9088 18884 9094 18896
rect 15672 18884 15700 18924
rect 9088 18856 15700 18884
rect 15740 18887 15798 18893
rect 9088 18844 9094 18856
rect 15740 18853 15752 18887
rect 15786 18884 15798 18887
rect 15838 18884 15844 18896
rect 15786 18856 15844 18884
rect 15786 18853 15798 18856
rect 15740 18847 15798 18853
rect 15838 18844 15844 18856
rect 15896 18844 15902 18896
rect 16960 18884 16988 18924
rect 17034 18912 17040 18964
rect 17092 18952 17098 18964
rect 17313 18955 17371 18961
rect 17313 18952 17325 18955
rect 17092 18924 17325 18952
rect 17092 18912 17098 18924
rect 17313 18921 17325 18924
rect 17359 18921 17371 18955
rect 17313 18915 17371 18921
rect 17678 18912 17684 18964
rect 17736 18952 17742 18964
rect 17865 18955 17923 18961
rect 17865 18952 17877 18955
rect 17736 18924 17877 18952
rect 17736 18912 17742 18924
rect 17865 18921 17877 18924
rect 17911 18921 17923 18955
rect 17865 18915 17923 18921
rect 18049 18955 18107 18961
rect 18049 18921 18061 18955
rect 18095 18952 18107 18955
rect 20530 18952 20536 18964
rect 18095 18924 20536 18952
rect 18095 18921 18107 18924
rect 18049 18915 18107 18921
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 18966 18884 18972 18896
rect 16960 18856 18972 18884
rect 18966 18844 18972 18856
rect 19024 18844 19030 18896
rect 19153 18887 19211 18893
rect 19153 18853 19165 18887
rect 19199 18884 19211 18887
rect 20346 18884 20352 18896
rect 19199 18856 20352 18884
rect 19199 18853 19211 18856
rect 19153 18847 19211 18853
rect 20346 18844 20352 18856
rect 20404 18844 20410 18896
rect 2498 18776 2504 18828
rect 2556 18816 2562 18828
rect 8849 18819 8907 18825
rect 8849 18816 8861 18819
rect 2556 18788 8861 18816
rect 2556 18776 2562 18788
rect 8849 18785 8861 18788
rect 8895 18785 8907 18819
rect 8849 18779 8907 18785
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 8260 18720 8616 18748
rect 8260 18708 8266 18720
rect 3050 18572 3056 18624
rect 3108 18612 3114 18624
rect 7650 18612 7656 18624
rect 3108 18584 7656 18612
rect 3108 18572 3114 18584
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 8202 18612 8208 18624
rect 8163 18584 8208 18612
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 8478 18612 8484 18624
rect 8439 18584 8484 18612
rect 8478 18572 8484 18584
rect 8536 18572 8542 18624
rect 8588 18612 8616 18720
rect 8864 18680 8892 18779
rect 9214 18776 9220 18828
rect 9272 18816 9278 18828
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 9272 18788 9689 18816
rect 9272 18776 9278 18788
rect 9677 18785 9689 18788
rect 9723 18816 9735 18819
rect 9766 18816 9772 18828
rect 9723 18788 9772 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 9766 18776 9772 18788
rect 9824 18776 9830 18828
rect 9944 18819 10002 18825
rect 9944 18785 9956 18819
rect 9990 18816 10002 18819
rect 11238 18816 11244 18828
rect 9990 18788 11244 18816
rect 9990 18785 10002 18788
rect 9944 18779 10002 18785
rect 11238 18776 11244 18788
rect 11296 18776 11302 18828
rect 11701 18819 11759 18825
rect 11701 18785 11713 18819
rect 11747 18785 11759 18819
rect 13354 18816 13360 18828
rect 11701 18779 11759 18785
rect 11900 18788 12940 18816
rect 13315 18788 13360 18816
rect 8938 18708 8944 18760
rect 8996 18748 9002 18760
rect 9398 18748 9404 18760
rect 8996 18720 9404 18748
rect 8996 18708 9002 18720
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 11146 18708 11152 18760
rect 11204 18748 11210 18760
rect 11716 18748 11744 18779
rect 11204 18720 11744 18748
rect 11204 18708 11210 18720
rect 11790 18708 11796 18760
rect 11848 18748 11854 18760
rect 11900 18757 11928 18788
rect 11885 18751 11943 18757
rect 11885 18748 11897 18751
rect 11848 18720 11897 18748
rect 11848 18708 11854 18720
rect 11885 18717 11897 18720
rect 11931 18717 11943 18751
rect 11885 18711 11943 18717
rect 12158 18708 12164 18760
rect 12216 18748 12222 18760
rect 12802 18748 12808 18760
rect 12216 18720 12808 18748
rect 12216 18708 12222 18720
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 12912 18757 12940 18788
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 13998 18776 14004 18828
rect 14056 18816 14062 18828
rect 14458 18816 14464 18828
rect 14056 18788 14464 18816
rect 14056 18776 14062 18788
rect 14458 18776 14464 18788
rect 14516 18816 14522 18828
rect 14553 18819 14611 18825
rect 14553 18816 14565 18819
rect 14516 18788 14565 18816
rect 14516 18776 14522 18788
rect 14553 18785 14565 18788
rect 14599 18785 14611 18819
rect 14553 18779 14611 18785
rect 14918 18776 14924 18828
rect 14976 18816 14982 18828
rect 17129 18819 17187 18825
rect 17129 18816 17141 18819
rect 14976 18788 17141 18816
rect 14976 18776 14982 18788
rect 17129 18785 17141 18788
rect 17175 18785 17187 18819
rect 17678 18816 17684 18828
rect 17639 18788 17684 18816
rect 17129 18779 17187 18785
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 18233 18819 18291 18825
rect 18233 18785 18245 18819
rect 18279 18816 18291 18819
rect 20254 18816 20260 18828
rect 18279 18788 20116 18816
rect 20215 18788 20260 18816
rect 18279 18785 18291 18788
rect 18233 18779 18291 18785
rect 12897 18751 12955 18757
rect 12897 18717 12909 18751
rect 12943 18717 12955 18751
rect 12897 18711 12955 18717
rect 14829 18751 14887 18757
rect 14829 18717 14841 18751
rect 14875 18748 14887 18751
rect 15194 18748 15200 18760
rect 14875 18720 15200 18748
rect 14875 18717 14887 18720
rect 14829 18711 14887 18717
rect 15194 18708 15200 18720
rect 15252 18708 15258 18760
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 11333 18683 11391 18689
rect 8864 18652 9720 18680
rect 8846 18612 8852 18624
rect 8588 18584 8852 18612
rect 8846 18572 8852 18584
rect 8904 18572 8910 18624
rect 9306 18612 9312 18624
rect 9267 18584 9312 18612
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 9692 18612 9720 18652
rect 11333 18649 11345 18683
rect 11379 18680 11391 18683
rect 14185 18683 14243 18689
rect 11379 18652 12572 18680
rect 11379 18649 11391 18652
rect 11333 18643 11391 18649
rect 11698 18612 11704 18624
rect 9692 18584 11704 18612
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 12345 18615 12403 18621
rect 12345 18581 12357 18615
rect 12391 18612 12403 18615
rect 12434 18612 12440 18624
rect 12391 18584 12440 18612
rect 12391 18581 12403 18584
rect 12345 18575 12403 18581
rect 12434 18572 12440 18584
rect 12492 18572 12498 18624
rect 12544 18612 12572 18652
rect 14185 18649 14197 18683
rect 14231 18680 14243 18683
rect 15378 18680 15384 18692
rect 14231 18652 15384 18680
rect 14231 18649 14243 18652
rect 14185 18643 14243 18649
rect 15378 18640 15384 18652
rect 15436 18640 15442 18692
rect 12894 18612 12900 18624
rect 12544 18584 12900 18612
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 14090 18572 14096 18624
rect 14148 18612 14154 18624
rect 15488 18612 15516 18711
rect 18138 18708 18144 18760
rect 18196 18748 18202 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 18196 18720 19257 18748
rect 18196 18708 18202 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 16482 18640 16488 18692
rect 16540 18680 16546 18692
rect 18049 18683 18107 18689
rect 18049 18680 18061 18683
rect 16540 18652 18061 18680
rect 16540 18640 16546 18652
rect 18049 18649 18061 18652
rect 18095 18649 18107 18683
rect 19260 18680 19288 18711
rect 19426 18708 19432 18760
rect 19484 18748 19490 18760
rect 20088 18748 20116 18788
rect 20254 18776 20260 18788
rect 20312 18776 20318 18828
rect 20901 18819 20959 18825
rect 20901 18785 20913 18819
rect 20947 18816 20959 18819
rect 21358 18816 21364 18828
rect 20947 18788 21364 18816
rect 20947 18785 20959 18788
rect 20901 18779 20959 18785
rect 21358 18776 21364 18788
rect 21416 18776 21422 18828
rect 21082 18748 21088 18760
rect 19484 18720 19529 18748
rect 20088 18720 21088 18748
rect 19484 18708 19490 18720
rect 21082 18708 21088 18720
rect 21140 18708 21146 18760
rect 19797 18683 19855 18689
rect 19797 18680 19809 18683
rect 19260 18652 19809 18680
rect 18049 18643 18107 18649
rect 19797 18649 19809 18652
rect 19843 18649 19855 18683
rect 19797 18643 19855 18649
rect 15746 18612 15752 18624
rect 14148 18584 15752 18612
rect 14148 18572 14154 18584
rect 15746 18572 15752 18584
rect 15804 18572 15810 18624
rect 16574 18572 16580 18624
rect 16632 18612 16638 18624
rect 16853 18615 16911 18621
rect 16853 18612 16865 18615
rect 16632 18584 16865 18612
rect 16632 18572 16638 18584
rect 16853 18581 16865 18584
rect 16899 18581 16911 18615
rect 16853 18575 16911 18581
rect 18417 18615 18475 18621
rect 18417 18581 18429 18615
rect 18463 18612 18475 18615
rect 18690 18612 18696 18624
rect 18463 18584 18696 18612
rect 18463 18581 18475 18584
rect 18417 18575 18475 18581
rect 18690 18572 18696 18584
rect 18748 18572 18754 18624
rect 18785 18615 18843 18621
rect 18785 18581 18797 18615
rect 18831 18612 18843 18615
rect 20070 18612 20076 18624
rect 18831 18584 20076 18612
rect 18831 18581 18843 18584
rect 18785 18575 18843 18581
rect 20070 18572 20076 18584
rect 20128 18572 20134 18624
rect 20438 18612 20444 18624
rect 20399 18584 20444 18612
rect 20438 18572 20444 18584
rect 20496 18572 20502 18624
rect 21085 18615 21143 18621
rect 21085 18581 21097 18615
rect 21131 18612 21143 18615
rect 21174 18612 21180 18624
rect 21131 18584 21180 18612
rect 21131 18581 21143 18584
rect 21085 18575 21143 18581
rect 21174 18572 21180 18584
rect 21232 18572 21238 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 7006 18368 7012 18420
rect 7064 18408 7070 18420
rect 7101 18411 7159 18417
rect 7101 18408 7113 18411
rect 7064 18380 7113 18408
rect 7064 18368 7070 18380
rect 7101 18377 7113 18380
rect 7147 18377 7159 18411
rect 7101 18371 7159 18377
rect 3602 18300 3608 18352
rect 3660 18340 3666 18352
rect 6546 18340 6552 18352
rect 3660 18312 6552 18340
rect 3660 18300 3666 18312
rect 6546 18300 6552 18312
rect 6604 18300 6610 18352
rect 1946 18232 1952 18284
rect 2004 18272 2010 18284
rect 7006 18272 7012 18284
rect 2004 18244 7012 18272
rect 2004 18232 2010 18244
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 5258 18164 5264 18216
rect 5316 18204 5322 18216
rect 6914 18204 6920 18216
rect 5316 18176 6920 18204
rect 5316 18164 5322 18176
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 7116 18204 7144 18371
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 8202 18408 8208 18420
rect 7616 18380 8208 18408
rect 7616 18368 7622 18380
rect 8202 18368 8208 18380
rect 8260 18408 8266 18420
rect 11146 18408 11152 18420
rect 8260 18380 11152 18408
rect 8260 18368 8266 18380
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 12069 18411 12127 18417
rect 12069 18377 12081 18411
rect 12115 18408 12127 18411
rect 12158 18408 12164 18420
rect 12115 18380 12164 18408
rect 12115 18377 12127 18380
rect 12069 18371 12127 18377
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 12253 18411 12311 18417
rect 12253 18377 12265 18411
rect 12299 18408 12311 18411
rect 13998 18408 14004 18420
rect 12299 18380 14004 18408
rect 12299 18377 12311 18380
rect 12253 18371 12311 18377
rect 13998 18368 14004 18380
rect 14056 18368 14062 18420
rect 14185 18411 14243 18417
rect 14185 18377 14197 18411
rect 14231 18408 14243 18411
rect 15657 18411 15715 18417
rect 14231 18380 15240 18408
rect 14231 18377 14243 18380
rect 14185 18371 14243 18377
rect 7469 18343 7527 18349
rect 7469 18309 7481 18343
rect 7515 18340 7527 18343
rect 8662 18340 8668 18352
rect 7515 18312 8668 18340
rect 7515 18309 7527 18312
rect 7469 18303 7527 18309
rect 8662 18300 8668 18312
rect 8720 18300 8726 18352
rect 10045 18343 10103 18349
rect 10045 18309 10057 18343
rect 10091 18340 10103 18343
rect 11238 18340 11244 18352
rect 10091 18312 11244 18340
rect 10091 18309 10103 18312
rect 10045 18303 10103 18309
rect 11238 18300 11244 18312
rect 11296 18300 11302 18352
rect 11790 18300 11796 18352
rect 11848 18340 11854 18352
rect 13906 18340 13912 18352
rect 11848 18312 13768 18340
rect 13867 18312 13912 18340
rect 11848 18300 11854 18312
rect 8113 18275 8171 18281
rect 8113 18241 8125 18275
rect 8159 18272 8171 18275
rect 8202 18272 8208 18284
rect 8159 18244 8208 18272
rect 8159 18241 8171 18244
rect 8113 18235 8171 18241
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 10060 18244 12265 18272
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 7116 18176 7849 18204
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 8665 18207 8723 18213
rect 8665 18173 8677 18207
rect 8711 18204 8723 18207
rect 9214 18204 9220 18216
rect 8711 18176 9220 18204
rect 8711 18173 8723 18176
rect 8665 18167 8723 18173
rect 9214 18164 9220 18176
rect 9272 18164 9278 18216
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 10060 18204 10088 18244
rect 12253 18241 12265 18244
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 12989 18275 13047 18281
rect 12989 18272 13001 18275
rect 12584 18244 13001 18272
rect 12584 18232 12590 18244
rect 12989 18241 13001 18244
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 9456 18176 10088 18204
rect 9456 18164 9462 18176
rect 10318 18164 10324 18216
rect 10376 18204 10382 18216
rect 10594 18204 10600 18216
rect 10376 18176 10600 18204
rect 10376 18164 10382 18176
rect 10594 18164 10600 18176
rect 10652 18164 10658 18216
rect 11241 18207 11299 18213
rect 11241 18173 11253 18207
rect 11287 18204 11299 18207
rect 12802 18204 12808 18216
rect 11287 18176 12725 18204
rect 12763 18176 12808 18204
rect 11287 18173 11299 18176
rect 11241 18167 11299 18173
rect 5810 18096 5816 18148
rect 5868 18136 5874 18148
rect 7098 18136 7104 18148
rect 5868 18108 7104 18136
rect 5868 18096 5874 18108
rect 7098 18096 7104 18108
rect 7156 18136 7162 18148
rect 7929 18139 7987 18145
rect 7929 18136 7941 18139
rect 7156 18108 7941 18136
rect 7156 18096 7162 18108
rect 7929 18105 7941 18108
rect 7975 18105 7987 18139
rect 7929 18099 7987 18105
rect 8932 18139 8990 18145
rect 8932 18105 8944 18139
rect 8978 18136 8990 18139
rect 9030 18136 9036 18148
rect 8978 18108 9036 18136
rect 8978 18105 8990 18108
rect 8932 18099 8990 18105
rect 9030 18096 9036 18108
rect 9088 18096 9094 18148
rect 9582 18096 9588 18148
rect 9640 18136 9646 18148
rect 9858 18136 9864 18148
rect 9640 18108 9864 18136
rect 9640 18096 9646 18108
rect 9858 18096 9864 18108
rect 9916 18096 9922 18148
rect 10226 18096 10232 18148
rect 10284 18136 10290 18148
rect 11517 18139 11575 18145
rect 10284 18108 10456 18136
rect 10284 18096 10290 18108
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 6178 18068 6184 18080
rect 4856 18040 6184 18068
rect 4856 18028 4862 18040
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 6362 18028 6368 18080
rect 6420 18068 6426 18080
rect 10134 18068 10140 18080
rect 6420 18040 10140 18068
rect 6420 18028 6426 18040
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 10318 18068 10324 18080
rect 10279 18040 10324 18068
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 10428 18068 10456 18108
rect 11517 18105 11529 18139
rect 11563 18136 11575 18139
rect 12697 18136 12725 18176
rect 12802 18164 12808 18176
rect 12860 18164 12866 18216
rect 12894 18164 12900 18216
rect 12952 18204 12958 18216
rect 13740 18213 13768 18312
rect 13906 18300 13912 18312
rect 13964 18300 13970 18352
rect 15212 18340 15240 18380
rect 15657 18377 15669 18411
rect 15703 18408 15715 18411
rect 15838 18408 15844 18420
rect 15703 18380 15844 18408
rect 15703 18377 15715 18380
rect 15657 18371 15715 18377
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 16209 18411 16267 18417
rect 16209 18377 16221 18411
rect 16255 18408 16267 18411
rect 20530 18408 20536 18420
rect 16255 18380 20536 18408
rect 16255 18377 16267 18380
rect 16209 18371 16267 18377
rect 20530 18368 20536 18380
rect 20588 18368 20594 18420
rect 16482 18340 16488 18352
rect 15212 18312 16488 18340
rect 16482 18300 16488 18312
rect 16540 18300 16546 18352
rect 16577 18343 16635 18349
rect 16577 18309 16589 18343
rect 16623 18340 16635 18343
rect 18046 18340 18052 18352
rect 16623 18312 18052 18340
rect 16623 18309 16635 18312
rect 16577 18303 16635 18309
rect 18046 18300 18052 18312
rect 18104 18300 18110 18352
rect 19705 18343 19763 18349
rect 19705 18309 19717 18343
rect 19751 18340 19763 18343
rect 20898 18340 20904 18352
rect 19751 18312 20904 18340
rect 19751 18309 19763 18312
rect 19705 18303 19763 18309
rect 20898 18300 20904 18312
rect 20956 18300 20962 18352
rect 17218 18272 17224 18284
rect 17179 18244 17224 18272
rect 17218 18232 17224 18244
rect 17276 18232 17282 18284
rect 19058 18232 19064 18284
rect 19116 18272 19122 18284
rect 19334 18272 19340 18284
rect 19116 18244 19340 18272
rect 19116 18232 19122 18244
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 20257 18275 20315 18281
rect 20257 18272 20269 18275
rect 19484 18244 20269 18272
rect 19484 18232 19490 18244
rect 20257 18241 20269 18244
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 13725 18207 13783 18213
rect 12952 18176 12997 18204
rect 12952 18164 12958 18176
rect 13725 18173 13737 18207
rect 13771 18173 13783 18207
rect 13725 18167 13783 18173
rect 13814 18164 13820 18216
rect 13872 18204 13878 18216
rect 14090 18204 14096 18216
rect 13872 18176 14096 18204
rect 13872 18164 13878 18176
rect 14090 18164 14096 18176
rect 14148 18204 14154 18216
rect 14277 18207 14335 18213
rect 14277 18204 14289 18207
rect 14148 18176 14289 18204
rect 14148 18164 14154 18176
rect 14277 18173 14289 18176
rect 14323 18173 14335 18207
rect 16025 18207 16083 18213
rect 16025 18204 16037 18207
rect 14277 18167 14335 18173
rect 14476 18176 16037 18204
rect 13170 18136 13176 18148
rect 11563 18108 12572 18136
rect 12697 18108 13176 18136
rect 11563 18105 11575 18108
rect 11517 18099 11575 18105
rect 10778 18068 10784 18080
rect 10428 18040 10784 18068
rect 10778 18028 10784 18040
rect 10836 18068 10842 18080
rect 10873 18071 10931 18077
rect 10873 18068 10885 18071
rect 10836 18040 10885 18068
rect 10836 18028 10842 18040
rect 10873 18037 10885 18040
rect 10919 18037 10931 18071
rect 10873 18031 10931 18037
rect 12158 18028 12164 18080
rect 12216 18068 12222 18080
rect 12437 18071 12495 18077
rect 12437 18068 12449 18071
rect 12216 18040 12449 18068
rect 12216 18028 12222 18040
rect 12437 18037 12449 18040
rect 12483 18037 12495 18071
rect 12544 18068 12572 18108
rect 13170 18096 13176 18108
rect 13228 18096 13234 18148
rect 13262 18096 13268 18148
rect 13320 18136 13326 18148
rect 14476 18136 14504 18176
rect 16025 18173 16037 18176
rect 16071 18173 16083 18207
rect 16025 18167 16083 18173
rect 13320 18108 14504 18136
rect 14544 18139 14602 18145
rect 13320 18096 13326 18108
rect 14544 18105 14556 18139
rect 14590 18136 14602 18139
rect 15194 18136 15200 18148
rect 14590 18108 15200 18136
rect 14590 18105 14602 18108
rect 14544 18099 14602 18105
rect 15194 18096 15200 18108
rect 15252 18096 15258 18148
rect 16040 18136 16068 18167
rect 16666 18164 16672 18216
rect 16724 18204 16730 18216
rect 16945 18207 17003 18213
rect 16945 18204 16957 18207
rect 16724 18176 16957 18204
rect 16724 18164 16730 18176
rect 16945 18173 16957 18176
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 17862 18164 17868 18216
rect 17920 18204 17926 18216
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 17920 18176 18061 18204
rect 17920 18164 17926 18176
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 18690 18164 18696 18216
rect 18748 18204 18754 18216
rect 20070 18204 20076 18216
rect 18748 18176 19196 18204
rect 20031 18176 20076 18204
rect 18748 18164 18754 18176
rect 17589 18139 17647 18145
rect 17589 18136 17601 18139
rect 16040 18108 17601 18136
rect 17589 18105 17601 18108
rect 17635 18136 17647 18139
rect 18138 18136 18144 18148
rect 17635 18108 18144 18136
rect 17635 18105 17647 18108
rect 17589 18099 17647 18105
rect 18138 18096 18144 18108
rect 18196 18096 18202 18148
rect 18316 18139 18374 18145
rect 18316 18105 18328 18139
rect 18362 18136 18374 18139
rect 19058 18136 19064 18148
rect 18362 18108 19064 18136
rect 18362 18105 18374 18108
rect 18316 18099 18374 18105
rect 19058 18096 19064 18108
rect 19116 18096 19122 18148
rect 19168 18136 19196 18176
rect 20070 18164 20076 18176
rect 20128 18164 20134 18216
rect 20806 18204 20812 18216
rect 20767 18176 20812 18204
rect 20806 18164 20812 18176
rect 20864 18164 20870 18216
rect 22094 18136 22100 18148
rect 19168 18108 22100 18136
rect 22094 18096 22100 18108
rect 22152 18096 22158 18148
rect 14185 18071 14243 18077
rect 14185 18068 14197 18071
rect 12544 18040 14197 18068
rect 12437 18031 12495 18037
rect 14185 18037 14197 18040
rect 14231 18037 14243 18071
rect 14185 18031 14243 18037
rect 17034 18028 17040 18080
rect 17092 18068 17098 18080
rect 19426 18068 19432 18080
rect 17092 18040 17137 18068
rect 19387 18040 19432 18068
rect 17092 18028 17098 18040
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 20162 18068 20168 18080
rect 20123 18040 20168 18068
rect 20162 18028 20168 18040
rect 20220 18028 20226 18080
rect 20990 18068 20996 18080
rect 20951 18040 20996 18068
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 7098 17864 7104 17876
rect 7059 17836 7104 17864
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 9030 17864 9036 17876
rect 8991 17836 9036 17864
rect 9030 17824 9036 17836
rect 9088 17824 9094 17876
rect 9677 17867 9735 17873
rect 9677 17833 9689 17867
rect 9723 17864 9735 17867
rect 11149 17867 11207 17873
rect 11149 17864 11161 17867
rect 9723 17836 11161 17864
rect 9723 17833 9735 17836
rect 9677 17827 9735 17833
rect 11149 17833 11161 17836
rect 11195 17833 11207 17867
rect 11149 17827 11207 17833
rect 11698 17824 11704 17876
rect 11756 17864 11762 17876
rect 13817 17867 13875 17873
rect 13817 17864 13829 17867
rect 11756 17836 13829 17864
rect 11756 17824 11762 17836
rect 13817 17833 13829 17836
rect 13863 17833 13875 17867
rect 16758 17864 16764 17876
rect 13817 17827 13875 17833
rect 14476 17836 16764 17864
rect 8662 17756 8668 17808
rect 8720 17796 8726 17808
rect 10137 17799 10195 17805
rect 10137 17796 10149 17799
rect 8720 17768 10149 17796
rect 8720 17756 8726 17768
rect 10137 17765 10149 17768
rect 10183 17765 10195 17799
rect 10137 17759 10195 17765
rect 13630 17756 13636 17808
rect 13688 17796 13694 17808
rect 13725 17799 13783 17805
rect 13725 17796 13737 17799
rect 13688 17768 13737 17796
rect 13688 17756 13694 17768
rect 13725 17765 13737 17768
rect 13771 17765 13783 17799
rect 14476 17796 14504 17836
rect 16758 17824 16764 17836
rect 16816 17824 16822 17876
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 17405 17867 17463 17873
rect 17405 17864 17417 17867
rect 17276 17836 17417 17864
rect 17276 17824 17282 17836
rect 17405 17833 17417 17836
rect 17451 17833 17463 17867
rect 17405 17827 17463 17833
rect 19337 17867 19395 17873
rect 19337 17833 19349 17867
rect 19383 17864 19395 17867
rect 20162 17864 20168 17876
rect 19383 17836 20168 17864
rect 19383 17833 19395 17836
rect 19337 17827 19395 17833
rect 16292 17799 16350 17805
rect 13725 17759 13783 17765
rect 13832 17768 14504 17796
rect 14568 17768 16252 17796
rect 7926 17737 7932 17740
rect 7920 17728 7932 17737
rect 7887 17700 7932 17728
rect 7920 17691 7932 17700
rect 7984 17728 7990 17740
rect 8202 17728 8208 17740
rect 7984 17700 8208 17728
rect 7926 17688 7932 17691
rect 7984 17688 7990 17700
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 8478 17688 8484 17740
rect 8536 17728 8542 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 8536 17700 10057 17728
rect 8536 17688 8542 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 11054 17728 11060 17740
rect 11015 17700 11060 17728
rect 10045 17691 10103 17697
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 12158 17728 12164 17740
rect 12119 17700 12164 17728
rect 12158 17688 12164 17700
rect 12216 17688 12222 17740
rect 12986 17688 12992 17740
rect 13044 17728 13050 17740
rect 13832 17728 13860 17768
rect 14568 17728 14596 17768
rect 13044 17700 13860 17728
rect 13924 17700 14596 17728
rect 13044 17688 13050 17700
rect 7653 17663 7711 17669
rect 7653 17629 7665 17663
rect 7699 17629 7711 17663
rect 7653 17623 7711 17629
rect 6270 17484 6276 17536
rect 6328 17524 6334 17536
rect 6733 17527 6791 17533
rect 6733 17524 6745 17527
rect 6328 17496 6745 17524
rect 6328 17484 6334 17496
rect 6733 17493 6745 17496
rect 6779 17493 6791 17527
rect 6733 17487 6791 17493
rect 7282 17484 7288 17536
rect 7340 17524 7346 17536
rect 7668 17524 7696 17623
rect 9030 17620 9036 17672
rect 9088 17660 9094 17672
rect 9582 17660 9588 17672
rect 9088 17632 9588 17660
rect 9088 17620 9094 17632
rect 9582 17620 9588 17632
rect 9640 17660 9646 17672
rect 10229 17663 10287 17669
rect 10229 17660 10241 17663
rect 9640 17632 10241 17660
rect 9640 17620 9646 17632
rect 10229 17629 10241 17632
rect 10275 17629 10287 17663
rect 11238 17660 11244 17672
rect 11199 17632 11244 17660
rect 10229 17623 10287 17629
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17660 12495 17663
rect 13924 17660 13952 17700
rect 14642 17688 14648 17740
rect 14700 17728 14706 17740
rect 15286 17728 15292 17740
rect 14700 17700 14745 17728
rect 15247 17700 15292 17728
rect 14700 17688 14706 17700
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 15746 17688 15752 17740
rect 15804 17728 15810 17740
rect 16025 17731 16083 17737
rect 16025 17728 16037 17731
rect 15804 17700 16037 17728
rect 15804 17688 15810 17700
rect 16025 17697 16037 17700
rect 16071 17697 16083 17731
rect 16224 17728 16252 17768
rect 16292 17765 16304 17799
rect 16338 17796 16350 17799
rect 16574 17796 16580 17808
rect 16338 17768 16580 17796
rect 16338 17765 16350 17768
rect 16292 17759 16350 17765
rect 16574 17756 16580 17768
rect 16632 17756 16638 17808
rect 17420 17796 17448 17827
rect 20162 17824 20168 17836
rect 20220 17824 20226 17876
rect 20346 17864 20352 17876
rect 20307 17836 20352 17864
rect 20346 17824 20352 17836
rect 20404 17824 20410 17876
rect 20806 17864 20812 17876
rect 20456 17836 20812 17864
rect 17926 17799 17984 17805
rect 17926 17796 17938 17799
rect 17420 17768 17938 17796
rect 17926 17765 17938 17768
rect 17972 17765 17984 17799
rect 20456 17796 20484 17836
rect 20806 17824 20812 17836
rect 20864 17824 20870 17876
rect 17926 17759 17984 17765
rect 18064 17768 20484 17796
rect 18064 17728 18092 17768
rect 20714 17756 20720 17808
rect 20772 17796 20778 17808
rect 21177 17799 21235 17805
rect 21177 17796 21189 17799
rect 20772 17768 21189 17796
rect 20772 17756 20778 17768
rect 21177 17765 21189 17768
rect 21223 17765 21235 17799
rect 21177 17759 21235 17765
rect 16224 17700 18092 17728
rect 16025 17691 16083 17697
rect 18230 17688 18236 17740
rect 18288 17728 18294 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 18288 17700 19717 17728
rect 18288 17688 18294 17700
rect 19705 17697 19717 17700
rect 19751 17697 19763 17731
rect 20898 17728 20904 17740
rect 20859 17700 20904 17728
rect 19705 17691 19763 17697
rect 20898 17688 20904 17700
rect 20956 17688 20962 17740
rect 12483 17632 13952 17660
rect 14001 17663 14059 17669
rect 12483 17629 12495 17632
rect 12437 17623 12495 17629
rect 14001 17629 14013 17663
rect 14047 17660 14059 17663
rect 14090 17660 14096 17672
rect 14047 17632 14096 17660
rect 14047 17629 14059 17632
rect 14001 17623 14059 17629
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 15562 17660 15568 17672
rect 15523 17632 15568 17660
rect 15562 17620 15568 17632
rect 15620 17620 15626 17672
rect 17586 17620 17592 17672
rect 17644 17660 17650 17672
rect 17681 17663 17739 17669
rect 17681 17660 17693 17663
rect 17644 17632 17693 17660
rect 17644 17620 17650 17632
rect 17681 17629 17693 17632
rect 17727 17629 17739 17663
rect 17681 17623 17739 17629
rect 18690 17620 18696 17672
rect 18748 17660 18754 17672
rect 19797 17663 19855 17669
rect 19797 17660 19809 17663
rect 18748 17632 19809 17660
rect 18748 17620 18754 17632
rect 19797 17629 19809 17632
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 19889 17663 19947 17669
rect 19889 17629 19901 17663
rect 19935 17629 19947 17663
rect 19889 17623 19947 17629
rect 9306 17552 9312 17604
rect 9364 17592 9370 17604
rect 19058 17592 19064 17604
rect 9364 17564 16068 17592
rect 18971 17564 19064 17592
rect 9364 17552 9370 17564
rect 9214 17524 9220 17536
rect 7340 17496 9220 17524
rect 7340 17484 7346 17496
rect 9214 17484 9220 17496
rect 9272 17484 9278 17536
rect 10502 17484 10508 17536
rect 10560 17524 10566 17536
rect 10689 17527 10747 17533
rect 10689 17524 10701 17527
rect 10560 17496 10701 17524
rect 10560 17484 10566 17496
rect 10689 17493 10701 17496
rect 10735 17493 10747 17527
rect 11790 17524 11796 17536
rect 11751 17496 11796 17524
rect 10689 17487 10747 17493
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 13078 17524 13084 17536
rect 13039 17496 13084 17524
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 13357 17527 13415 17533
rect 13357 17493 13369 17527
rect 13403 17524 13415 17527
rect 14550 17524 14556 17536
rect 13403 17496 14556 17524
rect 13403 17493 13415 17496
rect 13357 17487 13415 17493
rect 14550 17484 14556 17496
rect 14608 17484 14614 17536
rect 14826 17524 14832 17536
rect 14787 17496 14832 17524
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 16040 17524 16068 17564
rect 19058 17552 19064 17564
rect 19116 17592 19122 17604
rect 19904 17592 19932 17623
rect 19116 17564 19932 17592
rect 19116 17552 19122 17564
rect 17678 17524 17684 17536
rect 16040 17496 17684 17524
rect 17678 17484 17684 17496
rect 17736 17484 17742 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 7282 17320 7288 17332
rect 7024 17292 7288 17320
rect 7024 17193 7052 17292
rect 7282 17280 7288 17292
rect 7340 17280 7346 17332
rect 7926 17280 7932 17332
rect 7984 17320 7990 17332
rect 8389 17323 8447 17329
rect 8389 17320 8401 17323
rect 7984 17292 8401 17320
rect 7984 17280 7990 17292
rect 8389 17289 8401 17292
rect 8435 17289 8447 17323
rect 9125 17323 9183 17329
rect 9125 17320 9137 17323
rect 8389 17283 8447 17289
rect 8956 17292 9137 17320
rect 7009 17187 7067 17193
rect 7009 17153 7021 17187
rect 7055 17153 7067 17187
rect 7009 17147 7067 17153
rect 8386 17144 8392 17196
rect 8444 17184 8450 17196
rect 8956 17184 8984 17292
rect 9125 17289 9137 17292
rect 9171 17320 9183 17323
rect 9306 17320 9312 17332
rect 9171 17292 9312 17320
rect 9171 17289 9183 17292
rect 9125 17283 9183 17289
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 9493 17323 9551 17329
rect 9493 17289 9505 17323
rect 9539 17320 9551 17323
rect 11054 17320 11060 17332
rect 9539 17292 11060 17320
rect 9539 17289 9551 17292
rect 9493 17283 9551 17289
rect 11054 17280 11060 17292
rect 11112 17280 11118 17332
rect 11333 17323 11391 17329
rect 11333 17289 11345 17323
rect 11379 17320 11391 17323
rect 12437 17323 12495 17329
rect 11379 17292 12296 17320
rect 11379 17289 11391 17292
rect 11333 17283 11391 17289
rect 9030 17212 9036 17264
rect 9088 17252 9094 17264
rect 11698 17252 11704 17264
rect 9088 17224 11704 17252
rect 9088 17212 9094 17224
rect 11698 17212 11704 17224
rect 11756 17212 11762 17264
rect 12268 17252 12296 17292
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12894 17320 12900 17332
rect 12483 17292 12900 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12894 17280 12900 17292
rect 12952 17280 12958 17332
rect 13078 17280 13084 17332
rect 13136 17320 13142 17332
rect 14642 17320 14648 17332
rect 13136 17292 14648 17320
rect 13136 17280 13142 17292
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 16577 17323 16635 17329
rect 15620 17292 16252 17320
rect 15620 17280 15626 17292
rect 12618 17252 12624 17264
rect 11808 17224 12204 17252
rect 12268 17224 12624 17252
rect 8444 17156 8984 17184
rect 8444 17144 8450 17156
rect 9582 17144 9588 17196
rect 9640 17184 9646 17196
rect 11808 17193 11836 17224
rect 10045 17187 10103 17193
rect 10045 17184 10057 17187
rect 9640 17156 10057 17184
rect 9640 17144 9646 17156
rect 10045 17153 10057 17156
rect 10091 17153 10103 17187
rect 10045 17147 10103 17153
rect 11793 17187 11851 17193
rect 11793 17153 11805 17187
rect 11839 17153 11851 17187
rect 11974 17184 11980 17196
rect 11935 17156 11980 17184
rect 11793 17147 11851 17153
rect 11974 17144 11980 17156
rect 12032 17144 12038 17196
rect 12176 17184 12204 17224
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 14277 17255 14335 17261
rect 14277 17221 14289 17255
rect 14323 17221 14335 17255
rect 14277 17215 14335 17221
rect 12176 17156 12296 17184
rect 5902 17076 5908 17128
rect 5960 17116 5966 17128
rect 6638 17116 6644 17128
rect 5960 17088 6644 17116
rect 5960 17076 5966 17088
rect 6638 17076 6644 17088
rect 6696 17116 6702 17128
rect 7742 17116 7748 17128
rect 6696 17088 7748 17116
rect 6696 17076 6702 17088
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 9306 17076 9312 17128
rect 9364 17116 9370 17128
rect 9861 17119 9919 17125
rect 9364 17088 9812 17116
rect 9364 17076 9370 17088
rect 7276 17051 7334 17057
rect 7276 17017 7288 17051
rect 7322 17048 7334 17051
rect 9490 17048 9496 17060
rect 7322 17020 9496 17048
rect 7322 17017 7334 17020
rect 7276 17011 7334 17017
rect 9490 17008 9496 17020
rect 9548 17008 9554 17060
rect 9784 17048 9812 17088
rect 9861 17085 9873 17119
rect 9907 17116 9919 17119
rect 10318 17116 10324 17128
rect 9907 17088 10324 17116
rect 9907 17085 9919 17088
rect 9861 17079 9919 17085
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 10502 17116 10508 17128
rect 10463 17088 10508 17116
rect 10502 17076 10508 17088
rect 10560 17076 10566 17128
rect 11701 17119 11759 17125
rect 11701 17085 11713 17119
rect 11747 17116 11759 17119
rect 12161 17119 12219 17125
rect 12161 17116 12173 17119
rect 11747 17088 12173 17116
rect 11747 17085 11759 17088
rect 11701 17079 11759 17085
rect 12161 17085 12173 17088
rect 12207 17085 12219 17119
rect 12268 17116 12296 17156
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12897 17187 12955 17193
rect 12897 17184 12909 17187
rect 12492 17156 12909 17184
rect 12492 17144 12498 17156
rect 12897 17153 12909 17156
rect 12943 17153 12955 17187
rect 14292 17184 14320 17215
rect 14366 17212 14372 17264
rect 14424 17252 14430 17264
rect 14553 17255 14611 17261
rect 14553 17252 14565 17255
rect 14424 17224 14565 17252
rect 14424 17212 14430 17224
rect 14553 17221 14565 17224
rect 14599 17221 14611 17255
rect 14734 17252 14740 17264
rect 14647 17224 14740 17252
rect 14553 17215 14611 17221
rect 14660 17184 14688 17224
rect 14734 17212 14740 17224
rect 14792 17252 14798 17264
rect 16224 17252 16252 17292
rect 16577 17289 16589 17323
rect 16623 17320 16635 17323
rect 16666 17320 16672 17332
rect 16623 17292 16672 17320
rect 16623 17289 16635 17292
rect 16577 17283 16635 17289
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 21358 17320 21364 17332
rect 16776 17292 21364 17320
rect 16776 17252 16804 17292
rect 21358 17280 21364 17292
rect 21416 17280 21422 17332
rect 14792 17224 16160 17252
rect 16224 17224 16804 17252
rect 16960 17224 17172 17252
rect 14792 17212 14798 17224
rect 15194 17184 15200 17196
rect 14292 17156 14688 17184
rect 15107 17156 15200 17184
rect 12897 17147 12955 17153
rect 15194 17144 15200 17156
rect 15252 17184 15258 17196
rect 15838 17184 15844 17196
rect 15252 17156 15844 17184
rect 15252 17144 15258 17156
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 16132 17193 16160 17224
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 16960 17184 16988 17224
rect 17144 17193 17172 17224
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 18230 17252 18236 17264
rect 18012 17224 18236 17252
rect 18012 17212 18018 17224
rect 18230 17212 18236 17224
rect 18288 17212 18294 17264
rect 16632 17156 16988 17184
rect 17129 17187 17187 17193
rect 16632 17144 16638 17156
rect 17129 17153 17141 17187
rect 17175 17184 17187 17187
rect 17218 17184 17224 17196
rect 17175 17156 17224 17184
rect 17175 17153 17187 17156
rect 17129 17147 17187 17153
rect 17218 17144 17224 17156
rect 17276 17144 17282 17196
rect 17862 17144 17868 17196
rect 17920 17184 17926 17196
rect 18325 17187 18383 17193
rect 18325 17184 18337 17187
rect 17920 17156 18337 17184
rect 17920 17144 17926 17156
rect 18325 17153 18337 17156
rect 18371 17153 18383 17187
rect 20254 17184 20260 17196
rect 20215 17156 20260 17184
rect 18325 17147 18383 17153
rect 20254 17144 20260 17156
rect 20312 17144 20318 17196
rect 21082 17184 21088 17196
rect 21043 17156 21088 17184
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 12526 17116 12532 17128
rect 12268 17088 12532 17116
rect 12161 17079 12219 17085
rect 12526 17076 12532 17088
rect 12584 17076 12590 17128
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17116 12679 17119
rect 12986 17116 12992 17128
rect 12667 17088 12992 17116
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 12986 17076 12992 17088
rect 13044 17076 13050 17128
rect 13164 17119 13222 17125
rect 13164 17085 13176 17119
rect 13210 17116 13222 17119
rect 14090 17116 14096 17128
rect 13210 17088 14096 17116
rect 13210 17085 13222 17088
rect 13164 17079 13222 17085
rect 14090 17076 14096 17088
rect 14148 17076 14154 17128
rect 17954 17116 17960 17128
rect 14568 17088 17960 17116
rect 9953 17051 10011 17057
rect 9953 17048 9965 17051
rect 9784 17020 9965 17048
rect 9953 17017 9965 17020
rect 9999 17017 10011 17051
rect 9953 17011 10011 17017
rect 10781 17051 10839 17057
rect 10781 17017 10793 17051
rect 10827 17048 10839 17051
rect 14568 17048 14596 17088
rect 17954 17076 17960 17088
rect 18012 17076 18018 17128
rect 18592 17119 18650 17125
rect 18592 17085 18604 17119
rect 18638 17116 18650 17119
rect 19426 17116 19432 17128
rect 18638 17088 19432 17116
rect 18638 17085 18650 17088
rect 18592 17079 18650 17085
rect 19426 17076 19432 17088
rect 19484 17076 19490 17128
rect 20073 17119 20131 17125
rect 20073 17085 20085 17119
rect 20119 17085 20131 17119
rect 20073 17079 20131 17085
rect 10827 17020 14596 17048
rect 10827 17017 10839 17020
rect 10781 17011 10839 17017
rect 14642 17008 14648 17060
rect 14700 17048 14706 17060
rect 15013 17051 15071 17057
rect 15013 17048 15025 17051
rect 14700 17020 15025 17048
rect 14700 17008 14706 17020
rect 15013 17017 15025 17020
rect 15059 17017 15071 17051
rect 15013 17011 15071 17017
rect 18046 17008 18052 17060
rect 18104 17048 18110 17060
rect 20088 17048 20116 17079
rect 20346 17076 20352 17128
rect 20404 17116 20410 17128
rect 20809 17119 20867 17125
rect 20809 17116 20821 17119
rect 20404 17088 20821 17116
rect 20404 17076 20410 17088
rect 20809 17085 20821 17088
rect 20855 17085 20867 17119
rect 20809 17079 20867 17085
rect 18104 17020 20116 17048
rect 18104 17008 18110 17020
rect 6457 16983 6515 16989
rect 6457 16949 6469 16983
rect 6503 16980 6515 16983
rect 7190 16980 7196 16992
rect 6503 16952 7196 16980
rect 6503 16949 6515 16952
rect 6457 16943 6515 16949
rect 7190 16940 7196 16952
rect 7248 16980 7254 16992
rect 8478 16980 8484 16992
rect 7248 16952 8484 16980
rect 7248 16940 7254 16952
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 8754 16940 8760 16992
rect 8812 16980 8818 16992
rect 8849 16983 8907 16989
rect 8849 16980 8861 16983
rect 8812 16952 8861 16980
rect 8812 16940 8818 16952
rect 8849 16949 8861 16952
rect 8895 16980 8907 16983
rect 9030 16980 9036 16992
rect 8895 16952 9036 16980
rect 8895 16949 8907 16952
rect 8849 16943 8907 16949
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 12161 16983 12219 16989
rect 12161 16949 12173 16983
rect 12207 16980 12219 16983
rect 12802 16980 12808 16992
rect 12207 16952 12808 16980
rect 12207 16949 12219 16952
rect 12161 16943 12219 16949
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 13446 16940 13452 16992
rect 13504 16980 13510 16992
rect 13814 16980 13820 16992
rect 13504 16952 13820 16980
rect 13504 16940 13510 16952
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 13998 16940 14004 16992
rect 14056 16980 14062 16992
rect 14458 16980 14464 16992
rect 14056 16952 14464 16980
rect 14056 16940 14062 16952
rect 14458 16940 14464 16952
rect 14516 16980 14522 16992
rect 14921 16983 14979 16989
rect 14921 16980 14933 16983
rect 14516 16952 14933 16980
rect 14516 16940 14522 16952
rect 14921 16949 14933 16952
rect 14967 16949 14979 16983
rect 15562 16980 15568 16992
rect 15523 16952 15568 16980
rect 14921 16943 14979 16949
rect 15562 16940 15568 16952
rect 15620 16940 15626 16992
rect 15930 16980 15936 16992
rect 15891 16952 15936 16980
rect 15930 16940 15936 16952
rect 15988 16940 15994 16992
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 16942 16980 16948 16992
rect 16080 16952 16125 16980
rect 16903 16952 16948 16980
rect 16080 16940 16086 16952
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17037 16983 17095 16989
rect 17037 16949 17049 16983
rect 17083 16980 17095 16983
rect 17126 16980 17132 16992
rect 17083 16952 17132 16980
rect 17083 16949 17095 16952
rect 17037 16943 17095 16949
rect 17126 16940 17132 16952
rect 17184 16980 17190 16992
rect 17589 16983 17647 16989
rect 17589 16980 17601 16983
rect 17184 16952 17601 16980
rect 17184 16940 17190 16952
rect 17589 16949 17601 16952
rect 17635 16949 17647 16983
rect 17589 16943 17647 16949
rect 17678 16940 17684 16992
rect 17736 16980 17742 16992
rect 19334 16980 19340 16992
rect 17736 16952 19340 16980
rect 17736 16940 17742 16952
rect 19334 16940 19340 16952
rect 19392 16940 19398 16992
rect 19702 16980 19708 16992
rect 19663 16952 19708 16980
rect 19702 16940 19708 16952
rect 19760 16940 19766 16992
rect 20254 16940 20260 16992
rect 20312 16980 20318 16992
rect 21450 16980 21456 16992
rect 20312 16952 21456 16980
rect 20312 16940 20318 16952
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 5902 16776 5908 16788
rect 5863 16748 5908 16776
rect 5902 16736 5908 16748
rect 5960 16736 5966 16788
rect 7009 16779 7067 16785
rect 7009 16745 7021 16779
rect 7055 16776 7067 16779
rect 7742 16776 7748 16788
rect 7055 16748 7748 16776
rect 7055 16745 7067 16748
rect 7009 16739 7067 16745
rect 7742 16736 7748 16748
rect 7800 16776 7806 16788
rect 8938 16776 8944 16788
rect 7800 16748 8944 16776
rect 7800 16736 7806 16748
rect 8938 16736 8944 16748
rect 8996 16736 9002 16788
rect 9214 16736 9220 16788
rect 9272 16776 9278 16788
rect 10321 16779 10379 16785
rect 10321 16776 10333 16779
rect 9272 16748 10333 16776
rect 9272 16736 9278 16748
rect 10321 16745 10333 16748
rect 10367 16776 10379 16779
rect 10367 16748 10824 16776
rect 10367 16745 10379 16748
rect 10321 16739 10379 16745
rect 6641 16711 6699 16717
rect 6641 16677 6653 16711
rect 6687 16708 6699 16711
rect 7466 16708 7472 16720
rect 6687 16680 7472 16708
rect 6687 16677 6699 16680
rect 6641 16671 6699 16677
rect 7466 16668 7472 16680
rect 7524 16708 7530 16720
rect 10796 16708 10824 16748
rect 10870 16736 10876 16788
rect 10928 16776 10934 16788
rect 11146 16776 11152 16788
rect 10928 16748 11152 16776
rect 10928 16736 10934 16748
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 11974 16736 11980 16788
rect 12032 16776 12038 16788
rect 12161 16779 12219 16785
rect 12161 16776 12173 16779
rect 12032 16748 12173 16776
rect 12032 16736 12038 16748
rect 12161 16745 12173 16748
rect 12207 16745 12219 16779
rect 12161 16739 12219 16745
rect 12176 16708 12204 16739
rect 12894 16736 12900 16788
rect 12952 16776 12958 16788
rect 13446 16776 13452 16788
rect 12952 16748 13452 16776
rect 12952 16736 12958 16748
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 13817 16779 13875 16785
rect 13817 16745 13829 16779
rect 13863 16776 13875 16779
rect 14093 16779 14151 16785
rect 13863 16748 14044 16776
rect 13863 16745 13875 16748
rect 13817 16739 13875 16745
rect 12682 16711 12740 16717
rect 12682 16708 12694 16711
rect 7524 16680 8248 16708
rect 7524 16668 7530 16680
rect 7282 16640 7288 16652
rect 7243 16612 7288 16640
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 7552 16643 7610 16649
rect 7552 16609 7564 16643
rect 7598 16640 7610 16643
rect 8110 16640 8116 16652
rect 7598 16612 8116 16640
rect 7598 16609 7610 16612
rect 7552 16603 7610 16609
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 8220 16640 8248 16680
rect 10796 16680 11192 16708
rect 12176 16680 12694 16708
rect 8220 16612 8340 16640
rect 8312 16504 8340 16612
rect 8846 16600 8852 16652
rect 8904 16640 8910 16652
rect 9306 16640 9312 16652
rect 8904 16612 9312 16640
rect 8904 16600 8910 16612
rect 9306 16600 9312 16612
rect 9364 16640 9370 16652
rect 10318 16640 10324 16652
rect 9364 16612 10324 16640
rect 9364 16600 9370 16612
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10502 16640 10508 16652
rect 10463 16612 10508 16640
rect 10502 16600 10508 16612
rect 10560 16600 10566 16652
rect 10796 16649 10824 16680
rect 11054 16649 11060 16652
rect 10781 16643 10839 16649
rect 10781 16609 10793 16643
rect 10827 16609 10839 16643
rect 11048 16640 11060 16649
rect 11015 16612 11060 16640
rect 10781 16603 10839 16609
rect 11048 16603 11060 16612
rect 11054 16600 11060 16603
rect 11112 16600 11118 16652
rect 11164 16640 11192 16680
rect 12682 16677 12694 16680
rect 12728 16677 12740 16711
rect 12682 16671 12740 16677
rect 14016 16640 14044 16748
rect 14093 16745 14105 16779
rect 14139 16745 14151 16779
rect 14093 16739 14151 16745
rect 14108 16708 14136 16739
rect 14366 16736 14372 16788
rect 14424 16776 14430 16788
rect 14461 16779 14519 16785
rect 14461 16776 14473 16779
rect 14424 16748 14473 16776
rect 14424 16736 14430 16748
rect 14461 16745 14473 16748
rect 14507 16745 14519 16779
rect 14461 16739 14519 16745
rect 14550 16736 14556 16788
rect 14608 16776 14614 16788
rect 15289 16779 15347 16785
rect 14608 16748 14653 16776
rect 14608 16736 14614 16748
rect 15289 16745 15301 16779
rect 15335 16776 15347 16779
rect 16022 16776 16028 16788
rect 15335 16748 16028 16776
rect 15335 16745 15347 16748
rect 15289 16739 15347 16745
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 17126 16776 17132 16788
rect 17087 16748 17132 16776
rect 17126 16736 17132 16748
rect 17184 16736 17190 16788
rect 18138 16776 18144 16788
rect 18099 16748 18144 16776
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 18509 16779 18567 16785
rect 18509 16745 18521 16779
rect 18555 16745 18567 16779
rect 18509 16739 18567 16745
rect 15378 16708 15384 16720
rect 14108 16680 15384 16708
rect 15378 16668 15384 16680
rect 15436 16668 15442 16720
rect 15657 16711 15715 16717
rect 15657 16677 15669 16711
rect 15703 16677 15715 16711
rect 18524 16708 18552 16739
rect 18690 16736 18696 16788
rect 18748 16776 18754 16788
rect 21082 16776 21088 16788
rect 18748 16748 20300 16776
rect 21043 16748 21088 16776
rect 18748 16736 18754 16748
rect 20272 16717 20300 16748
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 20257 16711 20315 16717
rect 18524 16680 20024 16708
rect 15657 16671 15715 16677
rect 14090 16640 14096 16652
rect 11164 16612 12480 16640
rect 14003 16612 14096 16640
rect 12452 16584 12480 16612
rect 14090 16600 14096 16612
rect 14148 16640 14154 16652
rect 15194 16640 15200 16652
rect 14148 16612 15200 16640
rect 14148 16600 14154 16612
rect 15194 16600 15200 16612
rect 15252 16600 15258 16652
rect 15672 16640 15700 16671
rect 15580 16612 15700 16640
rect 16117 16643 16175 16649
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 14734 16572 14740 16584
rect 12492 16544 12537 16572
rect 14695 16544 14740 16572
rect 12492 16532 12498 16544
rect 14734 16532 14740 16544
rect 14792 16532 14798 16584
rect 8312 16476 10824 16504
rect 6270 16436 6276 16448
rect 6231 16408 6276 16436
rect 6270 16396 6276 16408
rect 6328 16396 6334 16448
rect 8665 16439 8723 16445
rect 8665 16405 8677 16439
rect 8711 16436 8723 16439
rect 8754 16436 8760 16448
rect 8711 16408 8760 16436
rect 8711 16405 8723 16408
rect 8665 16399 8723 16405
rect 8754 16396 8760 16408
rect 8812 16396 8818 16448
rect 9306 16436 9312 16448
rect 9267 16408 9312 16436
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 9858 16396 9864 16448
rect 9916 16436 9922 16448
rect 9953 16439 10011 16445
rect 9953 16436 9965 16439
rect 9916 16408 9965 16436
rect 9916 16396 9922 16408
rect 9953 16405 9965 16408
rect 9999 16405 10011 16439
rect 10796 16436 10824 16476
rect 13538 16464 13544 16516
rect 13596 16504 13602 16516
rect 15470 16504 15476 16516
rect 13596 16476 15476 16504
rect 13596 16464 13602 16476
rect 15470 16464 15476 16476
rect 15528 16464 15534 16516
rect 15580 16504 15608 16612
rect 16117 16609 16129 16643
rect 16163 16640 16175 16643
rect 17037 16643 17095 16649
rect 17037 16640 17049 16643
rect 16163 16612 17049 16640
rect 16163 16609 16175 16612
rect 16117 16603 16175 16609
rect 17037 16609 17049 16612
rect 17083 16609 17095 16643
rect 17037 16603 17095 16609
rect 17957 16643 18015 16649
rect 17957 16609 17969 16643
rect 18003 16640 18015 16643
rect 18690 16640 18696 16652
rect 18003 16612 18696 16640
rect 18003 16609 18015 16612
rect 17957 16603 18015 16609
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 18874 16640 18880 16652
rect 18835 16612 18880 16640
rect 18874 16600 18880 16612
rect 18932 16600 18938 16652
rect 19996 16649 20024 16680
rect 20257 16677 20269 16711
rect 20303 16677 20315 16711
rect 20257 16671 20315 16677
rect 19981 16643 20039 16649
rect 19981 16609 19993 16643
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 20714 16600 20720 16652
rect 20772 16640 20778 16652
rect 20901 16643 20959 16649
rect 20901 16640 20913 16643
rect 20772 16612 20913 16640
rect 20772 16600 20778 16612
rect 20901 16609 20913 16612
rect 20947 16609 20959 16643
rect 20901 16603 20959 16609
rect 15746 16572 15752 16584
rect 15707 16544 15752 16572
rect 15746 16532 15752 16544
rect 15804 16532 15810 16584
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 17218 16572 17224 16584
rect 15896 16544 15941 16572
rect 17179 16544 17224 16572
rect 15896 16532 15902 16544
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 18966 16572 18972 16584
rect 18927 16544 18972 16572
rect 18966 16532 18972 16544
rect 19024 16532 19030 16584
rect 19058 16532 19064 16584
rect 19116 16572 19122 16584
rect 19518 16572 19524 16584
rect 19116 16544 19161 16572
rect 19479 16544 19524 16572
rect 19116 16532 19122 16544
rect 19518 16532 19524 16544
rect 19576 16532 19582 16584
rect 15654 16504 15660 16516
rect 15580 16476 15660 16504
rect 15654 16464 15660 16476
rect 15712 16464 15718 16516
rect 16022 16464 16028 16516
rect 16080 16504 16086 16516
rect 19610 16504 19616 16516
rect 16080 16476 19616 16504
rect 16080 16464 16086 16476
rect 19610 16464 19616 16476
rect 19668 16464 19674 16516
rect 16114 16436 16120 16448
rect 10796 16408 16120 16436
rect 9953 16399 10011 16405
rect 16114 16396 16120 16408
rect 16172 16396 16178 16448
rect 16298 16436 16304 16448
rect 16259 16408 16304 16436
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 16669 16439 16727 16445
rect 16669 16405 16681 16439
rect 16715 16436 16727 16439
rect 17034 16436 17040 16448
rect 16715 16408 17040 16436
rect 16715 16405 16727 16408
rect 16669 16399 16727 16405
rect 17034 16396 17040 16408
rect 17092 16396 17098 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 8110 16192 8116 16244
rect 8168 16232 8174 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 8168 16204 8217 16232
rect 8168 16192 8174 16204
rect 8205 16201 8217 16204
rect 8251 16201 8263 16235
rect 9214 16232 9220 16244
rect 8205 16195 8263 16201
rect 8496 16204 9220 16232
rect 8496 16105 8524 16204
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 9490 16192 9496 16244
rect 9548 16232 9554 16244
rect 9861 16235 9919 16241
rect 9861 16232 9873 16235
rect 9548 16204 9873 16232
rect 9548 16192 9554 16204
rect 9861 16201 9873 16204
rect 9907 16201 9919 16235
rect 9861 16195 9919 16201
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 12526 16232 12532 16244
rect 12483 16204 12532 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 12526 16192 12532 16204
rect 12584 16192 12590 16244
rect 12802 16192 12808 16244
rect 12860 16232 12866 16244
rect 13078 16232 13084 16244
rect 12860 16204 13084 16232
rect 12860 16192 12866 16204
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 15105 16235 15163 16241
rect 15105 16201 15117 16235
rect 15151 16232 15163 16235
rect 15930 16232 15936 16244
rect 15151 16204 15936 16232
rect 15151 16201 15163 16204
rect 15105 16195 15163 16201
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 18693 16235 18751 16241
rect 18693 16201 18705 16235
rect 18739 16232 18751 16235
rect 18874 16232 18880 16244
rect 18739 16204 18880 16232
rect 18739 16201 18751 16204
rect 18693 16195 18751 16201
rect 18874 16192 18880 16204
rect 18932 16192 18938 16244
rect 19889 16235 19947 16241
rect 19889 16201 19901 16235
rect 19935 16232 19947 16235
rect 20346 16232 20352 16244
rect 19935 16204 20352 16232
rect 19935 16201 19947 16204
rect 19889 16195 19947 16201
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 11514 16164 11520 16176
rect 11427 16136 11520 16164
rect 11514 16124 11520 16136
rect 11572 16164 11578 16176
rect 11572 16136 13124 16164
rect 11572 16124 11578 16136
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 12069 16099 12127 16105
rect 12069 16065 12081 16099
rect 12115 16096 12127 16099
rect 12342 16096 12348 16108
rect 12115 16068 12348 16096
rect 12115 16065 12127 16068
rect 12069 16059 12127 16065
rect 12342 16056 12348 16068
rect 12400 16056 12406 16108
rect 13096 16105 13124 16136
rect 15378 16124 15384 16176
rect 15436 16164 15442 16176
rect 16117 16167 16175 16173
rect 15436 16136 15976 16164
rect 15436 16124 15442 16136
rect 13081 16099 13139 16105
rect 13081 16065 13093 16099
rect 13127 16065 13139 16099
rect 13081 16059 13139 16065
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7374 16028 7380 16040
rect 6871 16000 7380 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 8754 16037 8760 16040
rect 8748 16028 8760 16037
rect 8715 16000 8760 16028
rect 8748 15991 8760 16000
rect 8754 15988 8760 15991
rect 8812 15988 8818 16040
rect 9030 15988 9036 16040
rect 9088 16028 9094 16040
rect 9214 16028 9220 16040
rect 9088 16000 9220 16028
rect 9088 15988 9094 16000
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 9766 15988 9772 16040
rect 9824 16028 9830 16040
rect 10137 16031 10195 16037
rect 10137 16028 10149 16031
rect 9824 16000 10149 16028
rect 9824 15988 9830 16000
rect 10137 15997 10149 16000
rect 10183 15997 10195 16031
rect 10137 15991 10195 15997
rect 10336 16000 13032 16028
rect 7092 15963 7150 15969
rect 7092 15929 7104 15963
rect 7138 15960 7150 15963
rect 10336 15960 10364 16000
rect 7138 15932 10364 15960
rect 10404 15963 10462 15969
rect 7138 15929 7150 15932
rect 7092 15923 7150 15929
rect 10404 15929 10416 15963
rect 10450 15960 10462 15963
rect 10778 15960 10784 15972
rect 10450 15932 10784 15960
rect 10450 15929 10462 15932
rect 10404 15923 10462 15929
rect 10778 15920 10784 15932
rect 10836 15920 10842 15972
rect 10870 15920 10876 15972
rect 10928 15960 10934 15972
rect 12897 15963 12955 15969
rect 12897 15960 12909 15963
rect 10928 15932 12909 15960
rect 10928 15920 10934 15932
rect 12897 15929 12909 15932
rect 12943 15929 12955 15963
rect 12897 15923 12955 15929
rect 6454 15892 6460 15904
rect 6367 15864 6460 15892
rect 6454 15852 6460 15864
rect 6512 15892 6518 15904
rect 8938 15892 8944 15904
rect 6512 15864 8944 15892
rect 6512 15852 6518 15864
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 12066 15852 12072 15904
rect 12124 15892 12130 15904
rect 12805 15895 12863 15901
rect 12805 15892 12817 15895
rect 12124 15864 12817 15892
rect 12124 15852 12130 15864
rect 12805 15861 12817 15864
rect 12851 15861 12863 15895
rect 13004 15892 13032 16000
rect 13096 15960 13124 16059
rect 13446 16056 13452 16108
rect 13504 16096 13510 16108
rect 15749 16099 15807 16105
rect 13504 16068 13549 16096
rect 13504 16056 13510 16068
rect 15749 16065 15761 16099
rect 15795 16096 15807 16099
rect 15838 16096 15844 16108
rect 15795 16068 15844 16096
rect 15795 16065 15807 16068
rect 15749 16059 15807 16065
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 15948 16096 15976 16136
rect 16117 16133 16129 16167
rect 16163 16164 16175 16167
rect 16163 16136 17172 16164
rect 16163 16133 16175 16136
rect 16117 16127 16175 16133
rect 16577 16099 16635 16105
rect 16577 16096 16589 16099
rect 15948 16068 16589 16096
rect 16577 16065 16589 16068
rect 16623 16065 16635 16099
rect 16577 16059 16635 16065
rect 16669 16099 16727 16105
rect 16669 16065 16681 16099
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 13716 16031 13774 16037
rect 13716 15997 13728 16031
rect 13762 16028 13774 16031
rect 14734 16028 14740 16040
rect 13762 16000 14740 16028
rect 13762 15997 13774 16000
rect 13716 15991 13774 15997
rect 14734 15988 14740 16000
rect 14792 15988 14798 16040
rect 15562 15988 15568 16040
rect 15620 16028 15626 16040
rect 16485 16031 16543 16037
rect 16485 16028 16497 16031
rect 15620 16000 16497 16028
rect 15620 15988 15626 16000
rect 16485 15997 16497 16000
rect 16531 15997 16543 16031
rect 16485 15991 16543 15997
rect 13814 15960 13820 15972
rect 13096 15932 13820 15960
rect 13814 15920 13820 15932
rect 13872 15920 13878 15972
rect 16675 15960 16703 16059
rect 17144 16037 17172 16136
rect 19426 16124 19432 16176
rect 19484 16164 19490 16176
rect 19484 16136 20484 16164
rect 19484 16124 19490 16136
rect 19150 16096 19156 16108
rect 19111 16068 19156 16096
rect 19150 16056 19156 16068
rect 19208 16056 19214 16108
rect 19337 16099 19395 16105
rect 19337 16065 19349 16099
rect 19383 16096 19395 16099
rect 19702 16096 19708 16108
rect 19383 16068 19708 16096
rect 19383 16065 19395 16068
rect 19337 16059 19395 16065
rect 19702 16056 19708 16068
rect 19760 16056 19766 16108
rect 20456 16105 20484 16136
rect 20441 16099 20499 16105
rect 20441 16065 20453 16099
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 17129 16031 17187 16037
rect 17129 15997 17141 16031
rect 17175 15997 17187 16031
rect 17129 15991 17187 15997
rect 17954 15988 17960 16040
rect 18012 16028 18018 16040
rect 18141 16031 18199 16037
rect 18141 16028 18153 16031
rect 18012 16000 18153 16028
rect 18012 15988 18018 16000
rect 18141 15997 18153 16000
rect 18187 15997 18199 16031
rect 18141 15991 18199 15997
rect 19061 16031 19119 16037
rect 19061 15997 19073 16031
rect 19107 16028 19119 16031
rect 19518 16028 19524 16040
rect 19107 16000 19524 16028
rect 19107 15997 19119 16000
rect 19061 15991 19119 15997
rect 19518 15988 19524 16000
rect 19576 15988 19582 16040
rect 20901 16031 20959 16037
rect 20901 15997 20913 16031
rect 20947 15997 20959 16031
rect 20901 15991 20959 15997
rect 14844 15932 16703 15960
rect 17405 15963 17463 15969
rect 14844 15901 14872 15932
rect 17405 15929 17417 15963
rect 17451 15960 17463 15963
rect 20916 15960 20944 15991
rect 17451 15932 20944 15960
rect 17451 15929 17463 15932
rect 17405 15923 17463 15929
rect 14829 15895 14887 15901
rect 14829 15892 14841 15895
rect 13004 15864 14841 15892
rect 12805 15855 12863 15861
rect 14829 15861 14841 15864
rect 14875 15861 14887 15895
rect 14829 15855 14887 15861
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 15473 15895 15531 15901
rect 15473 15892 15485 15895
rect 15436 15864 15485 15892
rect 15436 15852 15442 15864
rect 15473 15861 15485 15864
rect 15519 15861 15531 15895
rect 15473 15855 15531 15861
rect 15562 15852 15568 15904
rect 15620 15892 15626 15904
rect 16390 15892 16396 15904
rect 15620 15864 16396 15892
rect 15620 15852 15626 15864
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 18322 15892 18328 15904
rect 18283 15864 18328 15892
rect 18322 15852 18328 15864
rect 18380 15852 18386 15904
rect 20070 15852 20076 15904
rect 20128 15892 20134 15904
rect 20257 15895 20315 15901
rect 20257 15892 20269 15895
rect 20128 15864 20269 15892
rect 20128 15852 20134 15864
rect 20257 15861 20269 15864
rect 20303 15861 20315 15895
rect 20257 15855 20315 15861
rect 20346 15852 20352 15904
rect 20404 15892 20410 15904
rect 20404 15864 20449 15892
rect 20404 15852 20410 15864
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 21085 15895 21143 15901
rect 21085 15892 21097 15895
rect 20680 15864 21097 15892
rect 20680 15852 20686 15864
rect 21085 15861 21097 15864
rect 21131 15861 21143 15895
rect 21085 15855 21143 15861
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 6178 15688 6184 15700
rect 6139 15660 6184 15688
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 6546 15688 6552 15700
rect 6507 15660 6552 15688
rect 6546 15648 6552 15660
rect 6604 15648 6610 15700
rect 6822 15648 6828 15700
rect 6880 15688 6886 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6880 15660 6929 15688
rect 6880 15648 6886 15660
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 6917 15651 6975 15657
rect 7285 15691 7343 15697
rect 7285 15657 7297 15691
rect 7331 15688 7343 15691
rect 8849 15691 8907 15697
rect 8849 15688 8861 15691
rect 7331 15660 8861 15688
rect 7331 15657 7343 15660
rect 7285 15651 7343 15657
rect 8849 15657 8861 15660
rect 8895 15657 8907 15691
rect 8849 15651 8907 15657
rect 10229 15691 10287 15697
rect 10229 15657 10241 15691
rect 10275 15688 10287 15691
rect 10870 15688 10876 15700
rect 10275 15660 10876 15688
rect 10275 15657 10287 15660
rect 10229 15651 10287 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 11241 15691 11299 15697
rect 11241 15657 11253 15691
rect 11287 15688 11299 15691
rect 12066 15688 12072 15700
rect 11287 15660 12072 15688
rect 11287 15657 11299 15660
rect 11241 15651 11299 15657
rect 12066 15648 12072 15660
rect 12124 15648 12130 15700
rect 12253 15691 12311 15697
rect 12253 15657 12265 15691
rect 12299 15657 12311 15691
rect 12253 15651 12311 15657
rect 6196 15620 6224 15648
rect 7745 15623 7803 15629
rect 7745 15620 7757 15623
rect 6196 15592 7757 15620
rect 7745 15589 7757 15592
rect 7791 15589 7803 15623
rect 10594 15620 10600 15632
rect 7745 15583 7803 15589
rect 7852 15592 10600 15620
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 7653 15555 7711 15561
rect 7653 15552 7665 15555
rect 6972 15524 7665 15552
rect 6972 15512 6978 15524
rect 7653 15521 7665 15524
rect 7699 15521 7711 15555
rect 7653 15515 7711 15521
rect 6546 15444 6552 15496
rect 6604 15484 6610 15496
rect 7852 15484 7880 15592
rect 10594 15580 10600 15592
rect 10652 15580 10658 15632
rect 12268 15620 12296 15651
rect 12802 15648 12808 15700
rect 12860 15688 12866 15700
rect 15378 15688 15384 15700
rect 12860 15660 15240 15688
rect 15339 15660 15384 15688
rect 12860 15648 12866 15660
rect 13633 15623 13691 15629
rect 13633 15620 13645 15623
rect 12268 15592 13645 15620
rect 13633 15589 13645 15592
rect 13679 15589 13691 15623
rect 15212 15620 15240 15660
rect 15378 15648 15384 15660
rect 15436 15648 15442 15700
rect 16114 15648 16120 15700
rect 16172 15688 16178 15700
rect 16393 15691 16451 15697
rect 16393 15688 16405 15691
rect 16172 15660 16405 15688
rect 16172 15648 16178 15660
rect 16393 15657 16405 15660
rect 16439 15657 16451 15691
rect 16942 15688 16948 15700
rect 16903 15660 16948 15688
rect 16393 15651 16451 15657
rect 16942 15648 16948 15660
rect 17000 15648 17006 15700
rect 18966 15648 18972 15700
rect 19024 15688 19030 15700
rect 19153 15691 19211 15697
rect 19153 15688 19165 15691
rect 19024 15660 19165 15688
rect 19024 15648 19030 15660
rect 19153 15657 19165 15660
rect 19199 15657 19211 15691
rect 19610 15688 19616 15700
rect 19571 15660 19616 15688
rect 19153 15651 19211 15657
rect 19610 15648 19616 15660
rect 19668 15648 19674 15700
rect 16301 15623 16359 15629
rect 16301 15620 16313 15623
rect 15212 15592 16313 15620
rect 13633 15583 13691 15589
rect 16301 15589 16313 15592
rect 16347 15620 16359 15623
rect 17034 15620 17040 15632
rect 16347 15592 17040 15620
rect 16347 15589 16359 15592
rect 16301 15583 16359 15589
rect 17034 15580 17040 15592
rect 17092 15580 17098 15632
rect 17764 15623 17822 15629
rect 17764 15589 17776 15623
rect 17810 15620 17822 15623
rect 19702 15620 19708 15632
rect 17810 15592 19708 15620
rect 17810 15589 17822 15592
rect 17764 15583 17822 15589
rect 19702 15580 19708 15592
rect 19760 15580 19766 15632
rect 20162 15580 20168 15632
rect 20220 15620 20226 15632
rect 20220 15592 20944 15620
rect 20220 15580 20226 15592
rect 8757 15555 8815 15561
rect 8757 15521 8769 15555
rect 8803 15552 8815 15555
rect 9030 15552 9036 15564
rect 8803 15524 9036 15552
rect 8803 15521 8815 15524
rect 8757 15515 8815 15521
rect 9030 15512 9036 15524
rect 9088 15512 9094 15564
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 11609 15555 11667 15561
rect 11609 15552 11621 15555
rect 11296 15524 11621 15552
rect 11296 15512 11302 15524
rect 11609 15521 11621 15524
rect 11655 15521 11667 15555
rect 11609 15515 11667 15521
rect 12621 15555 12679 15561
rect 12621 15521 12633 15555
rect 12667 15552 12679 15555
rect 14277 15555 14335 15561
rect 14277 15552 14289 15555
rect 12667 15524 14289 15552
rect 12667 15521 12679 15524
rect 12621 15515 12679 15521
rect 14277 15521 14289 15524
rect 14323 15521 14335 15555
rect 17052 15552 17080 15580
rect 20916 15561 20944 15592
rect 19521 15555 19579 15561
rect 19521 15552 19533 15555
rect 17052 15524 19533 15552
rect 14277 15515 14335 15521
rect 19521 15521 19533 15524
rect 19567 15521 19579 15555
rect 19521 15515 19579 15521
rect 20257 15555 20315 15561
rect 20257 15521 20269 15555
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 20901 15555 20959 15561
rect 20901 15521 20913 15555
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 6604 15456 7880 15484
rect 7929 15487 7987 15493
rect 6604 15444 6610 15456
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8202 15484 8208 15496
rect 7975 15456 8208 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 8846 15444 8852 15496
rect 8904 15484 8910 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8904 15456 8953 15484
rect 8904 15444 8910 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 9674 15484 9680 15496
rect 9635 15456 9680 15484
rect 8941 15447 8999 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 10689 15487 10747 15493
rect 10689 15453 10701 15487
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 6822 15376 6828 15428
rect 6880 15416 6886 15428
rect 10704 15416 10732 15447
rect 10778 15444 10784 15496
rect 10836 15484 10842 15496
rect 11698 15484 11704 15496
rect 10836 15456 10881 15484
rect 11659 15456 11704 15484
rect 10836 15444 10842 15456
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 11793 15487 11851 15493
rect 11793 15453 11805 15487
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 6880 15388 10732 15416
rect 10796 15416 10824 15444
rect 11808 15416 11836 15447
rect 12342 15444 12348 15496
rect 12400 15484 12406 15496
rect 12713 15487 12771 15493
rect 12713 15484 12725 15487
rect 12400 15456 12725 15484
rect 12400 15444 12406 15456
rect 12713 15453 12725 15456
rect 12759 15453 12771 15487
rect 12713 15447 12771 15453
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 12912 15416 12940 15447
rect 10796 15388 12940 15416
rect 6880 15376 6886 15388
rect 5905 15351 5963 15357
rect 5905 15317 5917 15351
rect 5951 15348 5963 15351
rect 7558 15348 7564 15360
rect 5951 15320 7564 15348
rect 5951 15317 5963 15320
rect 5905 15311 5963 15317
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 8389 15351 8447 15357
rect 8389 15317 8401 15351
rect 8435 15348 8447 15351
rect 8754 15348 8760 15360
rect 8435 15320 8760 15348
rect 8435 15317 8447 15320
rect 8389 15311 8447 15317
rect 8754 15308 8760 15320
rect 8812 15308 8818 15360
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 12802 15348 12808 15360
rect 8996 15320 12808 15348
rect 8996 15308 9002 15320
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 12912 15348 12940 15388
rect 13078 15376 13084 15428
rect 13136 15416 13142 15428
rect 13265 15419 13323 15425
rect 13265 15416 13277 15419
rect 13136 15388 13277 15416
rect 13136 15376 13142 15388
rect 13265 15385 13277 15388
rect 13311 15385 13323 15419
rect 13740 15416 13768 15447
rect 13814 15444 13820 15496
rect 13872 15484 13878 15496
rect 13872 15456 13917 15484
rect 13872 15444 13878 15456
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 14737 15487 14795 15493
rect 14737 15484 14749 15487
rect 14608 15456 14749 15484
rect 14608 15444 14614 15456
rect 14737 15453 14749 15456
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 16482 15444 16488 15496
rect 16540 15484 16546 15496
rect 17494 15484 17500 15496
rect 16540 15456 16585 15484
rect 17455 15456 17500 15484
rect 16540 15444 16546 15456
rect 17494 15444 17500 15456
rect 17552 15444 17558 15496
rect 19702 15484 19708 15496
rect 19663 15456 19708 15484
rect 19702 15444 19708 15456
rect 19760 15444 19766 15496
rect 15933 15419 15991 15425
rect 15933 15416 15945 15419
rect 13740 15388 15945 15416
rect 13265 15379 13323 15385
rect 15933 15385 15945 15388
rect 15979 15385 15991 15419
rect 15933 15379 15991 15385
rect 18877 15419 18935 15425
rect 18877 15385 18889 15419
rect 18923 15416 18935 15419
rect 19058 15416 19064 15428
rect 18923 15388 19064 15416
rect 18923 15385 18935 15388
rect 18877 15379 18935 15385
rect 19058 15376 19064 15388
rect 19116 15376 19122 15428
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 19610 15416 19616 15428
rect 19392 15388 19616 15416
rect 19392 15376 19398 15388
rect 19610 15376 19616 15388
rect 19668 15376 19674 15428
rect 16482 15348 16488 15360
rect 12912 15320 16488 15348
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 16574 15308 16580 15360
rect 16632 15348 16638 15360
rect 20272 15348 20300 15515
rect 20438 15348 20444 15360
rect 16632 15320 20300 15348
rect 20399 15320 20444 15348
rect 16632 15308 16638 15320
rect 20438 15308 20444 15320
rect 20496 15308 20502 15360
rect 20530 15308 20536 15360
rect 20588 15348 20594 15360
rect 21085 15351 21143 15357
rect 21085 15348 21097 15351
rect 20588 15320 21097 15348
rect 20588 15308 20594 15320
rect 21085 15317 21097 15320
rect 21131 15317 21143 15351
rect 21085 15311 21143 15317
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 6454 15144 6460 15156
rect 6415 15116 6460 15144
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 6914 15144 6920 15156
rect 6875 15116 6920 15144
rect 6914 15104 6920 15116
rect 6972 15144 6978 15156
rect 7282 15144 7288 15156
rect 6972 15116 7288 15144
rect 6972 15104 6978 15116
rect 7282 15104 7288 15116
rect 7340 15104 7346 15156
rect 7837 15147 7895 15153
rect 7837 15113 7849 15147
rect 7883 15144 7895 15147
rect 8938 15144 8944 15156
rect 7883 15116 8944 15144
rect 7883 15113 7895 15116
rect 7837 15107 7895 15113
rect 8938 15104 8944 15116
rect 8996 15104 9002 15156
rect 9030 15104 9036 15156
rect 9088 15144 9094 15156
rect 11698 15144 11704 15156
rect 9088 15116 11704 15144
rect 9088 15104 9094 15116
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 19981 15147 20039 15153
rect 19981 15144 19993 15147
rect 12492 15116 19993 15144
rect 12492 15104 12498 15116
rect 19981 15113 19993 15116
rect 20027 15113 20039 15147
rect 19981 15107 20039 15113
rect 20165 15147 20223 15153
rect 20165 15113 20177 15147
rect 20211 15144 20223 15147
rect 20346 15144 20352 15156
rect 20211 15116 20352 15144
rect 20211 15113 20223 15116
rect 20165 15107 20223 15113
rect 20346 15104 20352 15116
rect 20404 15104 20410 15156
rect 7650 15036 7656 15088
rect 7708 15076 7714 15088
rect 7708 15048 9720 15076
rect 7708 15036 7714 15048
rect 7469 15011 7527 15017
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 8386 15008 8392 15020
rect 7515 14980 8392 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 8846 14968 8852 15020
rect 8904 15008 8910 15020
rect 9033 15011 9091 15017
rect 9033 15008 9045 15011
rect 8904 14980 9045 15008
rect 8904 14968 8910 14980
rect 9033 14977 9045 14980
rect 9079 14977 9091 15011
rect 9033 14971 9091 14977
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 9493 14943 9551 14949
rect 9493 14940 9505 14943
rect 8352 14912 9505 14940
rect 8352 14900 8358 14912
rect 9493 14909 9505 14912
rect 9539 14909 9551 14943
rect 9692 14940 9720 15048
rect 9950 15036 9956 15088
rect 10008 15076 10014 15088
rect 10502 15076 10508 15088
rect 10008 15048 10508 15076
rect 10008 15036 10014 15048
rect 10502 15036 10508 15048
rect 10560 15076 10566 15088
rect 11425 15079 11483 15085
rect 11425 15076 11437 15079
rect 10560 15048 11437 15076
rect 10560 15036 10566 15048
rect 11425 15045 11437 15048
rect 11471 15045 11483 15079
rect 11425 15039 11483 15045
rect 11606 15036 11612 15088
rect 11664 15076 11670 15088
rect 11882 15076 11888 15088
rect 11664 15048 11888 15076
rect 11664 15036 11670 15048
rect 11882 15036 11888 15048
rect 11940 15036 11946 15088
rect 13357 15079 13415 15085
rect 13357 15045 13369 15079
rect 13403 15076 13415 15079
rect 14458 15076 14464 15088
rect 13403 15048 14464 15076
rect 13403 15045 13415 15048
rect 13357 15039 13415 15045
rect 14458 15036 14464 15048
rect 14516 15036 14522 15088
rect 16025 15079 16083 15085
rect 16025 15045 16037 15079
rect 16071 15076 16083 15079
rect 16482 15076 16488 15088
rect 16071 15048 16488 15076
rect 16071 15045 16083 15048
rect 16025 15039 16083 15045
rect 16482 15036 16488 15048
rect 16540 15036 16546 15088
rect 16666 15036 16672 15088
rect 16724 15076 16730 15088
rect 17313 15079 17371 15085
rect 17313 15076 17325 15079
rect 16724 15048 17325 15076
rect 16724 15036 16730 15048
rect 17313 15045 17325 15048
rect 17359 15045 17371 15079
rect 17313 15039 17371 15045
rect 9769 15011 9827 15017
rect 9769 14977 9781 15011
rect 9815 15008 9827 15011
rect 13906 15008 13912 15020
rect 9815 14980 13768 15008
rect 13867 14980 13912 15008
rect 9815 14977 9827 14980
rect 9769 14971 9827 14977
rect 9692 14912 9812 14940
rect 9493 14903 9551 14909
rect 8205 14875 8263 14881
rect 8205 14841 8217 14875
rect 8251 14872 8263 14875
rect 8849 14875 8907 14881
rect 8251 14844 8800 14872
rect 8251 14841 8263 14844
rect 8205 14835 8263 14841
rect 8481 14807 8539 14813
rect 8481 14773 8493 14807
rect 8527 14804 8539 14807
rect 8662 14804 8668 14816
rect 8527 14776 8668 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 8662 14764 8668 14776
rect 8720 14764 8726 14816
rect 8772 14804 8800 14844
rect 8849 14841 8861 14875
rect 8895 14872 8907 14875
rect 9674 14872 9680 14884
rect 8895 14844 9680 14872
rect 8895 14841 8907 14844
rect 8849 14835 8907 14841
rect 9674 14832 9680 14844
rect 9732 14832 9738 14884
rect 9784 14872 9812 14912
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10321 14943 10379 14949
rect 10321 14940 10333 14943
rect 10192 14912 10333 14940
rect 10192 14900 10198 14912
rect 10321 14909 10333 14912
rect 10367 14909 10379 14943
rect 10686 14940 10692 14952
rect 10647 14912 10692 14940
rect 10321 14903 10379 14909
rect 10686 14900 10692 14912
rect 10744 14940 10750 14952
rect 10870 14940 10876 14952
rect 10744 14912 10876 14940
rect 10744 14900 10750 14912
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 11609 14943 11667 14949
rect 11609 14909 11621 14943
rect 11655 14940 11667 14943
rect 12069 14943 12127 14949
rect 11655 14912 11928 14940
rect 11655 14909 11667 14912
rect 11609 14903 11667 14909
rect 10778 14872 10784 14884
rect 9784 14844 10784 14872
rect 10778 14832 10784 14844
rect 10836 14832 10842 14884
rect 8938 14804 8944 14816
rect 8772 14776 8944 14804
rect 8938 14764 8944 14776
rect 8996 14804 9002 14816
rect 10318 14804 10324 14816
rect 8996 14776 10324 14804
rect 8996 14764 9002 14776
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 11149 14807 11207 14813
rect 11149 14773 11161 14807
rect 11195 14804 11207 14807
rect 11238 14804 11244 14816
rect 11195 14776 11244 14804
rect 11195 14773 11207 14776
rect 11149 14767 11207 14773
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 11900 14813 11928 14912
rect 12069 14909 12081 14943
rect 12115 14909 12127 14943
rect 12069 14903 12127 14909
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14940 12495 14943
rect 12618 14940 12624 14952
rect 12483 14912 12624 14940
rect 12483 14909 12495 14912
rect 12437 14903 12495 14909
rect 12084 14872 12112 14903
rect 12618 14900 12624 14912
rect 12676 14900 12682 14952
rect 13740 14940 13768 14980
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 14424 14980 14657 15008
rect 14424 14968 14430 14980
rect 14645 14977 14657 14980
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 15654 14968 15660 15020
rect 15712 15008 15718 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 15712 14980 16865 15008
rect 15712 14968 15718 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 17328 15008 17356 15039
rect 20717 15011 20775 15017
rect 17328 14980 18276 15008
rect 16853 14971 16911 14977
rect 14274 14940 14280 14952
rect 13740 14912 14280 14940
rect 14274 14900 14280 14912
rect 14332 14900 14338 14952
rect 18248 14949 18276 14980
rect 20717 14977 20729 15011
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 17497 14943 17555 14949
rect 17497 14940 17509 14943
rect 14660 14912 17509 14940
rect 12526 14872 12532 14884
rect 12084 14844 12532 14872
rect 12526 14832 12532 14844
rect 12584 14832 12590 14884
rect 12710 14872 12716 14884
rect 12671 14844 12716 14872
rect 12710 14832 12716 14844
rect 12768 14832 12774 14884
rect 14660 14872 14688 14912
rect 17497 14909 17509 14912
rect 17543 14909 17555 14943
rect 17497 14903 17555 14909
rect 18233 14943 18291 14949
rect 18233 14909 18245 14943
rect 18279 14909 18291 14943
rect 18233 14903 18291 14909
rect 18509 14943 18567 14949
rect 18509 14909 18521 14943
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 18776 14943 18834 14949
rect 18776 14909 18788 14943
rect 18822 14940 18834 14943
rect 19058 14940 19064 14952
rect 18822 14912 19064 14940
rect 18822 14909 18834 14912
rect 18776 14903 18834 14909
rect 13556 14844 14688 14872
rect 11885 14807 11943 14813
rect 11885 14773 11897 14807
rect 11931 14804 11943 14807
rect 13556 14804 13584 14844
rect 14734 14832 14740 14884
rect 14792 14872 14798 14884
rect 14890 14875 14948 14881
rect 14890 14872 14902 14875
rect 14792 14844 14902 14872
rect 14792 14832 14798 14844
rect 14890 14841 14902 14844
rect 14936 14841 14948 14875
rect 14890 14835 14948 14841
rect 15378 14832 15384 14884
rect 15436 14872 15442 14884
rect 16669 14875 16727 14881
rect 16669 14872 16681 14875
rect 15436 14844 16681 14872
rect 15436 14832 15442 14844
rect 16669 14841 16681 14844
rect 16715 14841 16727 14875
rect 18524 14872 18552 14903
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 19981 14943 20039 14949
rect 19981 14909 19993 14943
rect 20027 14940 20039 14943
rect 20625 14943 20683 14949
rect 20625 14940 20637 14943
rect 20027 14912 20637 14940
rect 20027 14909 20039 14912
rect 19981 14903 20039 14909
rect 20625 14909 20637 14912
rect 20671 14909 20683 14943
rect 20625 14903 20683 14909
rect 16669 14835 16727 14841
rect 18064 14844 18552 14872
rect 18064 14816 18092 14844
rect 13722 14804 13728 14816
rect 11931 14776 13584 14804
rect 13683 14776 13728 14804
rect 11931 14773 11943 14776
rect 11885 14767 11943 14773
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 13872 14776 13917 14804
rect 13872 14764 13878 14776
rect 14090 14764 14096 14816
rect 14148 14804 14154 14816
rect 16301 14807 16359 14813
rect 16301 14804 16313 14807
rect 14148 14776 16313 14804
rect 14148 14764 14154 14776
rect 16301 14773 16313 14776
rect 16347 14773 16359 14807
rect 16758 14804 16764 14816
rect 16719 14776 16764 14804
rect 16301 14767 16359 14773
rect 16758 14764 16764 14776
rect 16816 14764 16822 14816
rect 18046 14804 18052 14816
rect 18007 14776 18052 14804
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18524 14804 18552 14844
rect 18598 14832 18604 14884
rect 18656 14872 18662 14884
rect 19242 14872 19248 14884
rect 18656 14844 19248 14872
rect 18656 14832 18662 14844
rect 19242 14832 19248 14844
rect 19300 14872 19306 14884
rect 20533 14875 20591 14881
rect 20533 14872 20545 14875
rect 19300 14844 20545 14872
rect 19300 14832 19306 14844
rect 20533 14841 20545 14844
rect 20579 14841 20591 14875
rect 20732 14872 20760 14971
rect 20533 14835 20591 14841
rect 20640 14844 20760 14872
rect 18874 14804 18880 14816
rect 18524 14776 18880 14804
rect 18874 14764 18880 14776
rect 18932 14764 18938 14816
rect 19886 14804 19892 14816
rect 19847 14776 19892 14804
rect 19886 14764 19892 14776
rect 19944 14804 19950 14816
rect 20640 14804 20668 14844
rect 21174 14804 21180 14816
rect 19944 14776 20668 14804
rect 21135 14776 21180 14804
rect 19944 14764 19950 14776
rect 21174 14764 21180 14776
rect 21232 14764 21238 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 6638 14560 6644 14612
rect 6696 14600 6702 14612
rect 6825 14603 6883 14609
rect 6825 14600 6837 14603
rect 6696 14572 6837 14600
rect 6696 14560 6702 14572
rect 6825 14569 6837 14572
rect 6871 14569 6883 14603
rect 6825 14563 6883 14569
rect 7285 14603 7343 14609
rect 7285 14569 7297 14603
rect 7331 14600 7343 14603
rect 7466 14600 7472 14612
rect 7331 14572 7472 14600
rect 7331 14569 7343 14572
rect 7285 14563 7343 14569
rect 7466 14560 7472 14572
rect 7524 14560 7530 14612
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 7708 14572 7941 14600
rect 7708 14560 7714 14572
rect 7929 14569 7941 14572
rect 7975 14569 7987 14603
rect 8294 14600 8300 14612
rect 8255 14572 8300 14600
rect 7929 14563 7987 14569
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 8662 14600 8668 14612
rect 8623 14572 8668 14600
rect 8662 14560 8668 14572
rect 8720 14560 8726 14612
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 8812 14572 8857 14600
rect 8812 14560 8818 14572
rect 8938 14560 8944 14612
rect 8996 14600 9002 14612
rect 11146 14600 11152 14612
rect 8996 14572 11152 14600
rect 8996 14560 9002 14572
rect 11146 14560 11152 14572
rect 11204 14600 11210 14612
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 11204 14572 11805 14600
rect 11204 14560 11210 14572
rect 11793 14569 11805 14572
rect 11839 14600 11851 14603
rect 11882 14600 11888 14612
rect 11839 14572 11888 14600
rect 11839 14569 11851 14572
rect 11793 14563 11851 14569
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 12529 14603 12587 14609
rect 12529 14569 12541 14603
rect 12575 14600 12587 14603
rect 13814 14600 13820 14612
rect 12575 14572 13820 14600
rect 12575 14569 12587 14572
rect 12529 14563 12587 14569
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 16574 14600 16580 14612
rect 13924 14572 16580 14600
rect 9944 14535 10002 14541
rect 9944 14501 9956 14535
rect 9990 14532 10002 14535
rect 12618 14532 12624 14544
rect 9990 14504 12624 14532
rect 9990 14501 10002 14504
rect 9944 14495 10002 14501
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 12710 14492 12716 14544
rect 12768 14532 12774 14544
rect 13924 14532 13952 14572
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 16666 14560 16672 14612
rect 16724 14600 16730 14612
rect 19426 14600 19432 14612
rect 16724 14572 19432 14600
rect 16724 14560 16730 14572
rect 19426 14560 19432 14572
rect 19484 14600 19490 14612
rect 19705 14603 19763 14609
rect 19705 14600 19717 14603
rect 19484 14572 19717 14600
rect 19484 14560 19490 14572
rect 19705 14569 19717 14572
rect 19751 14569 19763 14603
rect 19705 14563 19763 14569
rect 19797 14603 19855 14609
rect 19797 14569 19809 14603
rect 19843 14600 19855 14603
rect 20070 14600 20076 14612
rect 19843 14572 20076 14600
rect 19843 14569 19855 14572
rect 19797 14563 19855 14569
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 20165 14603 20223 14609
rect 20165 14569 20177 14603
rect 20211 14600 20223 14603
rect 21174 14600 21180 14612
rect 20211 14572 21180 14600
rect 20211 14569 20223 14572
rect 20165 14563 20223 14569
rect 21174 14560 21180 14572
rect 21232 14560 21238 14612
rect 12768 14504 13952 14532
rect 12768 14492 12774 14504
rect 14826 14492 14832 14544
rect 14884 14532 14890 14544
rect 14884 14504 15884 14532
rect 14884 14492 14890 14504
rect 7282 14424 7288 14476
rect 7340 14464 7346 14476
rect 8294 14464 8300 14476
rect 7340 14436 8300 14464
rect 7340 14424 7346 14436
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14464 9735 14467
rect 9766 14464 9772 14476
rect 9723 14436 9772 14464
rect 9723 14433 9735 14436
rect 9677 14427 9735 14433
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 11698 14464 11704 14476
rect 11611 14436 11704 14464
rect 11698 14424 11704 14436
rect 11756 14464 11762 14476
rect 12158 14464 12164 14476
rect 11756 14436 12164 14464
rect 11756 14424 11762 14436
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 12894 14464 12900 14476
rect 12855 14436 12900 14464
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 13814 14473 13820 14476
rect 13808 14464 13820 14473
rect 13775 14436 13820 14464
rect 13808 14427 13820 14436
rect 13814 14424 13820 14427
rect 13872 14424 13878 14476
rect 14274 14424 14280 14476
rect 14332 14464 14338 14476
rect 15654 14464 15660 14476
rect 14332 14436 14596 14464
rect 15615 14436 15660 14464
rect 14332 14424 14338 14436
rect 8941 14399 8999 14405
rect 8941 14365 8953 14399
rect 8987 14396 8999 14399
rect 9490 14396 9496 14408
rect 8987 14368 9496 14396
rect 8987 14365 8999 14368
rect 8941 14359 8999 14365
rect 9490 14356 9496 14368
rect 9548 14356 9554 14408
rect 11885 14399 11943 14405
rect 11885 14396 11897 14399
rect 11072 14368 11897 14396
rect 11072 14340 11100 14368
rect 11885 14365 11897 14368
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12989 14399 13047 14405
rect 12989 14396 13001 14399
rect 12492 14368 13001 14396
rect 12492 14356 12498 14368
rect 12989 14365 13001 14368
rect 13035 14365 13047 14399
rect 12989 14359 13047 14365
rect 13173 14399 13231 14405
rect 13173 14365 13185 14399
rect 13219 14365 13231 14399
rect 13538 14396 13544 14408
rect 13499 14368 13544 14396
rect 13173 14359 13231 14365
rect 11054 14328 11060 14340
rect 10967 14300 11060 14328
rect 11054 14288 11060 14300
rect 11112 14288 11118 14340
rect 12618 14328 12624 14340
rect 11256 14300 12020 14328
rect 7650 14260 7656 14272
rect 7611 14232 7656 14260
rect 7650 14220 7656 14232
rect 7708 14220 7714 14272
rect 8754 14220 8760 14272
rect 8812 14260 8818 14272
rect 10410 14260 10416 14272
rect 8812 14232 10416 14260
rect 8812 14220 8818 14232
rect 10410 14220 10416 14232
rect 10468 14260 10474 14272
rect 11256 14260 11284 14300
rect 10468 14232 11284 14260
rect 11333 14263 11391 14269
rect 10468 14220 10474 14232
rect 11333 14229 11345 14263
rect 11379 14260 11391 14263
rect 11882 14260 11888 14272
rect 11379 14232 11888 14260
rect 11379 14229 11391 14232
rect 11333 14223 11391 14229
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 11992 14260 12020 14300
rect 12360 14300 12624 14328
rect 12360 14260 12388 14300
rect 12618 14288 12624 14300
rect 12676 14288 12682 14340
rect 11992 14232 12388 14260
rect 12526 14220 12532 14272
rect 12584 14260 12590 14272
rect 13078 14260 13084 14272
rect 12584 14232 13084 14260
rect 12584 14220 12590 14232
rect 13078 14220 13084 14232
rect 13136 14220 13142 14272
rect 13188 14260 13216 14359
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 14568 14328 14596 14436
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 15194 14356 15200 14408
rect 15252 14396 15258 14408
rect 15856 14405 15884 14504
rect 15948 14504 18552 14532
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15252 14368 15761 14396
rect 15252 14356 15258 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 15948 14328 15976 14504
rect 16752 14467 16810 14473
rect 16752 14433 16764 14467
rect 16798 14464 16810 14467
rect 17770 14464 17776 14476
rect 16798 14436 17776 14464
rect 16798 14433 16810 14436
rect 16752 14427 16810 14433
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 17862 14424 17868 14476
rect 17920 14464 17926 14476
rect 18397 14467 18455 14473
rect 18397 14464 18409 14467
rect 17920 14436 18409 14464
rect 17920 14424 17926 14436
rect 18397 14433 18409 14436
rect 18443 14433 18455 14467
rect 18524 14464 18552 14504
rect 19518 14492 19524 14544
rect 19576 14532 19582 14544
rect 20254 14532 20260 14544
rect 19576 14504 20260 14532
rect 19576 14492 19582 14504
rect 20254 14492 20260 14504
rect 20312 14492 20318 14544
rect 20714 14464 20720 14476
rect 18524 14436 20720 14464
rect 18397 14427 18455 14433
rect 20714 14424 20720 14436
rect 20772 14424 20778 14476
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14464 20959 14467
rect 21174 14464 21180 14476
rect 20947 14436 21180 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 21174 14424 21180 14436
rect 21232 14424 21238 14476
rect 16485 14399 16543 14405
rect 16485 14396 16497 14399
rect 14568 14300 15976 14328
rect 16408 14368 16497 14396
rect 16408 14272 16436 14368
rect 16485 14365 16497 14368
rect 16531 14365 16543 14399
rect 16485 14359 16543 14365
rect 17494 14356 17500 14408
rect 17552 14396 17558 14408
rect 18046 14396 18052 14408
rect 17552 14368 18052 14396
rect 17552 14356 17558 14368
rect 18046 14356 18052 14368
rect 18104 14396 18110 14408
rect 18141 14399 18199 14405
rect 18141 14396 18153 14399
rect 18104 14368 18153 14396
rect 18104 14356 18110 14368
rect 18141 14365 18153 14368
rect 18187 14365 18199 14399
rect 18141 14359 18199 14365
rect 19886 14356 19892 14408
rect 19944 14396 19950 14408
rect 20349 14399 20407 14405
rect 20349 14396 20361 14399
rect 19944 14368 20361 14396
rect 19944 14356 19950 14368
rect 20349 14365 20361 14368
rect 20395 14365 20407 14399
rect 20349 14359 20407 14365
rect 14274 14260 14280 14272
rect 13188 14232 14280 14260
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 14734 14220 14740 14272
rect 14792 14260 14798 14272
rect 14921 14263 14979 14269
rect 14921 14260 14933 14263
rect 14792 14232 14933 14260
rect 14792 14220 14798 14232
rect 14921 14229 14933 14232
rect 14967 14229 14979 14263
rect 15286 14260 15292 14272
rect 15247 14232 15292 14260
rect 14921 14223 14979 14229
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 15746 14220 15752 14272
rect 15804 14260 15810 14272
rect 16390 14260 16396 14272
rect 15804 14232 16396 14260
rect 15804 14220 15810 14232
rect 16390 14220 16396 14232
rect 16448 14260 16454 14272
rect 17512 14260 17540 14356
rect 16448 14232 17540 14260
rect 16448 14220 16454 14232
rect 17678 14220 17684 14272
rect 17736 14260 17742 14272
rect 17862 14260 17868 14272
rect 17736 14232 17868 14260
rect 17736 14220 17742 14232
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 17954 14220 17960 14272
rect 18012 14260 18018 14272
rect 19521 14263 19579 14269
rect 19521 14260 19533 14263
rect 18012 14232 19533 14260
rect 18012 14220 18018 14232
rect 19521 14229 19533 14232
rect 19567 14229 19579 14263
rect 19521 14223 19579 14229
rect 19705 14263 19763 14269
rect 19705 14229 19717 14263
rect 19751 14260 19763 14263
rect 20346 14260 20352 14272
rect 19751 14232 20352 14260
rect 19751 14229 19763 14232
rect 19705 14223 19763 14229
rect 20346 14220 20352 14232
rect 20404 14220 20410 14272
rect 20622 14220 20628 14272
rect 20680 14260 20686 14272
rect 21085 14263 21143 14269
rect 21085 14260 21097 14263
rect 20680 14232 21097 14260
rect 20680 14220 20686 14232
rect 21085 14229 21097 14232
rect 21131 14229 21143 14263
rect 21085 14223 21143 14229
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 6454 14056 6460 14068
rect 6415 14028 6460 14056
rect 6454 14016 6460 14028
rect 6512 14016 6518 14068
rect 7285 14059 7343 14065
rect 7285 14025 7297 14059
rect 7331 14056 7343 14059
rect 7558 14056 7564 14068
rect 7331 14028 7564 14056
rect 7331 14025 7343 14028
rect 7285 14019 7343 14025
rect 7558 14016 7564 14028
rect 7616 14016 7622 14068
rect 7650 14016 7656 14068
rect 7708 14056 7714 14068
rect 8021 14059 8079 14065
rect 8021 14056 8033 14059
rect 7708 14028 8033 14056
rect 7708 14016 7714 14028
rect 8021 14025 8033 14028
rect 8067 14056 8079 14059
rect 8389 14059 8447 14065
rect 8389 14056 8401 14059
rect 8067 14028 8401 14056
rect 8067 14025 8079 14028
rect 8021 14019 8079 14025
rect 8389 14025 8401 14028
rect 8435 14056 8447 14059
rect 9030 14056 9036 14068
rect 8435 14028 9036 14056
rect 8435 14025 8447 14028
rect 8389 14019 8447 14025
rect 9030 14016 9036 14028
rect 9088 14016 9094 14068
rect 9766 14056 9772 14068
rect 9727 14028 9772 14056
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10870 14016 10876 14068
rect 10928 14056 10934 14068
rect 10928 14028 12296 14056
rect 10928 14016 10934 14028
rect 6917 13991 6975 13997
rect 6917 13957 6929 13991
rect 6963 13988 6975 13991
rect 7742 13988 7748 14000
rect 6963 13960 7748 13988
rect 6963 13957 6975 13960
rect 6917 13951 6975 13957
rect 7742 13948 7748 13960
rect 7800 13948 7806 14000
rect 8757 13991 8815 13997
rect 8757 13957 8769 13991
rect 8803 13988 8815 13991
rect 8938 13988 8944 14000
rect 8803 13960 8944 13988
rect 8803 13957 8815 13960
rect 8757 13951 8815 13957
rect 8938 13948 8944 13960
rect 8996 13948 9002 14000
rect 9784 13920 9812 14016
rect 12268 13988 12296 14028
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 13170 14056 13176 14068
rect 12492 14028 13176 14056
rect 12492 14016 12498 14028
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 14093 14059 14151 14065
rect 14093 14056 14105 14059
rect 13780 14028 14105 14056
rect 13780 14016 13786 14028
rect 14093 14025 14105 14028
rect 14139 14025 14151 14059
rect 14826 14056 14832 14068
rect 14093 14019 14151 14025
rect 14200 14028 14832 14056
rect 13814 13988 13820 14000
rect 12268 13960 12388 13988
rect 13727 13960 13820 13988
rect 10134 13920 10140 13932
rect 9784 13892 10140 13920
rect 10134 13880 10140 13892
rect 10192 13920 10198 13932
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 10192 13892 10241 13920
rect 10192 13880 10198 13892
rect 10229 13889 10241 13892
rect 10275 13889 10287 13923
rect 10229 13883 10287 13889
rect 11698 13880 11704 13932
rect 11756 13880 11762 13932
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 7561 13855 7619 13861
rect 7561 13852 7573 13855
rect 7340 13824 7573 13852
rect 7340 13812 7346 13824
rect 7561 13821 7573 13824
rect 7607 13821 7619 13855
rect 7561 13815 7619 13821
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 9033 13855 9091 13861
rect 9033 13852 9045 13855
rect 8812 13824 9045 13852
rect 8812 13812 8818 13824
rect 9033 13821 9045 13824
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13852 9551 13855
rect 9950 13852 9956 13864
rect 9539 13824 9812 13852
rect 9911 13824 9956 13852
rect 9539 13821 9551 13824
rect 9493 13815 9551 13821
rect 8938 13744 8944 13796
rect 8996 13784 9002 13796
rect 9398 13784 9404 13796
rect 8996 13756 9404 13784
rect 8996 13744 9002 13756
rect 9398 13744 9404 13756
rect 9456 13744 9462 13796
rect 9784 13784 9812 13824
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 10496 13855 10554 13861
rect 10496 13821 10508 13855
rect 10542 13852 10554 13855
rect 11054 13852 11060 13864
rect 10542 13824 11060 13852
rect 10542 13821 10554 13824
rect 10496 13815 10554 13821
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 11716 13784 11744 13880
rect 12250 13784 12256 13796
rect 9784 13756 12256 13784
rect 12250 13744 12256 13756
rect 12308 13744 12314 13796
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 11609 13719 11667 13725
rect 11609 13716 11621 13719
rect 11388 13688 11621 13716
rect 11388 13676 11394 13688
rect 11609 13685 11621 13688
rect 11655 13685 11667 13719
rect 11609 13679 11667 13685
rect 11698 13676 11704 13728
rect 11756 13716 11762 13728
rect 11885 13719 11943 13725
rect 11885 13716 11897 13719
rect 11756 13688 11897 13716
rect 11756 13676 11762 13688
rect 11885 13685 11897 13688
rect 11931 13685 11943 13719
rect 12360 13716 12388 13960
rect 13814 13948 13820 13960
rect 13872 13988 13878 14000
rect 14200 13988 14228 14028
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 15194 14056 15200 14068
rect 15155 14028 15200 14056
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 17681 14059 17739 14065
rect 15948 14028 17540 14056
rect 15746 13988 15752 14000
rect 13872 13960 14228 13988
rect 14476 13960 15752 13988
rect 13872 13948 13878 13960
rect 13538 13880 13544 13932
rect 13596 13920 13602 13932
rect 14476 13920 14504 13960
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 13596 13892 14504 13920
rect 14553 13923 14611 13929
rect 13596 13880 13602 13892
rect 14553 13889 14565 13923
rect 14599 13920 14611 13923
rect 14642 13920 14648 13932
rect 14599 13892 14648 13920
rect 14599 13889 14611 13892
rect 14553 13883 14611 13889
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13920 14795 13923
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 14783 13892 15853 13920
rect 14783 13889 14795 13892
rect 14737 13883 14795 13889
rect 15841 13889 15853 13892
rect 15887 13920 15899 13923
rect 15948 13920 15976 14028
rect 16577 13991 16635 13997
rect 16577 13957 16589 13991
rect 16623 13988 16635 13991
rect 17402 13988 17408 14000
rect 16623 13960 17408 13988
rect 16623 13957 16635 13960
rect 16577 13951 16635 13957
rect 17402 13948 17408 13960
rect 17460 13948 17466 14000
rect 17512 13988 17540 14028
rect 17681 14025 17693 14059
rect 17727 14056 17739 14059
rect 20438 14056 20444 14068
rect 17727 14028 20444 14056
rect 17727 14025 17739 14028
rect 17681 14019 17739 14025
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 17954 13988 17960 14000
rect 17512 13960 17960 13988
rect 17954 13948 17960 13960
rect 18012 13948 18018 14000
rect 20346 13948 20352 14000
rect 20404 13988 20410 14000
rect 20625 13991 20683 13997
rect 20625 13988 20637 13991
rect 20404 13960 20637 13988
rect 20404 13948 20410 13960
rect 20625 13957 20637 13960
rect 20671 13957 20683 13991
rect 20625 13951 20683 13957
rect 17034 13920 17040 13932
rect 15887 13892 15976 13920
rect 16995 13892 17040 13920
rect 15887 13889 15899 13892
rect 15841 13883 15899 13889
rect 12437 13855 12495 13861
rect 12437 13821 12449 13855
rect 12483 13852 12495 13855
rect 12526 13852 12532 13864
rect 12483 13824 12532 13852
rect 12483 13821 12495 13824
rect 12437 13815 12495 13821
rect 12526 13812 12532 13824
rect 12584 13812 12590 13864
rect 12704 13855 12762 13861
rect 12704 13821 12716 13855
rect 12750 13852 12762 13855
rect 14366 13852 14372 13864
rect 12750 13824 14372 13852
rect 12750 13821 12762 13824
rect 12704 13815 12762 13821
rect 14366 13812 14372 13824
rect 14424 13852 14430 13864
rect 14752 13852 14780 13883
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 17221 13923 17279 13929
rect 17221 13889 17233 13923
rect 17267 13920 17279 13923
rect 18690 13920 18696 13932
rect 17267 13892 18696 13920
rect 17267 13889 17279 13892
rect 17221 13883 17279 13889
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13920 21235 13923
rect 21542 13920 21548 13932
rect 21223 13892 21548 13920
rect 21223 13889 21235 13892
rect 21177 13883 21235 13889
rect 21542 13880 21548 13892
rect 21600 13880 21606 13932
rect 14424 13824 14780 13852
rect 14424 13812 14430 13824
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 15657 13855 15715 13861
rect 15657 13852 15669 13855
rect 15252 13824 15669 13852
rect 15252 13812 15258 13824
rect 15657 13821 15669 13824
rect 15703 13852 15715 13855
rect 15746 13852 15752 13864
rect 15703 13824 15752 13852
rect 15703 13821 15715 13824
rect 15657 13815 15715 13821
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 15930 13812 15936 13864
rect 15988 13852 15994 13864
rect 16209 13855 16267 13861
rect 16209 13852 16221 13855
rect 15988 13824 16221 13852
rect 15988 13812 15994 13824
rect 16209 13821 16221 13824
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 16574 13812 16580 13864
rect 16632 13852 16638 13864
rect 18509 13855 18567 13861
rect 18509 13852 18521 13855
rect 16632 13824 18521 13852
rect 16632 13812 16638 13824
rect 18509 13821 18521 13824
rect 18555 13821 18567 13855
rect 18509 13815 18567 13821
rect 18874 13812 18880 13864
rect 18932 13852 18938 13864
rect 19245 13855 19303 13861
rect 19245 13852 19257 13855
rect 18932 13824 19257 13852
rect 18932 13812 18938 13824
rect 19245 13821 19257 13824
rect 19291 13821 19303 13855
rect 19245 13815 19303 13821
rect 19512 13855 19570 13861
rect 19512 13821 19524 13855
rect 19558 13852 19570 13855
rect 19886 13852 19892 13864
rect 19558 13824 19892 13852
rect 19558 13821 19570 13824
rect 19512 13815 19570 13821
rect 19886 13812 19892 13824
rect 19944 13812 19950 13864
rect 20806 13812 20812 13864
rect 20864 13852 20870 13864
rect 20901 13855 20959 13861
rect 20901 13852 20913 13855
rect 20864 13824 20913 13852
rect 20864 13812 20870 13824
rect 20901 13821 20913 13824
rect 20947 13821 20959 13855
rect 20901 13815 20959 13821
rect 12618 13744 12624 13796
rect 12676 13784 12682 13796
rect 16945 13787 17003 13793
rect 16945 13784 16957 13787
rect 12676 13756 16957 13784
rect 12676 13744 12682 13756
rect 16945 13753 16957 13756
rect 16991 13753 17003 13787
rect 16945 13747 17003 13753
rect 17880 13756 20944 13784
rect 13538 13716 13544 13728
rect 12360 13688 13544 13716
rect 11885 13679 11943 13685
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 13998 13676 14004 13728
rect 14056 13716 14062 13728
rect 14461 13719 14519 13725
rect 14461 13716 14473 13719
rect 14056 13688 14473 13716
rect 14056 13676 14062 13688
rect 14461 13685 14473 13688
rect 14507 13685 14519 13719
rect 14461 13679 14519 13685
rect 15470 13676 15476 13728
rect 15528 13716 15534 13728
rect 15565 13719 15623 13725
rect 15565 13716 15577 13719
rect 15528 13688 15577 13716
rect 15528 13676 15534 13688
rect 15565 13685 15577 13688
rect 15611 13685 15623 13719
rect 15565 13679 15623 13685
rect 16206 13676 16212 13728
rect 16264 13716 16270 13728
rect 17880 13716 17908 13756
rect 20916 13728 20944 13756
rect 16264 13688 17908 13716
rect 16264 13676 16270 13688
rect 17954 13676 17960 13728
rect 18012 13716 18018 13728
rect 18049 13719 18107 13725
rect 18049 13716 18061 13719
rect 18012 13688 18061 13716
rect 18012 13676 18018 13688
rect 18049 13685 18061 13688
rect 18095 13685 18107 13719
rect 18414 13716 18420 13728
rect 18375 13688 18420 13716
rect 18049 13679 18107 13685
rect 18414 13676 18420 13688
rect 18472 13676 18478 13728
rect 20898 13676 20904 13728
rect 20956 13676 20962 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 7006 13472 7012 13524
rect 7064 13512 7070 13524
rect 8113 13515 8171 13521
rect 8113 13512 8125 13515
rect 7064 13484 8125 13512
rect 7064 13472 7070 13484
rect 8113 13481 8125 13484
rect 8159 13512 8171 13515
rect 8202 13512 8208 13524
rect 8159 13484 8208 13512
rect 8159 13481 8171 13484
rect 8113 13475 8171 13481
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 10686 13472 10692 13524
rect 10744 13512 10750 13524
rect 10870 13512 10876 13524
rect 10744 13484 10876 13512
rect 10744 13472 10750 13484
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 11425 13515 11483 13521
rect 11425 13481 11437 13515
rect 11471 13481 11483 13515
rect 11882 13512 11888 13524
rect 11843 13484 11888 13512
rect 11425 13475 11483 13481
rect 7466 13444 7472 13456
rect 7427 13416 7472 13444
rect 7466 13404 7472 13416
rect 7524 13404 7530 13456
rect 7650 13404 7656 13456
rect 7708 13444 7714 13456
rect 7745 13447 7803 13453
rect 7745 13444 7757 13447
rect 7708 13416 7757 13444
rect 7708 13404 7714 13416
rect 7745 13413 7757 13416
rect 7791 13413 7803 13447
rect 9122 13444 9128 13456
rect 9083 13416 9128 13444
rect 7745 13407 7803 13413
rect 9122 13404 9128 13416
rect 9180 13404 9186 13456
rect 9674 13444 9680 13456
rect 9600 13416 9680 13444
rect 8849 13379 8907 13385
rect 8849 13345 8861 13379
rect 8895 13376 8907 13379
rect 9600 13376 9628 13416
rect 9674 13404 9680 13416
rect 9732 13404 9738 13456
rect 10036 13447 10094 13453
rect 10036 13413 10048 13447
rect 10082 13444 10094 13447
rect 11330 13444 11336 13456
rect 10082 13416 11336 13444
rect 10082 13413 10094 13416
rect 10036 13407 10094 13413
rect 11330 13404 11336 13416
rect 11388 13404 11394 13456
rect 11440 13444 11468 13475
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 12897 13515 12955 13521
rect 12897 13512 12909 13515
rect 11992 13484 12909 13512
rect 11992 13444 12020 13484
rect 12897 13481 12909 13484
rect 12943 13481 12955 13515
rect 12897 13475 12955 13481
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 13722 13512 13728 13524
rect 13504 13484 13728 13512
rect 13504 13472 13510 13484
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 14550 13512 14556 13524
rect 14511 13484 14556 13512
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 15381 13515 15439 13521
rect 15381 13481 15393 13515
rect 15427 13481 15439 13515
rect 15381 13475 15439 13481
rect 15749 13515 15807 13521
rect 15749 13481 15761 13515
rect 15795 13512 15807 13515
rect 16942 13512 16948 13524
rect 15795 13484 16948 13512
rect 15795 13481 15807 13484
rect 15749 13475 15807 13481
rect 11440 13416 12020 13444
rect 12618 13404 12624 13456
rect 12676 13444 12682 13456
rect 13464 13444 13492 13472
rect 12676 13416 13492 13444
rect 12676 13404 12682 13416
rect 13538 13404 13544 13456
rect 13596 13444 13602 13456
rect 14645 13447 14703 13453
rect 14645 13444 14657 13447
rect 13596 13416 14657 13444
rect 13596 13404 13602 13416
rect 14645 13413 14657 13416
rect 14691 13413 14703 13447
rect 15396 13444 15424 13475
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 17770 13512 17776 13524
rect 17731 13484 17776 13512
rect 17770 13472 17776 13484
rect 17828 13472 17834 13524
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 20162 13512 20168 13524
rect 17920 13484 20168 13512
rect 17920 13472 17926 13484
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 21174 13444 21180 13456
rect 15396 13416 20944 13444
rect 21135 13416 21180 13444
rect 14645 13407 14703 13413
rect 9766 13376 9772 13388
rect 8895 13348 9628 13376
rect 9727 13348 9772 13376
rect 8895 13345 8907 13348
rect 8849 13339 8907 13345
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 11790 13376 11796 13388
rect 11751 13348 11796 13376
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 12066 13336 12072 13388
rect 12124 13376 12130 13388
rect 12805 13379 12863 13385
rect 12805 13376 12817 13379
rect 12124 13348 12817 13376
rect 12124 13336 12130 13348
rect 12805 13345 12817 13348
rect 12851 13345 12863 13379
rect 13446 13376 13452 13388
rect 13407 13348 13452 13376
rect 12805 13339 12863 13345
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 15194 13336 15200 13388
rect 15252 13376 15258 13388
rect 16390 13376 16396 13388
rect 15252 13348 16396 13376
rect 15252 13336 15258 13348
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 16660 13379 16718 13385
rect 16660 13345 16672 13379
rect 16706 13376 16718 13379
rect 16706 13348 18000 13376
rect 16706 13345 16718 13348
rect 16660 13339 16718 13345
rect 6270 13268 6276 13320
rect 6328 13308 6334 13320
rect 7101 13311 7159 13317
rect 7101 13308 7113 13311
rect 6328 13280 7113 13308
rect 6328 13268 6334 13280
rect 7101 13277 7113 13280
rect 7147 13308 7159 13311
rect 9490 13308 9496 13320
rect 7147 13280 9496 13308
rect 7147 13277 7159 13280
rect 7101 13271 7159 13277
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 11882 13308 11888 13320
rect 11388 13280 11888 13308
rect 11388 13268 11394 13280
rect 11882 13268 11888 13280
rect 11940 13308 11946 13320
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 11940 13280 11989 13308
rect 11940 13268 11946 13280
rect 11977 13277 11989 13280
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13277 13047 13311
rect 13630 13308 13636 13320
rect 13591 13280 13636 13308
rect 12989 13271 13047 13277
rect 6638 13200 6644 13252
rect 6696 13240 6702 13252
rect 9766 13240 9772 13252
rect 6696 13212 9772 13240
rect 6696 13200 6702 13212
rect 9766 13200 9772 13212
rect 9824 13200 9830 13252
rect 12434 13240 12440 13252
rect 12395 13212 12440 13240
rect 12434 13200 12440 13212
rect 12492 13200 12498 13252
rect 13004 13240 13032 13271
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 14366 13268 14372 13320
rect 14424 13308 14430 13320
rect 14737 13311 14795 13317
rect 14737 13308 14749 13311
rect 14424 13280 14749 13308
rect 14424 13268 14430 13280
rect 14737 13277 14749 13280
rect 14783 13277 14795 13311
rect 15838 13308 15844 13320
rect 15799 13280 15844 13308
rect 14737 13271 14795 13277
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 16025 13311 16083 13317
rect 16025 13277 16037 13311
rect 16071 13277 16083 13311
rect 16025 13271 16083 13277
rect 12544 13212 13032 13240
rect 14185 13243 14243 13249
rect 7466 13132 7472 13184
rect 7524 13172 7530 13184
rect 7742 13172 7748 13184
rect 7524 13144 7748 13172
rect 7524 13132 7530 13144
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 8573 13175 8631 13181
rect 8573 13141 8585 13175
rect 8619 13172 8631 13175
rect 8662 13172 8668 13184
rect 8619 13144 8668 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 11146 13172 11152 13184
rect 11059 13144 11152 13172
rect 11146 13132 11152 13144
rect 11204 13172 11210 13184
rect 12544 13172 12572 13212
rect 14185 13209 14197 13243
rect 14231 13240 14243 13243
rect 15654 13240 15660 13252
rect 14231 13212 15660 13240
rect 14231 13209 14243 13212
rect 14185 13203 14243 13209
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 11204 13144 12572 13172
rect 11204 13132 11210 13144
rect 12986 13132 12992 13184
rect 13044 13172 13050 13184
rect 13262 13172 13268 13184
rect 13044 13144 13268 13172
rect 13044 13132 13050 13144
rect 13262 13132 13268 13144
rect 13320 13132 13326 13184
rect 13630 13132 13636 13184
rect 13688 13172 13694 13184
rect 13998 13172 14004 13184
rect 13688 13144 14004 13172
rect 13688 13132 13694 13144
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 16040 13172 16068 13271
rect 17972 13240 18000 13348
rect 18322 13336 18328 13388
rect 18380 13376 18386 13388
rect 18417 13379 18475 13385
rect 18417 13376 18429 13379
rect 18380 13348 18429 13376
rect 18380 13336 18386 13348
rect 18417 13345 18429 13348
rect 18463 13345 18475 13379
rect 18417 13339 18475 13345
rect 18598 13336 18604 13388
rect 18656 13376 18662 13388
rect 19426 13385 19432 13388
rect 19409 13379 19432 13385
rect 19409 13376 19421 13379
rect 18656 13348 19421 13376
rect 18656 13336 18662 13348
rect 19409 13345 19421 13348
rect 19484 13376 19490 13388
rect 20916 13385 20944 13416
rect 21174 13404 21180 13416
rect 21232 13404 21238 13456
rect 20901 13379 20959 13385
rect 19484 13348 19557 13376
rect 19409 13339 19432 13345
rect 19426 13336 19432 13339
rect 19484 13336 19490 13348
rect 20901 13345 20913 13379
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 18506 13308 18512 13320
rect 18467 13280 18512 13308
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 18690 13308 18696 13320
rect 18651 13280 18696 13308
rect 18690 13268 18696 13280
rect 18748 13268 18754 13320
rect 18874 13268 18880 13320
rect 18932 13308 18938 13320
rect 19153 13311 19211 13317
rect 19153 13308 19165 13311
rect 18932 13280 19165 13308
rect 18932 13268 18938 13280
rect 19153 13277 19165 13280
rect 19199 13277 19211 13311
rect 19153 13271 19211 13277
rect 18708 13240 18736 13268
rect 17972 13212 18736 13240
rect 17678 13172 17684 13184
rect 16040 13144 17684 13172
rect 17678 13132 17684 13144
rect 17736 13132 17742 13184
rect 18046 13172 18052 13184
rect 18007 13144 18052 13172
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 18966 13132 18972 13184
rect 19024 13172 19030 13184
rect 20533 13175 20591 13181
rect 20533 13172 20545 13175
rect 19024 13144 20545 13172
rect 19024 13132 19030 13144
rect 20533 13141 20545 13144
rect 20579 13141 20591 13175
rect 20533 13135 20591 13141
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 7432 12940 7849 12968
rect 7432 12928 7438 12940
rect 7837 12937 7849 12940
rect 7883 12968 7895 12971
rect 9858 12968 9864 12980
rect 7883 12940 9864 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 9858 12928 9864 12940
rect 9916 12968 9922 12980
rect 10870 12968 10876 12980
rect 9916 12940 10876 12968
rect 9916 12928 9922 12940
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 11057 12971 11115 12977
rect 11057 12937 11069 12971
rect 11103 12968 11115 12971
rect 12066 12968 12072 12980
rect 11103 12940 12072 12968
rect 11103 12937 11115 12940
rect 11057 12931 11115 12937
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 13173 12971 13231 12977
rect 13173 12937 13185 12971
rect 13219 12968 13231 12971
rect 15746 12968 15752 12980
rect 13219 12940 15752 12968
rect 13219 12937 13231 12940
rect 13173 12931 13231 12937
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 16945 12971 17003 12977
rect 16945 12968 16957 12971
rect 15896 12940 16957 12968
rect 15896 12928 15902 12940
rect 16945 12937 16957 12940
rect 16991 12937 17003 12971
rect 16945 12931 17003 12937
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 18598 12968 18604 12980
rect 17184 12940 18604 12968
rect 17184 12928 17190 12940
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 18748 12940 20085 12968
rect 18748 12928 18754 12940
rect 20073 12937 20085 12940
rect 20119 12937 20131 12971
rect 20073 12931 20131 12937
rect 10045 12903 10103 12909
rect 10045 12869 10057 12903
rect 10091 12900 10103 12903
rect 13446 12900 13452 12912
rect 10091 12872 13452 12900
rect 10091 12869 10103 12872
rect 10045 12863 10103 12869
rect 13446 12860 13452 12872
rect 13504 12860 13510 12912
rect 16206 12900 16212 12912
rect 13740 12872 16212 12900
rect 6638 12792 6644 12844
rect 6696 12832 6702 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6696 12804 7389 12832
rect 6696 12792 6702 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 10502 12832 10508 12844
rect 10463 12804 10508 12832
rect 7377 12795 7435 12801
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 10689 12835 10747 12841
rect 10689 12801 10701 12835
rect 10735 12832 10747 12835
rect 11054 12832 11060 12844
rect 10735 12804 11060 12832
rect 10735 12801 10747 12804
rect 10689 12795 10747 12801
rect 11054 12792 11060 12804
rect 11112 12792 11118 12844
rect 11609 12835 11667 12841
rect 11609 12801 11621 12835
rect 11655 12832 11667 12835
rect 11882 12832 11888 12844
rect 11655 12804 11888 12832
rect 11655 12801 11667 12804
rect 11609 12795 11667 12801
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 12066 12792 12072 12844
rect 12124 12832 12130 12844
rect 12618 12832 12624 12844
rect 12124 12804 12624 12832
rect 12124 12792 12130 12804
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12832 12771 12835
rect 13740 12832 13768 12872
rect 16206 12860 16212 12872
rect 16264 12860 16270 12912
rect 20441 12903 20499 12909
rect 16316 12872 18276 12900
rect 12759 12804 13768 12832
rect 13817 12835 13875 12841
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 13817 12801 13829 12835
rect 13863 12832 13875 12835
rect 14366 12832 14372 12844
rect 13863 12804 14372 12832
rect 13863 12801 13875 12804
rect 13817 12795 13875 12801
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 14734 12832 14740 12844
rect 14695 12804 14740 12832
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 8113 12767 8171 12773
rect 8113 12733 8125 12767
rect 8159 12733 8171 12767
rect 8113 12727 8171 12733
rect 8380 12767 8438 12773
rect 8380 12733 8392 12767
rect 8426 12764 8438 12767
rect 11146 12764 11152 12776
rect 8426 12736 11152 12764
rect 8426 12733 8438 12736
rect 8380 12727 8438 12733
rect 8128 12696 8156 12727
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 11425 12767 11483 12773
rect 11425 12733 11437 12767
rect 11471 12764 11483 12767
rect 11698 12764 11704 12776
rect 11471 12736 11704 12764
rect 11471 12733 11483 12736
rect 11425 12727 11483 12733
rect 11698 12724 11704 12736
rect 11756 12724 11762 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 14090 12764 14096 12776
rect 12492 12736 12537 12764
rect 12636 12736 14096 12764
rect 12492 12724 12498 12736
rect 10134 12696 10140 12708
rect 8128 12668 10140 12696
rect 10134 12656 10140 12668
rect 10192 12656 10198 12708
rect 10413 12699 10471 12705
rect 10413 12665 10425 12699
rect 10459 12696 10471 12699
rect 12636 12696 12664 12736
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 16316 12773 16344 12872
rect 16577 12835 16635 12841
rect 16577 12801 16589 12835
rect 16623 12832 16635 12835
rect 17126 12832 17132 12844
rect 16623 12804 17132 12832
rect 16623 12801 16635 12804
rect 16577 12795 16635 12801
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12832 17647 12835
rect 17770 12832 17776 12844
rect 17635 12804 17776 12832
rect 17635 12801 17647 12804
rect 17589 12795 17647 12801
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 14200 12736 15209 12764
rect 13541 12699 13599 12705
rect 13541 12696 13553 12699
rect 10459 12668 12664 12696
rect 12820 12668 13553 12696
rect 10459 12665 10471 12668
rect 10413 12659 10471 12665
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 9493 12631 9551 12637
rect 9493 12628 9505 12631
rect 9456 12600 9505 12628
rect 9456 12588 9462 12600
rect 9493 12597 9505 12600
rect 9539 12597 9551 12631
rect 9493 12591 9551 12597
rect 9858 12588 9864 12640
rect 9916 12628 9922 12640
rect 10594 12628 10600 12640
rect 9916 12600 10600 12628
rect 9916 12588 9922 12600
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 11296 12600 11529 12628
rect 11296 12588 11302 12600
rect 11517 12597 11529 12600
rect 11563 12628 11575 12631
rect 11790 12628 11796 12640
rect 11563 12600 11796 12628
rect 11563 12597 11575 12600
rect 11517 12591 11575 12597
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 12250 12588 12256 12640
rect 12308 12628 12314 12640
rect 12618 12628 12624 12640
rect 12308 12600 12624 12628
rect 12308 12588 12314 12600
rect 12618 12588 12624 12600
rect 12676 12628 12682 12640
rect 12820 12628 12848 12668
rect 13541 12665 13553 12668
rect 13587 12665 13599 12699
rect 13541 12659 13599 12665
rect 13633 12699 13691 12705
rect 13633 12665 13645 12699
rect 13679 12696 13691 12699
rect 13722 12696 13728 12708
rect 13679 12668 13728 12696
rect 13679 12665 13691 12668
rect 13633 12659 13691 12665
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 14200 12637 14228 12736
rect 15197 12733 15209 12736
rect 15243 12733 15255 12767
rect 15197 12727 15255 12733
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12733 16359 12767
rect 16301 12727 16359 12733
rect 17405 12767 17463 12773
rect 17405 12733 17417 12767
rect 17451 12764 17463 12767
rect 18046 12764 18052 12776
rect 17451 12736 18052 12764
rect 17451 12733 17463 12736
rect 17405 12727 17463 12733
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 14553 12699 14611 12705
rect 14553 12665 14565 12699
rect 14599 12696 14611 12699
rect 15286 12696 15292 12708
rect 14599 12668 15292 12696
rect 14599 12665 14611 12668
rect 14553 12659 14611 12665
rect 15286 12656 15292 12668
rect 15344 12656 15350 12708
rect 15473 12699 15531 12705
rect 15473 12665 15485 12699
rect 15519 12696 15531 12699
rect 17313 12699 17371 12705
rect 15519 12668 17264 12696
rect 15519 12665 15531 12668
rect 15473 12659 15531 12665
rect 12676 12600 12848 12628
rect 14185 12631 14243 12637
rect 12676 12588 12682 12600
rect 14185 12597 14197 12631
rect 14231 12597 14243 12631
rect 14185 12591 14243 12597
rect 14458 12588 14464 12640
rect 14516 12628 14522 12640
rect 14645 12631 14703 12637
rect 14645 12628 14657 12631
rect 14516 12600 14657 12628
rect 14516 12588 14522 12600
rect 14645 12597 14657 12600
rect 14691 12597 14703 12631
rect 15930 12628 15936 12640
rect 15891 12600 15936 12628
rect 14645 12591 14703 12597
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 16022 12588 16028 12640
rect 16080 12628 16086 12640
rect 16298 12628 16304 12640
rect 16080 12600 16304 12628
rect 16080 12588 16086 12600
rect 16298 12588 16304 12600
rect 16356 12628 16362 12640
rect 16393 12631 16451 12637
rect 16393 12628 16405 12631
rect 16356 12600 16405 12628
rect 16356 12588 16362 12600
rect 16393 12597 16405 12600
rect 16439 12597 16451 12631
rect 17236 12628 17264 12668
rect 17313 12665 17325 12699
rect 17359 12696 17371 12699
rect 17954 12696 17960 12708
rect 17359 12668 17960 12696
rect 17359 12665 17371 12668
rect 17313 12659 17371 12665
rect 17954 12656 17960 12668
rect 18012 12656 18018 12708
rect 18248 12696 18276 12872
rect 20441 12869 20453 12903
rect 20487 12869 20499 12903
rect 20441 12863 20499 12869
rect 18598 12792 18604 12844
rect 18656 12832 18662 12844
rect 18693 12835 18751 12841
rect 18693 12832 18705 12835
rect 18656 12804 18705 12832
rect 18656 12792 18662 12804
rect 18693 12801 18705 12804
rect 18739 12801 18751 12835
rect 20456 12832 20484 12863
rect 18693 12795 18751 12801
rect 19720 12804 20484 12832
rect 18322 12724 18328 12776
rect 18380 12764 18386 12776
rect 18966 12773 18972 12776
rect 18960 12764 18972 12773
rect 18380 12736 18972 12764
rect 18380 12724 18386 12736
rect 18960 12727 18972 12736
rect 18966 12724 18972 12727
rect 19024 12724 19030 12776
rect 18248 12668 19003 12696
rect 17862 12628 17868 12640
rect 17236 12600 17868 12628
rect 16393 12591 16451 12597
rect 17862 12588 17868 12600
rect 17920 12588 17926 12640
rect 18049 12631 18107 12637
rect 18049 12597 18061 12631
rect 18095 12628 18107 12631
rect 18230 12628 18236 12640
rect 18095 12600 18236 12628
rect 18095 12597 18107 12600
rect 18049 12591 18107 12597
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 18598 12588 18604 12640
rect 18656 12628 18662 12640
rect 18874 12628 18880 12640
rect 18656 12600 18880 12628
rect 18656 12588 18662 12600
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 18975 12628 19003 12668
rect 19058 12656 19064 12708
rect 19116 12696 19122 12708
rect 19720 12696 19748 12804
rect 20622 12792 20628 12844
rect 20680 12832 20686 12844
rect 20993 12835 21051 12841
rect 20993 12832 21005 12835
rect 20680 12804 21005 12832
rect 20680 12792 20686 12804
rect 20993 12801 21005 12804
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 20438 12724 20444 12776
rect 20496 12764 20502 12776
rect 20809 12767 20867 12773
rect 20809 12764 20821 12767
rect 20496 12736 20821 12764
rect 20496 12724 20502 12736
rect 20809 12733 20821 12736
rect 20855 12733 20867 12767
rect 20809 12727 20867 12733
rect 19116 12668 19748 12696
rect 19116 12656 19122 12668
rect 20530 12656 20536 12708
rect 20588 12696 20594 12708
rect 20901 12699 20959 12705
rect 20901 12696 20913 12699
rect 20588 12668 20913 12696
rect 20588 12656 20594 12668
rect 20901 12665 20913 12668
rect 20947 12665 20959 12699
rect 20901 12659 20959 12665
rect 20714 12628 20720 12640
rect 18975 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 8113 12427 8171 12433
rect 8113 12424 8125 12427
rect 7340 12396 8125 12424
rect 7340 12384 7346 12396
rect 8113 12393 8125 12396
rect 8159 12424 8171 12427
rect 10137 12427 10195 12433
rect 10137 12424 10149 12427
rect 8159 12396 10149 12424
rect 8159 12393 8171 12396
rect 8113 12387 8171 12393
rect 10137 12393 10149 12396
rect 10183 12424 10195 12427
rect 14458 12424 14464 12436
rect 10183 12396 14464 12424
rect 10183 12393 10195 12396
rect 10137 12387 10195 12393
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 14553 12427 14611 12433
rect 14553 12393 14565 12427
rect 14599 12424 14611 12427
rect 15930 12424 15936 12436
rect 14599 12396 15936 12424
rect 14599 12393 14611 12396
rect 14553 12387 14611 12393
rect 15930 12384 15936 12396
rect 15988 12384 15994 12436
rect 16942 12424 16948 12436
rect 16903 12396 16948 12424
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 17402 12424 17408 12436
rect 17363 12396 17408 12424
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 18417 12427 18475 12433
rect 18417 12393 18429 12427
rect 18463 12424 18475 12427
rect 19150 12424 19156 12436
rect 18463 12396 19156 12424
rect 18463 12393 18475 12396
rect 18417 12387 18475 12393
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 20533 12427 20591 12433
rect 20533 12424 20545 12427
rect 19484 12396 20545 12424
rect 19484 12384 19490 12396
rect 20533 12393 20545 12396
rect 20579 12424 20591 12427
rect 20622 12424 20628 12436
rect 20579 12396 20628 12424
rect 20579 12393 20591 12396
rect 20533 12387 20591 12393
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 21085 12427 21143 12433
rect 21085 12393 21097 12427
rect 21131 12424 21143 12427
rect 21266 12424 21272 12436
rect 21131 12396 21272 12424
rect 21131 12393 21143 12396
rect 21085 12387 21143 12393
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 8481 12359 8539 12365
rect 8481 12325 8493 12359
rect 8527 12356 8539 12359
rect 8662 12356 8668 12368
rect 8527 12328 8668 12356
rect 8527 12325 8539 12328
rect 8481 12319 8539 12325
rect 8662 12316 8668 12328
rect 8720 12356 8726 12368
rect 9766 12356 9772 12368
rect 8720 12328 9772 12356
rect 8720 12316 8726 12328
rect 9766 12316 9772 12328
rect 9824 12356 9830 12368
rect 9950 12356 9956 12368
rect 9824 12328 9956 12356
rect 9824 12316 9830 12328
rect 9950 12316 9956 12328
rect 10008 12316 10014 12368
rect 11048 12359 11106 12365
rect 11048 12325 11060 12359
rect 11094 12356 11106 12359
rect 11238 12356 11244 12368
rect 11094 12328 11244 12356
rect 11094 12325 11106 12328
rect 11048 12319 11106 12325
rect 11238 12316 11244 12328
rect 11296 12316 11302 12368
rect 12526 12356 12532 12368
rect 11348 12328 12532 12356
rect 9214 12248 9220 12300
rect 9272 12288 9278 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 9272 12260 10057 12288
rect 9272 12248 9278 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 11348 12288 11376 12328
rect 12526 12316 12532 12328
rect 12584 12316 12590 12368
rect 13354 12316 13360 12368
rect 13412 12356 13418 12368
rect 13725 12359 13783 12365
rect 13725 12356 13737 12359
rect 13412 12328 13737 12356
rect 13412 12316 13418 12328
rect 13725 12325 13737 12328
rect 13771 12325 13783 12359
rect 13725 12319 13783 12325
rect 17313 12359 17371 12365
rect 17313 12325 17325 12359
rect 17359 12356 17371 12359
rect 18230 12356 18236 12368
rect 17359 12328 18236 12356
rect 17359 12325 17371 12328
rect 17313 12319 17371 12325
rect 18230 12316 18236 12328
rect 18288 12316 18294 12368
rect 18506 12356 18512 12368
rect 18467 12328 18512 12356
rect 18506 12316 18512 12328
rect 18564 12316 18570 12368
rect 18598 12316 18604 12368
rect 18656 12316 18662 12368
rect 18874 12316 18880 12368
rect 18932 12356 18938 12368
rect 19242 12356 19248 12368
rect 18932 12328 19248 12356
rect 18932 12316 18938 12328
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 10045 12251 10103 12257
rect 10796 12260 11376 12288
rect 10796 12232 10824 12260
rect 12342 12248 12348 12300
rect 12400 12288 12406 12300
rect 12805 12291 12863 12297
rect 12805 12288 12817 12291
rect 12400 12260 12817 12288
rect 12400 12248 12406 12260
rect 12805 12257 12817 12260
rect 12851 12257 12863 12291
rect 12805 12251 12863 12257
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12288 13507 12291
rect 14550 12288 14556 12300
rect 13495 12260 14556 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15562 12297 15568 12300
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 15252 12260 15301 12288
rect 15252 12248 15258 12260
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 15556 12288 15568 12297
rect 15523 12260 15568 12288
rect 15289 12251 15347 12257
rect 15556 12251 15568 12260
rect 15562 12248 15568 12251
rect 15620 12248 15626 12300
rect 18616 12288 18644 12316
rect 19153 12291 19211 12297
rect 19153 12288 19165 12291
rect 18616 12260 19165 12288
rect 19153 12257 19165 12260
rect 19199 12257 19211 12291
rect 19153 12251 19211 12257
rect 19420 12291 19478 12297
rect 19420 12257 19432 12291
rect 19466 12288 19478 12291
rect 20162 12288 20168 12300
rect 19466 12260 20168 12288
rect 19466 12257 19478 12260
rect 19420 12251 19478 12257
rect 20162 12248 20168 12260
rect 20220 12248 20226 12300
rect 20898 12288 20904 12300
rect 20859 12260 20904 12288
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 9122 12220 9128 12232
rect 9083 12192 9128 12220
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10778 12220 10784 12232
rect 10739 12192 10784 12220
rect 10229 12183 10287 12189
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 9582 12152 9588 12164
rect 9456 12124 9588 12152
rect 9456 12112 9462 12124
rect 9582 12112 9588 12124
rect 9640 12152 9646 12164
rect 10244 12152 10272 12183
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 12897 12223 12955 12229
rect 12897 12220 12909 12223
rect 11940 12192 12909 12220
rect 11940 12180 11946 12192
rect 12897 12189 12909 12192
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 14642 12220 14648 12232
rect 14603 12192 14648 12220
rect 12989 12183 13047 12189
rect 13004 12152 13032 12183
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12220 14887 12223
rect 17589 12223 17647 12229
rect 14875 12192 15332 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 9640 12124 10272 12152
rect 12176 12124 13032 12152
rect 9640 12112 9646 12124
rect 12176 12096 12204 12124
rect 8849 12087 8907 12093
rect 8849 12053 8861 12087
rect 8895 12084 8907 12087
rect 9214 12084 9220 12096
rect 8895 12056 9220 12084
rect 8895 12053 8907 12056
rect 8849 12047 8907 12053
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 9677 12087 9735 12093
rect 9677 12053 9689 12087
rect 9723 12084 9735 12087
rect 10134 12084 10140 12096
rect 9723 12056 10140 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 12158 12084 12164 12096
rect 12119 12056 12164 12084
rect 12158 12044 12164 12056
rect 12216 12044 12222 12096
rect 12434 12044 12440 12096
rect 12492 12084 12498 12096
rect 14182 12084 14188 12096
rect 12492 12056 12537 12084
rect 14143 12056 14188 12084
rect 12492 12044 12498 12056
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 15304 12084 15332 12192
rect 17589 12189 17601 12223
rect 17635 12220 17647 12223
rect 17770 12220 17776 12232
rect 17635 12192 17776 12220
rect 17635 12189 17647 12192
rect 17589 12183 17647 12189
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 18690 12220 18696 12232
rect 18651 12192 18696 12220
rect 18690 12180 18696 12192
rect 18748 12180 18754 12232
rect 18322 12152 18328 12164
rect 16224 12124 18328 12152
rect 16224 12084 16252 12124
rect 18322 12112 18328 12124
rect 18380 12112 18386 12164
rect 16666 12084 16672 12096
rect 15304 12056 16252 12084
rect 16627 12056 16672 12084
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 18049 12087 18107 12093
rect 18049 12084 18061 12087
rect 17368 12056 18061 12084
rect 17368 12044 17374 12056
rect 18049 12053 18061 12056
rect 18095 12053 18107 12087
rect 18049 12047 18107 12053
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 8846 11840 8852 11892
rect 8904 11880 8910 11892
rect 9306 11880 9312 11892
rect 8904 11852 9312 11880
rect 8904 11840 8910 11852
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11609 11883 11667 11889
rect 11609 11880 11621 11883
rect 11296 11852 11621 11880
rect 11296 11840 11302 11852
rect 11609 11849 11621 11852
rect 11655 11849 11667 11883
rect 17954 11880 17960 11892
rect 11609 11843 11667 11849
rect 14292 11852 17960 11880
rect 12342 11704 12348 11756
rect 12400 11744 12406 11756
rect 12437 11747 12495 11753
rect 12437 11744 12449 11747
rect 12400 11716 12449 11744
rect 12400 11704 12406 11716
rect 12437 11713 12449 11716
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 12526 11704 12532 11756
rect 12584 11744 12590 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12584 11716 13001 11744
rect 12584 11704 12590 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11645 8631 11679
rect 8573 11639 8631 11645
rect 8840 11679 8898 11685
rect 8840 11645 8852 11679
rect 8886 11676 8898 11679
rect 9582 11676 9588 11688
rect 8886 11648 9588 11676
rect 8886 11645 8898 11648
rect 8840 11639 8898 11645
rect 8588 11608 8616 11639
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 10226 11676 10232 11688
rect 9876 11648 10232 11676
rect 9876 11608 9904 11648
rect 10226 11636 10232 11648
rect 10284 11676 10290 11688
rect 10778 11676 10784 11688
rect 10284 11648 10784 11676
rect 10284 11636 10290 11648
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 10318 11608 10324 11620
rect 8588 11580 9904 11608
rect 9968 11580 10324 11608
rect 9968 11549 9996 11580
rect 10318 11568 10324 11580
rect 10376 11608 10382 11620
rect 10474 11611 10532 11617
rect 10474 11608 10486 11611
rect 10376 11580 10486 11608
rect 10376 11568 10382 11580
rect 10474 11577 10486 11580
rect 10520 11577 10532 11611
rect 10474 11571 10532 11577
rect 13256 11611 13314 11617
rect 13256 11577 13268 11611
rect 13302 11608 13314 11611
rect 13814 11608 13820 11620
rect 13302 11580 13820 11608
rect 13302 11577 13314 11580
rect 13256 11571 13314 11577
rect 13814 11568 13820 11580
rect 13872 11568 13878 11620
rect 9953 11543 10011 11549
rect 9953 11509 9965 11543
rect 9999 11509 10011 11543
rect 9953 11503 10011 11509
rect 11146 11500 11152 11552
rect 11204 11540 11210 11552
rect 11977 11543 12035 11549
rect 11977 11540 11989 11543
rect 11204 11512 11989 11540
rect 11204 11500 11210 11512
rect 11977 11509 11989 11512
rect 12023 11509 12035 11543
rect 11977 11503 12035 11509
rect 12342 11500 12348 11552
rect 12400 11540 12406 11552
rect 14292 11540 14320 11852
rect 17954 11840 17960 11852
rect 18012 11840 18018 11892
rect 18598 11840 18604 11892
rect 18656 11880 18662 11892
rect 19794 11880 19800 11892
rect 18656 11852 19800 11880
rect 18656 11840 18662 11852
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 20162 11880 20168 11892
rect 20123 11852 20168 11880
rect 20162 11840 20168 11852
rect 20220 11840 20226 11892
rect 20530 11880 20536 11892
rect 20491 11852 20536 11880
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 14366 11772 14372 11824
rect 14424 11812 14430 11824
rect 16945 11815 17003 11821
rect 14424 11784 14469 11812
rect 14424 11772 14430 11784
rect 16945 11781 16957 11815
rect 16991 11812 17003 11815
rect 16991 11784 18092 11812
rect 16991 11781 17003 11784
rect 16945 11775 17003 11781
rect 14384 11744 14412 11772
rect 17494 11744 17500 11756
rect 14384 11716 14780 11744
rect 14752 11688 14780 11716
rect 15672 11716 17500 11744
rect 14366 11636 14372 11688
rect 14424 11676 14430 11688
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 14424 11648 14657 11676
rect 14424 11636 14430 11648
rect 14645 11645 14657 11648
rect 14691 11645 14703 11679
rect 14645 11639 14703 11645
rect 14734 11636 14740 11688
rect 14792 11676 14798 11688
rect 14901 11679 14959 11685
rect 14901 11676 14913 11679
rect 14792 11648 14913 11676
rect 14792 11636 14798 11648
rect 14901 11645 14913 11648
rect 14947 11645 14959 11679
rect 14901 11639 14959 11645
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15672 11676 15700 11716
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 17589 11747 17647 11753
rect 17589 11713 17601 11747
rect 17635 11744 17647 11747
rect 17773 11747 17831 11753
rect 17773 11744 17785 11747
rect 17635 11716 17785 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 17773 11713 17785 11716
rect 17819 11713 17831 11747
rect 17773 11707 17831 11713
rect 15344 11648 15700 11676
rect 15344 11636 15350 11648
rect 16022 11636 16028 11688
rect 16080 11676 16086 11688
rect 16301 11679 16359 11685
rect 16301 11676 16313 11679
rect 16080 11648 16313 11676
rect 16080 11636 16086 11648
rect 16301 11645 16313 11648
rect 16347 11645 16359 11679
rect 17310 11676 17316 11688
rect 17271 11648 17316 11676
rect 16301 11639 16359 11645
rect 17310 11636 17316 11648
rect 17368 11636 17374 11688
rect 18064 11685 18092 11784
rect 18138 11704 18144 11756
rect 18196 11744 18202 11756
rect 18233 11747 18291 11753
rect 18233 11744 18245 11747
rect 18196 11716 18245 11744
rect 18196 11704 18202 11716
rect 18233 11713 18245 11716
rect 18279 11713 18291 11747
rect 18233 11707 18291 11713
rect 18322 11704 18328 11756
rect 18380 11744 18386 11756
rect 20180 11744 20208 11840
rect 21085 11747 21143 11753
rect 21085 11744 21097 11747
rect 18380 11716 18920 11744
rect 20180 11716 21097 11744
rect 18380 11704 18386 11716
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 18414 11636 18420 11688
rect 18472 11676 18478 11688
rect 18785 11679 18843 11685
rect 18785 11676 18797 11679
rect 18472 11648 18797 11676
rect 18472 11636 18478 11648
rect 18785 11645 18797 11648
rect 18831 11645 18843 11679
rect 18892 11676 18920 11716
rect 21085 11713 21097 11716
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 20806 11676 20812 11688
rect 18892 11648 20812 11676
rect 18785 11639 18843 11645
rect 20806 11636 20812 11648
rect 20864 11636 20870 11688
rect 17773 11611 17831 11617
rect 17773 11577 17785 11611
rect 17819 11608 17831 11611
rect 18966 11608 18972 11620
rect 17819 11580 18972 11608
rect 17819 11577 17831 11580
rect 17773 11571 17831 11577
rect 18966 11568 18972 11580
rect 19024 11617 19030 11620
rect 19024 11611 19088 11617
rect 19024 11577 19042 11611
rect 19076 11577 19088 11611
rect 19024 11571 19088 11577
rect 19024 11568 19030 11571
rect 20622 11568 20628 11620
rect 20680 11608 20686 11620
rect 20993 11611 21051 11617
rect 20993 11608 21005 11611
rect 20680 11580 21005 11608
rect 20680 11568 20686 11580
rect 20993 11577 21005 11580
rect 21039 11577 21051 11611
rect 20993 11571 21051 11577
rect 12400 11512 14320 11540
rect 12400 11500 12406 11512
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 15562 11540 15568 11552
rect 15252 11512 15568 11540
rect 15252 11500 15258 11512
rect 15562 11500 15568 11512
rect 15620 11540 15626 11552
rect 16025 11543 16083 11549
rect 16025 11540 16037 11543
rect 15620 11512 16037 11540
rect 15620 11500 15626 11512
rect 16025 11509 16037 11512
rect 16071 11509 16083 11543
rect 16025 11503 16083 11509
rect 17405 11543 17463 11549
rect 17405 11509 17417 11543
rect 17451 11540 17463 11543
rect 19242 11540 19248 11552
rect 17451 11512 19248 11540
rect 17451 11509 17463 11512
rect 17405 11503 17463 11509
rect 19242 11500 19248 11512
rect 19300 11500 19306 11552
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 20901 11543 20959 11549
rect 20901 11540 20913 11543
rect 20864 11512 20913 11540
rect 20864 11500 20870 11512
rect 20901 11509 20913 11512
rect 20947 11509 20959 11543
rect 20901 11503 20959 11509
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 7558 11296 7564 11348
rect 7616 11336 7622 11348
rect 8849 11339 8907 11345
rect 8849 11336 8861 11339
rect 7616 11308 8861 11336
rect 7616 11296 7622 11308
rect 8849 11305 8861 11308
rect 8895 11305 8907 11339
rect 9674 11336 9680 11348
rect 9635 11308 9680 11336
rect 8849 11299 8907 11305
rect 8864 11200 8892 11299
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10134 11336 10140 11348
rect 10095 11308 10140 11336
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11241 11339 11299 11345
rect 11241 11305 11253 11339
rect 11287 11336 11299 11339
rect 12986 11336 12992 11348
rect 11287 11308 12992 11336
rect 11287 11305 11299 11308
rect 11241 11299 11299 11305
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 13078 11296 13084 11348
rect 13136 11336 13142 11348
rect 14461 11339 14519 11345
rect 14461 11336 14473 11339
rect 13136 11308 14473 11336
rect 13136 11296 13142 11308
rect 14461 11305 14473 11308
rect 14507 11305 14519 11339
rect 14461 11299 14519 11305
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 15378 11336 15384 11348
rect 15335 11308 15384 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 18598 11336 18604 11348
rect 15528 11308 18604 11336
rect 15528 11296 15534 11308
rect 18598 11296 18604 11308
rect 18656 11296 18662 11348
rect 18966 11336 18972 11348
rect 18927 11308 18972 11336
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 19242 11336 19248 11348
rect 19203 11308 19248 11336
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 19610 11336 19616 11348
rect 19571 11308 19616 11336
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 20714 11296 20720 11348
rect 20772 11336 20778 11348
rect 20901 11339 20959 11345
rect 20901 11336 20913 11339
rect 20772 11308 20913 11336
rect 20772 11296 20778 11308
rect 20901 11305 20913 11308
rect 20947 11305 20959 11339
rect 20901 11299 20959 11305
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 10045 11271 10103 11277
rect 10045 11268 10057 11271
rect 9180 11240 10057 11268
rect 9180 11228 9186 11240
rect 10045 11237 10057 11240
rect 10091 11237 10103 11271
rect 10045 11231 10103 11237
rect 11054 11228 11060 11280
rect 11112 11268 11118 11280
rect 16178 11271 16236 11277
rect 16178 11268 16190 11271
rect 11112 11240 16190 11268
rect 11112 11228 11118 11240
rect 16178 11237 16190 11240
rect 16224 11268 16236 11271
rect 16666 11268 16672 11280
rect 16224 11240 16672 11268
rect 16224 11237 16236 11240
rect 16178 11231 16236 11237
rect 16666 11228 16672 11240
rect 16724 11228 16730 11280
rect 19058 11268 19064 11280
rect 16776 11240 19064 11268
rect 11517 11203 11575 11209
rect 8864 11172 11100 11200
rect 11072 11144 11100 11172
rect 11517 11169 11529 11203
rect 11563 11200 11575 11203
rect 11606 11200 11612 11212
rect 11563 11172 11612 11200
rect 11563 11169 11575 11172
rect 11517 11163 11575 11169
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 11784 11203 11842 11209
rect 11784 11169 11796 11203
rect 11830 11200 11842 11203
rect 12066 11200 12072 11212
rect 11830 11172 12072 11200
rect 11830 11169 11842 11172
rect 11784 11163 11842 11169
rect 12066 11160 12072 11172
rect 12124 11160 12130 11212
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 10318 11132 10324 11144
rect 10279 11104 10324 11132
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 11054 11092 11060 11144
rect 11112 11092 11118 11144
rect 13188 11132 13216 11163
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 16776 11200 16804 11240
rect 19058 11228 19064 11240
rect 19116 11228 19122 11280
rect 14700 11172 16804 11200
rect 17856 11203 17914 11209
rect 14700 11160 14706 11172
rect 17856 11169 17868 11203
rect 17902 11200 17914 11203
rect 18690 11200 18696 11212
rect 17902 11172 18696 11200
rect 17902 11169 17914 11172
rect 17856 11163 17914 11169
rect 18690 11160 18696 11172
rect 18748 11200 18754 11212
rect 18748 11172 19932 11200
rect 18748 11160 18754 11172
rect 15470 11132 15476 11144
rect 13188 11104 15476 11132
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11101 15991 11135
rect 15933 11095 15991 11101
rect 10686 11064 10692 11076
rect 10647 11036 10692 11064
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 12897 11067 12955 11073
rect 12897 11033 12909 11067
rect 12943 11064 12955 11067
rect 13814 11064 13820 11076
rect 12943 11036 13820 11064
rect 12943 11033 12955 11036
rect 12897 11027 12955 11033
rect 13814 11024 13820 11036
rect 13872 11064 13878 11076
rect 14366 11064 14372 11076
rect 13872 11036 14372 11064
rect 13872 11024 13878 11036
rect 14366 11024 14372 11036
rect 14424 11024 14430 11076
rect 14458 11024 14464 11076
rect 14516 11064 14522 11076
rect 15948 11064 15976 11095
rect 17494 11092 17500 11144
rect 17552 11132 17558 11144
rect 17589 11135 17647 11141
rect 17589 11132 17601 11135
rect 17552 11104 17601 11132
rect 17552 11092 17558 11104
rect 17589 11101 17601 11104
rect 17635 11101 17647 11135
rect 17589 11095 17647 11101
rect 17604 11064 17632 11095
rect 18598 11092 18604 11144
rect 18656 11132 18662 11144
rect 19334 11132 19340 11144
rect 18656 11104 19340 11132
rect 18656 11092 18662 11104
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 19702 11132 19708 11144
rect 19663 11104 19708 11132
rect 19702 11092 19708 11104
rect 19760 11092 19766 11144
rect 19904 11141 19932 11172
rect 19889 11135 19947 11141
rect 19889 11101 19901 11135
rect 19935 11132 19947 11135
rect 20714 11132 20720 11144
rect 19935 11104 20720 11132
rect 19935 11101 19947 11104
rect 19889 11095 19947 11101
rect 20714 11092 20720 11104
rect 20772 11092 20778 11144
rect 14516 11036 15976 11064
rect 14516 11024 14522 11036
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 9217 10999 9275 11005
rect 9217 10996 9229 10999
rect 8536 10968 9229 10996
rect 8536 10956 8542 10968
rect 9217 10965 9229 10968
rect 9263 10965 9275 10999
rect 9217 10959 9275 10965
rect 10502 10956 10508 11008
rect 10560 10996 10566 11008
rect 13998 10996 14004 11008
rect 10560 10968 14004 10996
rect 10560 10956 10566 10968
rect 13998 10956 14004 10968
rect 14056 10956 14062 11008
rect 15948 10996 15976 11036
rect 16868 11036 17632 11064
rect 20533 11067 20591 11073
rect 16868 10996 16896 11036
rect 20533 11033 20545 11067
rect 20579 11064 20591 11067
rect 20622 11064 20628 11076
rect 20579 11036 20628 11064
rect 20579 11033 20591 11036
rect 20533 11027 20591 11033
rect 20622 11024 20628 11036
rect 20680 11024 20686 11076
rect 15948 10968 16896 10996
rect 17313 10999 17371 11005
rect 17313 10965 17325 10999
rect 17359 10996 17371 10999
rect 17770 10996 17776 11008
rect 17359 10968 17776 10996
rect 17359 10965 17371 10968
rect 17313 10959 17371 10965
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 8757 10795 8815 10801
rect 8757 10761 8769 10795
rect 8803 10792 8815 10795
rect 10502 10792 10508 10804
rect 8803 10764 10508 10792
rect 8803 10761 8815 10764
rect 8757 10755 8815 10761
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 10781 10795 10839 10801
rect 10781 10761 10793 10795
rect 10827 10792 10839 10795
rect 11882 10792 11888 10804
rect 10827 10764 11888 10792
rect 10827 10761 10839 10764
rect 10781 10755 10839 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 14550 10752 14556 10804
rect 14608 10792 14614 10804
rect 14737 10795 14795 10801
rect 14737 10792 14749 10795
rect 14608 10764 14749 10792
rect 14608 10752 14614 10764
rect 14737 10761 14749 10764
rect 14783 10761 14795 10795
rect 14737 10755 14795 10761
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 17862 10792 17868 10804
rect 16172 10764 17868 10792
rect 16172 10752 16178 10764
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 20714 10792 20720 10804
rect 20675 10764 20720 10792
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 9769 10727 9827 10733
rect 9769 10693 9781 10727
rect 9815 10693 9827 10727
rect 9769 10687 9827 10693
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10588 9091 10591
rect 9784 10588 9812 10687
rect 9950 10684 9956 10736
rect 10008 10724 10014 10736
rect 12802 10724 12808 10736
rect 10008 10696 12808 10724
rect 10008 10684 10014 10696
rect 12802 10684 12808 10696
rect 12860 10724 12866 10736
rect 12860 10696 13216 10724
rect 12860 10684 12866 10696
rect 10410 10656 10416 10668
rect 10371 10628 10416 10656
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 13188 10665 13216 10696
rect 14642 10684 14648 10736
rect 14700 10724 14706 10736
rect 15749 10727 15807 10733
rect 15749 10724 15761 10727
rect 14700 10696 15761 10724
rect 14700 10684 14706 10696
rect 15749 10693 15761 10696
rect 15795 10693 15807 10727
rect 15749 10687 15807 10693
rect 11333 10659 11391 10665
rect 11333 10656 11345 10659
rect 11296 10628 11345 10656
rect 11296 10616 11302 10628
rect 11333 10625 11345 10628
rect 11379 10625 11391 10659
rect 11333 10619 11391 10625
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 13357 10659 13415 10665
rect 13357 10625 13369 10659
rect 13403 10625 13415 10659
rect 13357 10619 13415 10625
rect 11974 10588 11980 10600
rect 9079 10560 9812 10588
rect 10060 10560 11980 10588
rect 9079 10557 9091 10560
rect 9033 10551 9091 10557
rect 9309 10523 9367 10529
rect 9309 10489 9321 10523
rect 9355 10520 9367 10523
rect 10060 10520 10088 10560
rect 11974 10548 11980 10560
rect 12032 10548 12038 10600
rect 12986 10548 12992 10600
rect 13044 10588 13050 10600
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 13044 10560 13093 10588
rect 13044 10548 13050 10560
rect 13081 10557 13093 10560
rect 13127 10557 13139 10591
rect 13372 10588 13400 10619
rect 13538 10616 13544 10668
rect 13596 10656 13602 10668
rect 14277 10659 14335 10665
rect 14277 10656 14289 10659
rect 13596 10628 14289 10656
rect 13596 10616 13602 10628
rect 14277 10625 14289 10628
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 14366 10616 14372 10668
rect 14424 10656 14430 10668
rect 15289 10659 15347 10665
rect 15289 10656 15301 10659
rect 14424 10628 15301 10656
rect 14424 10616 14430 10628
rect 15289 10625 15301 10628
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 17589 10659 17647 10665
rect 17589 10625 17601 10659
rect 17635 10656 17647 10659
rect 18046 10656 18052 10668
rect 17635 10628 18052 10656
rect 17635 10625 17647 10628
rect 17589 10619 17647 10625
rect 13722 10588 13728 10600
rect 13372 10560 13728 10588
rect 13081 10551 13139 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 13906 10548 13912 10600
rect 13964 10588 13970 10600
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 13964 10560 14197 10588
rect 13964 10548 13970 10560
rect 14185 10557 14197 10560
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 14734 10548 14740 10600
rect 14792 10588 14798 10600
rect 15838 10588 15844 10600
rect 14792 10560 15844 10588
rect 14792 10548 14798 10560
rect 15838 10548 15844 10560
rect 15896 10588 15902 10600
rect 16316 10588 16344 10619
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18690 10656 18696 10668
rect 18651 10628 18696 10656
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 19334 10656 19340 10668
rect 19295 10628 19340 10656
rect 19334 10616 19340 10628
rect 19392 10616 19398 10668
rect 15896 10560 16344 10588
rect 15896 10548 15902 10560
rect 9355 10492 10088 10520
rect 10137 10523 10195 10529
rect 9355 10489 9367 10492
rect 9309 10483 9367 10489
rect 10137 10489 10149 10523
rect 10183 10520 10195 10523
rect 10870 10520 10876 10532
rect 10183 10492 10876 10520
rect 10183 10489 10195 10492
rect 10137 10483 10195 10489
rect 10870 10480 10876 10492
rect 10928 10480 10934 10532
rect 11054 10480 11060 10532
rect 11112 10520 11118 10532
rect 11238 10520 11244 10532
rect 11112 10492 11244 10520
rect 11112 10480 11118 10492
rect 11238 10480 11244 10492
rect 11296 10480 11302 10532
rect 12069 10523 12127 10529
rect 12069 10489 12081 10523
rect 12115 10520 12127 10523
rect 13446 10520 13452 10532
rect 12115 10492 13452 10520
rect 12115 10489 12127 10492
rect 12069 10483 12127 10489
rect 13446 10480 13452 10492
rect 13504 10480 13510 10532
rect 15197 10523 15255 10529
rect 15197 10520 15209 10523
rect 13740 10492 15209 10520
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 10284 10424 10329 10452
rect 10284 10412 10290 10424
rect 10686 10412 10692 10464
rect 10744 10452 10750 10464
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 10744 10424 11161 10452
rect 10744 10412 10750 10424
rect 11149 10421 11161 10424
rect 11195 10421 11207 10455
rect 11149 10415 11207 10421
rect 11882 10412 11888 10464
rect 11940 10452 11946 10464
rect 13740 10461 13768 10492
rect 15197 10489 15209 10492
rect 15243 10489 15255 10523
rect 15197 10483 15255 10489
rect 16022 10480 16028 10532
rect 16080 10520 16086 10532
rect 19610 10529 19616 10532
rect 16209 10523 16267 10529
rect 16209 10520 16221 10523
rect 16080 10492 16221 10520
rect 16080 10480 16086 10492
rect 16209 10489 16221 10492
rect 16255 10489 16267 10523
rect 16209 10483 16267 10489
rect 17313 10523 17371 10529
rect 17313 10489 17325 10523
rect 17359 10520 17371 10523
rect 17359 10492 18092 10520
rect 17359 10489 17371 10492
rect 17313 10483 17371 10489
rect 12713 10455 12771 10461
rect 12713 10452 12725 10455
rect 11940 10424 12725 10452
rect 11940 10412 11946 10424
rect 12713 10421 12725 10424
rect 12759 10421 12771 10455
rect 12713 10415 12771 10421
rect 13725 10455 13783 10461
rect 13725 10421 13737 10455
rect 13771 10421 13783 10455
rect 13725 10415 13783 10421
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 14093 10455 14151 10461
rect 14093 10452 14105 10455
rect 13872 10424 14105 10452
rect 13872 10412 13878 10424
rect 14093 10421 14105 10424
rect 14139 10421 14151 10455
rect 14093 10415 14151 10421
rect 14366 10412 14372 10464
rect 14424 10452 14430 10464
rect 15105 10455 15163 10461
rect 15105 10452 15117 10455
rect 14424 10424 15117 10452
rect 14424 10412 14430 10424
rect 15105 10421 15117 10424
rect 15151 10421 15163 10455
rect 16114 10452 16120 10464
rect 16075 10424 16120 10452
rect 15105 10415 15163 10421
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 16298 10412 16304 10464
rect 16356 10452 16362 10464
rect 16945 10455 17003 10461
rect 16945 10452 16957 10455
rect 16356 10424 16957 10452
rect 16356 10412 16362 10424
rect 16945 10421 16957 10424
rect 16991 10421 17003 10455
rect 17402 10452 17408 10464
rect 17363 10424 17408 10452
rect 16945 10415 17003 10421
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 18064 10461 18092 10492
rect 19604 10483 19616 10529
rect 19668 10520 19674 10532
rect 19668 10492 19704 10520
rect 19610 10480 19616 10483
rect 19668 10480 19674 10492
rect 18049 10455 18107 10461
rect 18049 10421 18061 10455
rect 18095 10421 18107 10455
rect 18049 10415 18107 10421
rect 18138 10412 18144 10464
rect 18196 10452 18202 10464
rect 18417 10455 18475 10461
rect 18417 10452 18429 10455
rect 18196 10424 18429 10452
rect 18196 10412 18202 10424
rect 18417 10421 18429 10424
rect 18463 10421 18475 10455
rect 18417 10415 18475 10421
rect 18506 10412 18512 10464
rect 18564 10452 18570 10464
rect 19518 10452 19524 10464
rect 18564 10424 19524 10452
rect 18564 10412 18570 10424
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 21269 10455 21327 10461
rect 21269 10421 21281 10455
rect 21315 10452 21327 10455
rect 21358 10452 21364 10464
rect 21315 10424 21364 10452
rect 21315 10421 21327 10424
rect 21269 10415 21327 10421
rect 21358 10412 21364 10424
rect 21416 10412 21422 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 8570 10248 8576 10260
rect 8531 10220 8576 10248
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 8662 10208 8668 10260
rect 8720 10248 8726 10260
rect 8849 10251 8907 10257
rect 8849 10248 8861 10251
rect 8720 10220 8861 10248
rect 8720 10208 8726 10220
rect 8849 10217 8861 10220
rect 8895 10248 8907 10251
rect 9122 10248 9128 10260
rect 8895 10220 9128 10248
rect 8895 10217 8907 10220
rect 8849 10211 8907 10217
rect 9122 10208 9128 10220
rect 9180 10248 9186 10260
rect 11606 10248 11612 10260
rect 9180 10220 11612 10248
rect 9180 10208 9186 10220
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 13357 10251 13415 10257
rect 13357 10248 13369 10251
rect 12032 10220 13369 10248
rect 12032 10208 12038 10220
rect 13357 10217 13369 10220
rect 13403 10248 13415 10251
rect 13538 10248 13544 10260
rect 13403 10220 13544 10248
rect 13403 10217 13415 10220
rect 13357 10211 13415 10217
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10248 13691 10251
rect 13814 10248 13820 10260
rect 13679 10220 13820 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14001 10251 14059 10257
rect 14001 10217 14013 10251
rect 14047 10248 14059 10251
rect 14458 10248 14464 10260
rect 14047 10220 14464 10248
rect 14047 10217 14059 10220
rect 14001 10211 14059 10217
rect 14458 10208 14464 10220
rect 14516 10248 14522 10260
rect 15286 10248 15292 10260
rect 14516 10220 15292 10248
rect 14516 10208 14522 10220
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 15657 10251 15715 10257
rect 15657 10217 15669 10251
rect 15703 10248 15715 10251
rect 15746 10248 15752 10260
rect 15703 10220 15752 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 17129 10251 17187 10257
rect 17129 10217 17141 10251
rect 17175 10248 17187 10251
rect 18509 10251 18567 10257
rect 18509 10248 18521 10251
rect 17175 10220 18521 10248
rect 17175 10217 17187 10220
rect 17129 10211 17187 10217
rect 18509 10217 18521 10220
rect 18555 10217 18567 10251
rect 19150 10248 19156 10260
rect 19111 10220 19156 10248
rect 18509 10211 18567 10217
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 19702 10248 19708 10260
rect 19663 10220 19708 10248
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 10410 10140 10416 10192
rect 10468 10180 10474 10192
rect 10566 10183 10624 10189
rect 10566 10180 10578 10183
rect 10468 10152 10578 10180
rect 10468 10140 10474 10152
rect 10566 10149 10578 10152
rect 10612 10149 10624 10183
rect 10566 10143 10624 10149
rect 12526 10140 12532 10192
rect 12584 10180 12590 10192
rect 17497 10183 17555 10189
rect 17497 10180 17509 10183
rect 12584 10152 17509 10180
rect 12584 10140 12590 10152
rect 17497 10149 17509 10152
rect 17543 10149 17555 10183
rect 17497 10143 17555 10149
rect 17589 10183 17647 10189
rect 17589 10149 17601 10183
rect 17635 10180 17647 10183
rect 17678 10180 17684 10192
rect 17635 10152 17684 10180
rect 17635 10149 17647 10152
rect 17589 10143 17647 10149
rect 17678 10140 17684 10152
rect 17736 10140 17742 10192
rect 20165 10183 20223 10189
rect 20165 10149 20177 10183
rect 20211 10180 20223 10183
rect 20254 10180 20260 10192
rect 20211 10152 20260 10180
rect 20211 10149 20223 10152
rect 20165 10143 20223 10149
rect 20254 10140 20260 10152
rect 20312 10140 20318 10192
rect 11698 10112 11704 10124
rect 10336 10084 11704 10112
rect 9306 10004 9312 10056
rect 9364 10044 9370 10056
rect 10336 10053 10364 10084
rect 11698 10072 11704 10084
rect 11756 10112 11762 10124
rect 11977 10115 12035 10121
rect 11977 10112 11989 10115
rect 11756 10084 11989 10112
rect 11756 10072 11762 10084
rect 11977 10081 11989 10084
rect 12023 10081 12035 10115
rect 12244 10115 12302 10121
rect 12244 10112 12256 10115
rect 11977 10075 12035 10081
rect 12084 10084 12256 10112
rect 10321 10047 10379 10053
rect 10321 10044 10333 10047
rect 9364 10016 10333 10044
rect 9364 10004 9370 10016
rect 10321 10013 10333 10016
rect 10367 10013 10379 10047
rect 12084 10044 12112 10084
rect 12244 10081 12256 10084
rect 12290 10112 12302 10115
rect 12290 10084 13032 10112
rect 12290 10081 12302 10084
rect 12244 10075 12302 10081
rect 10321 10007 10379 10013
rect 11716 10016 12112 10044
rect 6914 9936 6920 9988
rect 6972 9976 6978 9988
rect 9217 9979 9275 9985
rect 9217 9976 9229 9979
rect 6972 9948 9229 9976
rect 6972 9936 6978 9948
rect 9217 9945 9229 9948
rect 9263 9976 9275 9979
rect 9950 9976 9956 9988
rect 9263 9948 9956 9976
rect 9263 9945 9275 9948
rect 9217 9939 9275 9945
rect 9950 9936 9956 9948
rect 10008 9936 10014 9988
rect 11716 9985 11744 10016
rect 11701 9979 11759 9985
rect 11701 9945 11713 9979
rect 11747 9945 11759 9979
rect 13004 9976 13032 10084
rect 13538 10072 13544 10124
rect 13596 10112 13602 10124
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 13596 10084 15761 10112
rect 13596 10072 13602 10084
rect 15749 10081 15761 10084
rect 15795 10081 15807 10115
rect 16298 10112 16304 10124
rect 16259 10084 16304 10112
rect 15749 10075 15807 10081
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 16577 10115 16635 10121
rect 16577 10081 16589 10115
rect 16623 10112 16635 10115
rect 17218 10112 17224 10124
rect 16623 10084 17224 10112
rect 16623 10081 16635 10084
rect 16577 10075 16635 10081
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 20073 10115 20131 10121
rect 20073 10081 20085 10115
rect 20119 10112 20131 10115
rect 21358 10112 21364 10124
rect 20119 10084 21364 10112
rect 20119 10081 20131 10084
rect 20073 10075 20131 10081
rect 21358 10072 21364 10084
rect 21416 10072 21422 10124
rect 14090 10004 14096 10056
rect 14148 10044 14154 10056
rect 14277 10047 14335 10053
rect 14148 10016 14193 10044
rect 14148 10004 14154 10016
rect 14277 10013 14289 10047
rect 14323 10013 14335 10047
rect 14734 10044 14740 10056
rect 14695 10016 14740 10044
rect 14277 10007 14335 10013
rect 13722 9976 13728 9988
rect 13004 9948 13728 9976
rect 11701 9939 11759 9945
rect 13722 9936 13728 9948
rect 13780 9976 13786 9988
rect 14292 9976 14320 10007
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 15838 10004 15844 10056
rect 15896 10044 15902 10056
rect 17770 10044 17776 10056
rect 15896 10016 15941 10044
rect 17731 10016 17776 10044
rect 15896 10004 15902 10016
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 18598 10044 18604 10056
rect 18559 10016 18604 10044
rect 18598 10004 18604 10016
rect 18656 10004 18662 10056
rect 18690 10004 18696 10056
rect 18748 10044 18754 10056
rect 20257 10047 20315 10053
rect 18748 10016 18793 10044
rect 18748 10004 18754 10016
rect 20257 10013 20269 10047
rect 20303 10013 20315 10047
rect 20257 10007 20315 10013
rect 13780 9948 14320 9976
rect 13780 9936 13786 9948
rect 17402 9936 17408 9988
rect 17460 9976 17466 9988
rect 18141 9979 18199 9985
rect 18141 9976 18153 9979
rect 17460 9948 18153 9976
rect 17460 9936 17466 9948
rect 18141 9945 18153 9948
rect 18187 9945 18199 9979
rect 18141 9939 18199 9945
rect 19610 9936 19616 9988
rect 19668 9976 19674 9988
rect 20272 9976 20300 10007
rect 21358 9976 21364 9988
rect 19668 9948 20300 9976
rect 21319 9948 21364 9976
rect 19668 9936 19674 9948
rect 21358 9936 21364 9948
rect 21416 9936 21422 9988
rect 10042 9908 10048 9920
rect 10003 9880 10048 9908
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 12894 9868 12900 9920
rect 12952 9908 12958 9920
rect 14182 9908 14188 9920
rect 12952 9880 14188 9908
rect 12952 9868 12958 9880
rect 14182 9868 14188 9880
rect 14240 9908 14246 9920
rect 14458 9908 14464 9920
rect 14240 9880 14464 9908
rect 14240 9868 14246 9880
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 15289 9911 15347 9917
rect 15289 9908 15301 9911
rect 14792 9880 15301 9908
rect 14792 9868 14798 9880
rect 15289 9877 15301 9880
rect 15335 9877 15347 9911
rect 15289 9871 15347 9877
rect 17494 9868 17500 9920
rect 17552 9908 17558 9920
rect 18966 9908 18972 9920
rect 17552 9880 18972 9908
rect 17552 9868 17558 9880
rect 18966 9868 18972 9880
rect 19024 9868 19030 9920
rect 20990 9908 20996 9920
rect 20951 9880 20996 9908
rect 20990 9868 20996 9880
rect 21048 9868 21054 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 8570 9704 8576 9716
rect 8531 9676 8576 9704
rect 8570 9664 8576 9676
rect 8628 9664 8634 9716
rect 9232 9676 10180 9704
rect 8757 9639 8815 9645
rect 8757 9605 8769 9639
rect 8803 9636 8815 9639
rect 9232 9636 9260 9676
rect 8803 9608 9260 9636
rect 10152 9636 10180 9676
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 10597 9707 10655 9713
rect 10597 9704 10609 9707
rect 10468 9676 10609 9704
rect 10468 9664 10474 9676
rect 10597 9673 10609 9676
rect 10643 9673 10655 9707
rect 10870 9704 10876 9716
rect 10831 9676 10876 9704
rect 10597 9667 10655 9673
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 11885 9707 11943 9713
rect 11885 9704 11897 9707
rect 11756 9676 11897 9704
rect 11756 9664 11762 9676
rect 11885 9673 11897 9676
rect 11931 9673 11943 9707
rect 11885 9667 11943 9673
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 14366 9704 14372 9716
rect 12584 9676 14372 9704
rect 12584 9664 12590 9676
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 18690 9704 18696 9716
rect 18064 9676 18696 9704
rect 12437 9639 12495 9645
rect 10152 9608 11560 9636
rect 8803 9605 8815 9608
rect 8757 9599 8815 9605
rect 11348 9577 11376 9608
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9537 11391 9571
rect 11333 9531 11391 9537
rect 11425 9571 11483 9577
rect 11425 9537 11437 9571
rect 11471 9537 11483 9571
rect 11532 9568 11560 9608
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 12894 9636 12900 9648
rect 12483 9608 12900 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 13265 9639 13323 9645
rect 13265 9605 13277 9639
rect 13311 9636 13323 9639
rect 13906 9636 13912 9648
rect 13311 9608 13912 9636
rect 13311 9605 13323 9608
rect 13265 9599 13323 9605
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 14090 9596 14096 9648
rect 14148 9636 14154 9648
rect 14277 9639 14335 9645
rect 14277 9636 14289 9639
rect 14148 9608 14289 9636
rect 14148 9596 14154 9608
rect 14277 9605 14289 9608
rect 14323 9636 14335 9639
rect 14550 9636 14556 9648
rect 14323 9608 14556 9636
rect 14323 9605 14335 9608
rect 14277 9599 14335 9605
rect 14550 9596 14556 9608
rect 14608 9636 14614 9648
rect 17681 9639 17739 9645
rect 14608 9608 16252 9636
rect 14608 9596 14614 9608
rect 12710 9568 12716 9580
rect 11532 9540 12716 9568
rect 11425 9531 11483 9537
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9306 9500 9312 9512
rect 9263 9472 9312 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 9484 9503 9542 9509
rect 9484 9469 9496 9503
rect 9530 9500 9542 9503
rect 10962 9500 10968 9512
rect 9530 9472 10968 9500
rect 9530 9469 9542 9472
rect 9484 9463 9542 9469
rect 10962 9460 10968 9472
rect 11020 9500 11026 9512
rect 11440 9500 11468 9531
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 12912 9540 13676 9568
rect 12066 9500 12072 9512
rect 11020 9472 11468 9500
rect 12027 9472 12072 9500
rect 11020 9460 11026 9472
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 12912 9500 12940 9540
rect 12268 9472 12940 9500
rect 12989 9503 13047 9509
rect 3418 9392 3424 9444
rect 3476 9432 3482 9444
rect 3476 9404 8984 9432
rect 3476 9392 3482 9404
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 7800 9336 8769 9364
rect 7800 9324 7806 9336
rect 8757 9333 8769 9336
rect 8803 9364 8815 9367
rect 8849 9367 8907 9373
rect 8849 9364 8861 9367
rect 8803 9336 8861 9364
rect 8803 9333 8815 9336
rect 8757 9327 8815 9333
rect 8849 9333 8861 9336
rect 8895 9333 8907 9367
rect 8956 9364 8984 9404
rect 9950 9392 9956 9444
rect 10008 9432 10014 9444
rect 11241 9435 11299 9441
rect 11241 9432 11253 9435
rect 10008 9404 11253 9432
rect 10008 9392 10014 9404
rect 11241 9401 11253 9404
rect 11287 9401 11299 9435
rect 11241 9395 11299 9401
rect 12268 9364 12296 9472
rect 12989 9469 13001 9503
rect 13035 9500 13047 9503
rect 13078 9500 13084 9512
rect 13035 9472 13084 9500
rect 13035 9469 13047 9472
rect 12989 9463 13047 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 13648 9500 13676 9540
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 13817 9571 13875 9577
rect 13817 9568 13829 9571
rect 13780 9540 13829 9568
rect 13780 9528 13786 9540
rect 13817 9537 13829 9540
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 14458 9528 14464 9580
rect 14516 9568 14522 9580
rect 15197 9571 15255 9577
rect 15197 9568 15209 9571
rect 14516 9540 15209 9568
rect 14516 9528 14522 9540
rect 15197 9537 15209 9540
rect 15243 9537 15255 9571
rect 15197 9531 15255 9537
rect 16224 9500 16252 9608
rect 17681 9605 17693 9639
rect 17727 9636 17739 9639
rect 17954 9636 17960 9648
rect 17727 9608 17960 9636
rect 17727 9605 17739 9608
rect 17681 9599 17739 9605
rect 17954 9596 17960 9608
rect 18012 9636 18018 9648
rect 18064 9636 18092 9676
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 19610 9664 19616 9716
rect 19668 9704 19674 9716
rect 19705 9707 19763 9713
rect 19705 9704 19717 9707
rect 19668 9676 19717 9704
rect 19668 9664 19674 9676
rect 19705 9673 19717 9676
rect 19751 9673 19763 9707
rect 19705 9667 19763 9673
rect 19886 9664 19892 9716
rect 19944 9704 19950 9716
rect 20438 9704 20444 9716
rect 19944 9676 20444 9704
rect 19944 9664 19950 9676
rect 20438 9664 20444 9676
rect 20496 9664 20502 9716
rect 18012 9608 18092 9636
rect 18012 9596 18018 9608
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9568 16359 9571
rect 16347 9540 16436 9568
rect 16347 9537 16359 9540
rect 16301 9531 16359 9537
rect 16408 9512 16436 9540
rect 17310 9528 17316 9580
rect 17368 9568 17374 9580
rect 17368 9540 18368 9568
rect 17368 9528 17374 9540
rect 13648 9472 16160 9500
rect 16224 9472 16344 9500
rect 13538 9392 13544 9444
rect 13596 9432 13602 9444
rect 13725 9435 13783 9441
rect 13725 9432 13737 9435
rect 13596 9404 13737 9432
rect 13596 9392 13602 9404
rect 13725 9401 13737 9404
rect 13771 9401 13783 9435
rect 13725 9395 13783 9401
rect 15013 9435 15071 9441
rect 15013 9401 15025 9435
rect 15059 9432 15071 9435
rect 15657 9435 15715 9441
rect 15657 9432 15669 9435
rect 15059 9404 15669 9432
rect 15059 9401 15071 9404
rect 15013 9395 15071 9401
rect 15657 9401 15669 9404
rect 15703 9401 15715 9435
rect 16132 9432 16160 9472
rect 16316 9432 16344 9472
rect 16390 9460 16396 9512
rect 16448 9460 16454 9512
rect 16568 9503 16626 9509
rect 16568 9469 16580 9503
rect 16614 9500 16626 9503
rect 17770 9500 17776 9512
rect 16614 9472 17776 9500
rect 16614 9469 16626 9472
rect 16568 9463 16626 9469
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 18230 9500 18236 9512
rect 17880 9472 18236 9500
rect 17880 9432 17908 9472
rect 18230 9460 18236 9472
rect 18288 9460 18294 9512
rect 18340 9509 18368 9540
rect 20438 9528 20444 9580
rect 20496 9568 20502 9580
rect 20901 9571 20959 9577
rect 20901 9568 20913 9571
rect 20496 9540 20913 9568
rect 20496 9528 20502 9540
rect 20901 9537 20913 9540
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 18325 9503 18383 9509
rect 18325 9469 18337 9503
rect 18371 9500 18383 9503
rect 19334 9500 19340 9512
rect 18371 9472 19340 9500
rect 18371 9469 18383 9472
rect 18325 9463 18383 9469
rect 19334 9460 19340 9472
rect 19392 9460 19398 9512
rect 20809 9503 20867 9509
rect 20809 9469 20821 9503
rect 20855 9500 20867 9503
rect 21358 9500 21364 9512
rect 20855 9472 21364 9500
rect 20855 9469 20867 9472
rect 20809 9463 20867 9469
rect 21358 9460 21364 9472
rect 21416 9460 21422 9512
rect 16132 9404 16252 9432
rect 16316 9404 17908 9432
rect 15657 9395 15715 9401
rect 12802 9364 12808 9376
rect 8956 9336 12296 9364
rect 12763 9336 12808 9364
rect 8849 9327 8907 9333
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 13633 9367 13691 9373
rect 13633 9364 13645 9367
rect 13504 9336 13645 9364
rect 13504 9324 13510 9336
rect 13633 9333 13645 9336
rect 13679 9333 13691 9367
rect 14642 9364 14648 9376
rect 14603 9336 14648 9364
rect 13633 9327 13691 9333
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 15105 9367 15163 9373
rect 15105 9333 15117 9367
rect 15151 9364 15163 9367
rect 16114 9364 16120 9376
rect 15151 9336 16120 9364
rect 15151 9333 15163 9336
rect 15105 9327 15163 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16224 9364 16252 9404
rect 18046 9392 18052 9444
rect 18104 9432 18110 9444
rect 18506 9432 18512 9444
rect 18104 9404 18512 9432
rect 18104 9392 18110 9404
rect 18506 9392 18512 9404
rect 18564 9441 18570 9444
rect 18564 9435 18628 9441
rect 18564 9401 18582 9435
rect 18616 9401 18628 9435
rect 18564 9395 18628 9401
rect 18564 9392 18570 9395
rect 19242 9364 19248 9376
rect 16224 9336 19248 9364
rect 19242 9324 19248 9336
rect 19300 9364 19306 9376
rect 19981 9367 20039 9373
rect 19981 9364 19993 9367
rect 19300 9336 19993 9364
rect 19300 9324 19306 9336
rect 19981 9333 19993 9336
rect 20027 9333 20039 9367
rect 20346 9364 20352 9376
rect 20307 9336 20352 9364
rect 19981 9327 20039 9333
rect 20346 9324 20352 9336
rect 20404 9324 20410 9376
rect 20714 9364 20720 9376
rect 20675 9336 20720 9364
rect 20714 9324 20720 9336
rect 20772 9324 20778 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 9950 9160 9956 9172
rect 9911 9132 9956 9160
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 10226 9120 10232 9172
rect 10284 9160 10290 9172
rect 10413 9163 10471 9169
rect 10413 9160 10425 9163
rect 10284 9132 10425 9160
rect 10284 9120 10290 9132
rect 10413 9129 10425 9132
rect 10459 9129 10471 9163
rect 10413 9123 10471 9129
rect 10502 9120 10508 9172
rect 10560 9160 10566 9172
rect 10778 9160 10784 9172
rect 10560 9132 10784 9160
rect 10560 9120 10566 9132
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 11882 9160 11888 9172
rect 11843 9132 11888 9160
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 13357 9163 13415 9169
rect 13357 9129 13369 9163
rect 13403 9160 13415 9163
rect 13909 9163 13967 9169
rect 13909 9160 13921 9163
rect 13403 9132 13921 9160
rect 13403 9129 13415 9132
rect 13357 9123 13415 9129
rect 13909 9129 13921 9132
rect 13955 9129 13967 9163
rect 13909 9123 13967 9129
rect 14277 9163 14335 9169
rect 14277 9129 14289 9163
rect 14323 9160 14335 9163
rect 15289 9163 15347 9169
rect 15289 9160 15301 9163
rect 14323 9132 15301 9160
rect 14323 9129 14335 9132
rect 14277 9123 14335 9129
rect 15289 9129 15301 9132
rect 15335 9129 15347 9163
rect 15289 9123 15347 9129
rect 16390 9120 16396 9172
rect 16448 9160 16454 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 16448 9132 16681 9160
rect 16448 9120 16454 9132
rect 16669 9129 16681 9132
rect 16715 9160 16727 9163
rect 17310 9160 17316 9172
rect 16715 9132 17316 9160
rect 16715 9129 16727 9132
rect 16669 9123 16727 9129
rect 9309 9095 9367 9101
rect 9309 9061 9321 9095
rect 9355 9092 9367 9095
rect 10042 9092 10048 9104
rect 9355 9064 10048 9092
rect 9355 9061 9367 9064
rect 9309 9055 9367 9061
rect 10042 9052 10048 9064
rect 10100 9092 10106 9104
rect 11606 9092 11612 9104
rect 10100 9064 11612 9092
rect 10100 9052 10106 9064
rect 11606 9052 11612 9064
rect 11664 9052 11670 9104
rect 11793 9095 11851 9101
rect 11793 9061 11805 9095
rect 11839 9092 11851 9095
rect 13170 9092 13176 9104
rect 11839 9064 13176 9092
rect 11839 9061 11851 9064
rect 11793 9055 11851 9061
rect 13170 9052 13176 9064
rect 13228 9052 13234 9104
rect 13265 9095 13323 9101
rect 13265 9061 13277 9095
rect 13311 9092 13323 9095
rect 14642 9092 14648 9104
rect 13311 9064 14648 9092
rect 13311 9061 13323 9064
rect 13265 9055 13323 9061
rect 14642 9052 14648 9064
rect 14700 9052 14706 9104
rect 16758 9052 16764 9104
rect 16816 9092 16822 9104
rect 16816 9064 16896 9092
rect 16816 9052 16822 9064
rect 8941 9027 8999 9033
rect 8941 8993 8953 9027
rect 8987 9024 8999 9027
rect 10134 9024 10140 9036
rect 8987 8996 10140 9024
rect 8987 8993 8999 8996
rect 8941 8987 8999 8993
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10226 8984 10232 9036
rect 10284 9024 10290 9036
rect 10781 9027 10839 9033
rect 10781 9024 10793 9027
rect 10284 8996 10793 9024
rect 10284 8984 10290 8996
rect 10781 8993 10793 8996
rect 10827 8993 10839 9027
rect 10781 8987 10839 8993
rect 10873 9027 10931 9033
rect 10873 8993 10885 9027
rect 10919 9024 10931 9027
rect 11054 9024 11060 9036
rect 10919 8996 11060 9024
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 12621 9027 12679 9033
rect 12621 8993 12633 9027
rect 12667 9024 12679 9027
rect 12802 9024 12808 9036
rect 12667 8996 12808 9024
rect 12667 8993 12679 8996
rect 12621 8987 12679 8993
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 9024 15715 9027
rect 16022 9024 16028 9036
rect 15703 8996 16028 9024
rect 15703 8993 15715 8996
rect 15657 8987 15715 8993
rect 16022 8984 16028 8996
rect 16080 9024 16086 9036
rect 16868 9033 16896 9064
rect 17144 9033 17172 9132
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 17770 9120 17776 9172
rect 17828 9160 17834 9172
rect 18506 9160 18512 9172
rect 17828 9132 18092 9160
rect 18467 9132 18512 9160
rect 17828 9120 17834 9132
rect 17396 9095 17454 9101
rect 17396 9061 17408 9095
rect 17442 9092 17454 9095
rect 17954 9092 17960 9104
rect 17442 9064 17960 9092
rect 17442 9061 17454 9064
rect 17396 9055 17454 9061
rect 17954 9052 17960 9064
rect 18012 9052 18018 9104
rect 18064 9092 18092 9132
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 18598 9120 18604 9172
rect 18656 9160 18662 9172
rect 18785 9163 18843 9169
rect 18785 9160 18797 9163
rect 18656 9132 18797 9160
rect 18656 9120 18662 9132
rect 18785 9129 18797 9132
rect 18831 9129 18843 9163
rect 19150 9160 19156 9172
rect 19111 9132 19156 9160
rect 18785 9123 18843 9129
rect 19150 9120 19156 9132
rect 19208 9120 19214 9172
rect 20714 9120 20720 9172
rect 20772 9160 20778 9172
rect 20901 9163 20959 9169
rect 20901 9160 20913 9163
rect 20772 9132 20913 9160
rect 20772 9120 20778 9132
rect 20901 9129 20913 9132
rect 20947 9129 20959 9163
rect 20901 9123 20959 9129
rect 20165 9095 20223 9101
rect 18064 9064 19288 9092
rect 16117 9027 16175 9033
rect 16117 9024 16129 9027
rect 16080 8996 16129 9024
rect 16080 8984 16086 8996
rect 16117 8993 16129 8996
rect 16163 8993 16175 9027
rect 16117 8987 16175 8993
rect 16861 9027 16919 9033
rect 16861 8993 16873 9027
rect 16907 8993 16919 9027
rect 16861 8987 16919 8993
rect 17129 9027 17187 9033
rect 17129 8993 17141 9027
rect 17175 8993 17187 9027
rect 19260 9024 19288 9064
rect 20165 9061 20177 9095
rect 20211 9092 20223 9095
rect 20254 9092 20260 9104
rect 20211 9064 20260 9092
rect 20211 9061 20223 9064
rect 20165 9055 20223 9061
rect 19260 8996 19380 9024
rect 17129 8987 17187 8993
rect 10962 8956 10968 8968
rect 10923 8928 10968 8956
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11974 8956 11980 8968
rect 11935 8928 11980 8956
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 13541 8959 13599 8965
rect 13541 8925 13553 8959
rect 13587 8956 13599 8959
rect 13722 8956 13728 8968
rect 13587 8928 13728 8956
rect 13587 8925 13599 8928
rect 13541 8919 13599 8925
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 14366 8956 14372 8968
rect 14327 8928 14372 8956
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 14458 8916 14464 8968
rect 14516 8956 14522 8968
rect 15749 8959 15807 8965
rect 14516 8928 14561 8956
rect 14516 8916 14522 8928
rect 15749 8925 15761 8959
rect 15795 8956 15807 8959
rect 15838 8956 15844 8968
rect 15795 8928 15844 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8956 15991 8959
rect 16666 8956 16672 8968
rect 15979 8928 16672 8956
rect 15979 8925 15991 8928
rect 15933 8919 15991 8925
rect 16666 8916 16672 8928
rect 16724 8916 16730 8968
rect 18690 8916 18696 8968
rect 18748 8956 18754 8968
rect 19352 8965 19380 8996
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 18748 8928 19257 8956
rect 18748 8916 18754 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 19337 8959 19395 8965
rect 19337 8925 19349 8959
rect 19383 8925 19395 8959
rect 19337 8919 19395 8925
rect 11425 8891 11483 8897
rect 11425 8857 11437 8891
rect 11471 8888 11483 8891
rect 12526 8888 12532 8900
rect 11471 8860 12532 8888
rect 11471 8857 11483 8860
rect 11425 8851 11483 8857
rect 12526 8848 12532 8860
rect 12584 8848 12590 8900
rect 12805 8891 12863 8897
rect 12805 8857 12817 8891
rect 12851 8888 12863 8891
rect 16850 8888 16856 8900
rect 12851 8860 16856 8888
rect 12851 8857 12863 8860
rect 12805 8851 12863 8857
rect 16850 8848 16856 8860
rect 16908 8848 16914 8900
rect 18322 8848 18328 8900
rect 18380 8888 18386 8900
rect 20180 8888 20208 9055
rect 20254 9052 20260 9064
rect 20312 9052 20318 9104
rect 20257 8959 20315 8965
rect 20257 8925 20269 8959
rect 20303 8925 20315 8959
rect 20438 8956 20444 8968
rect 20399 8928 20444 8956
rect 20257 8919 20315 8925
rect 18380 8860 20208 8888
rect 18380 8848 18386 8860
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10778 8820 10784 8832
rect 9824 8792 10784 8820
rect 9824 8780 9830 8792
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 11882 8780 11888 8832
rect 11940 8820 11946 8832
rect 12066 8820 12072 8832
rect 11940 8792 12072 8820
rect 11940 8780 11946 8792
rect 12066 8780 12072 8792
rect 12124 8820 12130 8832
rect 12437 8823 12495 8829
rect 12437 8820 12449 8823
rect 12124 8792 12449 8820
rect 12124 8780 12130 8792
rect 12437 8789 12449 8792
rect 12483 8789 12495 8823
rect 12437 8783 12495 8789
rect 12710 8780 12716 8832
rect 12768 8820 12774 8832
rect 12897 8823 12955 8829
rect 12897 8820 12909 8823
rect 12768 8792 12909 8820
rect 12768 8780 12774 8792
rect 12897 8789 12909 8792
rect 12943 8789 12955 8823
rect 12897 8783 12955 8789
rect 16117 8823 16175 8829
rect 16117 8789 16129 8823
rect 16163 8820 16175 8823
rect 16393 8823 16451 8829
rect 16393 8820 16405 8823
rect 16163 8792 16405 8820
rect 16163 8789 16175 8792
rect 16117 8783 16175 8789
rect 16393 8789 16405 8792
rect 16439 8820 16451 8823
rect 18598 8820 18604 8832
rect 16439 8792 18604 8820
rect 16439 8789 16451 8792
rect 16393 8783 16451 8789
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 19794 8820 19800 8832
rect 19755 8792 19800 8820
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 20162 8780 20168 8832
rect 20220 8820 20226 8832
rect 20272 8820 20300 8919
rect 20438 8916 20444 8928
rect 20496 8916 20502 8968
rect 20220 8792 20300 8820
rect 20220 8780 20226 8792
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 8389 8619 8447 8625
rect 8389 8585 8401 8619
rect 8435 8616 8447 8619
rect 10042 8616 10048 8628
rect 8435 8588 10048 8616
rect 8435 8585 8447 8588
rect 8389 8579 8447 8585
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10962 8616 10968 8628
rect 10827 8588 10968 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 11756 8588 12204 8616
rect 11756 8576 11762 8588
rect 11348 8520 11744 8548
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 9364 8452 9413 8480
rect 9364 8440 9370 8452
rect 9401 8449 9413 8452
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 11348 8424 11376 8520
rect 11716 8489 11744 8520
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 12176 8480 12204 8588
rect 12250 8576 12256 8628
rect 12308 8616 12314 8628
rect 12434 8616 12440 8628
rect 12308 8588 12440 8616
rect 12308 8576 12314 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 14366 8576 14372 8628
rect 14424 8616 14430 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 14424 8588 16037 8616
rect 14424 8576 14430 8588
rect 16025 8585 16037 8588
rect 16071 8585 16083 8619
rect 16025 8579 16083 8585
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 17037 8619 17095 8625
rect 17037 8616 17049 8619
rect 16816 8588 17049 8616
rect 16816 8576 16822 8588
rect 17037 8585 17049 8588
rect 17083 8585 17095 8619
rect 17037 8579 17095 8585
rect 19242 8576 19248 8628
rect 19300 8616 19306 8628
rect 21085 8619 21143 8625
rect 21085 8616 21097 8619
rect 19300 8588 21097 8616
rect 19300 8576 19306 8588
rect 21085 8585 21097 8588
rect 21131 8585 21143 8619
rect 21085 8579 21143 8585
rect 13722 8508 13728 8560
rect 13780 8548 13786 8560
rect 13817 8551 13875 8557
rect 13817 8548 13829 8551
rect 13780 8520 13829 8548
rect 13780 8508 13786 8520
rect 13817 8517 13829 8520
rect 13863 8517 13875 8551
rect 15746 8548 15752 8560
rect 15707 8520 15752 8548
rect 13817 8511 13875 8517
rect 15746 8508 15752 8520
rect 15804 8508 15810 8560
rect 16114 8508 16120 8560
rect 16172 8548 16178 8560
rect 17497 8551 17555 8557
rect 17497 8548 17509 8551
rect 16172 8520 17509 8548
rect 16172 8508 16178 8520
rect 17497 8517 17509 8520
rect 17543 8517 17555 8551
rect 17497 8511 17555 8517
rect 18693 8551 18751 8557
rect 18693 8517 18705 8551
rect 18739 8548 18751 8551
rect 19334 8548 19340 8560
rect 18739 8520 19340 8548
rect 18739 8517 18751 8520
rect 18693 8511 18751 8517
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 12250 8480 12256 8492
rect 12163 8452 12256 8480
rect 11701 8443 11759 8449
rect 12250 8440 12256 8452
rect 12308 8480 12314 8492
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 12308 8452 12449 8480
rect 12308 8440 12314 8452
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 16482 8480 16488 8492
rect 16443 8452 16488 8480
rect 12437 8443 12495 8449
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8412 8815 8415
rect 8846 8412 8852 8424
rect 8803 8384 8852 8412
rect 8803 8381 8815 8384
rect 8757 8375 8815 8381
rect 8846 8372 8852 8384
rect 8904 8372 8910 8424
rect 9668 8415 9726 8421
rect 9668 8381 9680 8415
rect 9714 8412 9726 8415
rect 11330 8412 11336 8424
rect 9714 8384 11336 8412
rect 9714 8381 9726 8384
rect 9668 8375 9726 8381
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8412 11575 8415
rect 11974 8412 11980 8424
rect 11563 8384 11980 8412
rect 11563 8381 11575 8384
rect 11517 8375 11575 8381
rect 11974 8372 11980 8384
rect 12032 8412 12038 8424
rect 12342 8412 12348 8424
rect 12032 8384 12348 8412
rect 12032 8372 12038 8384
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 12452 8412 12480 8443
rect 16482 8440 16488 8452
rect 16540 8440 16546 8492
rect 16666 8480 16672 8492
rect 16627 8452 16672 8480
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8480 18107 8483
rect 18138 8480 18144 8492
rect 18095 8452 18144 8480
rect 18095 8449 18107 8452
rect 18049 8443 18107 8449
rect 18138 8440 18144 8452
rect 18196 8440 18202 8492
rect 19242 8480 19248 8492
rect 19203 8452 19248 8480
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 19426 8440 19432 8492
rect 19484 8480 19490 8492
rect 19705 8483 19763 8489
rect 19705 8480 19717 8483
rect 19484 8452 19717 8480
rect 19484 8440 19490 8452
rect 19705 8449 19717 8452
rect 19751 8449 19763 8483
rect 19705 8443 19763 8449
rect 14369 8415 14427 8421
rect 14369 8412 14381 8415
rect 12452 8384 14381 8412
rect 14369 8381 14381 8384
rect 14415 8381 14427 8415
rect 14369 8375 14427 8381
rect 14636 8415 14694 8421
rect 14636 8381 14648 8415
rect 14682 8412 14694 8415
rect 16684 8412 16712 8440
rect 14682 8384 16712 8412
rect 14682 8381 14694 8384
rect 14636 8375 14694 8381
rect 16850 8372 16856 8424
rect 16908 8412 16914 8424
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 16908 8384 17233 8412
rect 16908 8372 16914 8384
rect 17221 8381 17233 8384
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 19153 8415 19211 8421
rect 19153 8381 19165 8415
rect 19199 8412 19211 8415
rect 19794 8412 19800 8424
rect 19199 8384 19800 8412
rect 19199 8381 19211 8384
rect 19153 8375 19211 8381
rect 19794 8372 19800 8384
rect 19852 8372 19858 8424
rect 19972 8415 20030 8421
rect 19972 8381 19984 8415
rect 20018 8412 20030 8415
rect 20438 8412 20444 8424
rect 20018 8384 20444 8412
rect 20018 8381 20030 8384
rect 19972 8375 20030 8381
rect 20438 8372 20444 8384
rect 20496 8372 20502 8424
rect 7650 8304 7656 8356
rect 7708 8344 7714 8356
rect 9033 8347 9091 8353
rect 9033 8344 9045 8347
rect 7708 8316 9045 8344
rect 7708 8304 7714 8316
rect 9033 8313 9045 8316
rect 9079 8344 9091 8347
rect 10502 8344 10508 8356
rect 9079 8316 10508 8344
rect 9079 8313 9091 8316
rect 9033 8307 9091 8313
rect 10502 8304 10508 8316
rect 10560 8344 10566 8356
rect 11425 8347 11483 8353
rect 11425 8344 11437 8347
rect 10560 8316 11437 8344
rect 10560 8304 10566 8316
rect 11425 8313 11437 8316
rect 11471 8313 11483 8347
rect 11425 8307 11483 8313
rect 12704 8347 12762 8353
rect 12704 8313 12716 8347
rect 12750 8344 12762 8347
rect 14458 8344 14464 8356
rect 12750 8316 14464 8344
rect 12750 8313 12762 8316
rect 12704 8307 12762 8313
rect 14458 8304 14464 8316
rect 14516 8344 14522 8356
rect 15746 8344 15752 8356
rect 14516 8316 15752 8344
rect 14516 8304 14522 8316
rect 15746 8304 15752 8316
rect 15804 8304 15810 8356
rect 16393 8347 16451 8353
rect 16393 8344 16405 8347
rect 15856 8316 16405 8344
rect 10226 8236 10232 8288
rect 10284 8276 10290 8288
rect 11057 8279 11115 8285
rect 11057 8276 11069 8279
rect 10284 8248 11069 8276
rect 10284 8236 10290 8248
rect 11057 8245 11069 8248
rect 11103 8245 11115 8279
rect 11057 8239 11115 8245
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 14366 8276 14372 8288
rect 13504 8248 14372 8276
rect 13504 8236 13510 8248
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 14642 8236 14648 8288
rect 14700 8276 14706 8288
rect 15856 8276 15884 8316
rect 16393 8313 16405 8316
rect 16439 8313 16451 8347
rect 16393 8307 16451 8313
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 18138 8344 18144 8356
rect 16632 8316 18144 8344
rect 16632 8304 16638 8316
rect 18138 8304 18144 8316
rect 18196 8304 18202 8356
rect 19061 8347 19119 8353
rect 19061 8313 19073 8347
rect 19107 8344 19119 8347
rect 20346 8344 20352 8356
rect 19107 8316 20352 8344
rect 19107 8313 19119 8316
rect 19061 8307 19119 8313
rect 20346 8304 20352 8316
rect 20404 8304 20410 8356
rect 14700 8248 15884 8276
rect 14700 8236 14706 8248
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9677 8075 9735 8081
rect 9677 8072 9689 8075
rect 9539 8044 9689 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9677 8041 9689 8044
rect 9723 8041 9735 8075
rect 11054 8072 11060 8084
rect 11015 8044 11060 8072
rect 9677 8035 9735 8041
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 13998 8032 14004 8084
rect 14056 8072 14062 8084
rect 14185 8075 14243 8081
rect 14185 8072 14197 8075
rect 14056 8044 14197 8072
rect 14056 8032 14062 8044
rect 14185 8041 14197 8044
rect 14231 8041 14243 8075
rect 14550 8072 14556 8084
rect 14511 8044 14556 8072
rect 14185 8035 14243 8041
rect 14550 8032 14556 8044
rect 14608 8032 14614 8084
rect 14645 8075 14703 8081
rect 14645 8041 14657 8075
rect 14691 8072 14703 8075
rect 14734 8072 14740 8084
rect 14691 8044 14740 8072
rect 14691 8041 14703 8044
rect 14645 8035 14703 8041
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 16666 8072 16672 8084
rect 16627 8044 16672 8072
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 17589 8075 17647 8081
rect 17589 8041 17601 8075
rect 17635 8072 17647 8075
rect 17678 8072 17684 8084
rect 17635 8044 17684 8072
rect 17635 8041 17647 8044
rect 17589 8035 17647 8041
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 18233 8075 18291 8081
rect 18233 8041 18245 8075
rect 18279 8072 18291 8075
rect 19150 8072 19156 8084
rect 18279 8044 19156 8072
rect 18279 8041 18291 8044
rect 18233 8035 18291 8041
rect 19150 8032 19156 8044
rect 19208 8032 19214 8084
rect 20438 8032 20444 8084
rect 20496 8072 20502 8084
rect 20533 8075 20591 8081
rect 20533 8072 20545 8075
rect 20496 8044 20545 8072
rect 20496 8032 20502 8044
rect 20533 8041 20545 8044
rect 20579 8041 20591 8075
rect 20533 8035 20591 8041
rect 8573 8007 8631 8013
rect 8573 7973 8585 8007
rect 8619 8004 8631 8007
rect 9766 8004 9772 8016
rect 8619 7976 9772 8004
rect 8619 7973 8631 7976
rect 8573 7967 8631 7973
rect 9766 7964 9772 7976
rect 9824 8004 9830 8016
rect 10781 8007 10839 8013
rect 9824 7976 10732 8004
rect 9824 7964 9830 7976
rect 8849 7939 8907 7945
rect 8849 7905 8861 7939
rect 8895 7936 8907 7939
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 8895 7908 9505 7936
rect 8895 7905 8907 7908
rect 8849 7899 8907 7905
rect 9493 7905 9505 7908
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 10045 7939 10103 7945
rect 10045 7905 10057 7939
rect 10091 7936 10103 7939
rect 10704 7936 10732 7976
rect 10781 7973 10793 8007
rect 10827 8004 10839 8007
rect 11517 8007 11575 8013
rect 11517 8004 11529 8007
rect 10827 7976 11529 8004
rect 10827 7973 10839 7976
rect 10781 7967 10839 7973
rect 11517 7973 11529 7976
rect 11563 8004 11575 8007
rect 12066 8004 12072 8016
rect 11563 7976 12072 8004
rect 11563 7973 11575 7976
rect 11517 7967 11575 7973
rect 12066 7964 12072 7976
rect 12124 7964 12130 8016
rect 12520 8007 12578 8013
rect 12520 7973 12532 8007
rect 12566 8004 12578 8007
rect 13722 8004 13728 8016
rect 12566 7976 13728 8004
rect 12566 7973 12578 7976
rect 12520 7967 12578 7973
rect 13722 7964 13728 7976
rect 13780 7964 13786 8016
rect 17954 8004 17960 8016
rect 14476 7976 17960 8004
rect 11425 7939 11483 7945
rect 11425 7936 11437 7939
rect 10091 7908 10456 7936
rect 10704 7908 11437 7936
rect 10091 7905 10103 7908
rect 10045 7899 10103 7905
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7868 9183 7871
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 9171 7840 9413 7868
rect 9171 7837 9183 7840
rect 9125 7831 9183 7837
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 9732 7840 10149 7868
rect 9732 7828 9738 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10318 7868 10324 7880
rect 10279 7840 10324 7868
rect 10137 7831 10195 7837
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 7558 7760 7564 7812
rect 7616 7800 7622 7812
rect 10428 7800 10456 7908
rect 11425 7905 11437 7908
rect 11471 7936 11483 7939
rect 12250 7936 12256 7948
rect 11471 7908 12112 7936
rect 12211 7908 12256 7936
rect 11471 7905 11483 7908
rect 11425 7899 11483 7905
rect 11330 7828 11336 7880
rect 11388 7868 11394 7880
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11388 7840 11621 7868
rect 11388 7828 11394 7840
rect 11609 7837 11621 7840
rect 11655 7837 11667 7871
rect 12084 7868 12112 7908
rect 12250 7896 12256 7908
rect 12308 7896 12314 7948
rect 14476 7936 14504 7976
rect 17954 7964 17960 7976
rect 18012 7964 18018 8016
rect 18325 8007 18383 8013
rect 18325 7973 18337 8007
rect 18371 8004 18383 8007
rect 18690 8004 18696 8016
rect 18371 7976 18696 8004
rect 18371 7973 18383 7976
rect 18325 7967 18383 7973
rect 18690 7964 18696 7976
rect 18748 7964 18754 8016
rect 12360 7908 14504 7936
rect 15556 7939 15614 7945
rect 12360 7868 12388 7908
rect 15556 7905 15568 7939
rect 15602 7936 15614 7939
rect 16298 7936 16304 7948
rect 15602 7908 16304 7936
rect 15602 7905 15614 7908
rect 15556 7899 15614 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 16758 7896 16764 7948
rect 16816 7936 16822 7948
rect 17129 7939 17187 7945
rect 17129 7936 17141 7939
rect 16816 7908 17141 7936
rect 16816 7896 16822 7908
rect 17129 7905 17141 7908
rect 17175 7905 17187 7939
rect 17129 7899 17187 7905
rect 19420 7939 19478 7945
rect 19420 7905 19432 7939
rect 19466 7936 19478 7939
rect 20530 7936 20536 7948
rect 19466 7908 20536 7936
rect 19466 7905 19478 7908
rect 19420 7899 19478 7905
rect 20530 7896 20536 7908
rect 20588 7896 20594 7948
rect 12084 7840 12388 7868
rect 14829 7871 14887 7877
rect 11609 7831 11667 7837
rect 14829 7837 14841 7871
rect 14875 7868 14887 7871
rect 15194 7868 15200 7880
rect 14875 7840 15200 7868
rect 14875 7837 14887 7840
rect 14829 7831 14887 7837
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7837 18475 7871
rect 18417 7831 18475 7837
rect 7616 7772 10456 7800
rect 7616 7760 7622 7772
rect 7282 7692 7288 7744
rect 7340 7732 7346 7744
rect 8113 7735 8171 7741
rect 8113 7732 8125 7735
rect 7340 7704 8125 7732
rect 7340 7692 7346 7704
rect 8113 7701 8125 7704
rect 8159 7732 8171 7735
rect 8202 7732 8208 7744
rect 8159 7704 8208 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 10870 7732 10876 7744
rect 9447 7704 10876 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 13630 7732 13636 7744
rect 13591 7704 13636 7732
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 15304 7732 15332 7831
rect 16482 7760 16488 7812
rect 16540 7800 16546 7812
rect 17865 7803 17923 7809
rect 17865 7800 17877 7803
rect 16540 7772 17877 7800
rect 16540 7760 16546 7772
rect 17865 7769 17877 7772
rect 17911 7769 17923 7803
rect 17865 7763 17923 7769
rect 17954 7760 17960 7812
rect 18012 7800 18018 7812
rect 18432 7800 18460 7831
rect 18598 7828 18604 7880
rect 18656 7868 18662 7880
rect 19153 7871 19211 7877
rect 19153 7868 19165 7871
rect 18656 7840 19165 7868
rect 18656 7828 18662 7840
rect 19153 7837 19165 7840
rect 19199 7837 19211 7871
rect 20898 7868 20904 7880
rect 20859 7840 20904 7868
rect 19153 7831 19211 7837
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 18012 7772 18460 7800
rect 18012 7760 18018 7772
rect 16945 7735 17003 7741
rect 16945 7732 16957 7735
rect 15304 7704 16957 7732
rect 16945 7701 16957 7704
rect 16991 7732 17003 7735
rect 17126 7732 17132 7744
rect 16991 7704 17132 7732
rect 16991 7701 17003 7704
rect 16945 7695 17003 7701
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 7466 7488 7472 7540
rect 7524 7528 7530 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 7524 7500 7665 7528
rect 7524 7488 7530 7500
rect 7653 7497 7665 7500
rect 7699 7528 7711 7531
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 7699 7500 8217 7528
rect 7699 7497 7711 7500
rect 7653 7491 7711 7497
rect 8205 7497 8217 7500
rect 8251 7497 8263 7531
rect 8205 7491 8263 7497
rect 8404 7500 11192 7528
rect 8113 7463 8171 7469
rect 8113 7429 8125 7463
rect 8159 7460 8171 7463
rect 8404 7460 8432 7500
rect 11164 7472 11192 7500
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11425 7531 11483 7537
rect 11425 7528 11437 7531
rect 11296 7500 11437 7528
rect 11296 7488 11302 7500
rect 11425 7497 11437 7500
rect 11471 7497 11483 7531
rect 11974 7528 11980 7540
rect 11935 7500 11980 7528
rect 11425 7491 11483 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 14090 7488 14096 7540
rect 14148 7528 14154 7540
rect 14461 7531 14519 7537
rect 14461 7528 14473 7531
rect 14148 7500 14473 7528
rect 14148 7488 14154 7500
rect 14461 7497 14473 7500
rect 14507 7497 14519 7531
rect 16298 7528 16304 7540
rect 14461 7491 14519 7497
rect 14936 7500 16160 7528
rect 16259 7500 16304 7528
rect 8159 7432 8432 7460
rect 8159 7429 8171 7432
rect 8113 7423 8171 7429
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 14936 7460 14964 7500
rect 11204 7432 14964 7460
rect 16132 7460 16160 7500
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 20806 7460 20812 7472
rect 16132 7432 20812 7460
rect 11204 7420 11210 7432
rect 20806 7420 20812 7432
rect 20864 7420 20870 7472
rect 13630 7352 13636 7404
rect 13688 7392 13694 7404
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 13688 7364 14013 7392
rect 13688 7352 13694 7364
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 17589 7395 17647 7401
rect 17589 7361 17601 7395
rect 17635 7392 17647 7395
rect 17862 7392 17868 7404
rect 17635 7364 17868 7392
rect 17635 7361 17647 7364
rect 17589 7355 17647 7361
rect 17862 7352 17868 7364
rect 17920 7392 17926 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 17920 7364 18613 7392
rect 17920 7352 17926 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 20070 7392 20076 7404
rect 20031 7364 20076 7392
rect 18601 7355 18659 7361
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 21082 7392 21088 7404
rect 21043 7364 21088 7392
rect 21082 7352 21088 7364
rect 21140 7352 21146 7404
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 8260 7296 8401 7324
rect 8260 7284 8266 7296
rect 8389 7293 8401 7296
rect 8435 7324 8447 7327
rect 10045 7327 10103 7333
rect 10045 7324 10057 7327
rect 8435 7296 10057 7324
rect 8435 7293 8447 7296
rect 8389 7287 8447 7293
rect 10045 7293 10057 7296
rect 10091 7324 10103 7327
rect 10134 7324 10140 7336
rect 10091 7296 10140 7324
rect 10091 7293 10103 7296
rect 10045 7287 10103 7293
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10318 7333 10324 7336
rect 10312 7324 10324 7333
rect 10244 7296 10324 7324
rect 8662 7265 8668 7268
rect 8656 7256 8668 7265
rect 8623 7228 8668 7256
rect 8656 7219 8668 7228
rect 8662 7216 8668 7219
rect 8720 7216 8726 7268
rect 8205 7191 8263 7197
rect 8205 7157 8217 7191
rect 8251 7188 8263 7191
rect 8386 7188 8392 7200
rect 8251 7160 8392 7188
rect 8251 7157 8263 7160
rect 8205 7151 8263 7157
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 9769 7191 9827 7197
rect 9769 7157 9781 7191
rect 9815 7188 9827 7191
rect 10244 7188 10272 7296
rect 10312 7287 10324 7296
rect 10318 7284 10324 7287
rect 10376 7284 10382 7336
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 13538 7324 13544 7336
rect 11204 7296 13544 7324
rect 11204 7284 11210 7296
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 13817 7327 13875 7333
rect 13817 7293 13829 7327
rect 13863 7324 13875 7327
rect 14090 7324 14096 7336
rect 13863 7296 14096 7324
rect 13863 7293 13875 7296
rect 13817 7287 13875 7293
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 17126 7324 17132 7336
rect 14967 7296 17132 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 17126 7284 17132 7296
rect 17184 7284 17190 7336
rect 17405 7327 17463 7333
rect 17405 7293 17417 7327
rect 17451 7324 17463 7327
rect 17678 7324 17684 7336
rect 17451 7296 17684 7324
rect 17451 7293 17463 7296
rect 17405 7287 17463 7293
rect 17678 7284 17684 7296
rect 17736 7284 17742 7336
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 17972 7296 18521 7324
rect 12250 7216 12256 7268
rect 12308 7256 12314 7268
rect 12618 7256 12624 7268
rect 12308 7228 12624 7256
rect 12308 7216 12314 7228
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 13173 7259 13231 7265
rect 13173 7225 13185 7259
rect 13219 7256 13231 7259
rect 13354 7256 13360 7268
rect 13219 7228 13360 7256
rect 13219 7225 13231 7228
rect 13173 7219 13231 7225
rect 13354 7216 13360 7228
rect 13412 7216 13418 7268
rect 14366 7216 14372 7268
rect 14424 7256 14430 7268
rect 15188 7259 15246 7265
rect 14424 7228 14596 7256
rect 14424 7216 14430 7228
rect 12526 7188 12532 7200
rect 9815 7160 10272 7188
rect 12487 7160 12532 7188
rect 9815 7157 9827 7160
rect 9769 7151 9827 7157
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 13446 7188 13452 7200
rect 13407 7160 13452 7188
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 13909 7191 13967 7197
rect 13909 7157 13921 7191
rect 13955 7188 13967 7191
rect 14458 7188 14464 7200
rect 13955 7160 14464 7188
rect 13955 7157 13967 7160
rect 13909 7151 13967 7157
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 14568 7188 14596 7228
rect 15188 7225 15200 7259
rect 15234 7256 15246 7259
rect 16390 7256 16396 7268
rect 15234 7228 16396 7256
rect 15234 7225 15246 7228
rect 15188 7219 15246 7225
rect 16390 7216 16396 7228
rect 16448 7216 16454 7268
rect 16669 7259 16727 7265
rect 16669 7225 16681 7259
rect 16715 7256 16727 7259
rect 17313 7259 17371 7265
rect 17313 7256 17325 7259
rect 16715 7228 17325 7256
rect 16715 7225 16727 7228
rect 16669 7219 16727 7225
rect 17313 7225 17325 7228
rect 17359 7225 17371 7259
rect 17972 7256 18000 7296
rect 18509 7293 18521 7296
rect 18555 7324 18567 7327
rect 18874 7324 18880 7336
rect 18555 7296 18880 7324
rect 18555 7293 18567 7296
rect 18509 7287 18567 7293
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 19153 7327 19211 7333
rect 19153 7293 19165 7327
rect 19199 7324 19211 7327
rect 19889 7327 19947 7333
rect 19199 7296 19840 7324
rect 19199 7293 19211 7296
rect 19153 7287 19211 7293
rect 17313 7219 17371 7225
rect 17420 7228 18000 7256
rect 18417 7259 18475 7265
rect 16684 7188 16712 7219
rect 14568 7160 16712 7188
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 16945 7191 17003 7197
rect 16945 7188 16957 7191
rect 16816 7160 16957 7188
rect 16816 7148 16822 7160
rect 16945 7157 16957 7160
rect 16991 7157 17003 7191
rect 16945 7151 17003 7157
rect 17218 7148 17224 7200
rect 17276 7188 17282 7200
rect 17420 7188 17448 7228
rect 18417 7225 18429 7259
rect 18463 7256 18475 7259
rect 19242 7256 19248 7268
rect 18463 7228 19248 7256
rect 18463 7225 18475 7228
rect 18417 7219 18475 7225
rect 19242 7216 19248 7228
rect 19300 7216 19306 7268
rect 19812 7256 19840 7296
rect 19889 7293 19901 7327
rect 19935 7324 19947 7327
rect 20898 7324 20904 7336
rect 19935 7296 20904 7324
rect 19935 7293 19947 7296
rect 19889 7287 19947 7293
rect 20898 7284 20904 7296
rect 20956 7284 20962 7336
rect 20622 7256 20628 7268
rect 19812 7228 20628 7256
rect 20622 7216 20628 7228
rect 20680 7256 20686 7268
rect 20993 7259 21051 7265
rect 20993 7256 21005 7259
rect 20680 7228 21005 7256
rect 20680 7216 20686 7228
rect 20993 7225 21005 7228
rect 21039 7225 21051 7259
rect 20993 7219 21051 7225
rect 17276 7160 17448 7188
rect 17276 7148 17282 7160
rect 17494 7148 17500 7200
rect 17552 7188 17558 7200
rect 18049 7191 18107 7197
rect 18049 7188 18061 7191
rect 17552 7160 18061 7188
rect 17552 7148 17558 7160
rect 18049 7157 18061 7160
rect 18095 7157 18107 7191
rect 19518 7188 19524 7200
rect 19479 7160 19524 7188
rect 18049 7151 18107 7157
rect 19518 7148 19524 7160
rect 19576 7148 19582 7200
rect 19886 7148 19892 7200
rect 19944 7188 19950 7200
rect 19981 7191 20039 7197
rect 19981 7188 19993 7191
rect 19944 7160 19993 7188
rect 19944 7148 19950 7160
rect 19981 7157 19993 7160
rect 20027 7157 20039 7191
rect 19981 7151 20039 7157
rect 20162 7148 20168 7200
rect 20220 7188 20226 7200
rect 20533 7191 20591 7197
rect 20533 7188 20545 7191
rect 20220 7160 20545 7188
rect 20220 7148 20226 7160
rect 20533 7157 20545 7160
rect 20579 7157 20591 7191
rect 20533 7151 20591 7157
rect 20806 7148 20812 7200
rect 20864 7188 20870 7200
rect 20901 7191 20959 7197
rect 20901 7188 20913 7191
rect 20864 7160 20913 7188
rect 20864 7148 20870 7160
rect 20901 7157 20913 7160
rect 20947 7157 20959 7191
rect 20901 7151 20959 7157
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 7558 6984 7564 6996
rect 7519 6956 7564 6984
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 8938 6984 8944 6996
rect 8899 6956 8944 6984
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 9674 6984 9680 6996
rect 9635 6956 9680 6984
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 10137 6987 10195 6993
rect 10137 6953 10149 6987
rect 10183 6984 10195 6987
rect 10689 6987 10747 6993
rect 10689 6984 10701 6987
rect 10183 6956 10701 6984
rect 10183 6953 10195 6956
rect 10137 6947 10195 6953
rect 10689 6953 10701 6956
rect 10735 6953 10747 6987
rect 10689 6947 10747 6953
rect 11057 6987 11115 6993
rect 11057 6953 11069 6987
rect 11103 6984 11115 6987
rect 12526 6984 12532 6996
rect 11103 6956 12532 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 12526 6944 12532 6956
rect 12584 6984 12590 6996
rect 13262 6984 13268 6996
rect 12584 6956 13268 6984
rect 12584 6944 12590 6956
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 13354 6944 13360 6996
rect 13412 6984 13418 6996
rect 15838 6984 15844 6996
rect 13412 6956 15844 6984
rect 13412 6944 13418 6956
rect 15838 6944 15844 6956
rect 15896 6944 15902 6996
rect 16482 6984 16488 6996
rect 16443 6956 16488 6984
rect 16482 6944 16488 6956
rect 16540 6944 16546 6996
rect 16577 6987 16635 6993
rect 16577 6953 16589 6987
rect 16623 6984 16635 6987
rect 17494 6984 17500 6996
rect 16623 6956 17500 6984
rect 16623 6953 16635 6956
rect 16577 6947 16635 6953
rect 17494 6944 17500 6956
rect 17552 6944 17558 6996
rect 18877 6987 18935 6993
rect 18877 6953 18889 6987
rect 18923 6984 18935 6987
rect 19150 6984 19156 6996
rect 18923 6956 19156 6984
rect 18923 6953 18935 6956
rect 18877 6947 18935 6953
rect 19150 6944 19156 6956
rect 19208 6944 19214 6996
rect 20530 6984 20536 6996
rect 20491 6956 20536 6984
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 7929 6919 7987 6925
rect 7929 6885 7941 6919
rect 7975 6916 7987 6919
rect 9582 6916 9588 6928
rect 7975 6888 9588 6916
rect 7975 6885 7987 6888
rect 7929 6879 7987 6885
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 11146 6916 11152 6928
rect 9876 6888 11152 6916
rect 7190 6808 7196 6860
rect 7248 6848 7254 6860
rect 8754 6848 8760 6860
rect 7248 6820 8760 6848
rect 7248 6808 7254 6820
rect 8754 6808 8760 6820
rect 8812 6848 8818 6860
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 8812 6820 9045 6848
rect 8812 6808 8818 6820
rect 9033 6817 9045 6820
rect 9079 6817 9091 6851
rect 9033 6811 9091 6817
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 9876 6848 9904 6888
rect 11146 6876 11152 6888
rect 11204 6876 11210 6928
rect 12704 6919 12762 6925
rect 12704 6885 12716 6919
rect 12750 6916 12762 6919
rect 13630 6916 13636 6928
rect 12750 6888 13636 6916
rect 12750 6885 12762 6888
rect 12704 6879 12762 6885
rect 13630 6876 13636 6888
rect 13688 6916 13694 6928
rect 13688 6888 14688 6916
rect 13688 6876 13694 6888
rect 10042 6848 10048 6860
rect 9548 6820 9904 6848
rect 10003 6820 10048 6848
rect 9548 6808 9554 6820
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 11882 6848 11888 6860
rect 11843 6820 11888 6848
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 14366 6808 14372 6860
rect 14424 6848 14430 6860
rect 14461 6851 14519 6857
rect 14461 6848 14473 6851
rect 14424 6820 14473 6848
rect 14424 6808 14430 6820
rect 14461 6817 14473 6820
rect 14507 6817 14519 6851
rect 14461 6811 14519 6817
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 8662 6780 8668 6792
rect 8251 6752 8668 6780
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 6917 6715 6975 6721
rect 6917 6681 6929 6715
rect 6963 6712 6975 6715
rect 8036 6712 8064 6743
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8956 6752 9137 6780
rect 8573 6715 8631 6721
rect 8573 6712 8585 6715
rect 6963 6684 7972 6712
rect 8036 6684 8585 6712
rect 6963 6681 6975 6684
rect 6917 6675 6975 6681
rect 7190 6644 7196 6656
rect 7151 6616 7196 6644
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7944 6644 7972 6684
rect 8573 6681 8585 6684
rect 8619 6681 8631 6715
rect 8573 6675 8631 6681
rect 8754 6672 8760 6724
rect 8812 6712 8818 6724
rect 8956 6712 8984 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 9364 6752 10241 6780
rect 9364 6740 9370 6752
rect 10229 6749 10241 6752
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 10870 6740 10876 6792
rect 10928 6780 10934 6792
rect 11241 6783 11299 6789
rect 11241 6780 11253 6783
rect 10928 6752 11253 6780
rect 10928 6740 10934 6752
rect 11241 6749 11253 6752
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 8812 6684 8984 6712
rect 8812 6672 8818 6684
rect 12452 6656 12480 6743
rect 14182 6740 14188 6792
rect 14240 6780 14246 6792
rect 14660 6789 14688 6888
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 17218 6916 17224 6928
rect 14792 6888 17224 6916
rect 14792 6876 14798 6888
rect 17218 6876 17224 6888
rect 17276 6876 17282 6928
rect 17396 6919 17454 6925
rect 17396 6885 17408 6919
rect 17442 6916 17454 6919
rect 17862 6916 17868 6928
rect 17442 6888 17868 6916
rect 17442 6885 17454 6888
rect 17396 6879 17454 6885
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 19420 6919 19478 6925
rect 19420 6885 19432 6919
rect 19466 6916 19478 6919
rect 20070 6916 20076 6928
rect 19466 6888 20076 6916
rect 19466 6885 19478 6888
rect 19420 6879 19478 6885
rect 20070 6876 20076 6888
rect 20128 6876 20134 6928
rect 15749 6851 15807 6857
rect 15749 6817 15761 6851
rect 15795 6848 15807 6851
rect 16114 6848 16120 6860
rect 15795 6820 16120 6848
rect 15795 6817 15807 6820
rect 15749 6811 15807 6817
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 17126 6848 17132 6860
rect 17039 6820 17132 6848
rect 17126 6808 17132 6820
rect 17184 6848 17190 6860
rect 18598 6848 18604 6860
rect 17184 6820 18604 6848
rect 17184 6808 17190 6820
rect 18598 6808 18604 6820
rect 18656 6848 18662 6860
rect 19153 6851 19211 6857
rect 19153 6848 19165 6851
rect 18656 6820 19165 6848
rect 18656 6808 18662 6820
rect 19153 6817 19165 6820
rect 19199 6817 19211 6851
rect 19153 6811 19211 6817
rect 19702 6808 19708 6860
rect 19760 6848 19766 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 19760 6820 20913 6848
rect 19760 6808 19766 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 14240 6752 14565 6780
rect 14240 6740 14246 6752
rect 14553 6749 14565 6752
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 14568 6712 14596 6743
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 16669 6783 16727 6789
rect 16669 6780 16681 6783
rect 16448 6752 16681 6780
rect 16448 6740 16454 6752
rect 16669 6749 16681 6752
rect 16715 6749 16727 6783
rect 16669 6743 16727 6749
rect 15289 6715 15347 6721
rect 15289 6712 15301 6715
rect 14568 6684 15301 6712
rect 15289 6681 15301 6684
rect 15335 6681 15347 6715
rect 15289 6675 15347 6681
rect 8662 6644 8668 6656
rect 7944 6616 8668 6644
rect 8662 6604 8668 6616
rect 8720 6644 8726 6656
rect 9490 6644 9496 6656
rect 8720 6616 9496 6644
rect 8720 6604 8726 6616
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 10192 6616 11713 6644
rect 10192 6604 10198 6616
rect 11701 6613 11713 6616
rect 11747 6644 11759 6647
rect 12434 6644 12440 6656
rect 11747 6616 12440 6644
rect 11747 6613 11759 6616
rect 11701 6607 11759 6613
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 13722 6604 13728 6656
rect 13780 6644 13786 6656
rect 13817 6647 13875 6653
rect 13817 6644 13829 6647
rect 13780 6616 13829 6644
rect 13780 6604 13786 6616
rect 13817 6613 13829 6616
rect 13863 6613 13875 6647
rect 13817 6607 13875 6613
rect 14093 6647 14151 6653
rect 14093 6613 14105 6647
rect 14139 6644 14151 6647
rect 14550 6644 14556 6656
rect 14139 6616 14556 6644
rect 14139 6613 14151 6616
rect 14093 6607 14151 6613
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 15746 6604 15752 6656
rect 15804 6644 15810 6656
rect 16117 6647 16175 6653
rect 16117 6644 16129 6647
rect 15804 6616 16129 6644
rect 15804 6604 15810 6616
rect 16117 6613 16129 6616
rect 16163 6613 16175 6647
rect 16684 6644 16712 6743
rect 18966 6672 18972 6724
rect 19024 6712 19030 6724
rect 19150 6712 19156 6724
rect 19024 6684 19156 6712
rect 19024 6672 19030 6684
rect 19150 6672 19156 6684
rect 19208 6672 19214 6724
rect 18509 6647 18567 6653
rect 18509 6644 18521 6647
rect 16684 6616 18521 6644
rect 16117 6607 16175 6613
rect 18509 6613 18521 6616
rect 18555 6613 18567 6647
rect 18509 6607 18567 6613
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 7193 6443 7251 6449
rect 7193 6440 7205 6443
rect 7156 6412 7205 6440
rect 7156 6400 7162 6412
rect 7193 6409 7205 6412
rect 7239 6409 7251 6443
rect 8202 6440 8208 6452
rect 7193 6403 7251 6409
rect 7944 6412 8208 6440
rect 6822 6196 6828 6248
rect 6880 6236 6886 6248
rect 7944 6245 7972 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 9122 6440 9128 6452
rect 8720 6412 9128 6440
rect 8720 6400 8726 6412
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 9306 6440 9312 6452
rect 9267 6412 9312 6440
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 10100 6412 10333 6440
rect 10100 6400 10106 6412
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 14366 6440 14372 6452
rect 10321 6403 10379 6409
rect 11256 6412 13216 6440
rect 14327 6412 14372 6440
rect 9858 6332 9864 6384
rect 9916 6372 9922 6384
rect 11256 6372 11284 6412
rect 9916 6344 11284 6372
rect 11333 6375 11391 6381
rect 9916 6332 9922 6344
rect 11333 6341 11345 6375
rect 11379 6372 11391 6375
rect 12161 6375 12219 6381
rect 12161 6372 12173 6375
rect 11379 6344 12173 6372
rect 11379 6341 11391 6344
rect 11333 6335 11391 6341
rect 12161 6341 12173 6344
rect 12207 6341 12219 6375
rect 13078 6372 13084 6384
rect 12161 6335 12219 6341
rect 12268 6344 13084 6372
rect 9582 6304 9588 6316
rect 9543 6276 9588 6304
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 10870 6304 10876 6316
rect 10783 6276 10876 6304
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 11054 6264 11060 6316
rect 11112 6304 11118 6316
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 11112 6276 11989 6304
rect 11112 6264 11118 6276
rect 11977 6273 11989 6276
rect 12023 6304 12035 6307
rect 12268 6304 12296 6344
rect 13078 6332 13084 6344
rect 13136 6332 13142 6384
rect 12023 6276 12296 6304
rect 13188 6304 13216 6412
rect 14366 6400 14372 6412
rect 14424 6400 14430 6452
rect 16117 6443 16175 6449
rect 16117 6409 16129 6443
rect 16163 6440 16175 6443
rect 16301 6443 16359 6449
rect 16301 6440 16313 6443
rect 16163 6412 16313 6440
rect 16163 6409 16175 6412
rect 16117 6403 16175 6409
rect 16301 6409 16313 6412
rect 16347 6409 16359 6443
rect 16301 6403 16359 6409
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 16908 6412 17448 6440
rect 16908 6400 16914 6412
rect 17420 6384 17448 6412
rect 17678 6400 17684 6452
rect 17736 6440 17742 6452
rect 18417 6443 18475 6449
rect 18417 6440 18429 6443
rect 17736 6412 18429 6440
rect 17736 6400 17742 6412
rect 18417 6409 18429 6412
rect 18463 6409 18475 6443
rect 18417 6403 18475 6409
rect 18966 6400 18972 6452
rect 19024 6440 19030 6452
rect 19024 6412 19840 6440
rect 19024 6400 19030 6412
rect 13538 6332 13544 6384
rect 13596 6372 13602 6384
rect 15289 6375 15347 6381
rect 15289 6372 15301 6375
rect 13596 6344 15301 6372
rect 13596 6332 13602 6344
rect 15289 6341 15301 6344
rect 15335 6341 15347 6375
rect 15289 6335 15347 6341
rect 16390 6332 16396 6384
rect 16448 6372 16454 6384
rect 16448 6344 16896 6372
rect 16448 6332 16454 6344
rect 13188 6276 13553 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 8202 6245 8208 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 6880 6208 7941 6236
rect 6880 6196 6886 6208
rect 7929 6205 7941 6208
rect 7975 6205 7987 6239
rect 8196 6236 8208 6245
rect 8115 6208 8208 6236
rect 7929 6199 7987 6205
rect 8196 6199 8208 6208
rect 8260 6236 8266 6248
rect 8754 6236 8760 6248
rect 8260 6208 8760 6236
rect 8202 6196 8208 6199
rect 8260 6196 8266 6208
rect 8754 6196 8760 6208
rect 8812 6236 8818 6248
rect 10888 6236 10916 6264
rect 12529 6239 12587 6245
rect 12529 6236 12541 6239
rect 8812 6208 10916 6236
rect 11532 6208 12541 6236
rect 8812 6196 8818 6208
rect 10042 6128 10048 6180
rect 10100 6168 10106 6180
rect 10781 6171 10839 6177
rect 10781 6168 10793 6171
rect 10100 6140 10793 6168
rect 10100 6128 10106 6140
rect 10781 6137 10793 6140
rect 10827 6168 10839 6171
rect 10870 6168 10876 6180
rect 10827 6140 10876 6168
rect 10827 6137 10839 6140
rect 10781 6131 10839 6137
rect 10870 6128 10876 6140
rect 10928 6128 10934 6180
rect 7653 6103 7711 6109
rect 7653 6069 7665 6103
rect 7699 6100 7711 6103
rect 9950 6100 9956 6112
rect 7699 6072 9956 6100
rect 7699 6069 7711 6072
rect 7653 6063 7711 6069
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 10689 6103 10747 6109
rect 10689 6069 10701 6103
rect 10735 6100 10747 6103
rect 11532 6100 11560 6208
rect 12529 6205 12541 6208
rect 12575 6236 12587 6239
rect 13525 6236 13553 6276
rect 13630 6264 13636 6316
rect 13688 6304 13694 6316
rect 13909 6307 13967 6313
rect 13909 6304 13921 6307
rect 13688 6276 13921 6304
rect 13688 6264 13694 6276
rect 13909 6273 13921 6276
rect 13955 6273 13967 6307
rect 15746 6304 15752 6316
rect 15707 6276 15752 6304
rect 13909 6267 13967 6273
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16298 6304 16304 6316
rect 15979 6276 16304 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 16758 6304 16764 6316
rect 16719 6276 16764 6304
rect 16758 6264 16764 6276
rect 16816 6264 16822 6316
rect 16868 6313 16896 6344
rect 17402 6332 17408 6384
rect 17460 6372 17466 6384
rect 18049 6375 18107 6381
rect 18049 6372 18061 6375
rect 17460 6344 18061 6372
rect 17460 6332 17466 6344
rect 18049 6341 18061 6344
rect 18095 6341 18107 6375
rect 18049 6335 18107 6341
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6273 16911 6307
rect 19812 6304 19840 6412
rect 20901 6307 20959 6313
rect 20901 6304 20913 6307
rect 19812 6276 20913 6304
rect 16853 6267 16911 6273
rect 20901 6273 20913 6276
rect 20947 6273 20959 6307
rect 21082 6304 21088 6316
rect 21043 6276 21088 6304
rect 20901 6267 20959 6273
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 13814 6236 13820 6248
rect 12575 6208 13492 6236
rect 13525 6208 13820 6236
rect 12575 6205 12587 6208
rect 12529 6199 12587 6205
rect 11793 6171 11851 6177
rect 11793 6137 11805 6171
rect 11839 6168 11851 6171
rect 12986 6168 12992 6180
rect 11839 6140 12992 6168
rect 11839 6137 11851 6140
rect 11793 6131 11851 6137
rect 12986 6128 12992 6140
rect 13044 6128 13050 6180
rect 13464 6168 13492 6208
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 15838 6196 15844 6248
rect 15896 6236 15902 6248
rect 18138 6236 18144 6248
rect 15896 6208 18144 6236
rect 15896 6196 15902 6208
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 18598 6196 18604 6248
rect 18656 6236 18662 6248
rect 18785 6239 18843 6245
rect 18785 6236 18797 6239
rect 18656 6208 18797 6236
rect 18656 6196 18662 6208
rect 18785 6205 18797 6208
rect 18831 6205 18843 6239
rect 18785 6199 18843 6205
rect 18874 6196 18880 6248
rect 18932 6236 18938 6248
rect 19052 6239 19110 6245
rect 19052 6236 19064 6239
rect 18932 6208 19064 6236
rect 18932 6196 18938 6208
rect 19052 6205 19064 6208
rect 19098 6236 19110 6239
rect 21100 6236 21128 6264
rect 19098 6208 21128 6236
rect 19098 6205 19110 6208
rect 19052 6199 19110 6205
rect 13464 6140 13584 6168
rect 11698 6100 11704 6112
rect 10735 6072 11560 6100
rect 11659 6072 11704 6100
rect 10735 6069 10747 6072
rect 10689 6063 10747 6069
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 12161 6103 12219 6109
rect 12161 6069 12173 6103
rect 12207 6100 12219 6103
rect 12618 6100 12624 6112
rect 12207 6072 12624 6100
rect 12207 6069 12219 6072
rect 12161 6063 12219 6069
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 12894 6100 12900 6112
rect 12855 6072 12900 6100
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13354 6100 13360 6112
rect 13315 6072 13360 6100
rect 13354 6060 13360 6072
rect 13412 6060 13418 6112
rect 13556 6100 13584 6140
rect 13630 6128 13636 6180
rect 13688 6168 13694 6180
rect 13725 6171 13783 6177
rect 13725 6168 13737 6171
rect 13688 6140 13737 6168
rect 13688 6128 13694 6140
rect 13725 6137 13737 6140
rect 13771 6137 13783 6171
rect 15657 6171 15715 6177
rect 13725 6131 13783 6137
rect 14200 6140 15608 6168
rect 14200 6100 14228 6140
rect 13556 6072 14228 6100
rect 14458 6060 14464 6112
rect 14516 6100 14522 6112
rect 14737 6103 14795 6109
rect 14737 6100 14749 6103
rect 14516 6072 14749 6100
rect 14516 6060 14522 6072
rect 14737 6069 14749 6072
rect 14783 6069 14795 6103
rect 15580 6100 15608 6140
rect 15657 6137 15669 6171
rect 15703 6168 15715 6171
rect 16117 6171 16175 6177
rect 16117 6168 16129 6171
rect 15703 6140 16129 6168
rect 15703 6137 15715 6140
rect 15657 6131 15715 6137
rect 16117 6137 16129 6140
rect 16163 6137 16175 6171
rect 16117 6131 16175 6137
rect 16669 6171 16727 6177
rect 16669 6137 16681 6171
rect 16715 6168 16727 6171
rect 17313 6171 17371 6177
rect 17313 6168 17325 6171
rect 16715 6140 17325 6168
rect 16715 6137 16727 6140
rect 16669 6131 16727 6137
rect 17313 6137 17325 6140
rect 17359 6137 17371 6171
rect 17313 6131 17371 6137
rect 17954 6128 17960 6180
rect 18012 6168 18018 6180
rect 20809 6171 20867 6177
rect 20809 6168 20821 6171
rect 18012 6140 20821 6168
rect 18012 6128 18018 6140
rect 20809 6137 20821 6140
rect 20855 6137 20867 6171
rect 20809 6131 20867 6137
rect 16850 6100 16856 6112
rect 15580 6072 16856 6100
rect 14737 6063 14795 6069
rect 16850 6060 16856 6072
rect 16908 6060 16914 6112
rect 20070 6060 20076 6112
rect 20128 6100 20134 6112
rect 20165 6103 20223 6109
rect 20165 6100 20177 6103
rect 20128 6072 20177 6100
rect 20128 6060 20134 6072
rect 20165 6069 20177 6072
rect 20211 6069 20223 6103
rect 20165 6063 20223 6069
rect 20254 6060 20260 6112
rect 20312 6100 20318 6112
rect 20441 6103 20499 6109
rect 20441 6100 20453 6103
rect 20312 6072 20453 6100
rect 20312 6060 20318 6072
rect 20441 6069 20453 6072
rect 20487 6069 20499 6103
rect 20441 6063 20499 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 8202 5896 8208 5908
rect 8163 5868 8208 5896
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 8938 5896 8944 5908
rect 8619 5868 8944 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 8938 5856 8944 5868
rect 8996 5856 9002 5908
rect 9030 5856 9036 5908
rect 9088 5896 9094 5908
rect 9217 5899 9275 5905
rect 9217 5896 9229 5899
rect 9088 5868 9229 5896
rect 9088 5856 9094 5868
rect 9217 5865 9229 5868
rect 9263 5896 9275 5899
rect 9490 5896 9496 5908
rect 9263 5868 9496 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 10042 5896 10048 5908
rect 10003 5868 10048 5896
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 10502 5856 10508 5908
rect 10560 5856 10566 5908
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 11756 5868 14105 5896
rect 11756 5856 11762 5868
rect 14093 5865 14105 5868
rect 14139 5865 14151 5899
rect 14550 5896 14556 5908
rect 14511 5868 14556 5896
rect 14093 5859 14151 5865
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 15289 5899 15347 5905
rect 15289 5865 15301 5899
rect 15335 5896 15347 5899
rect 16761 5899 16819 5905
rect 16761 5896 16773 5899
rect 15335 5868 16773 5896
rect 15335 5865 15347 5868
rect 15289 5859 15347 5865
rect 16761 5865 16773 5868
rect 16807 5865 16819 5899
rect 16761 5859 16819 5865
rect 18693 5899 18751 5905
rect 18693 5865 18705 5899
rect 18739 5896 18751 5899
rect 18874 5896 18880 5908
rect 18739 5868 18880 5896
rect 18739 5865 18751 5868
rect 18693 5859 18751 5865
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 19521 5899 19579 5905
rect 19521 5865 19533 5899
rect 19567 5896 19579 5899
rect 19886 5896 19892 5908
rect 19567 5868 19892 5896
rect 19567 5865 19579 5868
rect 19521 5859 19579 5865
rect 19886 5856 19892 5868
rect 19944 5856 19950 5908
rect 20254 5896 20260 5908
rect 20215 5868 20260 5896
rect 20254 5856 20260 5868
rect 20312 5856 20318 5908
rect 8849 5831 8907 5837
rect 8849 5797 8861 5831
rect 8895 5828 8907 5831
rect 9122 5828 9128 5840
rect 8895 5800 9128 5828
rect 8895 5797 8907 5800
rect 8849 5791 8907 5797
rect 9122 5788 9128 5800
rect 9180 5828 9186 5840
rect 10520 5828 10548 5856
rect 9180 5800 10548 5828
rect 9180 5788 9186 5800
rect 4062 5720 4068 5772
rect 4120 5760 4126 5772
rect 6457 5763 6515 5769
rect 6457 5760 6469 5763
rect 4120 5732 6469 5760
rect 4120 5720 4126 5732
rect 6457 5729 6469 5732
rect 6503 5760 6515 5763
rect 7081 5763 7139 5769
rect 7081 5760 7093 5763
rect 6503 5732 7093 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 7081 5729 7093 5732
rect 7127 5729 7139 5763
rect 7081 5723 7139 5729
rect 10134 5720 10140 5772
rect 10192 5760 10198 5772
rect 10321 5763 10379 5769
rect 10321 5760 10333 5763
rect 10192 5732 10333 5760
rect 10192 5720 10198 5732
rect 10321 5729 10333 5732
rect 10367 5729 10379 5763
rect 10520 5760 10548 5800
rect 10588 5831 10646 5837
rect 10588 5797 10600 5831
rect 10634 5828 10646 5831
rect 11054 5828 11060 5840
rect 10634 5800 11060 5828
rect 10634 5797 10646 5800
rect 10588 5791 10646 5797
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 12618 5788 12624 5840
rect 12676 5828 12682 5840
rect 12802 5828 12808 5840
rect 12676 5800 12808 5828
rect 12676 5788 12682 5800
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 12894 5788 12900 5840
rect 12952 5828 12958 5840
rect 14461 5831 14519 5837
rect 14461 5828 14473 5831
rect 12952 5800 14473 5828
rect 12952 5788 12958 5800
rect 14461 5797 14473 5800
rect 14507 5797 14519 5831
rect 14461 5791 14519 5797
rect 14826 5788 14832 5840
rect 14884 5828 14890 5840
rect 15657 5831 15715 5837
rect 15657 5828 15669 5831
rect 14884 5800 15669 5828
rect 14884 5788 14890 5800
rect 15657 5797 15669 5800
rect 15703 5828 15715 5831
rect 15703 5800 16804 5828
rect 15703 5797 15715 5800
rect 15657 5791 15715 5797
rect 11882 5760 11888 5772
rect 10520 5732 11888 5760
rect 10321 5723 10379 5729
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 12066 5760 12072 5772
rect 12027 5732 12072 5760
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12704 5763 12762 5769
rect 12492 5732 12537 5760
rect 12492 5720 12498 5732
rect 12704 5729 12716 5763
rect 12750 5760 12762 5763
rect 16666 5760 16672 5772
rect 12750 5732 13768 5760
rect 16627 5732 16672 5760
rect 12750 5729 12762 5732
rect 12704 5723 12762 5729
rect 13740 5704 13768 5732
rect 16666 5720 16672 5732
rect 16724 5720 16730 5772
rect 16776 5760 16804 5800
rect 17494 5788 17500 5840
rect 17552 5837 17558 5840
rect 17552 5831 17616 5837
rect 17552 5797 17570 5831
rect 17604 5797 17616 5831
rect 20162 5828 20168 5840
rect 20123 5800 20168 5828
rect 17552 5791 17616 5797
rect 17552 5788 17558 5791
rect 20162 5788 20168 5800
rect 20220 5788 20226 5840
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 16776 5732 20913 5760
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 6822 5692 6828 5704
rect 6783 5664 6828 5692
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 13722 5652 13728 5704
rect 13780 5692 13786 5704
rect 14645 5695 14703 5701
rect 14645 5692 14657 5695
rect 13780 5664 14657 5692
rect 13780 5652 13786 5664
rect 14645 5661 14657 5664
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 15562 5652 15568 5704
rect 15620 5692 15626 5704
rect 15749 5695 15807 5701
rect 15749 5692 15761 5695
rect 15620 5664 15761 5692
rect 15620 5652 15626 5664
rect 15749 5661 15761 5664
rect 15795 5661 15807 5695
rect 15749 5655 15807 5661
rect 15838 5652 15844 5704
rect 15896 5692 15902 5704
rect 15896 5664 15941 5692
rect 15896 5652 15902 5664
rect 16390 5652 16396 5704
rect 16448 5692 16454 5704
rect 16853 5695 16911 5701
rect 16853 5692 16865 5695
rect 16448 5664 16865 5692
rect 16448 5652 16454 5664
rect 16853 5661 16865 5664
rect 16899 5661 16911 5695
rect 16853 5655 16911 5661
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5692 17279 5695
rect 17313 5695 17371 5701
rect 17313 5692 17325 5695
rect 17267 5664 17325 5692
rect 17267 5661 17279 5664
rect 17221 5655 17279 5661
rect 17313 5661 17325 5664
rect 17359 5661 17371 5695
rect 17313 5655 17371 5661
rect 18969 5695 19027 5701
rect 18969 5661 18981 5695
rect 19015 5692 19027 5695
rect 19426 5692 19432 5704
rect 19015 5664 19432 5692
rect 19015 5661 19027 5664
rect 18969 5655 19027 5661
rect 19426 5652 19432 5664
rect 19484 5652 19490 5704
rect 20070 5652 20076 5704
rect 20128 5692 20134 5704
rect 20349 5695 20407 5701
rect 20349 5692 20361 5695
rect 20128 5664 20361 5692
rect 20128 5652 20134 5664
rect 20349 5661 20361 5664
rect 20395 5661 20407 5695
rect 20349 5655 20407 5661
rect 12342 5624 12348 5636
rect 11256 5596 12348 5624
rect 9950 5516 9956 5568
rect 10008 5556 10014 5568
rect 11256 5556 11284 5596
rect 12342 5584 12348 5596
rect 12400 5584 12406 5636
rect 13906 5584 13912 5636
rect 13964 5624 13970 5636
rect 13964 5596 17356 5624
rect 13964 5584 13970 5596
rect 10008 5528 11284 5556
rect 11701 5559 11759 5565
rect 10008 5516 10014 5528
rect 11701 5525 11713 5559
rect 11747 5556 11759 5559
rect 11882 5556 11888 5568
rect 11747 5528 11888 5556
rect 11747 5525 11759 5528
rect 11701 5519 11759 5525
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 13078 5516 13084 5568
rect 13136 5556 13142 5568
rect 13817 5559 13875 5565
rect 13817 5556 13829 5559
rect 13136 5528 13829 5556
rect 13136 5516 13142 5528
rect 13817 5525 13829 5528
rect 13863 5525 13875 5559
rect 13817 5519 13875 5525
rect 16022 5516 16028 5568
rect 16080 5556 16086 5568
rect 16301 5559 16359 5565
rect 16301 5556 16313 5559
rect 16080 5528 16313 5556
rect 16080 5516 16086 5528
rect 16301 5525 16313 5528
rect 16347 5525 16359 5559
rect 16301 5519 16359 5525
rect 16574 5516 16580 5568
rect 16632 5556 16638 5568
rect 17221 5559 17279 5565
rect 17221 5556 17233 5559
rect 16632 5528 17233 5556
rect 16632 5516 16638 5528
rect 17221 5525 17233 5528
rect 17267 5525 17279 5559
rect 17328 5556 17356 5596
rect 17954 5556 17960 5568
rect 17328 5528 17960 5556
rect 17221 5519 17279 5525
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 19794 5556 19800 5568
rect 19755 5528 19800 5556
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 21085 5559 21143 5565
rect 21085 5525 21097 5559
rect 21131 5556 21143 5559
rect 22094 5556 22100 5568
rect 21131 5528 22100 5556
rect 21131 5525 21143 5528
rect 21085 5519 21143 5525
rect 22094 5516 22100 5528
rect 22152 5516 22158 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8389 5355 8447 5361
rect 8389 5352 8401 5355
rect 8352 5324 8401 5352
rect 8352 5312 8358 5324
rect 8389 5321 8401 5324
rect 8435 5352 8447 5355
rect 8754 5352 8760 5364
rect 8435 5324 8760 5352
rect 8435 5321 8447 5324
rect 8389 5315 8447 5321
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 9122 5352 9128 5364
rect 9083 5324 9128 5352
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 9585 5355 9643 5361
rect 9585 5321 9597 5355
rect 9631 5352 9643 5355
rect 9766 5352 9772 5364
rect 9631 5324 9772 5352
rect 9631 5321 9643 5324
rect 9585 5315 9643 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 9953 5355 10011 5361
rect 9953 5321 9965 5355
rect 9999 5352 10011 5355
rect 10502 5352 10508 5364
rect 9999 5324 10508 5352
rect 9999 5321 10011 5324
rect 9953 5315 10011 5321
rect 10502 5312 10508 5324
rect 10560 5352 10566 5364
rect 10560 5324 11744 5352
rect 10560 5312 10566 5324
rect 8849 5287 8907 5293
rect 8849 5253 8861 5287
rect 8895 5284 8907 5287
rect 9858 5284 9864 5296
rect 8895 5256 9864 5284
rect 8895 5253 8907 5256
rect 8849 5247 8907 5253
rect 9858 5244 9864 5256
rect 9916 5244 9922 5296
rect 10229 5287 10287 5293
rect 10229 5253 10241 5287
rect 10275 5284 10287 5287
rect 11606 5284 11612 5296
rect 10275 5256 11612 5284
rect 10275 5253 10287 5256
rect 10229 5247 10287 5253
rect 11606 5244 11612 5256
rect 11664 5244 11670 5296
rect 11716 5284 11744 5324
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 12437 5355 12495 5361
rect 12437 5352 12449 5355
rect 12032 5324 12449 5352
rect 12032 5312 12038 5324
rect 12437 5321 12449 5324
rect 12483 5321 12495 5355
rect 12986 5352 12992 5364
rect 12947 5324 12992 5352
rect 12437 5315 12495 5321
rect 12986 5312 12992 5324
rect 13044 5312 13050 5364
rect 14458 5312 14464 5364
rect 14516 5352 14522 5364
rect 15841 5355 15899 5361
rect 14516 5324 15424 5352
rect 14516 5312 14522 5324
rect 14366 5284 14372 5296
rect 11716 5256 14372 5284
rect 14366 5244 14372 5256
rect 14424 5244 14430 5296
rect 15396 5284 15424 5324
rect 15841 5321 15853 5355
rect 15887 5352 15899 5355
rect 16390 5352 16396 5364
rect 15887 5324 16396 5352
rect 15887 5321 15899 5324
rect 15841 5315 15899 5321
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 17862 5312 17868 5364
rect 17920 5352 17926 5364
rect 19429 5355 19487 5361
rect 19429 5352 19441 5355
rect 17920 5324 19441 5352
rect 17920 5312 17926 5324
rect 19429 5321 19441 5324
rect 19475 5321 19487 5355
rect 19429 5315 19487 5321
rect 16114 5284 16120 5296
rect 15396 5256 16120 5284
rect 16114 5244 16120 5256
rect 16172 5244 16178 5296
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5216 10931 5219
rect 11054 5216 11060 5228
rect 10919 5188 11060 5216
rect 10919 5185 10931 5188
rect 10873 5179 10931 5185
rect 11054 5176 11060 5188
rect 11112 5216 11118 5228
rect 11793 5219 11851 5225
rect 11793 5216 11805 5219
rect 11112 5188 11805 5216
rect 11112 5176 11118 5188
rect 11793 5185 11805 5188
rect 11839 5216 11851 5219
rect 11882 5216 11888 5228
rect 11839 5188 11888 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 13354 5176 13360 5228
rect 13412 5216 13418 5228
rect 13449 5219 13507 5225
rect 13449 5216 13461 5219
rect 13412 5188 13461 5216
rect 13412 5176 13418 5188
rect 13449 5185 13461 5188
rect 13495 5185 13507 5219
rect 13449 5179 13507 5185
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 13722 5216 13728 5228
rect 13679 5188 13728 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 13722 5176 13728 5188
rect 13780 5176 13786 5228
rect 17954 5176 17960 5228
rect 18012 5216 18018 5228
rect 19521 5219 19579 5225
rect 18012 5188 18184 5216
rect 18012 5176 18018 5188
rect 18156 5160 18184 5188
rect 19521 5185 19533 5219
rect 19567 5216 19579 5219
rect 19705 5219 19763 5225
rect 19705 5216 19717 5219
rect 19567 5188 19717 5216
rect 19567 5185 19579 5188
rect 19521 5179 19579 5185
rect 19705 5185 19717 5188
rect 19751 5185 19763 5219
rect 19705 5179 19763 5185
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 11609 5151 11667 5157
rect 11609 5148 11621 5151
rect 9824 5120 11621 5148
rect 9824 5108 9830 5120
rect 11609 5117 11621 5120
rect 11655 5117 11667 5151
rect 14458 5148 14464 5160
rect 11609 5111 11667 5117
rect 12912 5120 14228 5148
rect 14419 5120 14464 5148
rect 9306 5040 9312 5092
rect 9364 5080 9370 5092
rect 10502 5080 10508 5092
rect 9364 5052 10508 5080
rect 9364 5040 9370 5052
rect 10502 5040 10508 5052
rect 10560 5080 10566 5092
rect 10597 5083 10655 5089
rect 10597 5080 10609 5083
rect 10560 5052 10609 5080
rect 10560 5040 10566 5052
rect 10597 5049 10609 5052
rect 10643 5049 10655 5083
rect 10597 5043 10655 5049
rect 10689 5083 10747 5089
rect 10689 5049 10701 5083
rect 10735 5080 10747 5083
rect 11701 5083 11759 5089
rect 10735 5052 11652 5080
rect 10735 5049 10747 5052
rect 10689 5043 10747 5049
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 10962 5012 10968 5024
rect 9548 4984 10968 5012
rect 9548 4972 9554 4984
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11238 5012 11244 5024
rect 11199 4984 11244 5012
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 11624 5012 11652 5052
rect 11701 5049 11713 5083
rect 11747 5080 11759 5083
rect 12066 5080 12072 5092
rect 11747 5052 12072 5080
rect 11747 5049 11759 5052
rect 11701 5043 11759 5049
rect 12066 5040 12072 5052
rect 12124 5040 12130 5092
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 12526 5080 12532 5092
rect 12400 5052 12532 5080
rect 12400 5040 12406 5052
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 11974 5012 11980 5024
rect 11624 4984 11980 5012
rect 11974 4972 11980 4984
rect 12032 4972 12038 5024
rect 12084 5012 12112 5040
rect 12912 5012 12940 5120
rect 13357 5083 13415 5089
rect 13357 5049 13369 5083
rect 13403 5080 13415 5083
rect 13446 5080 13452 5092
rect 13403 5052 13452 5080
rect 13403 5049 13415 5052
rect 13357 5043 13415 5049
rect 13446 5040 13452 5052
rect 13504 5040 13510 5092
rect 12084 4984 12940 5012
rect 13262 4972 13268 5024
rect 13320 5012 13326 5024
rect 14090 5012 14096 5024
rect 13320 4984 14096 5012
rect 13320 4972 13326 4984
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14200 5012 14228 5120
rect 14458 5108 14464 5120
rect 14516 5148 14522 5160
rect 16390 5157 16396 5160
rect 16117 5151 16175 5157
rect 16117 5148 16129 5151
rect 14516 5120 16129 5148
rect 14516 5108 14522 5120
rect 16117 5117 16129 5120
rect 16163 5117 16175 5151
rect 16384 5148 16396 5157
rect 16351 5120 16396 5148
rect 16117 5111 16175 5117
rect 16384 5111 16396 5120
rect 14728 5083 14786 5089
rect 14728 5049 14740 5083
rect 14774 5080 14786 5083
rect 15838 5080 15844 5092
rect 14774 5052 15844 5080
rect 14774 5049 14786 5052
rect 14728 5043 14786 5049
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 16132 5080 16160 5111
rect 16390 5108 16396 5111
rect 16448 5108 16454 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 16592 5120 18061 5148
rect 16592 5092 16620 5120
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 16574 5080 16580 5092
rect 16132 5052 16580 5080
rect 16574 5040 16580 5052
rect 16632 5040 16638 5092
rect 17954 5080 17960 5092
rect 17328 5052 17960 5080
rect 17328 5012 17356 5052
rect 17954 5040 17960 5052
rect 18012 5040 18018 5092
rect 18064 5080 18092 5111
rect 18138 5108 18144 5160
rect 18196 5108 18202 5160
rect 18598 5148 18604 5160
rect 18248 5120 18604 5148
rect 18248 5080 18276 5120
rect 18598 5108 18604 5120
rect 18656 5108 18662 5160
rect 18874 5108 18880 5160
rect 18932 5148 18938 5160
rect 22646 5148 22652 5160
rect 18932 5120 22652 5148
rect 18932 5108 18938 5120
rect 22646 5108 22652 5120
rect 22704 5108 22710 5160
rect 18064 5052 18276 5080
rect 18316 5083 18374 5089
rect 18316 5049 18328 5083
rect 18362 5080 18374 5083
rect 19972 5083 20030 5089
rect 18362 5052 19656 5080
rect 18362 5049 18374 5052
rect 18316 5043 18374 5049
rect 19628 5024 19656 5052
rect 19972 5049 19984 5083
rect 20018 5080 20030 5083
rect 20070 5080 20076 5092
rect 20018 5052 20076 5080
rect 20018 5049 20030 5052
rect 19972 5043 20030 5049
rect 20070 5040 20076 5052
rect 20128 5040 20134 5092
rect 17494 5012 17500 5024
rect 14200 4984 17356 5012
rect 17455 4984 17500 5012
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 18598 4972 18604 5024
rect 18656 5012 18662 5024
rect 19521 5015 19579 5021
rect 19521 5012 19533 5015
rect 18656 4984 19533 5012
rect 18656 4972 18662 4984
rect 19521 4981 19533 4984
rect 19567 4981 19579 5015
rect 19521 4975 19579 4981
rect 19610 4972 19616 5024
rect 19668 5012 19674 5024
rect 21085 5015 21143 5021
rect 21085 5012 21097 5015
rect 19668 4984 21097 5012
rect 19668 4972 19674 4984
rect 21085 4981 21097 4984
rect 21131 4981 21143 5015
rect 21085 4975 21143 4981
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 10134 4808 10140 4820
rect 9692 4780 10140 4808
rect 9692 4681 9720 4780
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 18233 4811 18291 4817
rect 11716 4780 16988 4808
rect 9944 4743 10002 4749
rect 9944 4709 9956 4743
rect 9990 4740 10002 4743
rect 11054 4740 11060 4752
rect 9990 4712 11060 4740
rect 9990 4709 10002 4712
rect 9944 4703 10002 4709
rect 11054 4700 11060 4712
rect 11112 4700 11118 4752
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 10226 4672 10232 4684
rect 9677 4635 9735 4641
rect 9784 4644 10232 4672
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 9309 4607 9367 4613
rect 9309 4604 9321 4607
rect 8987 4576 9321 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 9309 4573 9321 4576
rect 9355 4604 9367 4607
rect 9784 4604 9812 4644
rect 10226 4632 10232 4644
rect 10284 4672 10290 4684
rect 11716 4681 11744 4780
rect 12526 4700 12532 4752
rect 12584 4740 12590 4752
rect 14737 4743 14795 4749
rect 12584 4712 13308 4740
rect 12584 4700 12590 4712
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 10284 4644 11713 4672
rect 10284 4632 10290 4644
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 11701 4635 11759 4641
rect 11974 4632 11980 4684
rect 12032 4672 12038 4684
rect 13153 4675 13211 4681
rect 13153 4672 13165 4675
rect 12032 4644 13165 4672
rect 12032 4632 12038 4644
rect 13153 4641 13165 4644
rect 13199 4641 13211 4675
rect 13280 4672 13308 4712
rect 14737 4709 14749 4743
rect 14783 4740 14795 4743
rect 16669 4743 16727 4749
rect 16669 4740 16681 4743
rect 14783 4712 16681 4740
rect 14783 4709 14795 4712
rect 14737 4703 14795 4709
rect 16669 4709 16681 4712
rect 16715 4709 16727 4743
rect 16669 4703 16727 4709
rect 16761 4743 16819 4749
rect 16761 4709 16773 4743
rect 16807 4740 16819 4743
rect 16850 4740 16856 4752
rect 16807 4712 16856 4740
rect 16807 4709 16819 4712
rect 16761 4703 16819 4709
rect 16850 4700 16856 4712
rect 16908 4700 16914 4752
rect 13630 4672 13636 4684
rect 13280 4644 13636 4672
rect 13153 4635 13211 4641
rect 13630 4632 13636 4644
rect 13688 4672 13694 4684
rect 15470 4672 15476 4684
rect 13688 4644 15476 4672
rect 13688 4632 13694 4644
rect 15470 4632 15476 4644
rect 15528 4632 15534 4684
rect 15654 4672 15660 4684
rect 15615 4644 15660 4672
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 15749 4675 15807 4681
rect 15749 4641 15761 4675
rect 15795 4672 15807 4675
rect 15795 4644 16068 4672
rect 15795 4641 15807 4644
rect 15749 4635 15807 4641
rect 9355 4576 9812 4604
rect 11793 4607 11851 4613
rect 9355 4573 9367 4576
rect 9309 4567 9367 4573
rect 11793 4573 11805 4607
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 10778 4496 10784 4548
rect 10836 4536 10842 4548
rect 11808 4536 11836 4567
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 11940 4576 11985 4604
rect 11940 4564 11946 4576
rect 12066 4564 12072 4616
rect 12124 4604 12130 4616
rect 12345 4607 12403 4613
rect 12345 4604 12357 4607
rect 12124 4576 12357 4604
rect 12124 4564 12130 4576
rect 12345 4573 12357 4576
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12894 4604 12900 4616
rect 12492 4576 12900 4604
rect 12492 4564 12498 4576
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 14090 4564 14096 4616
rect 14148 4604 14154 4616
rect 15764 4604 15792 4635
rect 14148 4576 15792 4604
rect 14148 4564 14154 4576
rect 15838 4564 15844 4616
rect 15896 4604 15902 4616
rect 16040 4604 16068 4644
rect 16390 4632 16396 4684
rect 16448 4672 16454 4684
rect 16448 4644 16896 4672
rect 16448 4632 16454 4644
rect 16868 4613 16896 4644
rect 16853 4607 16911 4613
rect 15896 4576 15941 4604
rect 16040 4576 16804 4604
rect 15896 4564 15902 4576
rect 14277 4539 14335 4545
rect 10836 4508 11928 4536
rect 10836 4496 10842 4508
rect 8573 4471 8631 4477
rect 8573 4437 8585 4471
rect 8619 4468 8631 4471
rect 9582 4468 9588 4480
rect 8619 4440 9588 4468
rect 8619 4437 8631 4440
rect 8573 4431 8631 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 11054 4468 11060 4480
rect 11015 4440 11060 4468
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 11146 4428 11152 4480
rect 11204 4468 11210 4480
rect 11333 4471 11391 4477
rect 11333 4468 11345 4471
rect 11204 4440 11345 4468
rect 11204 4428 11210 4440
rect 11333 4437 11345 4440
rect 11379 4437 11391 4471
rect 11900 4468 11928 4508
rect 14277 4505 14289 4539
rect 14323 4536 14335 4539
rect 15856 4536 15884 4564
rect 16666 4536 16672 4548
rect 14323 4508 15884 4536
rect 15948 4508 16672 4536
rect 14323 4505 14335 4508
rect 14277 4499 14335 4505
rect 12618 4468 12624 4480
rect 11900 4440 12624 4468
rect 11333 4431 11391 4437
rect 12618 4428 12624 4440
rect 12676 4468 12682 4480
rect 13630 4468 13636 4480
rect 12676 4440 13636 4468
rect 12676 4428 12682 4440
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 14090 4428 14096 4480
rect 14148 4468 14154 4480
rect 14734 4468 14740 4480
rect 14148 4440 14740 4468
rect 14148 4428 14154 4440
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 15289 4471 15347 4477
rect 15289 4437 15301 4471
rect 15335 4468 15347 4471
rect 15948 4468 15976 4508
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 15335 4440 15976 4468
rect 15335 4437 15347 4440
rect 15289 4431 15347 4437
rect 16114 4428 16120 4480
rect 16172 4468 16178 4480
rect 16301 4471 16359 4477
rect 16301 4468 16313 4471
rect 16172 4440 16313 4468
rect 16172 4428 16178 4440
rect 16301 4437 16313 4440
rect 16347 4437 16359 4471
rect 16776 4468 16804 4576
rect 16853 4573 16865 4607
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 16960 4536 16988 4780
rect 18233 4777 18245 4811
rect 18279 4808 18291 4811
rect 18874 4808 18880 4820
rect 18279 4780 18880 4808
rect 18279 4777 18291 4780
rect 18233 4771 18291 4777
rect 18874 4768 18880 4780
rect 18932 4768 18938 4820
rect 18969 4811 19027 4817
rect 18969 4777 18981 4811
rect 19015 4808 19027 4811
rect 19702 4808 19708 4820
rect 19015 4780 19708 4808
rect 19015 4777 19027 4780
rect 18969 4771 19027 4777
rect 19702 4768 19708 4780
rect 19760 4768 19766 4820
rect 19794 4768 19800 4820
rect 19852 4808 19858 4820
rect 20073 4811 20131 4817
rect 20073 4808 20085 4811
rect 19852 4780 20085 4808
rect 19852 4768 19858 4780
rect 20073 4777 20085 4780
rect 20119 4777 20131 4811
rect 20073 4771 20131 4777
rect 19518 4700 19524 4752
rect 19576 4740 19582 4752
rect 19981 4743 20039 4749
rect 19981 4740 19993 4743
rect 19576 4712 19993 4740
rect 19576 4700 19582 4712
rect 19981 4709 19993 4712
rect 20027 4709 20039 4743
rect 19981 4703 20039 4709
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4672 18107 4675
rect 18138 4672 18144 4684
rect 18095 4644 18144 4672
rect 18095 4641 18107 4644
rect 18049 4635 18107 4641
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 18230 4632 18236 4684
rect 18288 4672 18294 4684
rect 18874 4672 18880 4684
rect 18288 4644 18880 4672
rect 18288 4632 18294 4644
rect 18874 4632 18880 4644
rect 18932 4632 18938 4684
rect 19061 4675 19119 4681
rect 19061 4641 19073 4675
rect 19107 4672 19119 4675
rect 19886 4672 19892 4684
rect 19107 4644 19892 4672
rect 19107 4641 19119 4644
rect 19061 4635 19119 4641
rect 19886 4632 19892 4644
rect 19944 4632 19950 4684
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4641 20959 4675
rect 20901 4635 20959 4641
rect 17310 4604 17316 4616
rect 17271 4576 17316 4604
rect 17310 4564 17316 4576
rect 17368 4564 17374 4616
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4604 19303 4607
rect 19610 4604 19616 4616
rect 19291 4576 19616 4604
rect 19291 4573 19303 4576
rect 19245 4567 19303 4573
rect 19610 4564 19616 4576
rect 19668 4564 19674 4616
rect 19702 4564 19708 4616
rect 19760 4604 19766 4616
rect 19978 4604 19984 4616
rect 19760 4576 19984 4604
rect 19760 4564 19766 4576
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 20257 4607 20315 4613
rect 20257 4573 20269 4607
rect 20303 4604 20315 4607
rect 20530 4604 20536 4616
rect 20303 4576 20536 4604
rect 20303 4573 20315 4576
rect 20257 4567 20315 4573
rect 20530 4564 20536 4576
rect 20588 4564 20594 4616
rect 20916 4536 20944 4635
rect 16960 4508 20944 4536
rect 17954 4468 17960 4480
rect 16776 4440 17960 4468
rect 16301 4431 16359 4437
rect 17954 4428 17960 4440
rect 18012 4428 18018 4480
rect 18601 4471 18659 4477
rect 18601 4437 18613 4471
rect 18647 4468 18659 4471
rect 19518 4468 19524 4480
rect 18647 4440 19524 4468
rect 18647 4437 18659 4440
rect 18601 4431 18659 4437
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 19613 4471 19671 4477
rect 19613 4437 19625 4471
rect 19659 4468 19671 4471
rect 19978 4468 19984 4480
rect 19659 4440 19984 4468
rect 19659 4437 19671 4440
rect 19613 4431 19671 4437
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 21542 4468 21548 4480
rect 21131 4440 21548 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 8849 4267 8907 4273
rect 8849 4264 8861 4267
rect 7156 4236 8861 4264
rect 7156 4224 7162 4236
rect 8849 4233 8861 4236
rect 8895 4233 8907 4267
rect 8849 4227 8907 4233
rect 9309 4267 9367 4273
rect 9309 4233 9321 4267
rect 9355 4264 9367 4267
rect 9858 4264 9864 4276
rect 9355 4236 9864 4264
rect 9355 4233 9367 4236
rect 9309 4227 9367 4233
rect 8864 4196 8892 4227
rect 9858 4224 9864 4236
rect 9916 4224 9922 4276
rect 11974 4264 11980 4276
rect 10244 4236 11980 4264
rect 10042 4196 10048 4208
rect 8864 4168 10048 4196
rect 10042 4156 10048 4168
rect 10100 4156 10106 4208
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 7374 4128 7380 4140
rect 4212 4100 7380 4128
rect 4212 4088 4218 4100
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 8938 4128 8944 4140
rect 7616 4100 8944 4128
rect 7616 4088 7622 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 10244 4137 10272 4236
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 17954 4224 17960 4276
rect 18012 4264 18018 4276
rect 18966 4264 18972 4276
rect 18012 4236 18972 4264
rect 18012 4224 18018 4236
rect 18966 4224 18972 4236
rect 19024 4224 19030 4276
rect 19886 4224 19892 4276
rect 19944 4264 19950 4276
rect 20257 4267 20315 4273
rect 20257 4264 20269 4267
rect 19944 4236 20269 4264
rect 19944 4224 19950 4236
rect 20257 4233 20269 4236
rect 20303 4233 20315 4267
rect 20257 4227 20315 4233
rect 17494 4196 17500 4208
rect 16224 4168 17500 4196
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 13170 4128 13176 4140
rect 13044 4100 13176 4128
rect 13044 4088 13050 4100
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 16022 4128 16028 4140
rect 15983 4100 16028 4128
rect 16022 4088 16028 4100
rect 16080 4088 16086 4140
rect 16224 4137 16252 4168
rect 17494 4156 17500 4168
rect 17552 4156 17558 4208
rect 19981 4199 20039 4205
rect 19981 4165 19993 4199
rect 20027 4196 20039 4199
rect 20070 4196 20076 4208
rect 20027 4168 20076 4196
rect 20027 4165 20039 4168
rect 19981 4159 20039 4165
rect 20070 4156 20076 4168
rect 20128 4156 20134 4208
rect 16209 4131 16267 4137
rect 16209 4097 16221 4131
rect 16255 4097 16267 4131
rect 20088 4128 20116 4156
rect 20809 4131 20867 4137
rect 20809 4128 20821 4131
rect 20088 4100 20821 4128
rect 16209 4091 16267 4097
rect 20809 4097 20821 4100
rect 20855 4097 20867 4131
rect 20809 4091 20867 4097
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 8478 4060 8484 4072
rect 5868 4032 8484 4060
rect 5868 4020 5874 4032
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 10192 4032 10609 4060
rect 10192 4020 10198 4032
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 12526 4060 12532 4072
rect 10597 4023 10655 4029
rect 10796 4032 11744 4060
rect 12487 4032 12532 4060
rect 3050 3952 3056 4004
rect 3108 3992 3114 4004
rect 7650 3992 7656 4004
rect 3108 3964 7656 3992
rect 3108 3952 3114 3964
rect 7650 3952 7656 3964
rect 7708 3952 7714 4004
rect 7742 3952 7748 4004
rect 7800 3992 7806 4004
rect 8202 3992 8208 4004
rect 7800 3964 8208 3992
rect 7800 3952 7806 3964
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 8573 3995 8631 4001
rect 8573 3961 8585 3995
rect 8619 3992 8631 3995
rect 10796 3992 10824 4032
rect 8619 3964 10824 3992
rect 10864 3995 10922 4001
rect 8619 3961 8631 3964
rect 8573 3955 8631 3961
rect 10864 3961 10876 3995
rect 10910 3992 10922 3995
rect 11054 3992 11060 4004
rect 10910 3964 11060 3992
rect 10910 3961 10922 3964
rect 10864 3955 10922 3961
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 11146 3952 11152 4004
rect 11204 3992 11210 4004
rect 11514 3992 11520 4004
rect 11204 3964 11520 3992
rect 11204 3952 11210 3964
rect 11514 3952 11520 3964
rect 11572 3952 11578 4004
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 7190 3924 7196 3936
rect 2004 3896 7196 3924
rect 2004 3884 2010 3896
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 9585 3927 9643 3933
rect 9585 3893 9597 3927
rect 9631 3924 9643 3927
rect 9766 3924 9772 3936
rect 9631 3896 9772 3924
rect 9631 3893 9643 3896
rect 9585 3887 9643 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 9950 3924 9956 3936
rect 9911 3896 9956 3924
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 10594 3924 10600 3936
rect 10091 3896 10600 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11716 3924 11744 4032
rect 12526 4020 12532 4032
rect 12584 4020 12590 4072
rect 12894 4020 12900 4072
rect 12952 4060 12958 4072
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 12952 4032 13277 4060
rect 12952 4020 12958 4032
rect 13265 4029 13277 4032
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 14921 4063 14979 4069
rect 14921 4060 14933 4063
rect 13872 4032 14933 4060
rect 13872 4020 13878 4032
rect 14921 4029 14933 4032
rect 14967 4029 14979 4063
rect 14921 4023 14979 4029
rect 15933 4063 15991 4069
rect 15933 4029 15945 4063
rect 15979 4060 15991 4063
rect 16114 4060 16120 4072
rect 15979 4032 16120 4060
rect 15979 4029 15991 4032
rect 15933 4023 15991 4029
rect 16114 4020 16120 4032
rect 16172 4020 16178 4072
rect 16577 4063 16635 4069
rect 16577 4060 16589 4063
rect 16224 4032 16589 4060
rect 13446 3952 13452 4004
rect 13504 4001 13510 4004
rect 13504 3995 13568 4001
rect 13504 3961 13522 3995
rect 13556 3961 13568 3995
rect 13504 3955 13568 3961
rect 13504 3952 13510 3955
rect 13630 3952 13636 4004
rect 13688 3992 13694 4004
rect 16224 3992 16252 4032
rect 16577 4029 16589 4032
rect 16623 4029 16635 4063
rect 17126 4060 17132 4072
rect 17087 4032 17132 4060
rect 16577 4023 16635 4029
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 17954 4020 17960 4072
rect 18012 4060 18018 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 18012 4032 18061 4060
rect 18012 4020 18018 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 18138 4020 18144 4072
rect 18196 4060 18202 4072
rect 18601 4063 18659 4069
rect 18601 4060 18613 4063
rect 18196 4032 18613 4060
rect 18196 4020 18202 4032
rect 18601 4029 18613 4032
rect 18647 4029 18659 4063
rect 18601 4023 18659 4029
rect 18690 4020 18696 4072
rect 18748 4060 18754 4072
rect 21266 4060 21272 4072
rect 18748 4032 21272 4060
rect 18748 4020 18754 4032
rect 21266 4020 21272 4032
rect 21324 4020 21330 4072
rect 13688 3964 16252 3992
rect 13688 3952 13694 3964
rect 16390 3952 16396 4004
rect 16448 3992 16454 4004
rect 16448 3964 17356 3992
rect 16448 3952 16454 3964
rect 12434 3924 12440 3936
rect 11716 3896 12440 3924
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 12713 3927 12771 3933
rect 12713 3924 12725 3927
rect 12676 3896 12725 3924
rect 12676 3884 12682 3896
rect 12713 3893 12725 3896
rect 12759 3893 12771 3927
rect 12713 3887 12771 3893
rect 14645 3927 14703 3933
rect 14645 3893 14657 3927
rect 14691 3924 14703 3927
rect 14734 3924 14740 3936
rect 14691 3896 14740 3924
rect 14691 3893 14703 3896
rect 14645 3887 14703 3893
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 15105 3927 15163 3933
rect 15105 3893 15117 3927
rect 15151 3924 15163 3927
rect 15378 3924 15384 3936
rect 15151 3896 15384 3924
rect 15151 3893 15163 3896
rect 15105 3887 15163 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 15565 3927 15623 3933
rect 15565 3893 15577 3927
rect 15611 3924 15623 3927
rect 15746 3924 15752 3936
rect 15611 3896 15752 3924
rect 15611 3893 15623 3896
rect 15565 3887 15623 3893
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 15930 3884 15936 3936
rect 15988 3924 15994 3936
rect 17328 3933 17356 3964
rect 17402 3952 17408 4004
rect 17460 3992 17466 4004
rect 18868 3995 18926 4001
rect 17460 3964 18368 3992
rect 17460 3952 17466 3964
rect 16761 3927 16819 3933
rect 16761 3924 16773 3927
rect 15988 3896 16773 3924
rect 15988 3884 15994 3896
rect 16761 3893 16773 3896
rect 16807 3893 16819 3927
rect 16761 3887 16819 3893
rect 17313 3927 17371 3933
rect 17313 3893 17325 3927
rect 17359 3893 17371 3927
rect 17313 3887 17371 3893
rect 17678 3884 17684 3936
rect 17736 3924 17742 3936
rect 18233 3927 18291 3933
rect 18233 3924 18245 3927
rect 17736 3896 18245 3924
rect 17736 3884 17742 3896
rect 18233 3893 18245 3896
rect 18279 3893 18291 3927
rect 18340 3924 18368 3964
rect 18868 3961 18880 3995
rect 18914 3992 18926 3995
rect 19702 3992 19708 4004
rect 18914 3964 19708 3992
rect 18914 3961 18926 3964
rect 18868 3955 18926 3961
rect 19702 3952 19708 3964
rect 19760 3952 19766 4004
rect 20625 3927 20683 3933
rect 20625 3924 20637 3927
rect 18340 3896 20637 3924
rect 18233 3887 18291 3893
rect 20625 3893 20637 3896
rect 20671 3893 20683 3927
rect 20625 3887 20683 3893
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 20772 3896 20817 3924
rect 20772 3884 20778 3896
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 5258 3680 5264 3732
rect 5316 3720 5322 3732
rect 8662 3720 8668 3732
rect 5316 3692 8668 3720
rect 5316 3680 5322 3692
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 9309 3723 9367 3729
rect 9309 3689 9321 3723
rect 9355 3720 9367 3723
rect 9398 3720 9404 3732
rect 9355 3692 9404 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 10045 3723 10103 3729
rect 10045 3720 10057 3723
rect 9916 3692 10057 3720
rect 9916 3680 9922 3692
rect 10045 3689 10057 3692
rect 10091 3689 10103 3723
rect 10045 3683 10103 3689
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 10781 3723 10839 3729
rect 10781 3720 10793 3723
rect 10652 3692 10793 3720
rect 10652 3680 10658 3692
rect 10781 3689 10793 3692
rect 10827 3689 10839 3723
rect 12894 3720 12900 3732
rect 10781 3683 10839 3689
rect 12084 3692 12900 3720
rect 6454 3612 6460 3664
rect 6512 3652 6518 3664
rect 11974 3652 11980 3664
rect 6512 3624 11980 3652
rect 6512 3612 6518 3624
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 3602 3544 3608 3596
rect 3660 3584 3666 3596
rect 6914 3584 6920 3596
rect 3660 3556 6920 3584
rect 3660 3544 3666 3556
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 7006 3544 7012 3596
rect 7064 3584 7070 3596
rect 10686 3584 10692 3596
rect 7064 3556 10692 3584
rect 7064 3544 7070 3556
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 11146 3584 11152 3596
rect 11107 3556 11152 3584
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3584 11299 3587
rect 11514 3584 11520 3596
rect 11287 3556 11520 3584
rect 11287 3553 11299 3556
rect 11241 3547 11299 3553
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 12084 3593 12112 3692
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 14185 3723 14243 3729
rect 14185 3689 14197 3723
rect 14231 3720 14243 3723
rect 14274 3720 14280 3732
rect 14231 3692 14280 3720
rect 14231 3689 14243 3692
rect 14185 3683 14243 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 17402 3720 17408 3732
rect 15580 3692 17408 3720
rect 12158 3612 12164 3664
rect 12216 3652 12222 3664
rect 12314 3655 12372 3661
rect 12314 3652 12326 3655
rect 12216 3624 12326 3652
rect 12216 3612 12222 3624
rect 12314 3621 12326 3624
rect 12360 3621 12372 3655
rect 13906 3652 13912 3664
rect 13819 3624 13912 3652
rect 12314 3615 12372 3621
rect 13906 3612 13912 3624
rect 13964 3652 13970 3664
rect 15580 3652 15608 3692
rect 17402 3680 17408 3692
rect 17460 3680 17466 3732
rect 18049 3723 18107 3729
rect 18049 3689 18061 3723
rect 18095 3689 18107 3723
rect 19702 3720 19708 3732
rect 19663 3692 19708 3720
rect 18049 3683 18107 3689
rect 13964 3624 15608 3652
rect 16025 3655 16083 3661
rect 13964 3612 13970 3624
rect 16025 3621 16037 3655
rect 16071 3652 16083 3655
rect 17126 3652 17132 3664
rect 16071 3624 17132 3652
rect 16071 3621 16083 3624
rect 16025 3615 16083 3621
rect 17126 3612 17132 3624
rect 17184 3612 17190 3664
rect 18064 3652 18092 3683
rect 19702 3680 19708 3692
rect 19760 3680 19766 3732
rect 18598 3661 18604 3664
rect 18570 3655 18604 3661
rect 18570 3652 18582 3655
rect 18064 3624 18582 3652
rect 18570 3621 18582 3624
rect 18656 3652 18662 3664
rect 18656 3624 18718 3652
rect 18570 3615 18604 3621
rect 18598 3612 18604 3615
rect 18656 3612 18662 3624
rect 12069 3587 12127 3593
rect 12069 3553 12081 3587
rect 12115 3553 12127 3587
rect 12069 3547 12127 3553
rect 14553 3587 14611 3593
rect 14553 3553 14565 3587
rect 14599 3584 14611 3587
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 14599 3556 15301 3584
rect 14599 3553 14611 3556
rect 14553 3547 14611 3553
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 15746 3584 15752 3596
rect 15707 3556 15752 3584
rect 15289 3547 15347 3553
rect 15746 3544 15752 3556
rect 15804 3544 15810 3596
rect 16936 3587 16994 3593
rect 16936 3553 16948 3587
rect 16982 3584 16994 3587
rect 17494 3584 17500 3596
rect 16982 3556 17500 3584
rect 16982 3553 16994 3556
rect 16936 3547 16994 3553
rect 17494 3544 17500 3556
rect 17552 3544 17558 3596
rect 19978 3584 19984 3596
rect 19939 3556 19984 3584
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 20438 3544 20444 3596
rect 20496 3584 20502 3596
rect 20901 3587 20959 3593
rect 20901 3584 20913 3587
rect 20496 3556 20913 3584
rect 20496 3544 20502 3556
rect 20901 3553 20913 3556
rect 20947 3553 20959 3587
rect 20901 3547 20959 3553
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3516 9827 3519
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9815 3488 9873 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 9861 3485 9873 3488
rect 9907 3516 9919 3519
rect 10778 3516 10784 3528
rect 9907 3488 10784 3516
rect 9907 3485 9919 3488
rect 9861 3479 9919 3485
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 11330 3516 11336 3528
rect 11291 3488 11336 3516
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 14642 3516 14648 3528
rect 14603 3488 14648 3516
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 16666 3516 16672 3528
rect 14792 3488 14837 3516
rect 16627 3488 16672 3516
rect 14792 3476 14798 3488
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 18138 3476 18144 3528
rect 18196 3516 18202 3528
rect 18325 3519 18383 3525
rect 18325 3516 18337 3519
rect 18196 3488 18337 3516
rect 18196 3476 18202 3488
rect 18325 3485 18337 3488
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 20165 3519 20223 3525
rect 20165 3516 20177 3519
rect 19576 3488 20177 3516
rect 19576 3476 19582 3488
rect 20165 3485 20177 3488
rect 20211 3485 20223 3519
rect 20165 3479 20223 3485
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 8720 3420 12112 3448
rect 8720 3408 8726 3420
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 9861 3383 9919 3389
rect 9861 3380 9873 3383
rect 9640 3352 9873 3380
rect 9640 3340 9646 3352
rect 9861 3349 9873 3352
rect 9907 3349 9919 3383
rect 10502 3380 10508 3392
rect 10463 3352 10508 3380
rect 9861 3343 9919 3349
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 11974 3380 11980 3392
rect 11204 3352 11980 3380
rect 11204 3340 11210 3352
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 12084 3380 12112 3420
rect 13722 3408 13728 3460
rect 13780 3448 13786 3460
rect 15838 3448 15844 3460
rect 13780 3420 15844 3448
rect 13780 3408 13786 3420
rect 15838 3408 15844 3420
rect 15896 3408 15902 3460
rect 12986 3380 12992 3392
rect 12084 3352 12992 3380
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 13446 3380 13452 3392
rect 13407 3352 13452 3380
rect 13446 3340 13452 3352
rect 13504 3340 13510 3392
rect 20990 3340 20996 3392
rect 21048 3380 21054 3392
rect 21085 3383 21143 3389
rect 21085 3380 21097 3383
rect 21048 3352 21097 3380
rect 21048 3340 21054 3352
rect 21085 3349 21097 3352
rect 21131 3349 21143 3383
rect 21085 3343 21143 3349
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 9217 3179 9275 3185
rect 9217 3145 9229 3179
rect 9263 3176 9275 3179
rect 9674 3176 9680 3188
rect 9263 3148 9680 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 9674 3136 9680 3148
rect 9732 3176 9738 3188
rect 9858 3176 9864 3188
rect 9732 3148 9864 3176
rect 9732 3136 9738 3148
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 10008 3148 10793 3176
rect 10008 3136 10014 3148
rect 10781 3145 10793 3148
rect 10827 3145 10839 3179
rect 10781 3139 10839 3145
rect 13449 3179 13507 3185
rect 13449 3145 13461 3179
rect 13495 3176 13507 3179
rect 14642 3176 14648 3188
rect 13495 3148 14648 3176
rect 13495 3145 13507 3148
rect 13449 3139 13507 3145
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 17494 3176 17500 3188
rect 17455 3148 17500 3176
rect 17494 3136 17500 3148
rect 17552 3136 17558 3188
rect 18782 3136 18788 3188
rect 18840 3176 18846 3188
rect 19061 3179 19119 3185
rect 19061 3176 19073 3179
rect 18840 3148 19073 3176
rect 18840 3136 18846 3148
rect 19061 3145 19073 3148
rect 19107 3145 19119 3179
rect 19061 3139 19119 3145
rect 2498 3068 2504 3120
rect 2556 3108 2562 3120
rect 10226 3108 10232 3120
rect 2556 3080 10232 3108
rect 2556 3068 2562 3080
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 10413 3111 10471 3117
rect 10413 3077 10425 3111
rect 10459 3108 10471 3111
rect 10686 3108 10692 3120
rect 10459 3080 10692 3108
rect 10459 3077 10471 3080
rect 10413 3071 10471 3077
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 12253 3111 12311 3117
rect 12253 3108 12265 3111
rect 10980 3080 12265 3108
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 9674 3040 9680 3052
rect 1452 3012 9680 3040
rect 1452 3000 1458 3012
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3040 10011 3043
rect 10980 3040 11008 3080
rect 12253 3077 12265 3080
rect 12299 3077 12311 3111
rect 12253 3071 12311 3077
rect 9999 3012 11008 3040
rect 9999 3009 10011 3012
rect 9953 3003 10011 3009
rect 4798 2932 4804 2984
rect 4856 2972 4862 2984
rect 9968 2972 9996 3003
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11333 3043 11391 3049
rect 11333 3040 11345 3043
rect 11112 3012 11345 3040
rect 11112 3000 11118 3012
rect 11333 3009 11345 3012
rect 11379 3009 11391 3043
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 11333 3003 11391 3009
rect 11808 3012 12725 3040
rect 4856 2944 9996 2972
rect 10229 2975 10287 2981
rect 4856 2932 4862 2944
rect 10229 2941 10241 2975
rect 10275 2972 10287 2975
rect 11422 2972 11428 2984
rect 10275 2944 11428 2972
rect 10275 2941 10287 2944
rect 10229 2935 10287 2941
rect 11422 2932 11428 2944
rect 11480 2932 11486 2984
rect 11808 2981 11836 3012
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 12713 3003 12771 3009
rect 13446 3000 13452 3052
rect 13504 3040 13510 3052
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13504 3012 14013 3040
rect 13504 3000 13510 3012
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 18598 3040 18604 3052
rect 18559 3012 18604 3040
rect 14001 3003 14059 3009
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 19702 3040 19708 3052
rect 19392 3012 19564 3040
rect 19663 3012 19708 3040
rect 19392 3000 19398 3012
rect 11793 2975 11851 2981
rect 11793 2941 11805 2975
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 12529 2975 12587 2981
rect 12529 2941 12541 2975
rect 12575 2972 12587 2975
rect 13538 2972 13544 2984
rect 12575 2944 13544 2972
rect 12575 2941 12587 2944
rect 12529 2935 12587 2941
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 14458 2972 14464 2984
rect 14371 2944 14464 2972
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 14734 2981 14740 2984
rect 14728 2972 14740 2981
rect 14695 2944 14740 2972
rect 14728 2935 14740 2944
rect 14734 2932 14740 2935
rect 14792 2932 14798 2984
rect 16117 2975 16175 2981
rect 16117 2972 16129 2975
rect 15764 2944 16129 2972
rect 8849 2907 8907 2913
rect 8849 2873 8861 2907
rect 8895 2904 8907 2907
rect 12253 2907 12311 2913
rect 8895 2876 12204 2904
rect 8895 2873 8907 2876
rect 8849 2867 8907 2873
rect 290 2796 296 2848
rect 348 2836 354 2848
rect 9306 2836 9312 2848
rect 348 2808 9312 2836
rect 348 2796 354 2808
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 9490 2836 9496 2848
rect 9451 2808 9496 2836
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 10962 2836 10968 2848
rect 9732 2808 10968 2836
rect 9732 2796 9738 2808
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11146 2836 11152 2848
rect 11107 2808 11152 2836
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 11241 2839 11299 2845
rect 11241 2805 11253 2839
rect 11287 2836 11299 2839
rect 11698 2836 11704 2848
rect 11287 2808 11704 2836
rect 11287 2805 11299 2808
rect 11241 2799 11299 2805
rect 11698 2796 11704 2808
rect 11756 2796 11762 2848
rect 11977 2839 12035 2845
rect 11977 2805 11989 2839
rect 12023 2836 12035 2839
rect 12066 2836 12072 2848
rect 12023 2808 12072 2836
rect 12023 2805 12035 2808
rect 11977 2799 12035 2805
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 12176 2836 12204 2876
rect 12253 2873 12265 2907
rect 12299 2904 12311 2907
rect 13817 2907 13875 2913
rect 13817 2904 13829 2907
rect 12299 2876 13829 2904
rect 12299 2873 12311 2876
rect 12253 2867 12311 2873
rect 13817 2873 13829 2876
rect 13863 2873 13875 2907
rect 14476 2904 14504 2932
rect 15764 2904 15792 2944
rect 16117 2941 16129 2944
rect 16163 2972 16175 2975
rect 16666 2972 16672 2984
rect 16163 2944 16672 2972
rect 16163 2941 16175 2944
rect 16117 2935 16175 2941
rect 16666 2932 16672 2944
rect 16724 2972 16730 2984
rect 18138 2972 18144 2984
rect 16724 2944 18144 2972
rect 16724 2932 16730 2944
rect 18138 2932 18144 2944
rect 18196 2932 18202 2984
rect 18414 2972 18420 2984
rect 18375 2944 18420 2972
rect 18414 2932 18420 2944
rect 18472 2932 18478 2984
rect 19426 2972 19432 2984
rect 19387 2944 19432 2972
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 19536 2972 19564 3012
rect 19702 3000 19708 3012
rect 19760 3000 19766 3052
rect 20438 3040 20444 3052
rect 20399 3012 20444 3040
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 20165 2975 20223 2981
rect 20165 2972 20177 2975
rect 19536 2944 20177 2972
rect 20165 2941 20177 2944
rect 20211 2941 20223 2975
rect 20898 2972 20904 2984
rect 20859 2944 20904 2972
rect 20165 2935 20223 2941
rect 20898 2932 20904 2944
rect 20956 2932 20962 2984
rect 16362 2907 16420 2913
rect 16362 2904 16374 2907
rect 14476 2876 15792 2904
rect 15856 2876 16374 2904
rect 13817 2867 13875 2873
rect 13909 2839 13967 2845
rect 13909 2836 13921 2839
rect 12176 2808 13921 2836
rect 13909 2805 13921 2808
rect 13955 2836 13967 2839
rect 14182 2836 14188 2848
rect 13955 2808 14188 2836
rect 13955 2805 13967 2808
rect 13909 2799 13967 2805
rect 14182 2796 14188 2808
rect 14240 2796 14246 2848
rect 15856 2845 15884 2876
rect 16362 2873 16374 2876
rect 16408 2904 16420 2907
rect 16482 2904 16488 2916
rect 16408 2876 16488 2904
rect 16408 2873 16420 2876
rect 16362 2867 16420 2873
rect 16482 2864 16488 2876
rect 16540 2864 16546 2916
rect 19521 2907 19579 2913
rect 19521 2904 19533 2907
rect 18064 2876 19533 2904
rect 18064 2845 18092 2876
rect 19521 2873 19533 2876
rect 19567 2873 19579 2907
rect 19521 2867 19579 2873
rect 15841 2839 15899 2845
rect 15841 2805 15853 2839
rect 15887 2805 15899 2839
rect 15841 2799 15899 2805
rect 18049 2839 18107 2845
rect 18049 2805 18061 2839
rect 18095 2805 18107 2839
rect 18049 2799 18107 2805
rect 18138 2796 18144 2848
rect 18196 2836 18202 2848
rect 18509 2839 18567 2845
rect 18509 2836 18521 2839
rect 18196 2808 18521 2836
rect 18196 2796 18202 2808
rect 18509 2805 18521 2808
rect 18555 2805 18567 2839
rect 18509 2799 18567 2805
rect 19886 2796 19892 2848
rect 19944 2836 19950 2848
rect 21085 2839 21143 2845
rect 21085 2836 21097 2839
rect 19944 2808 21097 2836
rect 19944 2796 19950 2808
rect 21085 2805 21097 2808
rect 21131 2805 21143 2839
rect 21085 2799 21143 2805
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 7282 2592 7288 2644
rect 7340 2632 7346 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 7340 2604 8953 2632
rect 7340 2592 7346 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 8956 2360 8984 2595
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10505 2635 10563 2641
rect 10505 2632 10517 2635
rect 10284 2604 10517 2632
rect 10284 2592 10290 2604
rect 10505 2601 10517 2604
rect 10551 2632 10563 2635
rect 16301 2635 16359 2641
rect 16301 2632 16313 2635
rect 10551 2604 16313 2632
rect 10551 2601 10563 2604
rect 10505 2595 10563 2601
rect 16301 2601 16313 2604
rect 16347 2601 16359 2635
rect 16942 2632 16948 2644
rect 16903 2604 16948 2632
rect 16301 2595 16359 2601
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 17310 2632 17316 2644
rect 17271 2604 17316 2632
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 21266 2632 21272 2644
rect 21227 2604 21272 2632
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 10873 2567 10931 2573
rect 10873 2533 10885 2567
rect 10919 2564 10931 2567
rect 10962 2564 10968 2576
rect 10919 2536 10968 2564
rect 10919 2533 10931 2536
rect 10873 2527 10931 2533
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 11422 2564 11428 2576
rect 11383 2536 11428 2564
rect 11422 2524 11428 2536
rect 11480 2524 11486 2576
rect 13633 2567 13691 2573
rect 13633 2564 13645 2567
rect 11992 2536 13645 2564
rect 9766 2456 9772 2508
rect 9824 2496 9830 2508
rect 11992 2505 12020 2536
rect 13633 2533 13645 2536
rect 13679 2533 13691 2567
rect 15654 2564 15660 2576
rect 15615 2536 15660 2564
rect 13633 2527 13691 2533
rect 15654 2524 15660 2536
rect 15712 2524 15718 2576
rect 16206 2524 16212 2576
rect 16264 2564 16270 2576
rect 16393 2567 16451 2573
rect 16393 2564 16405 2567
rect 16264 2536 16405 2564
rect 16264 2524 16270 2536
rect 16393 2533 16405 2536
rect 16439 2533 16451 2567
rect 16393 2527 16451 2533
rect 17236 2536 18368 2564
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 9824 2468 11161 2496
rect 9824 2456 9830 2468
rect 11149 2465 11161 2468
rect 11195 2465 11207 2499
rect 11149 2459 11207 2465
rect 11977 2499 12035 2505
rect 11977 2465 11989 2499
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 12710 2496 12716 2508
rect 12667 2468 12716 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 12710 2456 12716 2468
rect 12768 2456 12774 2508
rect 12894 2456 12900 2508
rect 12952 2496 12958 2508
rect 13357 2499 13415 2505
rect 13357 2496 13369 2499
rect 12952 2468 13369 2496
rect 12952 2456 12958 2468
rect 13357 2465 13369 2468
rect 13403 2465 13415 2499
rect 14090 2496 14096 2508
rect 14051 2468 14096 2496
rect 13357 2459 13415 2465
rect 14090 2456 14096 2468
rect 14148 2456 14154 2508
rect 14642 2496 14648 2508
rect 14603 2468 14648 2496
rect 14642 2456 14648 2468
rect 14700 2456 14706 2508
rect 15562 2456 15568 2508
rect 15620 2496 15626 2508
rect 17236 2496 17264 2536
rect 18340 2505 18368 2536
rect 17405 2499 17463 2505
rect 17405 2496 17417 2499
rect 15620 2468 17264 2496
rect 17328 2468 17417 2496
rect 15620 2456 15626 2468
rect 10134 2428 10140 2440
rect 10095 2400 10140 2428
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 12526 2388 12532 2440
rect 12584 2428 12590 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12584 2400 12817 2428
rect 12584 2388 12590 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 16482 2428 16488 2440
rect 16443 2400 16488 2428
rect 12805 2391 12863 2397
rect 16482 2388 16488 2400
rect 16540 2388 16546 2440
rect 14090 2360 14096 2372
rect 8444 2332 8892 2360
rect 8956 2332 14096 2360
rect 8444 2320 8450 2332
rect 8294 2292 8300 2304
rect 8255 2264 8300 2292
rect 8294 2252 8300 2264
rect 8352 2252 8358 2304
rect 8665 2295 8723 2301
rect 8665 2261 8677 2295
rect 8711 2292 8723 2295
rect 8754 2292 8760 2304
rect 8711 2264 8760 2292
rect 8711 2261 8723 2264
rect 8665 2255 8723 2261
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 8864 2292 8892 2332
rect 14090 2320 14096 2332
rect 14148 2320 14154 2372
rect 15933 2363 15991 2369
rect 15933 2329 15945 2363
rect 15979 2360 15991 2363
rect 17328 2360 17356 2468
rect 17405 2465 17417 2468
rect 17451 2465 17463 2499
rect 17405 2459 17463 2465
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2496 18935 2499
rect 19150 2496 19156 2508
rect 18923 2468 19156 2496
rect 18923 2465 18935 2468
rect 18877 2459 18935 2465
rect 19150 2456 19156 2468
rect 19208 2456 19214 2508
rect 19426 2496 19432 2508
rect 19387 2468 19432 2496
rect 19426 2456 19432 2468
rect 19484 2456 19490 2508
rect 19981 2499 20039 2505
rect 19981 2465 19993 2499
rect 20027 2465 20039 2499
rect 20530 2496 20536 2508
rect 20491 2468 20536 2496
rect 19981 2459 20039 2465
rect 17494 2428 17500 2440
rect 17455 2400 17500 2428
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 19242 2388 19248 2440
rect 19300 2428 19306 2440
rect 19996 2428 20024 2459
rect 20530 2456 20536 2468
rect 20588 2456 20594 2508
rect 19300 2400 20024 2428
rect 19300 2388 19306 2400
rect 15979 2332 17356 2360
rect 15979 2329 15991 2332
rect 15933 2323 15991 2329
rect 18138 2320 18144 2372
rect 18196 2360 18202 2372
rect 19061 2363 19119 2369
rect 19061 2360 19073 2363
rect 18196 2332 19073 2360
rect 18196 2320 18202 2332
rect 19061 2329 19073 2332
rect 19107 2329 19119 2363
rect 19061 2323 19119 2329
rect 19334 2320 19340 2372
rect 19392 2360 19398 2372
rect 20165 2363 20223 2369
rect 20165 2360 20177 2363
rect 19392 2332 20177 2360
rect 19392 2320 19398 2332
rect 20165 2329 20177 2332
rect 20211 2329 20223 2363
rect 20165 2323 20223 2329
rect 9398 2292 9404 2304
rect 8864 2264 9404 2292
rect 9398 2252 9404 2264
rect 9456 2252 9462 2304
rect 12161 2295 12219 2301
rect 12161 2261 12173 2295
rect 12207 2292 12219 2295
rect 13170 2292 13176 2304
rect 12207 2264 13176 2292
rect 12207 2261 12219 2264
rect 12161 2255 12219 2261
rect 13170 2252 13176 2264
rect 13228 2252 13234 2304
rect 13722 2252 13728 2304
rect 13780 2292 13786 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13780 2264 14289 2292
rect 13780 2252 13786 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14826 2292 14832 2304
rect 14787 2264 14832 2292
rect 14277 2255 14335 2261
rect 14826 2252 14832 2264
rect 14884 2252 14890 2304
rect 17034 2252 17040 2304
rect 17092 2292 17098 2304
rect 18509 2295 18567 2301
rect 18509 2292 18521 2295
rect 17092 2264 18521 2292
rect 17092 2252 17098 2264
rect 18509 2261 18521 2264
rect 18555 2261 18567 2295
rect 18509 2255 18567 2261
rect 18782 2252 18788 2304
rect 18840 2292 18846 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 18840 2264 19625 2292
rect 18840 2252 18846 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 20438 2252 20444 2304
rect 20496 2292 20502 2304
rect 20717 2295 20775 2301
rect 20717 2292 20729 2295
rect 20496 2264 20729 2292
rect 20496 2252 20502 2264
rect 20717 2261 20729 2264
rect 20763 2261 20775 2295
rect 20717 2255 20775 2261
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 8754 2048 8760 2100
rect 8812 2088 8818 2100
rect 15562 2088 15568 2100
rect 8812 2060 15568 2088
rect 8812 2048 8818 2060
rect 15562 2048 15568 2060
rect 15620 2048 15626 2100
rect 15657 2091 15715 2097
rect 15657 2057 15669 2091
rect 15703 2088 15715 2091
rect 19242 2088 19248 2100
rect 15703 2060 19248 2088
rect 15703 2057 15715 2060
rect 15657 2051 15715 2057
rect 19242 2048 19248 2060
rect 19300 2048 19306 2100
rect 9766 1980 9772 2032
rect 9824 2020 9830 2032
rect 12250 2020 12256 2032
rect 9824 1992 12256 2020
rect 9824 1980 9830 1992
rect 12250 1980 12256 1992
rect 12308 1980 12314 2032
rect 8294 1912 8300 1964
rect 8352 1952 8358 1964
rect 16206 1952 16212 1964
rect 8352 1924 16212 1952
rect 8352 1912 8358 1924
rect 16206 1912 16212 1924
rect 16264 1912 16270 1964
rect 9398 1844 9404 1896
rect 9456 1884 9462 1896
rect 15657 1887 15715 1893
rect 15657 1884 15669 1887
rect 9456 1856 15669 1884
rect 9456 1844 9462 1856
rect 15657 1853 15669 1856
rect 15703 1853 15715 1887
rect 15657 1847 15715 1853
rect 10686 1096 10692 1148
rect 10744 1136 10750 1148
rect 14274 1136 14280 1148
rect 10744 1108 14280 1136
rect 10744 1096 10750 1108
rect 14274 1096 14280 1108
rect 14332 1096 14338 1148
<< via1 >>
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 12072 20544 12124 20596
rect 12348 20544 12400 20596
rect 14832 20544 14884 20596
rect 16304 20544 16356 20596
rect 17776 20544 17828 20596
rect 18144 20544 18196 20596
rect 18604 20544 18656 20596
rect 19340 20587 19392 20596
rect 12624 20476 12676 20528
rect 15384 20476 15436 20528
rect 10692 20408 10744 20460
rect 10968 20383 11020 20392
rect 10968 20349 10977 20383
rect 10977 20349 11011 20383
rect 11011 20349 11020 20383
rect 10968 20340 11020 20349
rect 12072 20340 12124 20392
rect 13452 20340 13504 20392
rect 12256 20272 12308 20324
rect 15844 20340 15896 20392
rect 18788 20476 18840 20528
rect 19340 20553 19349 20587
rect 19349 20553 19383 20587
rect 19383 20553 19392 20587
rect 19340 20544 19392 20553
rect 19892 20587 19944 20596
rect 19892 20553 19901 20587
rect 19901 20553 19935 20587
rect 19935 20553 19944 20587
rect 19892 20544 19944 20553
rect 19432 20408 19484 20460
rect 17776 20340 17828 20392
rect 18420 20340 18472 20392
rect 18604 20383 18656 20392
rect 18604 20349 18613 20383
rect 18613 20349 18647 20383
rect 18647 20349 18656 20383
rect 18604 20340 18656 20349
rect 19156 20383 19208 20392
rect 19156 20349 19165 20383
rect 19165 20349 19199 20383
rect 19199 20349 19208 20383
rect 19156 20340 19208 20349
rect 19524 20340 19576 20392
rect 20536 20383 20588 20392
rect 20536 20349 20545 20383
rect 20545 20349 20579 20383
rect 20579 20349 20588 20383
rect 20536 20340 20588 20349
rect 7748 20204 7800 20256
rect 10416 20204 10468 20256
rect 10784 20204 10836 20256
rect 11980 20204 12032 20256
rect 12992 20204 13044 20256
rect 13452 20204 13504 20256
rect 13544 20247 13596 20256
rect 13544 20213 13553 20247
rect 13553 20213 13587 20247
rect 13587 20213 13596 20247
rect 13544 20204 13596 20213
rect 15752 20204 15804 20256
rect 16028 20204 16080 20256
rect 19800 20272 19852 20324
rect 17132 20204 17184 20256
rect 17960 20204 18012 20256
rect 18880 20204 18932 20256
rect 20628 20204 20680 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 11244 20000 11296 20052
rect 13820 20000 13872 20052
rect 14372 20000 14424 20052
rect 15936 20000 15988 20052
rect 16580 20000 16632 20052
rect 18696 20000 18748 20052
rect 18972 20043 19024 20052
rect 18972 20009 18981 20043
rect 18981 20009 19015 20043
rect 19015 20009 19024 20043
rect 18972 20000 19024 20009
rect 9128 19932 9180 19984
rect 11888 19932 11940 19984
rect 13728 19932 13780 19984
rect 9680 19864 9732 19916
rect 11244 19864 11296 19916
rect 11704 19864 11756 19916
rect 10600 19839 10652 19848
rect 10600 19805 10609 19839
rect 10609 19805 10643 19839
rect 10643 19805 10652 19839
rect 10600 19796 10652 19805
rect 12164 19796 12216 19848
rect 13820 19796 13872 19848
rect 14464 19932 14516 19984
rect 15752 19932 15804 19984
rect 20996 20000 21048 20052
rect 19156 19932 19208 19984
rect 15660 19907 15712 19916
rect 15660 19873 15669 19907
rect 15669 19873 15703 19907
rect 15703 19873 15712 19907
rect 15660 19864 15712 19873
rect 16396 19864 16448 19916
rect 17316 19864 17368 19916
rect 17868 19907 17920 19916
rect 17868 19873 17877 19907
rect 17877 19873 17911 19907
rect 17911 19873 17920 19907
rect 17868 19864 17920 19873
rect 18420 19907 18472 19916
rect 18420 19873 18429 19907
rect 18429 19873 18463 19907
rect 18463 19873 18472 19907
rect 18420 19864 18472 19873
rect 18788 19907 18840 19916
rect 18788 19873 18797 19907
rect 18797 19873 18831 19907
rect 18831 19873 18840 19907
rect 18788 19864 18840 19873
rect 15384 19796 15436 19848
rect 15844 19839 15896 19848
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 15844 19796 15896 19805
rect 16580 19796 16632 19848
rect 7564 19660 7616 19712
rect 8392 19660 8444 19712
rect 11152 19728 11204 19780
rect 9864 19703 9916 19712
rect 9864 19669 9873 19703
rect 9873 19669 9907 19703
rect 9907 19669 9916 19703
rect 9864 19660 9916 19669
rect 11796 19660 11848 19712
rect 11888 19660 11940 19712
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 14648 19660 14700 19712
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 20720 19864 20772 19916
rect 18972 19796 19024 19848
rect 21548 19796 21600 19848
rect 19248 19728 19300 19780
rect 19156 19660 19208 19712
rect 19892 19703 19944 19712
rect 19892 19669 19901 19703
rect 19901 19669 19935 19703
rect 19935 19669 19944 19703
rect 19892 19660 19944 19669
rect 19984 19660 20036 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 9496 19456 9548 19508
rect 11704 19456 11756 19508
rect 12440 19456 12492 19508
rect 13820 19499 13872 19508
rect 12348 19388 12400 19440
rect 13820 19465 13829 19499
rect 13829 19465 13863 19499
rect 13863 19465 13872 19499
rect 13820 19456 13872 19465
rect 15660 19456 15712 19508
rect 15936 19456 15988 19508
rect 21548 19456 21600 19508
rect 9588 19320 9640 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 13820 19320 13872 19372
rect 296 19252 348 19304
rect 8576 19252 8628 19304
rect 9220 19252 9272 19304
rect 9680 19295 9732 19304
rect 9680 19261 9689 19295
rect 9689 19261 9723 19295
rect 9723 19261 9732 19295
rect 9680 19252 9732 19261
rect 9772 19252 9824 19304
rect 11244 19252 11296 19304
rect 12532 19252 12584 19304
rect 14096 19295 14148 19304
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 15200 19320 15252 19372
rect 19156 19388 19208 19440
rect 17868 19320 17920 19372
rect 18788 19320 18840 19372
rect 16580 19252 16632 19304
rect 16856 19252 16908 19304
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 19524 19252 19576 19304
rect 10140 19184 10192 19236
rect 10508 19227 10560 19236
rect 10508 19193 10542 19227
rect 10542 19193 10560 19227
rect 10508 19184 10560 19193
rect 13912 19184 13964 19236
rect 4160 19116 4212 19168
rect 8944 19116 8996 19168
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 10784 19116 10836 19168
rect 14740 19116 14792 19168
rect 16028 19184 16080 19236
rect 18788 19184 18840 19236
rect 18972 19184 19024 19236
rect 19800 19184 19852 19236
rect 22652 19184 22704 19236
rect 21456 19116 21508 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 848 18912 900 18964
rect 6368 18912 6420 18964
rect 6460 18912 6512 18964
rect 9864 18912 9916 18964
rect 10048 18912 10100 18964
rect 10508 18912 10560 18964
rect 11796 18955 11848 18964
rect 11796 18921 11805 18955
rect 11805 18921 11839 18955
rect 11839 18921 11848 18955
rect 11796 18912 11848 18921
rect 11888 18912 11940 18964
rect 13176 18912 13228 18964
rect 14648 18955 14700 18964
rect 14648 18921 14657 18955
rect 14657 18921 14691 18955
rect 14691 18921 14700 18955
rect 14648 18912 14700 18921
rect 1400 18844 1452 18896
rect 6828 18844 6880 18896
rect 9036 18844 9088 18896
rect 15844 18844 15896 18896
rect 17040 18912 17092 18964
rect 17684 18912 17736 18964
rect 20536 18912 20588 18964
rect 18972 18844 19024 18896
rect 20352 18844 20404 18896
rect 2504 18776 2556 18828
rect 8208 18708 8260 18760
rect 3056 18572 3108 18624
rect 7656 18572 7708 18624
rect 8208 18615 8260 18624
rect 8208 18581 8217 18615
rect 8217 18581 8251 18615
rect 8251 18581 8260 18615
rect 8208 18572 8260 18581
rect 8484 18615 8536 18624
rect 8484 18581 8493 18615
rect 8493 18581 8527 18615
rect 8527 18581 8536 18615
rect 8484 18572 8536 18581
rect 9220 18776 9272 18828
rect 9772 18776 9824 18828
rect 11244 18776 11296 18828
rect 13360 18819 13412 18828
rect 8944 18708 8996 18760
rect 9404 18708 9456 18760
rect 11152 18708 11204 18760
rect 11796 18708 11848 18760
rect 12164 18708 12216 18760
rect 12808 18751 12860 18760
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 13360 18785 13369 18819
rect 13369 18785 13403 18819
rect 13403 18785 13412 18819
rect 13360 18776 13412 18785
rect 14004 18776 14056 18828
rect 14464 18776 14516 18828
rect 14924 18776 14976 18828
rect 17684 18819 17736 18828
rect 17684 18785 17693 18819
rect 17693 18785 17727 18819
rect 17727 18785 17736 18819
rect 17684 18776 17736 18785
rect 20260 18819 20312 18828
rect 15200 18708 15252 18760
rect 8852 18572 8904 18624
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9312 18572 9364 18581
rect 11704 18572 11756 18624
rect 12440 18572 12492 18624
rect 15384 18640 15436 18692
rect 12900 18572 12952 18624
rect 14096 18572 14148 18624
rect 18144 18708 18196 18760
rect 16488 18640 16540 18692
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 20260 18785 20269 18819
rect 20269 18785 20303 18819
rect 20303 18785 20312 18819
rect 20260 18776 20312 18785
rect 21364 18776 21416 18828
rect 19432 18708 19484 18717
rect 21088 18708 21140 18760
rect 15752 18572 15804 18624
rect 16580 18572 16632 18624
rect 18696 18572 18748 18624
rect 20076 18572 20128 18624
rect 20444 18615 20496 18624
rect 20444 18581 20453 18615
rect 20453 18581 20487 18615
rect 20487 18581 20496 18615
rect 20444 18572 20496 18581
rect 21180 18572 21232 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 7012 18368 7064 18420
rect 3608 18300 3660 18352
rect 6552 18300 6604 18352
rect 1952 18232 2004 18284
rect 7012 18232 7064 18284
rect 5264 18164 5316 18216
rect 6920 18164 6972 18216
rect 7564 18368 7616 18420
rect 8208 18368 8260 18420
rect 11152 18368 11204 18420
rect 12164 18368 12216 18420
rect 14004 18368 14056 18420
rect 8668 18300 8720 18352
rect 11244 18300 11296 18352
rect 11796 18300 11848 18352
rect 13912 18343 13964 18352
rect 8208 18232 8260 18284
rect 9220 18164 9272 18216
rect 9404 18164 9456 18216
rect 12532 18232 12584 18284
rect 10324 18164 10376 18216
rect 10600 18164 10652 18216
rect 12808 18207 12860 18216
rect 5816 18096 5868 18148
rect 7104 18096 7156 18148
rect 9036 18096 9088 18148
rect 9588 18096 9640 18148
rect 9864 18096 9916 18148
rect 10232 18096 10284 18148
rect 4804 18028 4856 18080
rect 6184 18028 6236 18080
rect 6368 18028 6420 18080
rect 10140 18028 10192 18080
rect 10324 18071 10376 18080
rect 10324 18037 10333 18071
rect 10333 18037 10367 18071
rect 10367 18037 10376 18071
rect 10324 18028 10376 18037
rect 12808 18173 12817 18207
rect 12817 18173 12851 18207
rect 12851 18173 12860 18207
rect 12808 18164 12860 18173
rect 12900 18207 12952 18216
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 13912 18309 13921 18343
rect 13921 18309 13955 18343
rect 13955 18309 13964 18343
rect 13912 18300 13964 18309
rect 15844 18368 15896 18420
rect 20536 18368 20588 18420
rect 16488 18300 16540 18352
rect 18052 18300 18104 18352
rect 20904 18300 20956 18352
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 19064 18232 19116 18284
rect 19340 18232 19392 18284
rect 19432 18232 19484 18284
rect 12900 18164 12952 18173
rect 13820 18164 13872 18216
rect 14096 18164 14148 18216
rect 10784 18028 10836 18080
rect 12164 18028 12216 18080
rect 13176 18096 13228 18148
rect 13268 18096 13320 18148
rect 15200 18096 15252 18148
rect 16672 18164 16724 18216
rect 17868 18164 17920 18216
rect 18696 18164 18748 18216
rect 20076 18207 20128 18216
rect 18144 18096 18196 18148
rect 19064 18096 19116 18148
rect 20076 18173 20085 18207
rect 20085 18173 20119 18207
rect 20119 18173 20128 18207
rect 20076 18164 20128 18173
rect 20812 18207 20864 18216
rect 20812 18173 20821 18207
rect 20821 18173 20855 18207
rect 20855 18173 20864 18207
rect 20812 18164 20864 18173
rect 22100 18096 22152 18148
rect 17040 18071 17092 18080
rect 17040 18037 17049 18071
rect 17049 18037 17083 18071
rect 17083 18037 17092 18071
rect 19432 18071 19484 18080
rect 17040 18028 17092 18037
rect 19432 18037 19441 18071
rect 19441 18037 19475 18071
rect 19475 18037 19484 18071
rect 19432 18028 19484 18037
rect 20168 18071 20220 18080
rect 20168 18037 20177 18071
rect 20177 18037 20211 18071
rect 20211 18037 20220 18071
rect 20168 18028 20220 18037
rect 20996 18071 21048 18080
rect 20996 18037 21005 18071
rect 21005 18037 21039 18071
rect 21039 18037 21048 18071
rect 20996 18028 21048 18037
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 7104 17867 7156 17876
rect 7104 17833 7113 17867
rect 7113 17833 7147 17867
rect 7147 17833 7156 17867
rect 7104 17824 7156 17833
rect 9036 17867 9088 17876
rect 9036 17833 9045 17867
rect 9045 17833 9079 17867
rect 9079 17833 9088 17867
rect 9036 17824 9088 17833
rect 11704 17824 11756 17876
rect 8668 17756 8720 17808
rect 13636 17756 13688 17808
rect 16764 17824 16816 17876
rect 17224 17824 17276 17876
rect 7932 17731 7984 17740
rect 7932 17697 7966 17731
rect 7966 17697 7984 17731
rect 7932 17688 7984 17697
rect 8208 17688 8260 17740
rect 8484 17688 8536 17740
rect 11060 17731 11112 17740
rect 11060 17697 11069 17731
rect 11069 17697 11103 17731
rect 11103 17697 11112 17731
rect 11060 17688 11112 17697
rect 12164 17731 12216 17740
rect 12164 17697 12173 17731
rect 12173 17697 12207 17731
rect 12207 17697 12216 17731
rect 12164 17688 12216 17697
rect 12992 17688 13044 17740
rect 6276 17484 6328 17536
rect 7288 17484 7340 17536
rect 9036 17620 9088 17672
rect 9588 17620 9640 17672
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 14648 17731 14700 17740
rect 14648 17697 14657 17731
rect 14657 17697 14691 17731
rect 14691 17697 14700 17731
rect 15292 17731 15344 17740
rect 14648 17688 14700 17697
rect 15292 17697 15301 17731
rect 15301 17697 15335 17731
rect 15335 17697 15344 17731
rect 15292 17688 15344 17697
rect 15752 17688 15804 17740
rect 16580 17756 16632 17808
rect 20168 17824 20220 17876
rect 20352 17867 20404 17876
rect 20352 17833 20361 17867
rect 20361 17833 20395 17867
rect 20395 17833 20404 17867
rect 20352 17824 20404 17833
rect 20812 17824 20864 17876
rect 20720 17756 20772 17808
rect 18236 17688 18288 17740
rect 20904 17731 20956 17740
rect 20904 17697 20913 17731
rect 20913 17697 20947 17731
rect 20947 17697 20956 17731
rect 20904 17688 20956 17697
rect 14096 17620 14148 17672
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 17592 17620 17644 17672
rect 18696 17620 18748 17672
rect 9312 17552 9364 17604
rect 19064 17595 19116 17604
rect 9220 17484 9272 17536
rect 10508 17484 10560 17536
rect 11796 17527 11848 17536
rect 11796 17493 11805 17527
rect 11805 17493 11839 17527
rect 11839 17493 11848 17527
rect 11796 17484 11848 17493
rect 13084 17527 13136 17536
rect 13084 17493 13093 17527
rect 13093 17493 13127 17527
rect 13127 17493 13136 17527
rect 13084 17484 13136 17493
rect 14556 17484 14608 17536
rect 14832 17527 14884 17536
rect 14832 17493 14841 17527
rect 14841 17493 14875 17527
rect 14875 17493 14884 17527
rect 14832 17484 14884 17493
rect 19064 17561 19073 17595
rect 19073 17561 19107 17595
rect 19107 17561 19116 17595
rect 19064 17552 19116 17561
rect 17684 17484 17736 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 7288 17280 7340 17332
rect 7932 17280 7984 17332
rect 8392 17144 8444 17196
rect 9312 17280 9364 17332
rect 11060 17280 11112 17332
rect 9036 17212 9088 17264
rect 11704 17212 11756 17264
rect 12900 17280 12952 17332
rect 13084 17280 13136 17332
rect 14648 17280 14700 17332
rect 15568 17280 15620 17332
rect 9588 17144 9640 17196
rect 11980 17187 12032 17196
rect 11980 17153 11989 17187
rect 11989 17153 12023 17187
rect 12023 17153 12032 17187
rect 11980 17144 12032 17153
rect 12624 17212 12676 17264
rect 5908 17076 5960 17128
rect 6644 17076 6696 17128
rect 7748 17076 7800 17128
rect 9312 17076 9364 17128
rect 9496 17008 9548 17060
rect 10324 17076 10376 17128
rect 10508 17119 10560 17128
rect 10508 17085 10517 17119
rect 10517 17085 10551 17119
rect 10551 17085 10560 17119
rect 10508 17076 10560 17085
rect 12440 17144 12492 17196
rect 14372 17212 14424 17264
rect 14740 17212 14792 17264
rect 16672 17280 16724 17332
rect 21364 17280 21416 17332
rect 15200 17187 15252 17196
rect 15200 17153 15209 17187
rect 15209 17153 15243 17187
rect 15243 17153 15252 17187
rect 15200 17144 15252 17153
rect 15844 17144 15896 17196
rect 16580 17144 16632 17196
rect 17960 17212 18012 17264
rect 18236 17212 18288 17264
rect 17224 17144 17276 17196
rect 17868 17144 17920 17196
rect 20260 17187 20312 17196
rect 20260 17153 20269 17187
rect 20269 17153 20303 17187
rect 20303 17153 20312 17187
rect 20260 17144 20312 17153
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 12532 17076 12584 17128
rect 12992 17076 13044 17128
rect 14096 17076 14148 17128
rect 17960 17076 18012 17128
rect 19432 17076 19484 17128
rect 14648 17008 14700 17060
rect 18052 17008 18104 17060
rect 20352 17076 20404 17128
rect 7196 16940 7248 16992
rect 8484 16940 8536 16992
rect 8760 16940 8812 16992
rect 9036 16940 9088 16992
rect 12808 16940 12860 16992
rect 13452 16940 13504 16992
rect 13820 16940 13872 16992
rect 14004 16940 14056 16992
rect 14464 16940 14516 16992
rect 15568 16983 15620 16992
rect 15568 16949 15577 16983
rect 15577 16949 15611 16983
rect 15611 16949 15620 16983
rect 15568 16940 15620 16949
rect 15936 16983 15988 16992
rect 15936 16949 15945 16983
rect 15945 16949 15979 16983
rect 15979 16949 15988 16983
rect 15936 16940 15988 16949
rect 16028 16983 16080 16992
rect 16028 16949 16037 16983
rect 16037 16949 16071 16983
rect 16071 16949 16080 16983
rect 16948 16983 17000 16992
rect 16028 16940 16080 16949
rect 16948 16949 16957 16983
rect 16957 16949 16991 16983
rect 16991 16949 17000 16983
rect 16948 16940 17000 16949
rect 17132 16940 17184 16992
rect 17684 16940 17736 16992
rect 19340 16940 19392 16992
rect 19708 16983 19760 16992
rect 19708 16949 19717 16983
rect 19717 16949 19751 16983
rect 19751 16949 19760 16983
rect 19708 16940 19760 16949
rect 20260 16940 20312 16992
rect 21456 16940 21508 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 5908 16779 5960 16788
rect 5908 16745 5917 16779
rect 5917 16745 5951 16779
rect 5951 16745 5960 16779
rect 5908 16736 5960 16745
rect 7748 16736 7800 16788
rect 8944 16736 8996 16788
rect 9220 16736 9272 16788
rect 7472 16668 7524 16720
rect 10876 16736 10928 16788
rect 11152 16736 11204 16788
rect 11980 16736 12032 16788
rect 12900 16736 12952 16788
rect 13452 16736 13504 16788
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 8116 16600 8168 16652
rect 8852 16600 8904 16652
rect 9312 16600 9364 16652
rect 10324 16600 10376 16652
rect 10508 16643 10560 16652
rect 10508 16609 10517 16643
rect 10517 16609 10551 16643
rect 10551 16609 10560 16643
rect 10508 16600 10560 16609
rect 11060 16643 11112 16652
rect 11060 16609 11094 16643
rect 11094 16609 11112 16643
rect 11060 16600 11112 16609
rect 14372 16736 14424 16788
rect 14556 16779 14608 16788
rect 14556 16745 14565 16779
rect 14565 16745 14599 16779
rect 14599 16745 14608 16779
rect 14556 16736 14608 16745
rect 16028 16736 16080 16788
rect 17132 16779 17184 16788
rect 17132 16745 17141 16779
rect 17141 16745 17175 16779
rect 17175 16745 17184 16779
rect 17132 16736 17184 16745
rect 18144 16779 18196 16788
rect 18144 16745 18153 16779
rect 18153 16745 18187 16779
rect 18187 16745 18196 16779
rect 18144 16736 18196 16745
rect 15384 16668 15436 16720
rect 18696 16736 18748 16788
rect 21088 16779 21140 16788
rect 21088 16745 21097 16779
rect 21097 16745 21131 16779
rect 21131 16745 21140 16779
rect 21088 16736 21140 16745
rect 14096 16600 14148 16652
rect 15200 16600 15252 16652
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 14740 16575 14792 16584
rect 12440 16532 12492 16541
rect 14740 16541 14749 16575
rect 14749 16541 14783 16575
rect 14783 16541 14792 16575
rect 14740 16532 14792 16541
rect 6276 16439 6328 16448
rect 6276 16405 6285 16439
rect 6285 16405 6319 16439
rect 6319 16405 6328 16439
rect 6276 16396 6328 16405
rect 8760 16396 8812 16448
rect 9312 16439 9364 16448
rect 9312 16405 9321 16439
rect 9321 16405 9355 16439
rect 9355 16405 9364 16439
rect 9312 16396 9364 16405
rect 9864 16396 9916 16448
rect 13544 16464 13596 16516
rect 15476 16464 15528 16516
rect 18696 16600 18748 16652
rect 18880 16643 18932 16652
rect 18880 16609 18889 16643
rect 18889 16609 18923 16643
rect 18923 16609 18932 16643
rect 18880 16600 18932 16609
rect 20720 16600 20772 16652
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 17224 16575 17276 16584
rect 15844 16532 15896 16541
rect 17224 16541 17233 16575
rect 17233 16541 17267 16575
rect 17267 16541 17276 16575
rect 17224 16532 17276 16541
rect 18972 16575 19024 16584
rect 18972 16541 18981 16575
rect 18981 16541 19015 16575
rect 19015 16541 19024 16575
rect 18972 16532 19024 16541
rect 19064 16575 19116 16584
rect 19064 16541 19073 16575
rect 19073 16541 19107 16575
rect 19107 16541 19116 16575
rect 19524 16575 19576 16584
rect 19064 16532 19116 16541
rect 19524 16541 19533 16575
rect 19533 16541 19567 16575
rect 19567 16541 19576 16575
rect 19524 16532 19576 16541
rect 15660 16464 15712 16516
rect 16028 16464 16080 16516
rect 19616 16464 19668 16516
rect 16120 16439 16172 16448
rect 16120 16405 16129 16439
rect 16129 16405 16163 16439
rect 16163 16405 16172 16439
rect 16120 16396 16172 16405
rect 16304 16439 16356 16448
rect 16304 16405 16313 16439
rect 16313 16405 16347 16439
rect 16347 16405 16356 16439
rect 16304 16396 16356 16405
rect 17040 16396 17092 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 8116 16192 8168 16244
rect 9220 16192 9272 16244
rect 9496 16192 9548 16244
rect 12532 16192 12584 16244
rect 12808 16192 12860 16244
rect 13084 16192 13136 16244
rect 15936 16192 15988 16244
rect 18880 16192 18932 16244
rect 20352 16192 20404 16244
rect 11520 16167 11572 16176
rect 11520 16133 11529 16167
rect 11529 16133 11563 16167
rect 11563 16133 11572 16167
rect 11520 16124 11572 16133
rect 12348 16056 12400 16108
rect 15384 16124 15436 16176
rect 7380 15988 7432 16040
rect 8760 16031 8812 16040
rect 8760 15997 8794 16031
rect 8794 15997 8812 16031
rect 8760 15988 8812 15997
rect 9036 15988 9088 16040
rect 9220 15988 9272 16040
rect 9772 15988 9824 16040
rect 10784 15920 10836 15972
rect 10876 15920 10928 15972
rect 6460 15895 6512 15904
rect 6460 15861 6469 15895
rect 6469 15861 6503 15895
rect 6503 15861 6512 15895
rect 6460 15852 6512 15861
rect 8944 15852 8996 15904
rect 12072 15852 12124 15904
rect 13452 16099 13504 16108
rect 13452 16065 13461 16099
rect 13461 16065 13495 16099
rect 13495 16065 13504 16099
rect 13452 16056 13504 16065
rect 15844 16056 15896 16108
rect 14740 15988 14792 16040
rect 15568 15988 15620 16040
rect 13820 15920 13872 15972
rect 19432 16124 19484 16176
rect 19156 16099 19208 16108
rect 19156 16065 19165 16099
rect 19165 16065 19199 16099
rect 19199 16065 19208 16099
rect 19156 16056 19208 16065
rect 19708 16056 19760 16108
rect 17960 15988 18012 16040
rect 19524 15988 19576 16040
rect 15384 15852 15436 15904
rect 15568 15895 15620 15904
rect 15568 15861 15577 15895
rect 15577 15861 15611 15895
rect 15611 15861 15620 15895
rect 15568 15852 15620 15861
rect 16396 15852 16448 15904
rect 18328 15895 18380 15904
rect 18328 15861 18337 15895
rect 18337 15861 18371 15895
rect 18371 15861 18380 15895
rect 18328 15852 18380 15861
rect 20076 15852 20128 15904
rect 20352 15895 20404 15904
rect 20352 15861 20361 15895
rect 20361 15861 20395 15895
rect 20395 15861 20404 15895
rect 20352 15852 20404 15861
rect 20628 15852 20680 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 6184 15691 6236 15700
rect 6184 15657 6193 15691
rect 6193 15657 6227 15691
rect 6227 15657 6236 15691
rect 6184 15648 6236 15657
rect 6552 15691 6604 15700
rect 6552 15657 6561 15691
rect 6561 15657 6595 15691
rect 6595 15657 6604 15691
rect 6552 15648 6604 15657
rect 6828 15648 6880 15700
rect 10876 15648 10928 15700
rect 12072 15648 12124 15700
rect 10600 15623 10652 15632
rect 6920 15512 6972 15564
rect 6552 15444 6604 15496
rect 10600 15589 10609 15623
rect 10609 15589 10643 15623
rect 10643 15589 10652 15623
rect 10600 15580 10652 15589
rect 12808 15648 12860 15700
rect 15384 15691 15436 15700
rect 15384 15657 15393 15691
rect 15393 15657 15427 15691
rect 15427 15657 15436 15691
rect 15384 15648 15436 15657
rect 16120 15648 16172 15700
rect 16948 15691 17000 15700
rect 16948 15657 16957 15691
rect 16957 15657 16991 15691
rect 16991 15657 17000 15691
rect 16948 15648 17000 15657
rect 18972 15648 19024 15700
rect 19616 15691 19668 15700
rect 19616 15657 19625 15691
rect 19625 15657 19659 15691
rect 19659 15657 19668 15691
rect 19616 15648 19668 15657
rect 17040 15580 17092 15632
rect 19708 15580 19760 15632
rect 20168 15580 20220 15632
rect 9036 15512 9088 15564
rect 11244 15512 11296 15564
rect 8208 15444 8260 15496
rect 8852 15444 8904 15496
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 6828 15376 6880 15428
rect 10784 15487 10836 15496
rect 10784 15453 10793 15487
rect 10793 15453 10827 15487
rect 10827 15453 10836 15487
rect 11704 15487 11756 15496
rect 10784 15444 10836 15453
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 12348 15444 12400 15496
rect 7564 15308 7616 15360
rect 8760 15308 8812 15360
rect 8944 15308 8996 15360
rect 12808 15308 12860 15360
rect 13084 15376 13136 15428
rect 13820 15487 13872 15496
rect 13820 15453 13829 15487
rect 13829 15453 13863 15487
rect 13863 15453 13872 15487
rect 13820 15444 13872 15453
rect 14556 15444 14608 15496
rect 16488 15487 16540 15496
rect 16488 15453 16497 15487
rect 16497 15453 16531 15487
rect 16531 15453 16540 15487
rect 17500 15487 17552 15496
rect 16488 15444 16540 15453
rect 17500 15453 17509 15487
rect 17509 15453 17543 15487
rect 17543 15453 17552 15487
rect 17500 15444 17552 15453
rect 19708 15487 19760 15496
rect 19708 15453 19717 15487
rect 19717 15453 19751 15487
rect 19751 15453 19760 15487
rect 19708 15444 19760 15453
rect 19064 15376 19116 15428
rect 19340 15376 19392 15428
rect 19616 15376 19668 15428
rect 16488 15308 16540 15360
rect 16580 15308 16632 15360
rect 20444 15351 20496 15360
rect 20444 15317 20453 15351
rect 20453 15317 20487 15351
rect 20487 15317 20496 15351
rect 20444 15308 20496 15317
rect 20536 15308 20588 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 6460 15147 6512 15156
rect 6460 15113 6469 15147
rect 6469 15113 6503 15147
rect 6503 15113 6512 15147
rect 6460 15104 6512 15113
rect 6920 15147 6972 15156
rect 6920 15113 6929 15147
rect 6929 15113 6963 15147
rect 6963 15113 6972 15147
rect 6920 15104 6972 15113
rect 7288 15104 7340 15156
rect 8944 15104 8996 15156
rect 9036 15104 9088 15156
rect 11704 15104 11756 15156
rect 12440 15104 12492 15156
rect 20352 15104 20404 15156
rect 7656 15036 7708 15088
rect 8392 14968 8444 15020
rect 8852 14968 8904 15020
rect 8300 14900 8352 14952
rect 9956 15036 10008 15088
rect 10508 15036 10560 15088
rect 11612 15036 11664 15088
rect 11888 15036 11940 15088
rect 14464 15036 14516 15088
rect 16488 15036 16540 15088
rect 16672 15036 16724 15088
rect 13912 15011 13964 15020
rect 8668 14764 8720 14816
rect 9680 14832 9732 14884
rect 10140 14900 10192 14952
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 10876 14900 10928 14952
rect 10784 14832 10836 14884
rect 8944 14807 8996 14816
rect 8944 14773 8953 14807
rect 8953 14773 8987 14807
rect 8987 14773 8996 14807
rect 8944 14764 8996 14773
rect 10324 14764 10376 14816
rect 11244 14764 11296 14816
rect 12624 14900 12676 14952
rect 13912 14977 13921 15011
rect 13921 14977 13955 15011
rect 13955 14977 13964 15011
rect 13912 14968 13964 14977
rect 14372 14968 14424 15020
rect 15660 14968 15712 15020
rect 14280 14900 14332 14952
rect 12532 14832 12584 14884
rect 12716 14875 12768 14884
rect 12716 14841 12725 14875
rect 12725 14841 12759 14875
rect 12759 14841 12768 14875
rect 12716 14832 12768 14841
rect 14740 14832 14792 14884
rect 15384 14832 15436 14884
rect 19064 14900 19116 14952
rect 13728 14807 13780 14816
rect 13728 14773 13737 14807
rect 13737 14773 13771 14807
rect 13771 14773 13780 14807
rect 13728 14764 13780 14773
rect 13820 14807 13872 14816
rect 13820 14773 13829 14807
rect 13829 14773 13863 14807
rect 13863 14773 13872 14807
rect 13820 14764 13872 14773
rect 14096 14764 14148 14816
rect 16764 14807 16816 14816
rect 16764 14773 16773 14807
rect 16773 14773 16807 14807
rect 16807 14773 16816 14807
rect 16764 14764 16816 14773
rect 18052 14807 18104 14816
rect 18052 14773 18061 14807
rect 18061 14773 18095 14807
rect 18095 14773 18104 14807
rect 18052 14764 18104 14773
rect 18604 14832 18656 14884
rect 19248 14832 19300 14884
rect 18880 14764 18932 14816
rect 19892 14807 19944 14816
rect 19892 14773 19901 14807
rect 19901 14773 19935 14807
rect 19935 14773 19944 14807
rect 21180 14807 21232 14816
rect 19892 14764 19944 14773
rect 21180 14773 21189 14807
rect 21189 14773 21223 14807
rect 21223 14773 21232 14807
rect 21180 14764 21232 14773
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 6644 14560 6696 14612
rect 7472 14560 7524 14612
rect 7656 14560 7708 14612
rect 8300 14603 8352 14612
rect 8300 14569 8309 14603
rect 8309 14569 8343 14603
rect 8343 14569 8352 14603
rect 8300 14560 8352 14569
rect 8668 14603 8720 14612
rect 8668 14569 8677 14603
rect 8677 14569 8711 14603
rect 8711 14569 8720 14603
rect 8668 14560 8720 14569
rect 8760 14603 8812 14612
rect 8760 14569 8769 14603
rect 8769 14569 8803 14603
rect 8803 14569 8812 14603
rect 8760 14560 8812 14569
rect 8944 14560 8996 14612
rect 11152 14560 11204 14612
rect 11888 14560 11940 14612
rect 13820 14560 13872 14612
rect 12624 14492 12676 14544
rect 12716 14492 12768 14544
rect 16580 14560 16632 14612
rect 16672 14560 16724 14612
rect 19432 14560 19484 14612
rect 20076 14560 20128 14612
rect 21180 14560 21232 14612
rect 14832 14492 14884 14544
rect 7288 14424 7340 14476
rect 8300 14424 8352 14476
rect 9772 14424 9824 14476
rect 11704 14467 11756 14476
rect 11704 14433 11713 14467
rect 11713 14433 11747 14467
rect 11747 14433 11756 14467
rect 11704 14424 11756 14433
rect 12164 14424 12216 14476
rect 12900 14467 12952 14476
rect 12900 14433 12909 14467
rect 12909 14433 12943 14467
rect 12943 14433 12952 14467
rect 12900 14424 12952 14433
rect 13820 14467 13872 14476
rect 13820 14433 13854 14467
rect 13854 14433 13872 14467
rect 13820 14424 13872 14433
rect 14280 14424 14332 14476
rect 15660 14467 15712 14476
rect 9496 14356 9548 14408
rect 12440 14356 12492 14408
rect 13544 14399 13596 14408
rect 11060 14331 11112 14340
rect 11060 14297 11069 14331
rect 11069 14297 11103 14331
rect 11103 14297 11112 14331
rect 11060 14288 11112 14297
rect 7656 14263 7708 14272
rect 7656 14229 7665 14263
rect 7665 14229 7699 14263
rect 7699 14229 7708 14263
rect 7656 14220 7708 14229
rect 8760 14220 8812 14272
rect 10416 14220 10468 14272
rect 11888 14220 11940 14272
rect 12624 14288 12676 14340
rect 12532 14220 12584 14272
rect 13084 14220 13136 14272
rect 13544 14365 13553 14399
rect 13553 14365 13587 14399
rect 13587 14365 13596 14399
rect 13544 14356 13596 14365
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 15200 14356 15252 14408
rect 17776 14424 17828 14476
rect 17868 14424 17920 14476
rect 19524 14492 19576 14544
rect 20260 14535 20312 14544
rect 20260 14501 20269 14535
rect 20269 14501 20303 14535
rect 20303 14501 20312 14535
rect 20260 14492 20312 14501
rect 20720 14424 20772 14476
rect 21180 14424 21232 14476
rect 17500 14356 17552 14408
rect 18052 14356 18104 14408
rect 19892 14356 19944 14408
rect 14280 14220 14332 14272
rect 14740 14220 14792 14272
rect 15292 14263 15344 14272
rect 15292 14229 15301 14263
rect 15301 14229 15335 14263
rect 15335 14229 15344 14263
rect 15292 14220 15344 14229
rect 15752 14220 15804 14272
rect 16396 14220 16448 14272
rect 17684 14220 17736 14272
rect 17868 14263 17920 14272
rect 17868 14229 17877 14263
rect 17877 14229 17911 14263
rect 17911 14229 17920 14263
rect 17868 14220 17920 14229
rect 17960 14220 18012 14272
rect 20352 14220 20404 14272
rect 20628 14220 20680 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 6460 14059 6512 14068
rect 6460 14025 6469 14059
rect 6469 14025 6503 14059
rect 6503 14025 6512 14059
rect 6460 14016 6512 14025
rect 7564 14016 7616 14068
rect 7656 14016 7708 14068
rect 9036 14016 9088 14068
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 10876 14016 10928 14068
rect 7748 13948 7800 14000
rect 8944 13948 8996 14000
rect 12440 14016 12492 14068
rect 13176 14016 13228 14068
rect 13728 14016 13780 14068
rect 13820 13991 13872 14000
rect 10140 13880 10192 13932
rect 11704 13880 11756 13932
rect 7288 13812 7340 13864
rect 8760 13812 8812 13864
rect 9956 13855 10008 13864
rect 8944 13744 8996 13796
rect 9404 13744 9456 13796
rect 9956 13821 9965 13855
rect 9965 13821 9999 13855
rect 9999 13821 10008 13855
rect 9956 13812 10008 13821
rect 11060 13812 11112 13864
rect 12256 13744 12308 13796
rect 11336 13676 11388 13728
rect 11704 13676 11756 13728
rect 13820 13957 13829 13991
rect 13829 13957 13863 13991
rect 13863 13957 13872 13991
rect 14832 14016 14884 14068
rect 15200 14059 15252 14068
rect 15200 14025 15209 14059
rect 15209 14025 15243 14059
rect 15243 14025 15252 14059
rect 15200 14016 15252 14025
rect 13820 13948 13872 13957
rect 13544 13880 13596 13932
rect 15752 13948 15804 14000
rect 14648 13880 14700 13932
rect 17408 13948 17460 14000
rect 20444 14016 20496 14068
rect 17960 13948 18012 14000
rect 20352 13948 20404 14000
rect 17040 13923 17092 13932
rect 12532 13812 12584 13864
rect 14372 13812 14424 13864
rect 17040 13889 17049 13923
rect 17049 13889 17083 13923
rect 17083 13889 17092 13923
rect 17040 13880 17092 13889
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 21548 13880 21600 13932
rect 15200 13812 15252 13864
rect 15752 13812 15804 13864
rect 15936 13812 15988 13864
rect 16580 13812 16632 13864
rect 18880 13812 18932 13864
rect 19892 13812 19944 13864
rect 20812 13812 20864 13864
rect 12624 13744 12676 13796
rect 13544 13676 13596 13728
rect 14004 13676 14056 13728
rect 15476 13676 15528 13728
rect 16212 13676 16264 13728
rect 17960 13676 18012 13728
rect 18420 13719 18472 13728
rect 18420 13685 18429 13719
rect 18429 13685 18463 13719
rect 18463 13685 18472 13719
rect 18420 13676 18472 13685
rect 20904 13676 20956 13728
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 7012 13472 7064 13524
rect 8208 13472 8260 13524
rect 10692 13472 10744 13524
rect 10876 13472 10928 13524
rect 11888 13515 11940 13524
rect 7472 13447 7524 13456
rect 7472 13413 7481 13447
rect 7481 13413 7515 13447
rect 7515 13413 7524 13447
rect 7472 13404 7524 13413
rect 7656 13404 7708 13456
rect 9128 13447 9180 13456
rect 9128 13413 9137 13447
rect 9137 13413 9171 13447
rect 9171 13413 9180 13447
rect 9128 13404 9180 13413
rect 9680 13404 9732 13456
rect 11336 13404 11388 13456
rect 11888 13481 11897 13515
rect 11897 13481 11931 13515
rect 11931 13481 11940 13515
rect 11888 13472 11940 13481
rect 13452 13472 13504 13524
rect 13728 13472 13780 13524
rect 14556 13515 14608 13524
rect 14556 13481 14565 13515
rect 14565 13481 14599 13515
rect 14599 13481 14608 13515
rect 14556 13472 14608 13481
rect 12624 13404 12676 13456
rect 13544 13404 13596 13456
rect 16948 13472 17000 13524
rect 17776 13515 17828 13524
rect 17776 13481 17785 13515
rect 17785 13481 17819 13515
rect 17819 13481 17828 13515
rect 17776 13472 17828 13481
rect 17868 13472 17920 13524
rect 20168 13472 20220 13524
rect 21180 13447 21232 13456
rect 9772 13379 9824 13388
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 9772 13336 9824 13345
rect 11796 13379 11848 13388
rect 11796 13345 11805 13379
rect 11805 13345 11839 13379
rect 11839 13345 11848 13379
rect 11796 13336 11848 13345
rect 12072 13336 12124 13388
rect 13452 13379 13504 13388
rect 13452 13345 13461 13379
rect 13461 13345 13495 13379
rect 13495 13345 13504 13379
rect 13452 13336 13504 13345
rect 15200 13336 15252 13388
rect 16396 13379 16448 13388
rect 16396 13345 16405 13379
rect 16405 13345 16439 13379
rect 16439 13345 16448 13379
rect 16396 13336 16448 13345
rect 6276 13268 6328 13320
rect 9496 13268 9548 13320
rect 11336 13268 11388 13320
rect 11888 13268 11940 13320
rect 13636 13311 13688 13320
rect 6644 13200 6696 13252
rect 9772 13200 9824 13252
rect 12440 13243 12492 13252
rect 12440 13209 12449 13243
rect 12449 13209 12483 13243
rect 12483 13209 12492 13243
rect 12440 13200 12492 13209
rect 13636 13277 13645 13311
rect 13645 13277 13679 13311
rect 13679 13277 13688 13311
rect 13636 13268 13688 13277
rect 14372 13268 14424 13320
rect 15844 13311 15896 13320
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 15844 13268 15896 13277
rect 7472 13132 7524 13184
rect 7748 13132 7800 13184
rect 8668 13132 8720 13184
rect 11152 13175 11204 13184
rect 11152 13141 11161 13175
rect 11161 13141 11195 13175
rect 11195 13141 11204 13175
rect 15660 13200 15712 13252
rect 11152 13132 11204 13141
rect 12992 13132 13044 13184
rect 13268 13132 13320 13184
rect 13636 13132 13688 13184
rect 14004 13132 14056 13184
rect 18328 13336 18380 13388
rect 18604 13336 18656 13388
rect 19432 13379 19484 13388
rect 19432 13345 19455 13379
rect 19455 13345 19484 13379
rect 21180 13413 21189 13447
rect 21189 13413 21223 13447
rect 21223 13413 21232 13447
rect 21180 13404 21232 13413
rect 19432 13336 19484 13345
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 18696 13311 18748 13320
rect 18696 13277 18705 13311
rect 18705 13277 18739 13311
rect 18739 13277 18748 13311
rect 18696 13268 18748 13277
rect 18880 13268 18932 13320
rect 17684 13132 17736 13184
rect 18052 13175 18104 13184
rect 18052 13141 18061 13175
rect 18061 13141 18095 13175
rect 18095 13141 18104 13175
rect 18052 13132 18104 13141
rect 18972 13132 19024 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 7380 12928 7432 12980
rect 9864 12928 9916 12980
rect 10876 12928 10928 12980
rect 12072 12928 12124 12980
rect 15752 12928 15804 12980
rect 15844 12928 15896 12980
rect 17132 12928 17184 12980
rect 18604 12928 18656 12980
rect 18696 12928 18748 12980
rect 13452 12860 13504 12912
rect 6644 12792 6696 12844
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 11060 12792 11112 12844
rect 11888 12792 11940 12844
rect 12072 12792 12124 12844
rect 12624 12792 12676 12844
rect 16212 12860 16264 12912
rect 14372 12792 14424 12844
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 14740 12792 14792 12801
rect 11152 12724 11204 12776
rect 11704 12724 11756 12776
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 10140 12656 10192 12708
rect 14096 12724 14148 12776
rect 17132 12792 17184 12844
rect 17776 12792 17828 12844
rect 9404 12588 9456 12640
rect 9864 12588 9916 12640
rect 10600 12588 10652 12640
rect 11244 12588 11296 12640
rect 11796 12588 11848 12640
rect 12256 12588 12308 12640
rect 12624 12588 12676 12640
rect 13728 12656 13780 12708
rect 18052 12724 18104 12776
rect 15292 12656 15344 12708
rect 14464 12588 14516 12640
rect 15936 12631 15988 12640
rect 15936 12597 15945 12631
rect 15945 12597 15979 12631
rect 15979 12597 15988 12631
rect 15936 12588 15988 12597
rect 16028 12588 16080 12640
rect 16304 12588 16356 12640
rect 17960 12656 18012 12708
rect 18604 12792 18656 12844
rect 18328 12724 18380 12776
rect 18972 12767 19024 12776
rect 18972 12733 19006 12767
rect 19006 12733 19024 12767
rect 18972 12724 19024 12733
rect 17868 12588 17920 12640
rect 18236 12588 18288 12640
rect 18604 12588 18656 12640
rect 18880 12588 18932 12640
rect 19064 12656 19116 12708
rect 20628 12792 20680 12844
rect 20444 12724 20496 12776
rect 20536 12656 20588 12708
rect 20720 12588 20772 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 7288 12384 7340 12436
rect 14464 12384 14516 12436
rect 15936 12384 15988 12436
rect 16948 12427 17000 12436
rect 16948 12393 16957 12427
rect 16957 12393 16991 12427
rect 16991 12393 17000 12427
rect 16948 12384 17000 12393
rect 17408 12427 17460 12436
rect 17408 12393 17417 12427
rect 17417 12393 17451 12427
rect 17451 12393 17460 12427
rect 17408 12384 17460 12393
rect 19156 12384 19208 12436
rect 19432 12384 19484 12436
rect 20628 12384 20680 12436
rect 21272 12384 21324 12436
rect 8668 12316 8720 12368
rect 9772 12316 9824 12368
rect 9956 12316 10008 12368
rect 11244 12316 11296 12368
rect 9220 12248 9272 12300
rect 12532 12316 12584 12368
rect 13360 12316 13412 12368
rect 18236 12316 18288 12368
rect 18512 12359 18564 12368
rect 18512 12325 18521 12359
rect 18521 12325 18555 12359
rect 18555 12325 18564 12359
rect 18512 12316 18564 12325
rect 18604 12316 18656 12368
rect 18880 12316 18932 12368
rect 19248 12316 19300 12368
rect 12348 12248 12400 12300
rect 14556 12248 14608 12300
rect 15200 12248 15252 12300
rect 15568 12291 15620 12300
rect 15568 12257 15602 12291
rect 15602 12257 15620 12291
rect 15568 12248 15620 12257
rect 20168 12248 20220 12300
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 10784 12223 10836 12232
rect 9404 12112 9456 12164
rect 9588 12112 9640 12164
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 11888 12180 11940 12232
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 9220 12044 9272 12096
rect 10140 12044 10192 12096
rect 12164 12087 12216 12096
rect 12164 12053 12173 12087
rect 12173 12053 12207 12087
rect 12207 12053 12216 12087
rect 12164 12044 12216 12053
rect 12440 12087 12492 12096
rect 12440 12053 12449 12087
rect 12449 12053 12483 12087
rect 12483 12053 12492 12087
rect 14188 12087 14240 12096
rect 12440 12044 12492 12053
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 17776 12180 17828 12232
rect 18696 12223 18748 12232
rect 18696 12189 18705 12223
rect 18705 12189 18739 12223
rect 18739 12189 18748 12223
rect 18696 12180 18748 12189
rect 18328 12112 18380 12164
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 17316 12044 17368 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 8852 11840 8904 11892
rect 9312 11840 9364 11892
rect 11244 11840 11296 11892
rect 12348 11704 12400 11756
rect 12532 11704 12584 11756
rect 9588 11636 9640 11688
rect 10232 11679 10284 11688
rect 10232 11645 10241 11679
rect 10241 11645 10275 11679
rect 10275 11645 10284 11679
rect 10232 11636 10284 11645
rect 10784 11636 10836 11688
rect 10324 11568 10376 11620
rect 13820 11568 13872 11620
rect 11152 11500 11204 11552
rect 12348 11500 12400 11552
rect 17960 11840 18012 11892
rect 18604 11840 18656 11892
rect 19800 11840 19852 11892
rect 20168 11883 20220 11892
rect 20168 11849 20177 11883
rect 20177 11849 20211 11883
rect 20211 11849 20220 11883
rect 20168 11840 20220 11849
rect 20536 11883 20588 11892
rect 20536 11849 20545 11883
rect 20545 11849 20579 11883
rect 20579 11849 20588 11883
rect 20536 11840 20588 11849
rect 14372 11815 14424 11824
rect 14372 11781 14381 11815
rect 14381 11781 14415 11815
rect 14415 11781 14424 11815
rect 14372 11772 14424 11781
rect 14372 11636 14424 11688
rect 14740 11636 14792 11688
rect 15292 11636 15344 11688
rect 17500 11704 17552 11756
rect 16028 11636 16080 11688
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 18144 11704 18196 11756
rect 18328 11704 18380 11756
rect 18420 11636 18472 11688
rect 20812 11636 20864 11688
rect 18972 11568 19024 11620
rect 20628 11568 20680 11620
rect 15200 11500 15252 11552
rect 15568 11500 15620 11552
rect 19248 11500 19300 11552
rect 20812 11500 20864 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 7564 11296 7616 11348
rect 9680 11339 9732 11348
rect 9680 11305 9689 11339
rect 9689 11305 9723 11339
rect 9723 11305 9732 11339
rect 9680 11296 9732 11305
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 12992 11296 13044 11348
rect 13084 11296 13136 11348
rect 15384 11296 15436 11348
rect 15476 11296 15528 11348
rect 18604 11296 18656 11348
rect 18972 11339 19024 11348
rect 18972 11305 18981 11339
rect 18981 11305 19015 11339
rect 19015 11305 19024 11339
rect 18972 11296 19024 11305
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 19616 11339 19668 11348
rect 19616 11305 19625 11339
rect 19625 11305 19659 11339
rect 19659 11305 19668 11339
rect 19616 11296 19668 11305
rect 20720 11296 20772 11348
rect 9128 11228 9180 11280
rect 11060 11228 11112 11280
rect 16672 11228 16724 11280
rect 11612 11160 11664 11212
rect 12072 11160 12124 11212
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 11060 11092 11112 11144
rect 14648 11160 14700 11212
rect 19064 11228 19116 11280
rect 18696 11160 18748 11212
rect 15476 11092 15528 11144
rect 10692 11067 10744 11076
rect 10692 11033 10701 11067
rect 10701 11033 10735 11067
rect 10735 11033 10744 11067
rect 10692 11024 10744 11033
rect 13820 11024 13872 11076
rect 14372 11024 14424 11076
rect 14464 11024 14516 11076
rect 17500 11092 17552 11144
rect 18604 11092 18656 11144
rect 19340 11092 19392 11144
rect 19708 11135 19760 11144
rect 19708 11101 19717 11135
rect 19717 11101 19751 11135
rect 19751 11101 19760 11135
rect 19708 11092 19760 11101
rect 20720 11092 20772 11144
rect 8484 10956 8536 11008
rect 10508 10956 10560 11008
rect 14004 10956 14056 11008
rect 20628 11024 20680 11076
rect 17776 10956 17828 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 10508 10752 10560 10804
rect 11888 10752 11940 10804
rect 14556 10752 14608 10804
rect 16120 10752 16172 10804
rect 17868 10752 17920 10804
rect 20720 10795 20772 10804
rect 20720 10761 20729 10795
rect 20729 10761 20763 10795
rect 20763 10761 20772 10795
rect 20720 10752 20772 10761
rect 9956 10684 10008 10736
rect 12808 10684 12860 10736
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 11244 10616 11296 10668
rect 14648 10684 14700 10736
rect 11980 10548 12032 10600
rect 12992 10548 13044 10600
rect 13544 10616 13596 10668
rect 14372 10616 14424 10668
rect 13728 10548 13780 10600
rect 13912 10548 13964 10600
rect 14740 10548 14792 10600
rect 15844 10548 15896 10600
rect 18052 10616 18104 10668
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 19340 10659 19392 10668
rect 19340 10625 19349 10659
rect 19349 10625 19383 10659
rect 19383 10625 19392 10659
rect 19340 10616 19392 10625
rect 10876 10480 10928 10532
rect 11060 10480 11112 10532
rect 11244 10523 11296 10532
rect 11244 10489 11253 10523
rect 11253 10489 11287 10523
rect 11287 10489 11296 10523
rect 11244 10480 11296 10489
rect 13452 10480 13504 10532
rect 10232 10455 10284 10464
rect 10232 10421 10241 10455
rect 10241 10421 10275 10455
rect 10275 10421 10284 10455
rect 10232 10412 10284 10421
rect 10692 10412 10744 10464
rect 11888 10412 11940 10464
rect 16028 10480 16080 10532
rect 13820 10412 13872 10464
rect 14372 10412 14424 10464
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 16304 10412 16356 10464
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 19616 10523 19668 10532
rect 19616 10489 19650 10523
rect 19650 10489 19668 10523
rect 19616 10480 19668 10489
rect 18144 10412 18196 10464
rect 18512 10455 18564 10464
rect 18512 10421 18521 10455
rect 18521 10421 18555 10455
rect 18555 10421 18564 10455
rect 18512 10412 18564 10421
rect 19524 10412 19576 10464
rect 21364 10412 21416 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 8576 10251 8628 10260
rect 8576 10217 8585 10251
rect 8585 10217 8619 10251
rect 8619 10217 8628 10251
rect 8576 10208 8628 10217
rect 8668 10208 8720 10260
rect 9128 10208 9180 10260
rect 11612 10208 11664 10260
rect 11980 10208 12032 10260
rect 13544 10208 13596 10260
rect 13820 10208 13872 10260
rect 14464 10208 14516 10260
rect 15292 10208 15344 10260
rect 15752 10208 15804 10260
rect 19156 10251 19208 10260
rect 19156 10217 19165 10251
rect 19165 10217 19199 10251
rect 19199 10217 19208 10251
rect 19156 10208 19208 10217
rect 19708 10251 19760 10260
rect 19708 10217 19717 10251
rect 19717 10217 19751 10251
rect 19751 10217 19760 10251
rect 19708 10208 19760 10217
rect 10416 10140 10468 10192
rect 12532 10140 12584 10192
rect 17684 10140 17736 10192
rect 20260 10140 20312 10192
rect 9312 10004 9364 10056
rect 11704 10072 11756 10124
rect 6920 9936 6972 9988
rect 9956 9936 10008 9988
rect 13544 10072 13596 10124
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 17224 10072 17276 10124
rect 21364 10072 21416 10124
rect 14096 10047 14148 10056
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 14096 10004 14148 10013
rect 14740 10047 14792 10056
rect 13728 9936 13780 9988
rect 14740 10013 14749 10047
rect 14749 10013 14783 10047
rect 14783 10013 14792 10047
rect 14740 10004 14792 10013
rect 15844 10047 15896 10056
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 17776 10047 17828 10056
rect 15844 10004 15896 10013
rect 17776 10013 17785 10047
rect 17785 10013 17819 10047
rect 17819 10013 17828 10047
rect 17776 10004 17828 10013
rect 18604 10047 18656 10056
rect 18604 10013 18613 10047
rect 18613 10013 18647 10047
rect 18647 10013 18656 10047
rect 18604 10004 18656 10013
rect 18696 10047 18748 10056
rect 18696 10013 18705 10047
rect 18705 10013 18739 10047
rect 18739 10013 18748 10047
rect 18696 10004 18748 10013
rect 17408 9936 17460 9988
rect 19616 9936 19668 9988
rect 21364 9979 21416 9988
rect 21364 9945 21373 9979
rect 21373 9945 21407 9979
rect 21407 9945 21416 9979
rect 21364 9936 21416 9945
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 12900 9868 12952 9920
rect 14188 9868 14240 9920
rect 14464 9868 14516 9920
rect 14740 9868 14792 9920
rect 17500 9868 17552 9920
rect 18972 9868 19024 9920
rect 20996 9911 21048 9920
rect 20996 9877 21005 9911
rect 21005 9877 21039 9911
rect 21039 9877 21048 9911
rect 20996 9868 21048 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 8576 9707 8628 9716
rect 8576 9673 8585 9707
rect 8585 9673 8619 9707
rect 8619 9673 8628 9707
rect 8576 9664 8628 9673
rect 10416 9664 10468 9716
rect 10876 9707 10928 9716
rect 10876 9673 10885 9707
rect 10885 9673 10919 9707
rect 10919 9673 10928 9707
rect 10876 9664 10928 9673
rect 11704 9664 11756 9716
rect 12532 9664 12584 9716
rect 14372 9664 14424 9716
rect 12900 9596 12952 9648
rect 13912 9596 13964 9648
rect 14096 9596 14148 9648
rect 14556 9596 14608 9648
rect 9312 9460 9364 9512
rect 10968 9460 11020 9512
rect 12716 9528 12768 9580
rect 12072 9503 12124 9512
rect 12072 9469 12081 9503
rect 12081 9469 12115 9503
rect 12115 9469 12124 9503
rect 12072 9460 12124 9469
rect 3424 9392 3476 9444
rect 7748 9324 7800 9376
rect 9956 9392 10008 9444
rect 13084 9460 13136 9512
rect 13728 9528 13780 9580
rect 14464 9528 14516 9580
rect 17960 9596 18012 9648
rect 18696 9664 18748 9716
rect 19616 9664 19668 9716
rect 19892 9664 19944 9716
rect 20444 9664 20496 9716
rect 17316 9528 17368 9580
rect 13544 9392 13596 9444
rect 16396 9460 16448 9512
rect 17776 9460 17828 9512
rect 18236 9460 18288 9512
rect 20444 9528 20496 9580
rect 19340 9460 19392 9512
rect 21364 9460 21416 9512
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 13452 9324 13504 9376
rect 14648 9367 14700 9376
rect 14648 9333 14657 9367
rect 14657 9333 14691 9367
rect 14691 9333 14700 9367
rect 14648 9324 14700 9333
rect 16120 9324 16172 9376
rect 18052 9392 18104 9444
rect 18512 9392 18564 9444
rect 19248 9324 19300 9376
rect 20352 9367 20404 9376
rect 20352 9333 20361 9367
rect 20361 9333 20395 9367
rect 20395 9333 20404 9367
rect 20352 9324 20404 9333
rect 20720 9367 20772 9376
rect 20720 9333 20729 9367
rect 20729 9333 20763 9367
rect 20763 9333 20772 9367
rect 20720 9324 20772 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 9956 9163 10008 9172
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 10232 9120 10284 9172
rect 10508 9120 10560 9172
rect 10784 9120 10836 9172
rect 11888 9163 11940 9172
rect 11888 9129 11897 9163
rect 11897 9129 11931 9163
rect 11931 9129 11940 9163
rect 11888 9120 11940 9129
rect 16396 9120 16448 9172
rect 10048 9052 10100 9104
rect 11612 9052 11664 9104
rect 13176 9052 13228 9104
rect 14648 9052 14700 9104
rect 16764 9052 16816 9104
rect 10140 8984 10192 9036
rect 10232 8984 10284 9036
rect 11060 8984 11112 9036
rect 12808 9027 12860 9036
rect 12808 8993 12817 9027
rect 12817 8993 12851 9027
rect 12851 8993 12860 9027
rect 12808 8984 12860 8993
rect 16028 8984 16080 9036
rect 17316 9120 17368 9172
rect 17776 9120 17828 9172
rect 18512 9163 18564 9172
rect 17960 9052 18012 9104
rect 18512 9129 18521 9163
rect 18521 9129 18555 9163
rect 18555 9129 18564 9163
rect 18512 9120 18564 9129
rect 18604 9120 18656 9172
rect 19156 9163 19208 9172
rect 19156 9129 19165 9163
rect 19165 9129 19199 9163
rect 19199 9129 19208 9163
rect 19156 9120 19208 9129
rect 20720 9120 20772 9172
rect 10968 8959 11020 8968
rect 10968 8925 10977 8959
rect 10977 8925 11011 8959
rect 11011 8925 11020 8959
rect 10968 8916 11020 8925
rect 11980 8959 12032 8968
rect 11980 8925 11989 8959
rect 11989 8925 12023 8959
rect 12023 8925 12032 8959
rect 11980 8916 12032 8925
rect 13728 8916 13780 8968
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 14372 8916 14424 8925
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 15844 8916 15896 8968
rect 16672 8916 16724 8968
rect 18696 8916 18748 8968
rect 12532 8848 12584 8900
rect 16856 8848 16908 8900
rect 18328 8848 18380 8900
rect 20260 9052 20312 9104
rect 20444 8959 20496 8968
rect 9772 8780 9824 8832
rect 10784 8780 10836 8832
rect 11888 8780 11940 8832
rect 12072 8780 12124 8832
rect 12716 8780 12768 8832
rect 18604 8780 18656 8832
rect 19800 8823 19852 8832
rect 19800 8789 19809 8823
rect 19809 8789 19843 8823
rect 19843 8789 19852 8823
rect 19800 8780 19852 8789
rect 20168 8780 20220 8832
rect 20444 8925 20453 8959
rect 20453 8925 20487 8959
rect 20487 8925 20496 8959
rect 20444 8916 20496 8925
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 10048 8576 10100 8628
rect 10968 8576 11020 8628
rect 11704 8576 11756 8628
rect 9312 8440 9364 8492
rect 12256 8576 12308 8628
rect 12440 8576 12492 8628
rect 14372 8576 14424 8628
rect 16764 8576 16816 8628
rect 19248 8576 19300 8628
rect 13728 8508 13780 8560
rect 15752 8551 15804 8560
rect 15752 8517 15761 8551
rect 15761 8517 15795 8551
rect 15795 8517 15804 8551
rect 15752 8508 15804 8517
rect 16120 8508 16172 8560
rect 19340 8508 19392 8560
rect 12256 8440 12308 8492
rect 16488 8483 16540 8492
rect 8852 8372 8904 8424
rect 11336 8372 11388 8424
rect 11980 8372 12032 8424
rect 12348 8372 12400 8424
rect 16488 8449 16497 8483
rect 16497 8449 16531 8483
rect 16531 8449 16540 8483
rect 16488 8440 16540 8449
rect 16672 8483 16724 8492
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 18144 8440 18196 8492
rect 19248 8483 19300 8492
rect 19248 8449 19257 8483
rect 19257 8449 19291 8483
rect 19291 8449 19300 8483
rect 19248 8440 19300 8449
rect 19432 8440 19484 8492
rect 16856 8372 16908 8424
rect 19800 8372 19852 8424
rect 20444 8372 20496 8424
rect 7656 8304 7708 8356
rect 10508 8304 10560 8356
rect 14464 8304 14516 8356
rect 15752 8304 15804 8356
rect 10232 8236 10284 8288
rect 13452 8236 13504 8288
rect 14372 8236 14424 8288
rect 14648 8236 14700 8288
rect 16580 8304 16632 8356
rect 18144 8304 18196 8356
rect 20352 8304 20404 8356
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 11060 8075 11112 8084
rect 11060 8041 11069 8075
rect 11069 8041 11103 8075
rect 11103 8041 11112 8075
rect 11060 8032 11112 8041
rect 14004 8032 14056 8084
rect 14556 8075 14608 8084
rect 14556 8041 14565 8075
rect 14565 8041 14599 8075
rect 14599 8041 14608 8075
rect 14556 8032 14608 8041
rect 14740 8032 14792 8084
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 17684 8032 17736 8084
rect 19156 8032 19208 8084
rect 20444 8032 20496 8084
rect 9772 7964 9824 8016
rect 12072 7964 12124 8016
rect 13728 7964 13780 8016
rect 9680 7828 9732 7880
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 7564 7760 7616 7812
rect 12256 7939 12308 7948
rect 11336 7828 11388 7880
rect 12256 7905 12265 7939
rect 12265 7905 12299 7939
rect 12299 7905 12308 7939
rect 12256 7896 12308 7905
rect 17960 7964 18012 8016
rect 18696 7964 18748 8016
rect 16304 7896 16356 7948
rect 16764 7896 16816 7948
rect 20536 7896 20588 7948
rect 15200 7828 15252 7880
rect 7288 7692 7340 7744
rect 8208 7692 8260 7744
rect 10876 7692 10928 7744
rect 13636 7735 13688 7744
rect 13636 7701 13645 7735
rect 13645 7701 13679 7735
rect 13679 7701 13688 7735
rect 13636 7692 13688 7701
rect 16488 7760 16540 7812
rect 17960 7760 18012 7812
rect 18604 7828 18656 7880
rect 20904 7871 20956 7880
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 17132 7692 17184 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 7472 7488 7524 7540
rect 11244 7488 11296 7540
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 14096 7488 14148 7540
rect 16304 7531 16356 7540
rect 11152 7420 11204 7472
rect 16304 7497 16313 7531
rect 16313 7497 16347 7531
rect 16347 7497 16356 7531
rect 16304 7488 16356 7497
rect 20812 7420 20864 7472
rect 13636 7352 13688 7404
rect 17868 7352 17920 7404
rect 20076 7395 20128 7404
rect 20076 7361 20085 7395
rect 20085 7361 20119 7395
rect 20119 7361 20128 7395
rect 20076 7352 20128 7361
rect 21088 7395 21140 7404
rect 21088 7361 21097 7395
rect 21097 7361 21131 7395
rect 21131 7361 21140 7395
rect 21088 7352 21140 7361
rect 8208 7284 8260 7336
rect 10140 7284 10192 7336
rect 10324 7327 10376 7336
rect 8668 7259 8720 7268
rect 8668 7225 8702 7259
rect 8702 7225 8720 7259
rect 8668 7216 8720 7225
rect 8392 7148 8444 7200
rect 10324 7293 10358 7327
rect 10358 7293 10376 7327
rect 10324 7284 10376 7293
rect 11152 7284 11204 7336
rect 13544 7284 13596 7336
rect 14096 7284 14148 7336
rect 17132 7284 17184 7336
rect 17684 7284 17736 7336
rect 12256 7216 12308 7268
rect 12624 7216 12676 7268
rect 13360 7216 13412 7268
rect 14372 7216 14424 7268
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 13452 7191 13504 7200
rect 13452 7157 13461 7191
rect 13461 7157 13495 7191
rect 13495 7157 13504 7191
rect 13452 7148 13504 7157
rect 14464 7148 14516 7200
rect 16396 7216 16448 7268
rect 18880 7284 18932 7336
rect 16764 7148 16816 7200
rect 17224 7148 17276 7200
rect 19248 7216 19300 7268
rect 20904 7284 20956 7336
rect 20628 7216 20680 7268
rect 17500 7148 17552 7200
rect 19524 7191 19576 7200
rect 19524 7157 19533 7191
rect 19533 7157 19567 7191
rect 19567 7157 19576 7191
rect 19524 7148 19576 7157
rect 19892 7148 19944 7200
rect 20168 7148 20220 7200
rect 20812 7148 20864 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 7564 6987 7616 6996
rect 7564 6953 7573 6987
rect 7573 6953 7607 6987
rect 7607 6953 7616 6987
rect 7564 6944 7616 6953
rect 8944 6987 8996 6996
rect 8944 6953 8953 6987
rect 8953 6953 8987 6987
rect 8987 6953 8996 6987
rect 8944 6944 8996 6953
rect 9680 6987 9732 6996
rect 9680 6953 9689 6987
rect 9689 6953 9723 6987
rect 9723 6953 9732 6987
rect 9680 6944 9732 6953
rect 12532 6944 12584 6996
rect 13268 6944 13320 6996
rect 13360 6944 13412 6996
rect 15844 6944 15896 6996
rect 16488 6987 16540 6996
rect 16488 6953 16497 6987
rect 16497 6953 16531 6987
rect 16531 6953 16540 6987
rect 16488 6944 16540 6953
rect 17500 6944 17552 6996
rect 19156 6944 19208 6996
rect 20536 6987 20588 6996
rect 20536 6953 20545 6987
rect 20545 6953 20579 6987
rect 20579 6953 20588 6987
rect 20536 6944 20588 6953
rect 9588 6876 9640 6928
rect 11152 6919 11204 6928
rect 7196 6808 7248 6860
rect 8760 6808 8812 6860
rect 9496 6808 9548 6860
rect 11152 6885 11161 6919
rect 11161 6885 11195 6919
rect 11195 6885 11204 6919
rect 11152 6876 11204 6885
rect 13636 6876 13688 6928
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 11888 6851 11940 6860
rect 11888 6817 11897 6851
rect 11897 6817 11931 6851
rect 11931 6817 11940 6851
rect 11888 6808 11940 6817
rect 14372 6808 14424 6860
rect 8668 6740 8720 6792
rect 7196 6647 7248 6656
rect 7196 6613 7205 6647
rect 7205 6613 7239 6647
rect 7239 6613 7248 6647
rect 7196 6604 7248 6613
rect 8760 6672 8812 6724
rect 9312 6740 9364 6792
rect 10876 6740 10928 6792
rect 14188 6740 14240 6792
rect 14740 6876 14792 6928
rect 17224 6876 17276 6928
rect 17868 6876 17920 6928
rect 20076 6876 20128 6928
rect 16120 6808 16172 6860
rect 17132 6851 17184 6860
rect 17132 6817 17141 6851
rect 17141 6817 17175 6851
rect 17175 6817 17184 6851
rect 17132 6808 17184 6817
rect 18604 6808 18656 6860
rect 19708 6808 19760 6860
rect 16396 6740 16448 6792
rect 8668 6604 8720 6656
rect 9496 6604 9548 6656
rect 10140 6604 10192 6656
rect 12440 6604 12492 6656
rect 13728 6604 13780 6656
rect 14556 6604 14608 6656
rect 15752 6604 15804 6656
rect 18972 6672 19024 6724
rect 19156 6672 19208 6724
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 7104 6400 7156 6452
rect 6828 6196 6880 6248
rect 8208 6400 8260 6452
rect 8668 6400 8720 6452
rect 9128 6400 9180 6452
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 10048 6400 10100 6452
rect 14372 6443 14424 6452
rect 9864 6332 9916 6384
rect 9588 6307 9640 6316
rect 9588 6273 9597 6307
rect 9597 6273 9631 6307
rect 9631 6273 9640 6307
rect 9588 6264 9640 6273
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 11060 6264 11112 6316
rect 13084 6332 13136 6384
rect 14372 6409 14381 6443
rect 14381 6409 14415 6443
rect 14415 6409 14424 6443
rect 14372 6400 14424 6409
rect 16856 6400 16908 6452
rect 17684 6400 17736 6452
rect 18972 6400 19024 6452
rect 13544 6332 13596 6384
rect 16396 6332 16448 6384
rect 8208 6239 8260 6248
rect 8208 6205 8242 6239
rect 8242 6205 8260 6239
rect 8208 6196 8260 6205
rect 8760 6196 8812 6248
rect 10048 6128 10100 6180
rect 10876 6128 10928 6180
rect 9956 6060 10008 6112
rect 13636 6264 13688 6316
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 16304 6264 16356 6316
rect 16764 6307 16816 6316
rect 16764 6273 16773 6307
rect 16773 6273 16807 6307
rect 16807 6273 16816 6307
rect 16764 6264 16816 6273
rect 17408 6332 17460 6384
rect 21088 6307 21140 6316
rect 21088 6273 21097 6307
rect 21097 6273 21131 6307
rect 21131 6273 21140 6307
rect 21088 6264 21140 6273
rect 13820 6239 13872 6248
rect 12992 6128 13044 6180
rect 13820 6205 13829 6239
rect 13829 6205 13863 6239
rect 13863 6205 13872 6239
rect 13820 6196 13872 6205
rect 15844 6196 15896 6248
rect 18144 6196 18196 6248
rect 18604 6196 18656 6248
rect 18880 6196 18932 6248
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 12624 6060 12676 6112
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 13360 6103 13412 6112
rect 13360 6069 13369 6103
rect 13369 6069 13403 6103
rect 13403 6069 13412 6103
rect 13360 6060 13412 6069
rect 13636 6128 13688 6180
rect 14464 6060 14516 6112
rect 17960 6128 18012 6180
rect 16856 6060 16908 6112
rect 20076 6060 20128 6112
rect 20260 6060 20312 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 8944 5856 8996 5908
rect 9036 5856 9088 5908
rect 9496 5856 9548 5908
rect 10048 5899 10100 5908
rect 10048 5865 10057 5899
rect 10057 5865 10091 5899
rect 10091 5865 10100 5899
rect 10048 5856 10100 5865
rect 10508 5856 10560 5908
rect 11704 5856 11756 5908
rect 14556 5899 14608 5908
rect 14556 5865 14565 5899
rect 14565 5865 14599 5899
rect 14599 5865 14608 5899
rect 14556 5856 14608 5865
rect 18880 5856 18932 5908
rect 19892 5856 19944 5908
rect 20260 5899 20312 5908
rect 20260 5865 20269 5899
rect 20269 5865 20303 5899
rect 20303 5865 20312 5899
rect 20260 5856 20312 5865
rect 9128 5788 9180 5840
rect 4068 5720 4120 5772
rect 10140 5720 10192 5772
rect 11060 5788 11112 5840
rect 12624 5788 12676 5840
rect 12808 5788 12860 5840
rect 12900 5788 12952 5840
rect 14832 5788 14884 5840
rect 11888 5720 11940 5772
rect 12072 5763 12124 5772
rect 12072 5729 12081 5763
rect 12081 5729 12115 5763
rect 12115 5729 12124 5763
rect 12072 5720 12124 5729
rect 12440 5763 12492 5772
rect 12440 5729 12449 5763
rect 12449 5729 12483 5763
rect 12483 5729 12492 5763
rect 12440 5720 12492 5729
rect 16672 5763 16724 5772
rect 16672 5729 16681 5763
rect 16681 5729 16715 5763
rect 16715 5729 16724 5763
rect 16672 5720 16724 5729
rect 17500 5788 17552 5840
rect 20168 5831 20220 5840
rect 20168 5797 20177 5831
rect 20177 5797 20211 5831
rect 20211 5797 20220 5831
rect 20168 5788 20220 5797
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 13728 5652 13780 5704
rect 15568 5652 15620 5704
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 16396 5652 16448 5704
rect 19432 5652 19484 5704
rect 20076 5652 20128 5704
rect 9956 5516 10008 5568
rect 12348 5584 12400 5636
rect 13912 5584 13964 5636
rect 11888 5516 11940 5568
rect 13084 5516 13136 5568
rect 16028 5516 16080 5568
rect 16580 5516 16632 5568
rect 17960 5516 18012 5568
rect 19800 5559 19852 5568
rect 19800 5525 19809 5559
rect 19809 5525 19843 5559
rect 19843 5525 19852 5559
rect 19800 5516 19852 5525
rect 22100 5516 22152 5568
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 8300 5312 8352 5364
rect 8760 5312 8812 5364
rect 9128 5355 9180 5364
rect 9128 5321 9137 5355
rect 9137 5321 9171 5355
rect 9171 5321 9180 5355
rect 9128 5312 9180 5321
rect 9772 5312 9824 5364
rect 10508 5312 10560 5364
rect 9864 5244 9916 5296
rect 11612 5244 11664 5296
rect 11980 5312 12032 5364
rect 12992 5355 13044 5364
rect 12992 5321 13001 5355
rect 13001 5321 13035 5355
rect 13035 5321 13044 5355
rect 12992 5312 13044 5321
rect 14464 5312 14516 5364
rect 14372 5244 14424 5296
rect 16396 5312 16448 5364
rect 17868 5312 17920 5364
rect 16120 5244 16172 5296
rect 11060 5176 11112 5228
rect 11888 5176 11940 5228
rect 13360 5176 13412 5228
rect 13728 5176 13780 5228
rect 17960 5176 18012 5228
rect 9772 5108 9824 5160
rect 14464 5151 14516 5160
rect 9312 5040 9364 5092
rect 10508 5040 10560 5092
rect 9496 4972 9548 5024
rect 10968 4972 11020 5024
rect 11244 5015 11296 5024
rect 11244 4981 11253 5015
rect 11253 4981 11287 5015
rect 11287 4981 11296 5015
rect 11244 4972 11296 4981
rect 12072 5040 12124 5092
rect 12348 5040 12400 5092
rect 12532 5040 12584 5092
rect 11980 4972 12032 5024
rect 13452 5040 13504 5092
rect 13268 4972 13320 5024
rect 14096 5015 14148 5024
rect 14096 4981 14105 5015
rect 14105 4981 14139 5015
rect 14139 4981 14148 5015
rect 14096 4972 14148 4981
rect 14464 5117 14473 5151
rect 14473 5117 14507 5151
rect 14507 5117 14516 5151
rect 14464 5108 14516 5117
rect 16396 5151 16448 5160
rect 16396 5117 16430 5151
rect 16430 5117 16448 5151
rect 15844 5040 15896 5092
rect 16396 5108 16448 5117
rect 16580 5040 16632 5092
rect 17960 5040 18012 5092
rect 18144 5108 18196 5160
rect 18604 5108 18656 5160
rect 18880 5108 18932 5160
rect 22652 5108 22704 5160
rect 20076 5040 20128 5092
rect 17500 5015 17552 5024
rect 17500 4981 17509 5015
rect 17509 4981 17543 5015
rect 17543 4981 17552 5015
rect 17500 4972 17552 4981
rect 18604 4972 18656 5024
rect 19616 4972 19668 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 10140 4768 10192 4820
rect 11060 4700 11112 4752
rect 10232 4632 10284 4684
rect 12532 4700 12584 4752
rect 11980 4632 12032 4684
rect 16856 4700 16908 4752
rect 13636 4632 13688 4684
rect 15476 4632 15528 4684
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 10784 4496 10836 4548
rect 11888 4607 11940 4616
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 11888 4564 11940 4573
rect 12072 4564 12124 4616
rect 12440 4564 12492 4616
rect 12900 4607 12952 4616
rect 12900 4573 12909 4607
rect 12909 4573 12943 4607
rect 12943 4573 12952 4607
rect 12900 4564 12952 4573
rect 14096 4564 14148 4616
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 16396 4632 16448 4684
rect 15844 4564 15896 4573
rect 9588 4428 9640 4480
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 11152 4428 11204 4480
rect 12624 4428 12676 4480
rect 13636 4428 13688 4480
rect 14096 4428 14148 4480
rect 14740 4428 14792 4480
rect 16672 4496 16724 4548
rect 16120 4428 16172 4480
rect 18880 4768 18932 4820
rect 19708 4768 19760 4820
rect 19800 4768 19852 4820
rect 19524 4700 19576 4752
rect 18144 4632 18196 4684
rect 18236 4632 18288 4684
rect 18880 4632 18932 4684
rect 19892 4632 19944 4684
rect 17316 4607 17368 4616
rect 17316 4573 17325 4607
rect 17325 4573 17359 4607
rect 17359 4573 17368 4607
rect 17316 4564 17368 4573
rect 19616 4564 19668 4616
rect 19708 4564 19760 4616
rect 19984 4564 20036 4616
rect 20536 4564 20588 4616
rect 17960 4428 18012 4480
rect 19524 4428 19576 4480
rect 19984 4428 20036 4480
rect 21548 4428 21600 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 7104 4224 7156 4276
rect 9864 4224 9916 4276
rect 11980 4267 12032 4276
rect 10048 4156 10100 4208
rect 4160 4088 4212 4140
rect 7380 4088 7432 4140
rect 7564 4088 7616 4140
rect 8944 4088 8996 4140
rect 11980 4233 11989 4267
rect 11989 4233 12023 4267
rect 12023 4233 12032 4267
rect 11980 4224 12032 4233
rect 17960 4224 18012 4276
rect 18972 4224 19024 4276
rect 19892 4224 19944 4276
rect 12992 4088 13044 4140
rect 13176 4088 13228 4140
rect 16028 4131 16080 4140
rect 16028 4097 16037 4131
rect 16037 4097 16071 4131
rect 16071 4097 16080 4131
rect 16028 4088 16080 4097
rect 17500 4156 17552 4208
rect 20076 4156 20128 4208
rect 5816 4020 5868 4072
rect 8484 4020 8536 4072
rect 10140 4020 10192 4072
rect 12532 4063 12584 4072
rect 3056 3952 3108 4004
rect 7656 3952 7708 4004
rect 7748 3952 7800 4004
rect 8208 3952 8260 4004
rect 11060 3952 11112 4004
rect 11152 3952 11204 4004
rect 11520 3952 11572 4004
rect 1952 3884 2004 3936
rect 7196 3884 7248 3936
rect 9772 3884 9824 3936
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 10600 3884 10652 3936
rect 12532 4029 12541 4063
rect 12541 4029 12575 4063
rect 12575 4029 12584 4063
rect 12532 4020 12584 4029
rect 12900 4020 12952 4072
rect 13820 4020 13872 4072
rect 16120 4020 16172 4072
rect 13452 3952 13504 4004
rect 13636 3952 13688 4004
rect 17132 4063 17184 4072
rect 17132 4029 17141 4063
rect 17141 4029 17175 4063
rect 17175 4029 17184 4063
rect 17132 4020 17184 4029
rect 17960 4020 18012 4072
rect 18144 4020 18196 4072
rect 18696 4020 18748 4072
rect 21272 4063 21324 4072
rect 21272 4029 21281 4063
rect 21281 4029 21315 4063
rect 21315 4029 21324 4063
rect 21272 4020 21324 4029
rect 16396 3952 16448 4004
rect 12440 3884 12492 3936
rect 12624 3884 12676 3936
rect 14740 3884 14792 3936
rect 15384 3884 15436 3936
rect 15752 3884 15804 3936
rect 15936 3884 15988 3936
rect 17408 3952 17460 4004
rect 17684 3884 17736 3936
rect 19708 3952 19760 4004
rect 20720 3927 20772 3936
rect 20720 3893 20729 3927
rect 20729 3893 20763 3927
rect 20763 3893 20772 3927
rect 20720 3884 20772 3893
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 5264 3680 5316 3732
rect 8668 3680 8720 3732
rect 9404 3680 9456 3732
rect 9864 3680 9916 3732
rect 10600 3680 10652 3732
rect 6460 3612 6512 3664
rect 11980 3612 12032 3664
rect 3608 3544 3660 3596
rect 6920 3544 6972 3596
rect 7012 3544 7064 3596
rect 10692 3544 10744 3596
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 11520 3544 11572 3596
rect 12900 3680 12952 3732
rect 14280 3680 14332 3732
rect 12164 3612 12216 3664
rect 13912 3655 13964 3664
rect 13912 3621 13921 3655
rect 13921 3621 13955 3655
rect 13955 3621 13964 3655
rect 17408 3680 17460 3732
rect 19708 3723 19760 3732
rect 13912 3612 13964 3621
rect 17132 3612 17184 3664
rect 19708 3689 19717 3723
rect 19717 3689 19751 3723
rect 19751 3689 19760 3723
rect 19708 3680 19760 3689
rect 18604 3655 18656 3664
rect 18604 3621 18616 3655
rect 18616 3621 18656 3655
rect 18604 3612 18656 3621
rect 15752 3587 15804 3596
rect 15752 3553 15761 3587
rect 15761 3553 15795 3587
rect 15795 3553 15804 3587
rect 15752 3544 15804 3553
rect 17500 3544 17552 3596
rect 19984 3587 20036 3596
rect 19984 3553 19993 3587
rect 19993 3553 20027 3587
rect 20027 3553 20036 3587
rect 19984 3544 20036 3553
rect 20444 3544 20496 3596
rect 10784 3476 10836 3528
rect 11336 3519 11388 3528
rect 11336 3485 11345 3519
rect 11345 3485 11379 3519
rect 11379 3485 11388 3519
rect 11336 3476 11388 3485
rect 14648 3519 14700 3528
rect 14648 3485 14657 3519
rect 14657 3485 14691 3519
rect 14691 3485 14700 3519
rect 14648 3476 14700 3485
rect 14740 3519 14792 3528
rect 14740 3485 14749 3519
rect 14749 3485 14783 3519
rect 14783 3485 14792 3519
rect 16672 3519 16724 3528
rect 14740 3476 14792 3485
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 18144 3476 18196 3528
rect 19524 3476 19576 3528
rect 8668 3408 8720 3460
rect 9588 3340 9640 3392
rect 10508 3383 10560 3392
rect 10508 3349 10517 3383
rect 10517 3349 10551 3383
rect 10551 3349 10560 3383
rect 10508 3340 10560 3349
rect 11152 3340 11204 3392
rect 11980 3340 12032 3392
rect 13728 3408 13780 3460
rect 15844 3408 15896 3460
rect 12992 3340 13044 3392
rect 13452 3383 13504 3392
rect 13452 3349 13461 3383
rect 13461 3349 13495 3383
rect 13495 3349 13504 3383
rect 13452 3340 13504 3349
rect 20996 3340 21048 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 9680 3136 9732 3188
rect 9864 3136 9916 3188
rect 9956 3136 10008 3188
rect 14648 3136 14700 3188
rect 17500 3179 17552 3188
rect 17500 3145 17509 3179
rect 17509 3145 17543 3179
rect 17543 3145 17552 3179
rect 17500 3136 17552 3145
rect 18788 3136 18840 3188
rect 2504 3068 2556 3120
rect 10232 3068 10284 3120
rect 10692 3068 10744 3120
rect 1400 3000 1452 3052
rect 9680 3000 9732 3052
rect 4804 2932 4856 2984
rect 11060 3000 11112 3052
rect 11428 2932 11480 2984
rect 13452 3000 13504 3052
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 19340 3000 19392 3052
rect 19708 3043 19760 3052
rect 13544 2932 13596 2984
rect 14464 2975 14516 2984
rect 14464 2941 14473 2975
rect 14473 2941 14507 2975
rect 14507 2941 14516 2975
rect 14464 2932 14516 2941
rect 14740 2975 14792 2984
rect 14740 2941 14774 2975
rect 14774 2941 14792 2975
rect 14740 2932 14792 2941
rect 296 2796 348 2848
rect 9312 2796 9364 2848
rect 9496 2839 9548 2848
rect 9496 2805 9505 2839
rect 9505 2805 9539 2839
rect 9539 2805 9548 2839
rect 9496 2796 9548 2805
rect 9680 2796 9732 2848
rect 10968 2796 11020 2848
rect 11152 2839 11204 2848
rect 11152 2805 11161 2839
rect 11161 2805 11195 2839
rect 11195 2805 11204 2839
rect 11152 2796 11204 2805
rect 11704 2796 11756 2848
rect 12072 2796 12124 2848
rect 16672 2932 16724 2984
rect 18144 2932 18196 2984
rect 18420 2975 18472 2984
rect 18420 2941 18429 2975
rect 18429 2941 18463 2975
rect 18463 2941 18472 2975
rect 18420 2932 18472 2941
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19432 2932 19484 2941
rect 19708 3009 19717 3043
rect 19717 3009 19751 3043
rect 19751 3009 19760 3043
rect 19708 3000 19760 3009
rect 20444 3043 20496 3052
rect 20444 3009 20453 3043
rect 20453 3009 20487 3043
rect 20487 3009 20496 3043
rect 20444 3000 20496 3009
rect 20904 2975 20956 2984
rect 20904 2941 20913 2975
rect 20913 2941 20947 2975
rect 20947 2941 20956 2975
rect 20904 2932 20956 2941
rect 14188 2796 14240 2848
rect 16488 2864 16540 2916
rect 18144 2796 18196 2848
rect 19892 2796 19944 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 7288 2592 7340 2644
rect 8392 2320 8444 2372
rect 10232 2592 10284 2644
rect 16948 2635 17000 2644
rect 16948 2601 16957 2635
rect 16957 2601 16991 2635
rect 16991 2601 17000 2635
rect 16948 2592 17000 2601
rect 17316 2635 17368 2644
rect 17316 2601 17325 2635
rect 17325 2601 17359 2635
rect 17359 2601 17368 2635
rect 17316 2592 17368 2601
rect 21272 2635 21324 2644
rect 21272 2601 21281 2635
rect 21281 2601 21315 2635
rect 21315 2601 21324 2635
rect 21272 2592 21324 2601
rect 10968 2524 11020 2576
rect 11428 2567 11480 2576
rect 11428 2533 11437 2567
rect 11437 2533 11471 2567
rect 11471 2533 11480 2567
rect 11428 2524 11480 2533
rect 9772 2456 9824 2508
rect 15660 2567 15712 2576
rect 15660 2533 15669 2567
rect 15669 2533 15703 2567
rect 15703 2533 15712 2567
rect 15660 2524 15712 2533
rect 16212 2524 16264 2576
rect 12716 2456 12768 2508
rect 12900 2456 12952 2508
rect 14096 2499 14148 2508
rect 14096 2465 14105 2499
rect 14105 2465 14139 2499
rect 14139 2465 14148 2499
rect 14096 2456 14148 2465
rect 14648 2499 14700 2508
rect 14648 2465 14657 2499
rect 14657 2465 14691 2499
rect 14691 2465 14700 2499
rect 14648 2456 14700 2465
rect 15568 2456 15620 2508
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 12532 2388 12584 2440
rect 16488 2431 16540 2440
rect 16488 2397 16497 2431
rect 16497 2397 16531 2431
rect 16531 2397 16540 2431
rect 16488 2388 16540 2397
rect 8300 2295 8352 2304
rect 8300 2261 8309 2295
rect 8309 2261 8343 2295
rect 8343 2261 8352 2295
rect 8300 2252 8352 2261
rect 8760 2252 8812 2304
rect 14096 2320 14148 2372
rect 19156 2456 19208 2508
rect 19432 2499 19484 2508
rect 19432 2465 19441 2499
rect 19441 2465 19475 2499
rect 19475 2465 19484 2499
rect 19432 2456 19484 2465
rect 20536 2499 20588 2508
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 19248 2388 19300 2440
rect 20536 2465 20545 2499
rect 20545 2465 20579 2499
rect 20579 2465 20588 2499
rect 20536 2456 20588 2465
rect 18144 2320 18196 2372
rect 19340 2320 19392 2372
rect 9404 2295 9456 2304
rect 9404 2261 9413 2295
rect 9413 2261 9447 2295
rect 9447 2261 9456 2295
rect 9404 2252 9456 2261
rect 13176 2252 13228 2304
rect 13728 2252 13780 2304
rect 14832 2295 14884 2304
rect 14832 2261 14841 2295
rect 14841 2261 14875 2295
rect 14875 2261 14884 2295
rect 14832 2252 14884 2261
rect 17040 2252 17092 2304
rect 18788 2252 18840 2304
rect 20444 2252 20496 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 8760 2048 8812 2100
rect 15568 2048 15620 2100
rect 19248 2048 19300 2100
rect 9772 1980 9824 2032
rect 12256 1980 12308 2032
rect 8300 1912 8352 1964
rect 16212 1912 16264 1964
rect 9404 1844 9456 1896
rect 10692 1096 10744 1148
rect 14280 1096 14332 1148
<< metal2 >>
rect 294 22200 350 23000
rect 846 22200 902 23000
rect 1398 22200 1454 23000
rect 1950 22200 2006 23000
rect 2502 22200 2558 23000
rect 3054 22200 3110 23000
rect 3606 22200 3662 23000
rect 4158 22200 4214 23000
rect 4710 22200 4766 23000
rect 5262 22200 5318 23000
rect 5814 22200 5870 23000
rect 6458 22200 6514 23000
rect 7010 22200 7066 23000
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10874 22200 10930 23000
rect 11426 22200 11482 23000
rect 12070 22200 12126 23000
rect 12622 22200 12678 23000
rect 13174 22200 13230 23000
rect 13726 22200 13782 23000
rect 14278 22200 14334 23000
rect 14830 22200 14886 23000
rect 15382 22200 15438 23000
rect 15934 22200 15990 23000
rect 16486 22200 16542 23000
rect 17038 22200 17094 23000
rect 17682 22200 17738 23000
rect 18234 22200 18290 23000
rect 18786 22200 18842 23000
rect 19062 22672 19118 22681
rect 19062 22607 19118 22616
rect 18878 22264 18934 22273
rect 308 19310 336 22200
rect 296 19304 348 19310
rect 296 19246 348 19252
rect 860 18970 888 22200
rect 848 18964 900 18970
rect 848 18906 900 18912
rect 1412 18902 1440 22200
rect 1400 18896 1452 18902
rect 1400 18838 1452 18844
rect 1964 18290 1992 22200
rect 2516 18834 2544 22200
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 3068 18630 3096 22200
rect 3056 18624 3108 18630
rect 3056 18566 3108 18572
rect 3620 18358 3648 22200
rect 4172 19174 4200 22200
rect 4724 20788 4752 22200
rect 4724 20760 4844 20788
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 3608 18352 3660 18358
rect 3608 18294 3660 18300
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 4816 18086 4844 20760
rect 5276 18222 5304 22200
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5828 18154 5856 22200
rect 6472 18970 6500 22200
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 6380 18086 6408 18906
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6552 18352 6604 18358
rect 6552 18294 6604 18300
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 3422 17232 3478 17241
rect 3422 17167 3478 17176
rect 3436 9450 3464 17167
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5920 16794 5948 17070
rect 5908 16788 5960 16794
rect 5908 16730 5960 16736
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 6196 15706 6224 18022
rect 6276 17536 6328 17542
rect 6276 17478 6328 17484
rect 6288 16454 6316 17478
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 6288 13326 6316 16390
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6472 15162 6500 15846
rect 6564 15706 6592 18294
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6564 15502 6592 15642
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6472 14074 6500 15098
rect 6656 14618 6684 17070
rect 6840 15706 6868 18838
rect 7024 18426 7052 22200
rect 7576 19718 7604 22200
rect 8128 20346 8156 22200
rect 8128 20318 8248 20346
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6840 15434 6868 15642
rect 6932 15570 6960 18158
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 6932 15162 6960 15506
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6656 13258 6684 14554
rect 7024 13530 7052 18226
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 7116 17882 7144 18090
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 6656 12850 6684 13194
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 4066 5808 4122 5817
rect 4066 5743 4068 5752
rect 4120 5743 4122 5752
rect 4068 5714 4120 5720
rect 6840 5710 6868 6190
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 846 3496 902 3505
rect 846 3431 902 3440
rect 296 2848 348 2854
rect 296 2790 348 2796
rect 308 800 336 2790
rect 860 800 888 3431
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1412 800 1440 2994
rect 1964 800 1992 3878
rect 2504 3120 2556 3126
rect 2504 3062 2556 3068
rect 2516 800 2544 3062
rect 3068 800 3096 3946
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3620 800 3648 3538
rect 4172 800 4200 4082
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4816 1442 4844 2926
rect 4724 1414 4844 1442
rect 4724 800 4752 1414
rect 5276 800 5304 3674
rect 5828 800 5856 4014
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6472 800 6500 3606
rect 6932 3602 6960 9930
rect 7116 6458 7144 17818
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7300 17338 7328 17478
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 7208 13852 7236 16934
rect 7300 16658 7328 17274
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7288 16652 7340 16658
rect 7340 16612 7420 16640
rect 7288 16594 7340 16600
rect 7392 16046 7420 16612
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7300 14482 7328 15098
rect 7484 14618 7512 16662
rect 7576 15366 7604 18362
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7288 13864 7340 13870
rect 7208 13824 7288 13852
rect 7288 13806 7340 13812
rect 7300 12442 7328 13806
rect 7484 13462 7512 14554
rect 7576 14074 7604 15302
rect 7668 15094 7696 18566
rect 7760 17134 7788 20198
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8220 18766 8248 20318
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8220 18426 8248 18566
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8220 17746 8248 18226
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 7944 17338 7972 17682
rect 8404 17626 8432 19654
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8496 17746 8524 18566
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8220 17598 8432 17626
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7668 14618 7696 15030
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7668 14074 7696 14214
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7472 13456 7524 13462
rect 7472 13398 7524 13404
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7208 6662 7236 6802
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7116 4282 7144 6394
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7208 3942 7236 6598
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7024 800 7052 3538
rect 7300 2650 7328 7686
rect 7392 4146 7420 12922
rect 7484 7546 7512 13126
rect 7576 11354 7604 14010
rect 7668 13462 7696 14010
rect 7760 14006 7788 16730
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8128 16250 8156 16594
rect 8220 16402 8248 17598
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8404 16810 8432 17138
rect 8496 16998 8524 17682
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8404 16782 8524 16810
rect 8220 16374 8340 16402
rect 8116 16244 8168 16250
rect 8168 16204 8248 16232
rect 8116 16186 8168 16192
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8220 15502 8248 16204
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8312 15314 8340 16374
rect 8390 15736 8446 15745
rect 8390 15671 8446 15680
rect 8220 15286 8340 15314
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 8220 13852 8248 15286
rect 8404 15026 8432 15671
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8312 14618 8340 14894
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7760 13824 8248 13852
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7760 13190 7788 13824
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7576 7002 7604 7754
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7576 800 7604 4082
rect 7668 4010 7696 8298
rect 7760 4010 7788 9318
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 8220 7750 8248 13466
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8220 6458 8248 7278
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 8220 5914 8248 6190
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8312 5370 8340 14418
rect 8496 11014 8524 16782
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8220 2564 8248 3946
rect 8128 2536 8248 2564
rect 8128 800 8156 2536
rect 8404 2378 8432 7142
rect 8496 4078 8524 10950
rect 8588 10266 8616 19246
rect 8680 18442 8708 22200
rect 9128 19984 9180 19990
rect 9128 19926 9180 19932
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 8956 18766 8984 19110
rect 9048 18902 9076 19110
rect 9036 18896 9088 18902
rect 9036 18838 9088 18844
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8680 18414 8800 18442
rect 8668 18352 8720 18358
rect 8668 18294 8720 18300
rect 8680 17814 8708 18294
rect 8668 17808 8720 17814
rect 8668 17750 8720 17756
rect 8772 17320 8800 18414
rect 8763 17292 8800 17320
rect 8763 17218 8791 17292
rect 8763 17190 8800 17218
rect 8772 16998 8800 17190
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8864 16658 8892 18566
rect 8956 16794 8984 18702
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 9048 17882 9076 18090
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 9048 17678 9076 17818
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 9036 17264 9088 17270
rect 9036 17206 9088 17212
rect 9048 16998 9076 17206
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8760 16448 8812 16454
rect 8760 16390 8812 16396
rect 8772 16046 8800 16390
rect 9048 16046 9076 16934
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 8772 15586 8800 15982
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8772 15558 8892 15586
rect 8864 15502 8892 15558
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8680 14618 8708 14758
rect 8772 14618 8800 15302
rect 8864 15026 8892 15438
rect 8956 15366 8984 15846
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8942 15192 8998 15201
rect 9048 15162 9076 15506
rect 8942 15127 8944 15136
rect 8996 15127 8998 15136
rect 9036 15156 9088 15162
rect 8944 15098 8996 15104
rect 9036 15098 9088 15104
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8944 14816 8996 14822
rect 8864 14776 8944 14804
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 13870 8800 14214
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8680 12374 8708 13126
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8666 12200 8722 12209
rect 8666 12135 8722 12144
rect 8680 10266 8708 12135
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8588 9722 8616 10202
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8588 6610 8616 9658
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8680 6798 8708 7210
rect 8772 6866 8800 13806
rect 8864 12481 8892 14776
rect 8944 14758 8996 14764
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8956 14006 8984 14554
rect 9048 14074 9076 15098
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 8850 12472 8906 12481
rect 8850 12407 8906 12416
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8864 8430 8892 11834
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8668 6792 8720 6798
rect 8666 6760 8668 6769
rect 8720 6760 8722 6769
rect 8666 6695 8722 6704
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8668 6656 8720 6662
rect 8588 6604 8668 6610
rect 8588 6598 8720 6604
rect 8588 6582 8708 6598
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8680 3738 8708 6394
rect 8772 6254 8800 6666
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 8312 1970 8340 2246
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 8680 800 8708 3402
rect 8772 2310 8800 5306
rect 8864 4049 8892 8366
rect 8956 7002 8984 13738
rect 9140 13462 9168 19926
rect 9232 19310 9260 22200
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9232 18222 9260 18770
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9232 17542 9260 18158
rect 9324 17610 9352 18566
rect 9416 18222 9444 18702
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9232 16794 9260 17478
rect 9324 17338 9352 17546
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9324 17134 9352 17274
rect 9508 17184 9536 19450
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9600 18154 9628 19314
rect 9692 19310 9720 19858
rect 9784 19802 9812 22200
rect 9784 19774 9996 19802
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9784 18834 9812 19246
rect 9876 18970 9904 19654
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9588 17672 9640 17678
rect 9876 17649 9904 18090
rect 9588 17614 9640 17620
rect 9862 17640 9918 17649
rect 9600 17202 9628 17614
rect 9862 17575 9918 17584
rect 9416 17156 9536 17184
rect 9588 17196 9640 17202
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 9232 16250 9260 16730
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9324 16454 9352 16594
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 9232 13308 9260 15982
rect 9140 13280 9260 13308
rect 9140 12424 9168 13280
rect 9048 12396 9168 12424
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8956 5914 8984 6938
rect 9048 5914 9076 12396
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9140 11286 9168 12174
rect 9232 12102 9260 12242
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9140 6458 9168 10202
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 8956 4146 8984 5850
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 9140 5370 9168 5782
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8850 4040 8906 4049
rect 8850 3975 8906 3984
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8772 2106 8800 2246
rect 8760 2100 8812 2106
rect 8760 2042 8812 2048
rect 9232 800 9260 12038
rect 9324 11898 9352 16390
rect 9416 13802 9444 17156
rect 9588 17138 9640 17144
rect 9496 17060 9548 17066
rect 9496 17002 9548 17008
rect 9508 16250 9536 17002
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9508 14414 9536 16186
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9692 14890 9720 15438
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9784 14482 9812 15982
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9784 14074 9812 14418
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9586 13560 9642 13569
rect 9586 13495 9642 13504
rect 9600 13444 9628 13495
rect 9508 13416 9628 13444
rect 9680 13456 9732 13462
rect 9508 13326 9536 13416
rect 9680 13398 9732 13404
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9416 12170 9444 12582
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9324 9518 9352 9998
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9324 8498 9352 9454
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9508 6984 9536 13262
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9600 11694 9628 12106
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9692 11354 9720 13398
rect 9784 13394 9812 14010
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9770 13288 9826 13297
rect 9770 13223 9772 13232
rect 9824 13223 9826 13232
rect 9772 13194 9824 13200
rect 9876 12986 9904 16390
rect 9968 15201 9996 19774
rect 10138 19272 10194 19281
rect 10138 19207 10140 19216
rect 10192 19207 10194 19216
rect 10140 19178 10192 19184
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9954 15192 10010 15201
rect 9954 15127 10010 15136
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9968 13870 9996 15030
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9954 12744 10010 12753
rect 9954 12679 10010 12688
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9784 8838 9812 12310
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9692 7002 9720 7822
rect 9416 6956 9536 6984
rect 9680 6996 9732 7002
rect 9312 6792 9364 6798
rect 9310 6760 9312 6769
rect 9364 6760 9366 6769
rect 9310 6695 9366 6704
rect 9324 6458 9352 6695
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9324 2854 9352 5034
rect 9416 3777 9444 6956
rect 9680 6938 9732 6944
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9678 6896 9734 6905
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9508 6662 9536 6802
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9600 6322 9628 6870
rect 9678 6831 9734 6840
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9508 5030 9536 5850
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9402 3768 9458 3777
rect 9402 3703 9404 3712
rect 9456 3703 9458 3712
rect 9404 3674 9456 3680
rect 9416 3643 9444 3674
rect 9508 2854 9536 4966
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9600 3398 9628 4422
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9692 3194 9720 6831
rect 9784 5370 9812 7958
rect 9876 6390 9904 12582
rect 9968 12374 9996 12679
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 9968 9994 9996 10678
rect 10060 10146 10088 18906
rect 10336 18222 10364 22200
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10152 14958 10180 18022
rect 10244 15042 10272 18090
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10336 17134 10364 18022
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10322 16688 10378 16697
rect 10322 16623 10324 16632
rect 10376 16623 10378 16632
rect 10324 16594 10376 16600
rect 10244 15014 10364 15042
rect 10140 14952 10192 14958
rect 10138 14920 10140 14929
rect 10192 14920 10194 14929
rect 10138 14855 10194 14864
rect 10336 14822 10364 15014
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10428 14278 10456 20198
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10612 19258 10640 19790
rect 10520 19242 10640 19258
rect 10508 19236 10640 19242
rect 10560 19230 10640 19236
rect 10508 19178 10560 19184
rect 10520 18970 10548 19178
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 17134 10548 17478
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10520 15094 10548 16594
rect 10612 15745 10640 18158
rect 10598 15736 10654 15745
rect 10598 15671 10654 15680
rect 10600 15632 10652 15638
rect 10600 15574 10652 15580
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10152 12714 10180 13874
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 10152 12186 10180 12650
rect 10152 12158 10272 12186
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10152 11354 10180 12038
rect 10244 11694 10272 12158
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10336 11150 10364 11562
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10520 11014 10548 12786
rect 10612 12646 10640 15574
rect 10704 14958 10732 20402
rect 10784 20256 10836 20262
rect 10782 20224 10784 20233
rect 10836 20224 10838 20233
rect 10782 20159 10838 20168
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10796 18086 10824 19110
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10888 16794 10916 22200
rect 11440 20788 11468 22200
rect 11256 20760 11468 20788
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10796 15502 10824 15914
rect 10888 15706 10916 15914
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10796 13977 10824 14826
rect 10888 14074 10916 14894
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10782 13968 10838 13977
rect 10782 13903 10838 13912
rect 10888 13530 10916 14010
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10598 12336 10654 12345
rect 10598 12271 10654 12280
rect 10508 11008 10560 11014
rect 10322 10976 10378 10985
rect 10508 10950 10560 10956
rect 10322 10911 10378 10920
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10060 10118 10180 10146
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 9968 9178 9996 9386
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10060 9110 10088 9862
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 10152 9042 10180 10118
rect 10244 9178 10272 10406
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10046 8936 10102 8945
rect 10046 8871 10102 8880
rect 10060 8634 10088 8871
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10060 7041 10088 8570
rect 10152 7449 10180 8978
rect 10244 8294 10272 8978
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10336 7970 10364 10911
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10428 10198 10456 10610
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10428 9722 10456 10134
rect 10520 10033 10548 10746
rect 10506 10024 10562 10033
rect 10506 9959 10562 9968
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10520 9330 10548 9959
rect 10244 7942 10364 7970
rect 10428 9302 10548 9330
rect 10138 7440 10194 7449
rect 10138 7375 10194 7384
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10046 7032 10102 7041
rect 10046 6967 10102 6976
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6458 10088 6802
rect 10152 6662 10180 7278
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9784 5166 9812 5306
rect 9876 5302 9904 6326
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9968 5574 9996 6054
rect 10060 5914 10088 6122
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10152 5778 10180 6598
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9876 4282 9904 5238
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9968 4026 9996 5510
rect 10152 4826 10180 5714
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10048 4208 10100 4214
rect 10046 4176 10048 4185
rect 10100 4176 10102 4185
rect 10046 4111 10102 4120
rect 10152 4078 10180 4762
rect 10244 4690 10272 7942
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10336 7342 10364 7822
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 9876 3998 9996 4026
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9692 2854 9720 2994
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9784 2514 9812 3878
rect 9876 3738 9904 3998
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9968 3194 9996 3878
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9956 3188 10008 3194
rect 10428 3176 10456 9302
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10520 8362 10548 9114
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10508 5908 10560 5914
rect 10612 5896 10640 12271
rect 10704 11234 10732 13466
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10888 12889 10916 12922
rect 10874 12880 10930 12889
rect 10874 12815 10930 12824
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10796 11694 10824 12174
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10704 11206 10824 11234
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10704 10470 10732 11018
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10560 5868 10640 5896
rect 10508 5850 10560 5856
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10520 5098 10548 5306
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10506 4040 10562 4049
rect 10506 3975 10562 3984
rect 10520 3398 10548 3975
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3738 10640 3878
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10704 3602 10732 10406
rect 10796 9178 10824 11206
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10888 9722 10916 10474
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10980 9602 11008 20334
rect 11256 20058 11284 20760
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 12084 20602 12112 22200
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 11888 19984 11940 19990
rect 11888 19926 11940 19932
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11704 19916 11756 19922
rect 11704 19858 11756 19864
rect 11150 19816 11206 19825
rect 11150 19751 11152 19760
rect 11204 19751 11206 19760
rect 11152 19722 11204 19728
rect 11256 19310 11284 19858
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11716 19514 11744 19858
rect 11900 19718 11928 19926
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11244 18828 11296 18834
rect 11244 18770 11296 18776
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11164 18426 11192 18702
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 11072 17338 11100 17682
rect 11164 17524 11192 18362
rect 11256 18358 11284 18770
rect 11716 18748 11744 19450
rect 11808 18970 11836 19654
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11900 18970 11928 19314
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11886 18864 11942 18873
rect 11992 18850 12020 20198
rect 11942 18822 12020 18850
rect 11886 18799 11942 18808
rect 11796 18760 11848 18766
rect 11716 18720 11796 18748
rect 11796 18702 11848 18708
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11244 18352 11296 18358
rect 11244 18294 11296 18300
rect 11256 17678 11284 18294
rect 11716 17882 11744 18566
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11808 17542 11836 18294
rect 11796 17536 11848 17542
rect 11164 17496 11284 17524
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 11072 16153 11100 16594
rect 11058 16144 11114 16153
rect 11058 16079 11114 16088
rect 11164 14618 11192 16730
rect 11256 15570 11284 17496
rect 11796 17478 11848 17484
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11704 17264 11756 17270
rect 11702 17232 11704 17241
rect 11756 17232 11758 17241
rect 11702 17167 11758 17176
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11520 16176 11572 16182
rect 11518 16144 11520 16153
rect 11572 16144 11574 16153
rect 11518 16079 11574 16088
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11716 15162 11744 15438
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11060 14340 11112 14346
rect 11060 14282 11112 14288
rect 11072 13870 11100 14282
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 11072 11286 11100 12786
rect 11164 12782 11192 13126
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11256 12646 11284 14758
rect 11624 14362 11652 15030
rect 11716 14482 11744 15098
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11624 14334 11744 14362
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11716 13938 11744 14334
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11348 13462 11376 13670
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 11348 13326 11376 13398
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11716 12782 11744 13670
rect 11808 13394 11836 17478
rect 11900 15094 11928 18799
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11992 16794 12020 17138
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 12084 15994 12112 20334
rect 12256 20324 12308 20330
rect 12256 20266 12308 20272
rect 12164 19848 12216 19854
rect 12162 19816 12164 19825
rect 12216 19816 12218 19825
rect 12162 19751 12218 19760
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12176 18426 12204 18702
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12176 17746 12204 18022
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12268 16096 12296 20266
rect 12360 19446 12388 20538
rect 12636 20534 12664 22200
rect 12624 20528 12676 20534
rect 12624 20470 12676 20476
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12452 18873 12480 19450
rect 12544 19310 12572 19654
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12438 18864 12494 18873
rect 12438 18799 12494 18808
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12452 18170 12480 18566
rect 12544 18290 12572 19246
rect 12808 18760 12860 18766
rect 12806 18728 12808 18737
rect 12860 18728 12862 18737
rect 12806 18663 12862 18672
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12912 18222 12940 18566
rect 12808 18216 12860 18222
rect 12452 18164 12808 18170
rect 12452 18158 12860 18164
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12452 18142 12848 18158
rect 13004 18068 13032 20198
rect 13188 18970 13216 22200
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13464 20262 13492 20334
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 19961 13584 20198
rect 13740 20074 13768 22200
rect 14292 20074 14320 22200
rect 14844 20602 14872 22200
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 15396 20534 15424 22200
rect 15384 20528 15436 20534
rect 15384 20470 15436 20476
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15752 20256 15804 20262
rect 14462 20224 14518 20233
rect 15752 20198 15804 20204
rect 14462 20159 14518 20168
rect 13740 20058 13860 20074
rect 14292 20058 14412 20074
rect 13740 20052 13872 20058
rect 13740 20046 13820 20052
rect 14292 20052 14424 20058
rect 14292 20046 14372 20052
rect 13820 19994 13872 20000
rect 14372 19994 14424 20000
rect 14476 19990 14504 20159
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15764 19990 15792 20198
rect 13728 19984 13780 19990
rect 13542 19952 13598 19961
rect 13728 19926 13780 19932
rect 14464 19984 14516 19990
rect 14464 19926 14516 19932
rect 15752 19984 15804 19990
rect 15752 19926 15804 19932
rect 15856 19938 15884 20334
rect 15948 20058 15976 22200
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 13542 19887 13598 19896
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 12728 18040 13032 18068
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12452 16590 12480 17138
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12544 16250 12572 17070
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12348 16108 12400 16114
rect 12268 16068 12348 16096
rect 12348 16050 12400 16056
rect 11992 15966 12112 15994
rect 11888 15088 11940 15094
rect 11888 15030 11940 15036
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11900 14521 11928 14554
rect 11886 14512 11942 14521
rect 11886 14447 11942 14456
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11900 13530 11928 14214
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11704 12776 11756 12782
rect 11808 12753 11836 13330
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11900 12850 11928 13262
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11704 12718 11756 12724
rect 11794 12744 11850 12753
rect 11992 12730 12020 15966
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 12084 15706 12112 15846
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12360 15502 12388 16050
rect 12438 15736 12494 15745
rect 12438 15671 12494 15680
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12176 13433 12204 14418
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 12162 13424 12218 13433
rect 12072 13388 12124 13394
rect 12162 13359 12218 13368
rect 12072 13330 12124 13336
rect 12084 12986 12112 13330
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12070 12880 12126 12889
rect 12070 12815 12072 12824
rect 12124 12815 12126 12824
rect 12072 12786 12124 12792
rect 11794 12679 11850 12688
rect 11900 12702 12020 12730
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11256 11898 11284 12310
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10538 11100 11086
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 10888 9574 11008 9602
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 4842 10824 8774
rect 10888 7750 10916 9574
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10980 8974 11008 9454
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10980 8634 11008 8910
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11072 8090 11100 8978
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 11164 7478 11192 11494
rect 11256 10674 11284 11834
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11624 11098 11652 11154
rect 11624 11070 11744 11098
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11242 10568 11298 10577
rect 11242 10503 11244 10512
rect 11296 10503 11298 10512
rect 11244 10474 11296 10480
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11624 10169 11652 10202
rect 11610 10160 11666 10169
rect 11716 10130 11744 11070
rect 11610 10095 11666 10104
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11716 9722 11744 10066
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11610 9480 11666 9489
rect 11610 9415 11666 9424
rect 11624 9110 11652 9415
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11716 8634 11744 9658
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11348 7886 11376 8366
rect 11336 7880 11388 7886
rect 11256 7840 11336 7868
rect 11256 7546 11284 7840
rect 11336 7822 11388 7828
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11164 6934 11192 7278
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10888 6322 10916 6734
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 10874 6216 10930 6225
rect 10874 6151 10876 6160
rect 10928 6151 10930 6160
rect 10876 6122 10928 6128
rect 11072 5846 11100 6258
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11716 5914 11744 6054
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10966 5128 11022 5137
rect 10966 5063 11022 5072
rect 10980 5030 11008 5063
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10796 4814 11008 4842
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10796 3534 10824 4490
rect 10980 3924 11008 4814
rect 11072 4758 11100 5170
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11072 4010 11100 4422
rect 11164 4010 11192 4422
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 10888 3896 11008 3924
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 9956 3130 10008 3136
rect 10336 3148 10456 3176
rect 9876 2961 9904 3130
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 9862 2952 9918 2961
rect 9862 2887 9918 2896
rect 10244 2650 10272 3062
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 10140 2440 10192 2446
rect 10138 2408 10140 2417
rect 10192 2408 10194 2417
rect 10138 2343 10194 2352
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9416 1902 9444 2246
rect 9772 2032 9824 2038
rect 9772 1974 9824 1980
rect 9404 1896 9456 1902
rect 9404 1838 9456 1844
rect 9784 800 9812 1974
rect 10336 800 10364 3148
rect 10520 3097 10548 3334
rect 10692 3120 10744 3126
rect 10506 3088 10562 3097
rect 10692 3062 10744 3068
rect 10506 3023 10562 3032
rect 10704 1154 10732 3062
rect 10692 1148 10744 1154
rect 10692 1090 10744 1096
rect 10888 800 10916 3896
rect 11072 3482 11100 3946
rect 11256 3618 11284 4966
rect 11624 4468 11652 5238
rect 11624 4440 11744 4468
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 11164 3602 11284 3618
rect 11532 3602 11560 3946
rect 11152 3596 11284 3602
rect 11204 3590 11284 3596
rect 11520 3596 11572 3602
rect 11152 3538 11204 3544
rect 11520 3538 11572 3544
rect 11336 3528 11388 3534
rect 11072 3476 11336 3482
rect 11072 3470 11388 3476
rect 11072 3454 11376 3470
rect 11072 3058 11100 3454
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10966 2952 11022 2961
rect 10966 2887 11022 2896
rect 10980 2854 11008 2887
rect 11164 2854 11192 3334
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 10980 2582 11008 2790
rect 11440 2582 11468 2926
rect 11716 2854 11744 4440
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 11428 2576 11480 2582
rect 11428 2518 11480 2524
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11808 2088 11836 12582
rect 11900 12322 11928 12702
rect 12268 12646 12296 13738
rect 12360 12889 12388 15438
rect 12452 15162 12480 15671
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12636 14958 12664 17206
rect 12728 15178 12756 18040
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12820 16250 12848 16934
rect 12912 16794 12940 17274
rect 13004 17134 13032 17682
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13096 17338 13124 17478
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 13096 16402 13124 17274
rect 13004 16374 13124 16402
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12820 15366 12848 15642
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12728 15150 12848 15178
rect 12624 14952 12676 14958
rect 12438 14920 12494 14929
rect 12624 14894 12676 14900
rect 12438 14855 12494 14864
rect 12532 14884 12584 14890
rect 12452 14414 12480 14855
rect 12532 14826 12584 14832
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12544 14278 12572 14826
rect 12728 14550 12756 14826
rect 12624 14544 12676 14550
rect 12622 14512 12624 14521
rect 12716 14544 12768 14550
rect 12676 14512 12678 14521
rect 12716 14486 12768 14492
rect 12622 14447 12678 14456
rect 12820 14396 12848 15150
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12728 14368 12848 14396
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12452 13258 12480 14010
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12346 12880 12402 12889
rect 12346 12815 12402 12824
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12254 12472 12310 12481
rect 12254 12407 12310 12416
rect 11900 12294 12020 12322
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11900 10810 11928 12174
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11992 10606 12020 12294
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11888 10464 11940 10470
rect 12084 10418 12112 11154
rect 11888 10406 11940 10412
rect 11900 9178 11928 10406
rect 11992 10390 12112 10418
rect 11992 10266 12020 10390
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11992 8974 12020 10202
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 12084 8838 12112 9454
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 11900 6866 11928 8774
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11992 7546 12020 8366
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11886 5808 11942 5817
rect 11886 5743 11888 5752
rect 11940 5743 11942 5752
rect 11888 5714 11940 5720
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11900 5234 11928 5510
rect 11992 5370 12020 7482
rect 12084 5778 12112 7958
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11900 4622 11928 5170
rect 11992 5030 12020 5306
rect 12084 5098 12112 5714
rect 12072 5092 12124 5098
rect 12072 5034 12124 5040
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11992 4282 12020 4626
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11980 3664 12032 3670
rect 11978 3632 11980 3641
rect 12032 3632 12034 3641
rect 11978 3567 12034 3576
rect 12084 3482 12112 4558
rect 12176 3670 12204 12038
rect 12268 8634 12296 12407
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12360 11762 12388 12242
rect 12452 12102 12480 12718
rect 12544 12374 12572 13806
rect 12636 13802 12664 14282
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12636 12850 12664 13398
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12544 11762 12572 12310
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12268 7954 12296 8434
rect 12360 8430 12388 11494
rect 12532 10192 12584 10198
rect 12530 10160 12532 10169
rect 12584 10160 12586 10169
rect 12530 10095 12586 10104
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12544 8906 12572 9658
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12346 8256 12402 8265
rect 12346 8191 12402 8200
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 12164 3664 12216 3670
rect 12164 3606 12216 3612
rect 11992 3454 12112 3482
rect 11992 3398 12020 3454
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 11440 2060 11836 2088
rect 11440 800 11468 2060
rect 12084 800 12112 2790
rect 12268 2038 12296 7210
rect 12360 5681 12388 8191
rect 12452 6882 12480 8570
rect 12636 7274 12664 12582
rect 12728 9586 12756 14368
rect 12912 13977 12940 14418
rect 12898 13968 12954 13977
rect 12898 13903 12954 13912
rect 13004 13512 13032 16374
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13096 15434 13124 16186
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 12912 13484 13032 13512
rect 12806 12880 12862 12889
rect 12806 12815 12862 12824
rect 12820 10742 12848 12815
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12912 10033 12940 13484
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13004 11354 13032 13126
rect 13096 11354 13124 14214
rect 13188 14074 13216 18090
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13174 13968 13230 13977
rect 13174 13903 13230 13912
rect 13188 13002 13216 13903
rect 13280 13190 13308 18090
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13188 12974 13308 13002
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13004 10606 13032 11290
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 12898 10024 12954 10033
rect 12898 9959 12954 9968
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9654 12940 9862
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12820 9042 12848 9318
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 13004 8956 13032 10542
rect 13096 9518 13124 11290
rect 13174 10160 13230 10169
rect 13174 10095 13230 10104
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13188 9110 13216 10095
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13004 8928 13216 8956
rect 13280 8945 13308 12974
rect 13372 12374 13400 18770
rect 13636 17808 13688 17814
rect 13636 17750 13688 17756
rect 13648 17649 13676 17750
rect 13634 17640 13690 17649
rect 13634 17575 13690 17584
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16794 13492 16934
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13464 16114 13492 16730
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13464 15065 13492 16050
rect 13450 15056 13506 15065
rect 13450 14991 13506 15000
rect 13556 14498 13584 16458
rect 13740 14940 13768 19926
rect 15660 19916 15712 19922
rect 15856 19910 15976 19938
rect 15660 19858 15712 19864
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 13832 19514 13860 19790
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13832 19378 13860 19450
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14186 19272 14242 19281
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13924 18358 13952 19178
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 14016 18426 14044 18770
rect 14108 18630 14136 19246
rect 14186 19207 14242 19216
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 14108 18222 14136 18566
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 13832 16998 13860 18158
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14108 17134 14136 17614
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13832 15502 13860 15914
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13464 14470 13584 14498
rect 13648 14912 13768 14940
rect 13464 13530 13492 14470
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13556 13938 13584 14350
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13556 13462 13584 13670
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13464 12918 13492 13330
rect 13648 13326 13676 14912
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13740 14074 13768 14758
rect 13832 14618 13860 14758
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13924 14498 13952 14962
rect 13832 14482 13952 14498
rect 13820 14476 13952 14482
rect 13872 14470 13952 14476
rect 13820 14418 13872 14424
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13832 14006 13860 14418
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 14016 13734 14044 16934
rect 14108 16658 14136 17070
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13464 9382 13492 10474
rect 13556 10266 13584 10610
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13556 9450 13584 10066
rect 13648 9466 13676 13126
rect 13740 12714 13768 13466
rect 14016 13190 14044 13670
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14108 12782 14136 14758
rect 14200 14090 14228 19207
rect 14660 18970 14688 19654
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14752 18850 14780 19110
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 14752 18834 14964 18850
rect 14464 18828 14516 18834
rect 14752 18828 14976 18834
rect 14752 18822 14924 18828
rect 14464 18770 14516 18776
rect 14924 18770 14976 18776
rect 14372 17264 14424 17270
rect 14372 17206 14424 17212
rect 14384 16794 14412 17206
rect 14476 16998 14504 18770
rect 15212 18766 15240 19314
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15212 18154 15240 18702
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 14830 17776 14886 17785
rect 14648 17740 14700 17746
rect 15304 17746 15332 19654
rect 15396 18698 15424 19790
rect 15672 19514 15700 19858
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15856 18902 15884 19790
rect 15948 19514 15976 19910
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 16040 19242 16068 20198
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15764 17921 15792 18566
rect 15856 18426 15884 18838
rect 16316 18737 16344 20538
rect 16394 20496 16450 20505
rect 16394 20431 16450 20440
rect 16408 19922 16436 20431
rect 16500 20074 16528 22200
rect 16500 20058 16620 20074
rect 16500 20052 16632 20058
rect 16500 20046 16580 20052
rect 16580 19994 16632 20000
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16302 18728 16358 18737
rect 16302 18663 16358 18672
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15750 17912 15806 17921
rect 15750 17847 15806 17856
rect 15764 17746 15792 17847
rect 14830 17711 14886 17720
rect 15292 17740 15344 17746
rect 14648 17682 14700 17688
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14568 16794 14596 17478
rect 14660 17338 14688 17682
rect 14844 17542 14872 17711
rect 15292 17682 15344 17688
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15750 17640 15806 17649
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 15580 17338 15608 17614
rect 15750 17575 15806 17584
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 14740 17264 14792 17270
rect 14740 17206 14792 17212
rect 14648 17060 14700 17066
rect 14648 17002 14700 17008
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14464 15088 14516 15094
rect 14370 15056 14426 15065
rect 14464 15030 14516 15036
rect 14370 14991 14372 15000
rect 14424 14991 14426 15000
rect 14372 14962 14424 14968
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14292 14482 14320 14894
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14280 14272 14332 14278
rect 14332 14220 14412 14226
rect 14280 14214 14412 14220
rect 14292 14198 14412 14214
rect 14200 14062 14320 14090
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11801 14228 12038
rect 14186 11792 14242 11801
rect 14186 11727 14242 11736
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13832 11082 13860 11562
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13740 9994 13768 10542
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 10266 13860 10406
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13740 9586 13768 9930
rect 13924 9654 13952 10542
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13544 9444 13596 9450
rect 13648 9438 13952 9466
rect 13544 9386 13596 9392
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 7002 12572 7142
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12452 6854 12572 6882
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12452 5778 12480 6598
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12346 5672 12402 5681
rect 12346 5607 12348 5616
rect 12400 5607 12402 5616
rect 12348 5578 12400 5584
rect 12360 5547 12388 5578
rect 12346 5128 12402 5137
rect 12346 5063 12348 5072
rect 12400 5063 12402 5072
rect 12348 5034 12400 5040
rect 12452 4622 12480 5714
rect 12544 5692 12572 6854
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12636 5846 12664 6054
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12544 5664 12664 5692
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12544 4758 12572 5034
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12636 4486 12664 5664
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12532 4072 12584 4078
rect 12438 4040 12494 4049
rect 12532 4014 12584 4020
rect 12438 3975 12494 3984
rect 12452 3942 12480 3975
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12544 2446 12572 4014
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12256 2032 12308 2038
rect 12256 1974 12308 1980
rect 12636 800 12664 3878
rect 12728 2514 12756 8774
rect 13084 6384 13136 6390
rect 13084 6326 13136 6332
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12912 5846 12940 6054
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12820 2530 12848 5782
rect 13004 5370 13032 6122
rect 13096 5574 13124 6326
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12912 4078 12940 4558
rect 13188 4146 13216 8928
rect 13266 8936 13322 8945
rect 13266 8871 13322 8880
rect 13464 8294 13492 9318
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13556 7342 13584 9386
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13740 8566 13768 8910
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13740 8022 13768 8502
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13648 7410 13676 7686
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13372 7002 13400 7210
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13280 5030 13308 6938
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13372 5234 13400 6054
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13464 5098 13492 7142
rect 13648 6934 13676 7346
rect 13636 6928 13688 6934
rect 13636 6870 13688 6876
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12912 3738 12940 4014
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 13004 3398 13032 4082
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13464 3398 13492 3946
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13464 3058 13492 3334
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13556 2990 13584 6326
rect 13648 6322 13676 6870
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13924 6610 13952 9438
rect 14016 8090 14044 10950
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14108 9897 14136 9998
rect 14188 9920 14240 9926
rect 14094 9888 14150 9897
rect 14188 9862 14240 9868
rect 14094 9823 14150 9832
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 14108 7546 14136 9590
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14108 7342 14136 7482
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14200 6798 14228 9862
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13648 4690 13676 6122
rect 13740 5710 13768 6598
rect 13924 6582 14228 6610
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13740 5234 13768 5646
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13648 4010 13676 4422
rect 13832 4078 13860 6190
rect 13910 5672 13966 5681
rect 13910 5607 13912 5616
rect 13964 5607 13966 5616
rect 13912 5578 13964 5584
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14108 4622 14136 4966
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13912 3664 13964 3670
rect 13726 3632 13782 3641
rect 13912 3606 13964 3612
rect 13726 3567 13782 3576
rect 13740 3466 13768 3567
rect 13924 3505 13952 3606
rect 13910 3496 13966 3505
rect 13728 3460 13780 3466
rect 13910 3431 13966 3440
rect 13728 3402 13780 3408
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 12820 2514 12940 2530
rect 14108 2514 14136 4422
rect 14200 2854 14228 6582
rect 14292 3738 14320 14062
rect 14384 13870 14412 14198
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14384 13326 14412 13806
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14384 11830 14412 12786
rect 14476 12646 14504 15030
rect 14568 13530 14596 15438
rect 14660 13938 14688 17002
rect 14752 16590 14780 17206
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 15212 16658 15240 17138
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15384 16720 15436 16726
rect 15384 16662 15436 16668
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14752 16046 14780 16526
rect 15396 16182 15424 16662
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 15384 16176 15436 16182
rect 15384 16118 15436 16124
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 15384 15904 15436 15910
rect 15488 15892 15516 16458
rect 15580 16046 15608 16934
rect 15764 16590 15792 17575
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15856 16590 15884 17138
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15568 15904 15620 15910
rect 15488 15864 15568 15892
rect 15384 15846 15436 15852
rect 15568 15846 15620 15852
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15396 15706 15424 15846
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15672 15144 15700 16458
rect 15764 15416 15792 16526
rect 15856 16114 15884 16526
rect 15948 16250 15976 16934
rect 16040 16794 16068 16934
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 16040 15473 16068 16458
rect 16316 16454 16344 18663
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16132 15706 16160 16390
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16026 15464 16082 15473
rect 15764 15388 15884 15416
rect 16026 15399 16082 15408
rect 15488 15116 15700 15144
rect 15488 14929 15516 15116
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15474 14920 15530 14929
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 15384 14884 15436 14890
rect 15474 14855 15530 14864
rect 15384 14826 15436 14832
rect 14752 14278 14780 14826
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14832 14544 14884 14550
rect 14832 14486 14884 14492
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14660 12481 14688 13874
rect 14752 12850 14780 14214
rect 14844 14074 14872 14486
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15212 14074 15240 14350
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15200 13864 15252 13870
rect 15198 13832 15200 13841
rect 15252 13832 15254 13841
rect 15198 13767 15254 13776
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14646 12472 14702 12481
rect 14476 12442 14646 12458
rect 14464 12436 14646 12442
rect 14516 12430 14646 12436
rect 14817 12464 15113 12484
rect 14646 12407 14702 12416
rect 14464 12378 14516 12384
rect 15212 12306 15240 13330
rect 15304 12714 15332 14214
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14372 11688 14424 11694
rect 14372 11630 14424 11636
rect 14384 11234 14412 11630
rect 14384 11206 14504 11234
rect 14476 11082 14504 11206
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14384 10674 14412 11018
rect 14568 10810 14596 12242
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14660 11218 14688 12174
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14384 9722 14412 10406
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14476 9926 14504 10202
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14554 9888 14610 9897
rect 14554 9823 14610 9832
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14568 9654 14596 9823
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14476 8974 14504 9522
rect 14660 9466 14688 10678
rect 14752 10606 14780 11630
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 14738 10160 14794 10169
rect 14738 10095 14794 10104
rect 14752 10062 14780 10095
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14568 9438 14688 9466
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14384 8634 14412 8910
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14476 8362 14504 8910
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14372 8288 14424 8294
rect 14424 8236 14504 8242
rect 14372 8230 14504 8236
rect 14384 8214 14504 8230
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 14384 6866 14412 7210
rect 14476 7206 14504 8214
rect 14568 8090 14596 9438
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14660 9110 14688 9318
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14384 6458 14412 6802
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14384 5302 14412 6394
rect 14476 6118 14504 7142
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5370 14504 6054
rect 14568 5914 14596 6598
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14660 5794 14688 8230
rect 14752 8090 14780 9862
rect 14830 9752 14886 9761
rect 14830 9687 14886 9696
rect 14844 9625 14872 9687
rect 14830 9616 14886 9625
rect 14830 9551 14886 9560
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 15212 7886 15240 11494
rect 15304 10266 15332 11630
rect 15396 11354 15424 14826
rect 15488 13734 15516 14855
rect 15672 14600 15700 14962
rect 15580 14572 15700 14600
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13297 15516 13670
rect 15474 13288 15530 13297
rect 15474 13223 15530 13232
rect 15580 12306 15608 14572
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15672 13258 15700 14418
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15764 14006 15792 14214
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15752 13864 15804 13870
rect 15856 13852 15884 15388
rect 15804 13824 15884 13852
rect 15936 13864 15988 13870
rect 15752 13806 15804 13812
rect 16132 13841 16160 15642
rect 15936 13806 15988 13812
rect 16118 13832 16174 13841
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15750 13016 15806 13025
rect 15856 12986 15884 13262
rect 15750 12951 15752 12960
rect 15804 12951 15806 12960
rect 15844 12980 15896 12986
rect 15752 12922 15804 12928
rect 15844 12922 15896 12928
rect 15948 12730 15976 13806
rect 16118 13767 16174 13776
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 12918 16252 13670
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 15764 12702 15976 12730
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15580 11558 15608 12242
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15488 11150 15516 11290
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15764 10266 15792 12702
rect 16316 12646 16344 16390
rect 16408 15910 16436 19858
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16592 19310 16620 19790
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16488 18692 16540 18698
rect 16488 18634 16540 18640
rect 16500 18358 16528 18634
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16488 18352 16540 18358
rect 16488 18294 16540 18300
rect 16592 17814 16620 18566
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16580 17808 16632 17814
rect 16580 17750 16632 17756
rect 16592 17202 16620 17750
rect 16684 17338 16712 18158
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16776 16776 16804 17818
rect 16684 16748 16804 16776
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16500 15366 16528 15438
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16500 15094 16528 15302
rect 16488 15088 16540 15094
rect 16488 15030 16540 15036
rect 16592 14618 16620 15302
rect 16684 15094 16712 16748
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16684 14521 16712 14554
rect 16670 14512 16726 14521
rect 16670 14447 16726 14456
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 13394 16436 14214
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 15948 12442 15976 12582
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 16040 12322 16068 12582
rect 15948 12294 16068 12322
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15290 9616 15346 9625
rect 15290 9551 15346 9560
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14568 5766 14688 5794
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14476 2990 14504 5102
rect 14568 3097 14596 5766
rect 14752 4486 14780 6870
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14832 5840 14884 5846
rect 14830 5808 14832 5817
rect 14884 5808 14886 5817
rect 14830 5743 14886 5752
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14752 3534 14780 3878
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14660 3194 14688 3470
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 14554 3088 14610 3097
rect 14554 3023 14610 3032
rect 14752 2990 14780 3470
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 14646 2816 14702 2825
rect 12716 2508 12768 2514
rect 12820 2508 12952 2514
rect 12820 2502 12900 2508
rect 12716 2450 12768 2456
rect 12900 2450 12952 2456
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 14108 2378 14136 2450
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13188 800 13216 2246
rect 13740 800 13768 2246
rect 14200 1601 14228 2790
rect 14646 2751 14702 2760
rect 14660 2514 14688 2751
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14186 1592 14242 1601
rect 14186 1527 14242 1536
rect 14280 1148 14332 1154
rect 14280 1090 14332 1096
rect 14292 800 14320 1090
rect 14844 800 14872 2246
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13726 0 13782 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15304 649 15332 9551
rect 15764 8956 15792 10202
rect 15856 10062 15884 10542
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15844 8968 15896 8974
rect 15764 8928 15844 8956
rect 15844 8910 15896 8916
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15764 8362 15792 8502
rect 15752 8356 15804 8362
rect 15752 8298 15804 8304
rect 15658 7848 15714 7857
rect 15658 7783 15714 7792
rect 15672 6225 15700 7783
rect 15856 7002 15884 8910
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 6322 15792 6598
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15856 6254 15884 6938
rect 15844 6248 15896 6254
rect 15658 6216 15714 6225
rect 15844 6190 15896 6196
rect 15658 6151 15714 6160
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15488 4185 15516 4626
rect 15474 4176 15530 4185
rect 15474 4111 15530 4120
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15396 800 15424 3878
rect 15580 2514 15608 5646
rect 15672 4690 15700 6151
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15856 5098 15884 5646
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15672 2582 15700 4626
rect 15856 4622 15884 5034
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15948 4026 15976 12294
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16040 10538 16068 11630
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 16040 9042 16068 10474
rect 16132 10470 16160 10746
rect 16592 10577 16620 13806
rect 16776 13025 16804 14758
rect 16762 13016 16818 13025
rect 16762 12951 16818 12960
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 11286 16712 12038
rect 16672 11280 16724 11286
rect 16672 11222 16724 11228
rect 16578 10568 16634 10577
rect 16578 10503 16634 10512
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16132 9382 16160 10406
rect 16316 10130 16344 10406
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 16132 8566 16160 9318
rect 16408 9178 16436 9454
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16486 8936 16542 8945
rect 16486 8871 16542 8880
rect 16120 8560 16172 8566
rect 16120 8502 16172 8508
rect 16132 6866 16160 8502
rect 16500 8498 16528 8871
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16592 8362 16620 10503
rect 16868 9160 16896 19246
rect 17052 18970 17080 22200
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 15706 16988 16934
rect 17052 16454 17080 18022
rect 17144 16998 17172 20198
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17236 17882 17264 18226
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17144 16697 17172 16730
rect 17130 16688 17186 16697
rect 17130 16623 17186 16632
rect 17236 16590 17264 17138
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 17052 13938 17080 15574
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16960 12442 16988 13466
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 16868 9132 16988 9160
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16684 8498 16712 8910
rect 16776 8634 16804 9046
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16684 8090 16712 8434
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16776 7954 16804 8570
rect 16868 8430 16896 8842
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16316 7546 16344 7890
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16316 6322 16344 7482
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 16408 6798 16436 7210
rect 16500 7002 16528 7754
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16408 6390 16436 6734
rect 16396 6384 16448 6390
rect 16396 6326 16448 6332
rect 16776 6322 16804 7142
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16868 6118 16896 6394
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 16040 4146 16068 5510
rect 16408 5370 16436 5646
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16120 5296 16172 5302
rect 16118 5264 16120 5273
rect 16172 5264 16174 5273
rect 16118 5199 16174 5208
rect 16408 5166 16436 5306
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16408 4690 16436 5102
rect 16592 5098 16620 5510
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16684 4554 16712 5714
rect 16868 4758 16896 6054
rect 16856 4752 16908 4758
rect 16856 4694 16908 4700
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 16028 4140 16080 4146
rect 16028 4082 16080 4088
rect 16132 4078 16160 4422
rect 15856 3998 15976 4026
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16396 4004 16448 4010
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15764 3602 15792 3878
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15856 3466 15884 3998
rect 16396 3946 16448 3952
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15580 2106 15608 2450
rect 15568 2100 15620 2106
rect 15568 2042 15620 2048
rect 15948 800 15976 3878
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16224 2009 16252 2518
rect 16210 2000 16266 2009
rect 16408 1986 16436 3946
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16684 2990 16712 3470
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16500 2446 16528 2858
rect 16960 2650 16988 9132
rect 17052 4049 17080 13874
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17144 12850 17172 12922
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17328 12186 17356 19858
rect 17696 18970 17724 22200
rect 18248 20890 18276 22200
rect 18156 20862 18276 20890
rect 18156 20602 18184 20862
rect 18694 20768 18750 20777
rect 18282 20700 18578 20720
rect 18694 20703 18750 20712
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 17788 20398 17816 20538
rect 18616 20505 18644 20538
rect 18602 20496 18658 20505
rect 18602 20431 18658 20440
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17880 19378 17908 19858
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17590 17912 17646 17921
rect 17590 17847 17646 17856
rect 17604 17678 17632 17847
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17696 17542 17724 18770
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 17880 17921 17908 18158
rect 17866 17912 17922 17921
rect 17866 17847 17922 17856
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17696 16998 17724 17478
rect 17880 17202 17908 17847
rect 17972 17270 18000 20198
rect 18432 19922 18460 20334
rect 18420 19916 18472 19922
rect 18420 19858 18472 19864
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18052 19304 18104 19310
rect 18050 19272 18052 19281
rect 18104 19272 18106 19281
rect 18050 19207 18106 19216
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17972 16046 18000 17070
rect 18064 17066 18092 18294
rect 18156 18154 18184 18702
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18144 18148 18196 18154
rect 18144 18090 18196 18096
rect 18142 18048 18198 18057
rect 18142 17983 18198 17992
rect 18052 17060 18104 17066
rect 18052 17002 18104 17008
rect 18156 16794 18184 17983
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18248 17649 18276 17682
rect 18234 17640 18290 17649
rect 18234 17575 18290 17584
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18248 16538 18276 17206
rect 18156 16510 18276 16538
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17512 14414 17540 15438
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17420 12442 17448 13942
rect 17590 13832 17646 13841
rect 17590 13767 17646 13776
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17236 12158 17356 12186
rect 17236 10130 17264 12158
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11694 17356 12038
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17316 11688 17368 11694
rect 17512 11665 17540 11698
rect 17316 11630 17368 11636
rect 17498 11656 17554 11665
rect 17498 11591 17554 11600
rect 17498 11248 17554 11257
rect 17498 11183 17554 11192
rect 17512 11150 17540 11183
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17420 9994 17448 10406
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17328 9178 17356 9522
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17144 7342 17172 7686
rect 17132 7336 17184 7342
rect 17512 7290 17540 9862
rect 17132 7278 17184 7284
rect 17144 6866 17172 7278
rect 17420 7262 17540 7290
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17236 6934 17264 7142
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17420 6390 17448 7262
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17512 7002 17540 7142
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17408 6384 17460 6390
rect 17408 6326 17460 6332
rect 17500 5840 17552 5846
rect 17500 5782 17552 5788
rect 17512 5030 17540 5782
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17132 4072 17184 4078
rect 17038 4040 17094 4049
rect 17132 4014 17184 4020
rect 17038 3975 17094 3984
rect 17144 3670 17172 4014
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17328 2650 17356 4558
rect 17512 4214 17540 4966
rect 17500 4208 17552 4214
rect 17500 4150 17552 4156
rect 17408 4004 17460 4010
rect 17408 3946 17460 3952
rect 17420 3738 17448 3946
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17512 3194 17540 3538
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17512 2446 17540 3130
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 16408 1958 16528 1986
rect 16210 1935 16212 1944
rect 16264 1935 16266 1944
rect 16212 1906 16264 1912
rect 16224 1875 16252 1906
rect 16500 800 16528 1958
rect 17052 800 17080 2246
rect 17604 2009 17632 13767
rect 17696 13190 17724 14214
rect 17788 13530 17816 14418
rect 17880 14278 17908 14418
rect 18064 14414 18092 14758
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17972 14006 18000 14214
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17682 12880 17738 12889
rect 17788 12850 17816 13466
rect 17682 12815 17738 12824
rect 17776 12844 17828 12850
rect 17696 10198 17724 12815
rect 17776 12786 17828 12792
rect 17788 12238 17816 12786
rect 17880 12646 17908 13466
rect 17972 12714 18000 13670
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18064 12782 18092 13126
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17866 12336 17922 12345
rect 17866 12271 17922 12280
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17696 8090 17724 10134
rect 17788 10062 17816 10950
rect 17880 10810 17908 12271
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17972 11393 18000 11834
rect 18156 11762 18184 16510
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18328 15904 18380 15910
rect 18328 15846 18380 15852
rect 18340 15609 18368 15846
rect 18326 15600 18382 15609
rect 18326 15535 18382 15544
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18616 14929 18644 20334
rect 18708 20058 18736 20703
rect 18800 20534 18828 22200
rect 18878 22199 18934 22208
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18892 20262 18920 22199
rect 18970 20360 19026 20369
rect 18970 20295 19026 20304
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18984 20058 19012 20295
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18970 19952 19026 19961
rect 18788 19916 18840 19922
rect 18970 19887 19026 19896
rect 18788 19858 18840 19864
rect 18800 19378 18828 19858
rect 18984 19854 19012 19887
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18788 19236 18840 19242
rect 18788 19178 18840 19184
rect 18972 19236 19024 19242
rect 19076 19224 19104 22607
rect 19338 22200 19394 23000
rect 19890 22200 19946 23000
rect 20442 22200 20498 23000
rect 20994 22200 21050 23000
rect 21546 22200 21602 23000
rect 22098 22200 22154 23000
rect 22650 22200 22706 23000
rect 19352 21842 19380 22200
rect 19352 21814 19472 21842
rect 19338 21720 19394 21729
rect 19338 21655 19394 21664
rect 19352 20602 19380 21655
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19444 20466 19472 21814
rect 19904 21434 19932 22200
rect 19812 21406 19932 21434
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19168 19990 19196 20334
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 19168 19446 19196 19654
rect 19156 19440 19208 19446
rect 19156 19382 19208 19388
rect 19024 19196 19104 19224
rect 18972 19178 19024 19184
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18708 18465 18736 18566
rect 18694 18456 18750 18465
rect 18694 18391 18750 18400
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18708 17785 18736 18158
rect 18694 17776 18750 17785
rect 18694 17711 18750 17720
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18708 17241 18736 17614
rect 18694 17232 18750 17241
rect 18694 17167 18750 17176
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18708 16658 18736 16730
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18602 14920 18658 14929
rect 18602 14855 18604 14864
rect 18656 14855 18658 14864
rect 18604 14826 18656 14832
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18418 13832 18474 13841
rect 18418 13767 18474 13776
rect 18432 13734 18460 13767
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18328 13388 18380 13394
rect 18328 13330 18380 13336
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18340 13297 18368 13330
rect 18512 13320 18564 13326
rect 18326 13288 18382 13297
rect 18326 13223 18382 13232
rect 18510 13288 18512 13297
rect 18564 13288 18566 13297
rect 18510 13223 18566 13232
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18616 12986 18644 13330
rect 18708 13326 18736 13874
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18708 12986 18736 13262
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18510 12744 18566 12753
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18248 12374 18276 12582
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 18340 12170 18368 12718
rect 18510 12679 18566 12688
rect 18524 12374 18552 12679
rect 18616 12646 18644 12786
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18616 12374 18644 12582
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18328 12164 18380 12170
rect 18328 12106 18380 12112
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18326 11792 18382 11801
rect 18144 11756 18196 11762
rect 18326 11727 18328 11736
rect 18144 11698 18196 11704
rect 18380 11727 18382 11736
rect 18328 11698 18380 11704
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 17958 11384 18014 11393
rect 17958 11319 18014 11328
rect 18432 11257 18460 11630
rect 18616 11354 18644 11834
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18418 11248 18474 11257
rect 18474 11206 18644 11234
rect 18708 11218 18736 12174
rect 18418 11183 18474 11192
rect 18616 11150 18644 11206
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17866 10704 17922 10713
rect 17866 10639 17922 10648
rect 18052 10668 18104 10674
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17788 9518 17816 9998
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17788 9178 17816 9454
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17696 7342 17724 8026
rect 17880 7868 17908 10639
rect 18052 10610 18104 10616
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17972 9110 18000 9590
rect 18064 9450 18092 10610
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 18156 8498 18184 10406
rect 18524 10033 18552 10406
rect 18708 10062 18736 10610
rect 18604 10056 18656 10062
rect 18510 10024 18566 10033
rect 18604 9998 18656 10004
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18510 9959 18566 9968
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18326 9480 18382 9489
rect 18248 8945 18276 9454
rect 18326 9415 18382 9424
rect 18512 9444 18564 9450
rect 18234 8936 18290 8945
rect 18340 8906 18368 9415
rect 18512 9386 18564 9392
rect 18524 9178 18552 9386
rect 18616 9178 18644 9998
rect 18708 9722 18736 9998
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18602 9072 18658 9081
rect 18602 9007 18658 9016
rect 18234 8871 18290 8880
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18616 8838 18644 9007
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 17958 8120 18014 8129
rect 17958 8055 18014 8064
rect 17972 8022 18000 8055
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 17788 7840 17908 7868
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17696 6458 17724 7278
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17590 2000 17646 2009
rect 17590 1935 17646 1944
rect 17696 800 17724 3878
rect 15290 640 15346 649
rect 15290 575 15346 584
rect 15382 0 15438 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17682 0 17738 800
rect 17788 241 17816 7840
rect 17960 7812 18012 7818
rect 17880 7772 17960 7800
rect 17880 7410 17908 7772
rect 17960 7754 18012 7760
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17880 6934 17908 7346
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17880 5370 17908 6870
rect 18156 6338 18184 8298
rect 18708 8022 18736 8910
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18616 6866 18644 7822
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18156 6310 18276 6338
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17972 5574 18000 6122
rect 18156 5817 18184 6190
rect 18142 5808 18198 5817
rect 18142 5743 18198 5752
rect 18248 5658 18276 6310
rect 18616 6254 18644 6802
rect 18604 6248 18656 6254
rect 18708 6225 18736 7958
rect 18604 6190 18656 6196
rect 18694 6216 18750 6225
rect 18156 5630 18276 5658
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17972 5234 18000 5510
rect 18156 5250 18184 5630
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 17960 5228 18012 5234
rect 18156 5222 18276 5250
rect 17960 5170 18012 5176
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17972 4865 18000 5034
rect 17958 4856 18014 4865
rect 17958 4791 18014 4800
rect 18156 4690 18184 5102
rect 18248 4690 18276 5222
rect 18616 5166 18644 6190
rect 18694 6151 18750 6160
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18616 5030 18644 5102
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 17958 4584 18014 4593
rect 17958 4519 18014 4528
rect 17972 4486 18000 4519
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 17958 4312 18014 4321
rect 18282 4304 18578 4324
rect 17958 4247 17960 4256
rect 18012 4247 18014 4256
rect 17960 4218 18012 4224
rect 17972 4078 18000 4218
rect 18708 4078 18736 6151
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18050 3632 18106 3641
rect 18050 3567 18106 3576
rect 18064 2836 18092 3567
rect 18156 3534 18184 4014
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18156 2990 18184 3470
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18616 3058 18644 3606
rect 18800 3194 18828 19178
rect 18984 18902 19012 19178
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 19076 18154 19104 18226
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 19076 17610 19104 18090
rect 19064 17604 19116 17610
rect 19064 17546 19116 17552
rect 18880 16652 18932 16658
rect 18880 16594 18932 16600
rect 18892 16250 18920 16594
rect 18972 16584 19024 16590
rect 18972 16526 19024 16532
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 18984 15706 19012 16526
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 19076 15434 19104 16526
rect 19168 16114 19196 19382
rect 19260 17513 19288 19722
rect 19536 19310 19564 20334
rect 19812 20330 19840 21406
rect 19890 21312 19946 21321
rect 19890 21247 19946 21256
rect 19904 20602 19932 21247
rect 19892 20596 19944 20602
rect 19892 20538 19944 20544
rect 19800 20324 19852 20330
rect 19800 20266 19852 20272
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19904 19417 19932 19654
rect 19890 19408 19946 19417
rect 19890 19343 19946 19352
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 19800 19236 19852 19242
rect 19800 19178 19852 19184
rect 19432 18760 19484 18766
rect 19352 18720 19432 18748
rect 19352 18290 19380 18720
rect 19432 18702 19484 18708
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19444 18086 19472 18226
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19246 17504 19302 17513
rect 19246 17439 19302 17448
rect 19444 17134 19472 18022
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19352 15434 19380 16934
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19432 16176 19484 16182
rect 19432 16118 19484 16124
rect 19064 15428 19116 15434
rect 19064 15370 19116 15376
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19076 14958 19104 15370
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18892 13870 18920 14758
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18892 13326 18920 13806
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18892 12646 18920 13262
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18984 12782 19012 13126
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18892 11132 18920 12310
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18984 11354 19012 11562
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 19076 11286 19104 12650
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 18892 11104 19104 11132
rect 18970 10976 19026 10985
rect 18970 10911 19026 10920
rect 18878 10840 18934 10849
rect 18878 10775 18934 10784
rect 18892 7342 18920 10775
rect 18984 9926 19012 10911
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18970 9208 19026 9217
rect 18970 9143 19026 9152
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18984 6730 19012 9143
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18892 5914 18920 6190
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18880 5160 18932 5166
rect 18880 5102 18932 5108
rect 18892 4826 18920 5102
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18144 2984 18196 2990
rect 18420 2984 18472 2990
rect 18144 2926 18196 2932
rect 18418 2952 18420 2961
rect 18472 2952 18474 2961
rect 18418 2887 18474 2896
rect 18144 2848 18196 2854
rect 18064 2808 18144 2836
rect 18144 2790 18196 2796
rect 18156 2553 18184 2790
rect 18142 2544 18198 2553
rect 18142 2479 18198 2488
rect 18144 2372 18196 2378
rect 18144 2314 18196 2320
rect 18156 1170 18184 2314
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18156 1142 18276 1170
rect 18248 800 18276 1142
rect 18800 800 18828 2246
rect 18892 1057 18920 4626
rect 18984 4282 19012 6394
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 19076 3505 19104 11104
rect 19168 10266 19196 12378
rect 19260 12374 19288 14826
rect 19444 14618 19472 16118
rect 19536 16046 19564 16526
rect 19616 16516 19668 16522
rect 19616 16458 19668 16464
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19628 15706 19656 16458
rect 19720 16114 19748 16934
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19720 15638 19748 16050
rect 19708 15632 19760 15638
rect 19708 15574 19760 15580
rect 19720 15502 19748 15574
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19444 12442 19472 13330
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19260 11354 19288 11494
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19352 10674 19380 11086
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19352 9518 19380 10610
rect 19536 10470 19564 14486
rect 19628 11354 19656 15370
rect 19812 11898 19840 19178
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19904 14414 19932 14758
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19904 13870 19932 14350
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19616 10532 19668 10538
rect 19616 10474 19668 10480
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19628 9994 19656 10474
rect 19720 10266 19748 11086
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19616 9988 19668 9994
rect 19616 9930 19668 9936
rect 19628 9722 19656 9930
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 19892 9716 19944 9722
rect 19892 9658 19944 9664
rect 19340 9512 19392 9518
rect 19154 9480 19210 9489
rect 19340 9454 19392 9460
rect 19154 9415 19210 9424
rect 19168 9178 19196 9415
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19168 8090 19196 9114
rect 19260 8634 19288 9318
rect 19352 8650 19380 9454
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19248 8628 19300 8634
rect 19352 8622 19472 8650
rect 19248 8570 19300 8576
rect 19260 8498 19288 8570
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19168 7002 19196 8026
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 19062 3496 19118 3505
rect 19062 3431 19118 3440
rect 19168 2514 19196 6666
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 19168 2417 19196 2450
rect 19260 2446 19288 7210
rect 19352 3058 19380 8502
rect 19444 8498 19472 8622
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19812 8430 19840 8774
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19904 7206 19932 9658
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19444 2990 19472 5646
rect 19536 4758 19564 7142
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19616 5024 19668 5030
rect 19616 4966 19668 4972
rect 19524 4752 19576 4758
rect 19524 4694 19576 4700
rect 19628 4622 19656 4966
rect 19720 4826 19748 6802
rect 19904 5914 19932 7142
rect 19892 5908 19944 5914
rect 19892 5850 19944 5856
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19812 4826 19840 5510
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19708 4616 19760 4622
rect 19708 4558 19760 4564
rect 19524 4480 19576 4486
rect 19720 4434 19748 4558
rect 19576 4428 19748 4434
rect 19524 4422 19748 4428
rect 19536 4406 19748 4422
rect 19904 4282 19932 4626
rect 19996 4622 20024 19654
rect 20352 18896 20404 18902
rect 20352 18838 20404 18844
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 20088 18222 20116 18566
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20180 17882 20208 18022
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 20272 17202 20300 18770
rect 20364 17882 20392 18838
rect 20456 18714 20484 22200
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20548 18970 20576 20334
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20640 18873 20668 20198
rect 21008 20058 21036 22200
rect 20996 20052 21048 20058
rect 20996 19994 21048 20000
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20626 18864 20682 18873
rect 20626 18799 20682 18808
rect 20456 18686 20576 18714
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20352 17876 20404 17882
rect 20352 17818 20404 17824
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20352 17128 20404 17134
rect 20456 17105 20484 18566
rect 20548 18426 20576 18686
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20732 17814 20760 19858
rect 21560 19854 21588 22200
rect 21548 19848 21600 19854
rect 21270 19816 21326 19825
rect 21548 19790 21600 19796
rect 21270 19751 21326 19760
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 20904 18352 20956 18358
rect 20904 18294 20956 18300
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20824 17882 20852 18158
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 20720 17808 20772 17814
rect 20720 17750 20772 17756
rect 20916 17746 20944 18294
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20352 17070 20404 17076
rect 20442 17096 20498 17105
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 20088 14618 20116 15846
rect 20168 15632 20220 15638
rect 20168 15574 20220 15580
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20180 13530 20208 15574
rect 20272 14550 20300 16934
rect 20364 16250 20392 17070
rect 20442 17031 20498 17040
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20364 15162 20392 15846
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20260 14544 20312 14550
rect 20260 14486 20312 14492
rect 20352 14272 20404 14278
rect 20456 14249 20484 15302
rect 20352 14214 20404 14220
rect 20442 14240 20498 14249
rect 20364 14006 20392 14214
rect 20442 14175 20498 14184
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20352 14000 20404 14006
rect 20352 13942 20404 13948
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 20456 12782 20484 14010
rect 20548 13841 20576 15302
rect 20640 14657 20668 15846
rect 20626 14648 20682 14657
rect 20626 14583 20682 14592
rect 20732 14482 20760 16594
rect 21008 16153 21036 18022
rect 21100 17202 21128 18702
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 20994 16144 21050 16153
rect 20994 16079 21050 16088
rect 21100 15201 21128 16730
rect 21192 16561 21220 18566
rect 21178 16552 21234 16561
rect 21178 16487 21234 16496
rect 21086 15192 21142 15201
rect 21086 15127 21142 15136
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21192 14618 21220 14758
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20534 13832 20590 13841
rect 20534 13767 20590 13776
rect 20640 13297 20668 14214
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20626 13288 20682 13297
rect 20626 13223 20682 13232
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 20180 11898 20208 12242
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20456 10441 20484 12718
rect 20536 12708 20588 12714
rect 20536 12650 20588 12656
rect 20548 11898 20576 12650
rect 20640 12442 20668 12786
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20640 11082 20668 11562
rect 20732 11354 20760 12582
rect 20824 11694 20852 13806
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20916 12306 20944 13670
rect 21192 13462 21220 14418
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21284 12442 21312 19751
rect 21548 19508 21600 19514
rect 21548 19450 21600 19456
rect 21456 19168 21508 19174
rect 21456 19110 21508 19116
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21376 17338 21404 18770
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21468 16998 21496 19110
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21560 13938 21588 19450
rect 22112 18154 22140 22200
rect 22664 19242 22692 22200
rect 22652 19236 22704 19242
rect 22652 19178 22704 19184
rect 22100 18148 22152 18154
rect 22100 18090 22152 18096
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20442 10432 20498 10441
rect 20442 10367 20498 10376
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 20166 9208 20222 9217
rect 20166 9143 20222 9152
rect 20180 8838 20208 9143
rect 20272 9110 20300 10134
rect 20456 9722 20484 10367
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20260 9104 20312 9110
rect 20260 9046 20312 9052
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20088 6934 20116 7346
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 20088 6118 20116 6870
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 20088 5710 20116 6054
rect 20180 5846 20208 7142
rect 20272 6769 20300 9046
rect 20364 8362 20392 9318
rect 20456 8974 20484 9522
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20456 8430 20484 8910
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20352 8356 20404 8362
rect 20352 8298 20404 8304
rect 20456 8090 20484 8366
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 20548 7002 20576 7890
rect 20640 7274 20668 11018
rect 20732 10810 20760 11086
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20732 9178 20760 9318
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20824 7478 20852 11494
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 21376 10130 21404 10406
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21376 10033 21404 10066
rect 21362 10024 21418 10033
rect 21362 9959 21364 9968
rect 21416 9959 21418 9968
rect 21364 9930 21416 9936
rect 20996 9920 21048 9926
rect 20996 9862 21048 9868
rect 21008 9489 21036 9862
rect 21376 9518 21404 9930
rect 21364 9512 21416 9518
rect 20994 9480 21050 9489
rect 21364 9454 21416 9460
rect 20994 9415 21050 9424
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20258 6760 20314 6769
rect 20258 6695 20314 6704
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20272 5914 20300 6054
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20168 5840 20220 5846
rect 20168 5782 20220 5788
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 19708 4004 19760 4010
rect 19708 3946 19760 3952
rect 19720 3738 19748 3946
rect 19708 3732 19760 3738
rect 19708 3674 19760 3680
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19536 2836 19564 3470
rect 19720 3058 19748 3674
rect 19996 3602 20024 4422
rect 20088 4214 20116 5034
rect 20548 4622 20576 6938
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20076 4208 20128 4214
rect 20076 4150 20128 4156
rect 20534 4176 20590 4185
rect 20534 4111 20590 4120
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 20444 3596 20496 3602
rect 20444 3538 20496 3544
rect 20456 3058 20484 3538
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 19444 2808 19564 2836
rect 19892 2848 19944 2854
rect 19444 2514 19472 2808
rect 19892 2790 19944 2796
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19248 2440 19300 2446
rect 19154 2408 19210 2417
rect 19248 2382 19300 2388
rect 19154 2343 19210 2352
rect 19260 2106 19288 2382
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 19248 2100 19300 2106
rect 19248 2042 19300 2048
rect 18878 1048 18934 1057
rect 18878 983 18934 992
rect 19352 800 19380 2314
rect 19904 800 19932 2790
rect 20548 2514 20576 4111
rect 20640 3913 20668 7210
rect 20824 7206 20852 7414
rect 20916 7342 20944 7822
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 20812 7200 20864 7206
rect 20810 7168 20812 7177
rect 20864 7168 20866 7177
rect 20810 7103 20866 7112
rect 21100 6322 21128 7346
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21272 4072 21324 4078
rect 20718 4040 20774 4049
rect 21272 4014 21324 4020
rect 20718 3975 20774 3984
rect 20732 3942 20760 3975
rect 20720 3936 20772 3942
rect 20626 3904 20682 3913
rect 20720 3878 20772 3884
rect 20626 3839 20682 3848
rect 20732 2961 20760 3878
rect 20996 3392 21048 3398
rect 20996 3334 21048 3340
rect 20902 3088 20958 3097
rect 20902 3023 20958 3032
rect 20916 2990 20944 3023
rect 20904 2984 20956 2990
rect 20718 2952 20774 2961
rect 20904 2926 20956 2932
rect 20718 2887 20774 2896
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 20456 800 20484 2246
rect 21008 800 21036 3334
rect 21284 2650 21312 4014
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 21560 800 21588 4422
rect 22112 800 22140 5510
rect 22652 5160 22704 5166
rect 22652 5102 22704 5108
rect 22664 800 22692 5102
rect 17774 232 17830 241
rect 17774 167 17830 176
rect 18234 0 18290 800
rect 18786 0 18842 800
rect 19338 0 19394 800
rect 19890 0 19946 800
rect 20442 0 20498 800
rect 20994 0 21050 800
rect 21546 0 21602 800
rect 22098 0 22154 800
rect 22650 0 22706 800
<< via2 >>
rect 19062 22616 19118 22672
rect 18878 22208 18934 22264
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 3422 17176 3478 17232
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4066 5772 4122 5808
rect 4066 5752 4068 5772
rect 4068 5752 4120 5772
rect 4120 5752 4122 5772
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 846 3440 902 3496
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 8390 15680 8446 15736
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 8942 15156 8998 15192
rect 8942 15136 8944 15156
rect 8944 15136 8996 15156
rect 8996 15136 8998 15156
rect 8666 12144 8722 12200
rect 8850 12416 8906 12472
rect 8666 6740 8668 6760
rect 8668 6740 8720 6760
rect 8720 6740 8722 6760
rect 8666 6704 8722 6740
rect 9862 17584 9918 17640
rect 8850 3984 8906 4040
rect 9586 13504 9642 13560
rect 9770 13252 9826 13288
rect 9770 13232 9772 13252
rect 9772 13232 9824 13252
rect 9824 13232 9826 13252
rect 10138 19236 10194 19272
rect 10138 19216 10140 19236
rect 10140 19216 10192 19236
rect 10192 19216 10194 19236
rect 9954 15136 10010 15192
rect 9954 12688 10010 12744
rect 9310 6740 9312 6760
rect 9312 6740 9364 6760
rect 9364 6740 9366 6760
rect 9310 6704 9366 6740
rect 9678 6840 9734 6896
rect 9402 3732 9458 3768
rect 9402 3712 9404 3732
rect 9404 3712 9456 3732
rect 9456 3712 9458 3732
rect 10322 16652 10378 16688
rect 10322 16632 10324 16652
rect 10324 16632 10376 16652
rect 10376 16632 10378 16652
rect 10138 14900 10140 14920
rect 10140 14900 10192 14920
rect 10192 14900 10194 14920
rect 10138 14864 10194 14900
rect 10598 15680 10654 15736
rect 10782 20204 10784 20224
rect 10784 20204 10836 20224
rect 10836 20204 10838 20224
rect 10782 20168 10838 20204
rect 10782 13912 10838 13968
rect 10598 12280 10654 12336
rect 10322 10920 10378 10976
rect 10046 8880 10102 8936
rect 10506 9968 10562 10024
rect 10138 7384 10194 7440
rect 10046 6976 10102 7032
rect 10046 4156 10048 4176
rect 10048 4156 10100 4176
rect 10100 4156 10102 4176
rect 10046 4120 10102 4156
rect 10874 12824 10930 12880
rect 10506 3984 10562 4040
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11150 19780 11206 19816
rect 11150 19760 11152 19780
rect 11152 19760 11204 19780
rect 11204 19760 11206 19780
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11886 18808 11942 18864
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11058 16088 11114 16144
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11702 17212 11704 17232
rect 11704 17212 11756 17232
rect 11756 17212 11758 17232
rect 11702 17176 11758 17212
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11518 16124 11520 16144
rect 11520 16124 11572 16144
rect 11572 16124 11574 16144
rect 11518 16088 11574 16124
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 12162 19796 12164 19816
rect 12164 19796 12216 19816
rect 12216 19796 12218 19816
rect 12162 19760 12218 19796
rect 12438 18808 12494 18864
rect 12806 18708 12808 18728
rect 12808 18708 12860 18728
rect 12860 18708 12862 18728
rect 12806 18672 12862 18708
rect 14462 20168 14518 20224
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 13542 19896 13598 19952
rect 11886 14456 11942 14512
rect 11794 12688 11850 12744
rect 12438 15680 12494 15736
rect 12162 13368 12218 13424
rect 12070 12844 12126 12880
rect 12070 12824 12072 12844
rect 12072 12824 12124 12844
rect 12124 12824 12126 12844
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11242 10532 11298 10568
rect 11242 10512 11244 10532
rect 11244 10512 11296 10532
rect 11296 10512 11298 10532
rect 11610 10104 11666 10160
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11610 9424 11666 9480
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 10874 6180 10930 6216
rect 10874 6160 10876 6180
rect 10876 6160 10928 6180
rect 10928 6160 10930 6180
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 10966 5072 11022 5128
rect 9862 2896 9918 2952
rect 10138 2388 10140 2408
rect 10140 2388 10192 2408
rect 10192 2388 10194 2408
rect 10138 2352 10194 2388
rect 10506 3032 10562 3088
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 10966 2896 11022 2952
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12438 14864 12494 14920
rect 12622 14492 12624 14512
rect 12624 14492 12676 14512
rect 12676 14492 12678 14512
rect 12622 14456 12678 14492
rect 12346 12824 12402 12880
rect 12254 12416 12310 12472
rect 11886 5772 11942 5808
rect 11886 5752 11888 5772
rect 11888 5752 11940 5772
rect 11940 5752 11942 5772
rect 11978 3612 11980 3632
rect 11980 3612 12032 3632
rect 12032 3612 12034 3632
rect 11978 3576 12034 3612
rect 12530 10140 12532 10160
rect 12532 10140 12584 10160
rect 12584 10140 12586 10160
rect 12530 10104 12586 10140
rect 12346 8200 12402 8256
rect 12898 13912 12954 13968
rect 12806 12824 12862 12880
rect 13174 13912 13230 13968
rect 12898 9968 12954 10024
rect 13174 10104 13230 10160
rect 13634 17584 13690 17640
rect 13450 15000 13506 15056
rect 14186 19216 14242 19272
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14830 17720 14886 17776
rect 16394 20440 16450 20496
rect 16302 18672 16358 18728
rect 15750 17856 15806 17912
rect 15750 17584 15806 17640
rect 14370 15020 14426 15056
rect 14370 15000 14372 15020
rect 14372 15000 14424 15020
rect 14424 15000 14426 15020
rect 14186 11736 14242 11792
rect 12346 5636 12402 5672
rect 12346 5616 12348 5636
rect 12348 5616 12400 5636
rect 12400 5616 12402 5636
rect 12346 5092 12402 5128
rect 12346 5072 12348 5092
rect 12348 5072 12400 5092
rect 12400 5072 12402 5092
rect 12438 3984 12494 4040
rect 13266 8880 13322 8936
rect 14094 9832 14150 9888
rect 13910 5636 13966 5672
rect 13910 5616 13912 5636
rect 13912 5616 13964 5636
rect 13964 5616 13966 5636
rect 13726 3576 13782 3632
rect 13910 3440 13966 3496
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 16026 15408 16082 15464
rect 15474 14864 15530 14920
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 15198 13812 15200 13832
rect 15200 13812 15252 13832
rect 15252 13812 15254 13832
rect 15198 13776 15254 13812
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14646 12416 14702 12472
rect 14554 9832 14610 9888
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14738 10104 14794 10160
rect 14830 9696 14886 9752
rect 14830 9560 14886 9616
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 15474 13232 15530 13288
rect 15750 12980 15806 13016
rect 15750 12960 15752 12980
rect 15752 12960 15804 12980
rect 15804 12960 15806 12980
rect 16118 13776 16174 13832
rect 16670 14456 16726 14512
rect 15290 9560 15346 9616
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14830 5788 14832 5808
rect 14832 5788 14884 5808
rect 14884 5788 14886 5808
rect 14830 5752 14886 5788
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14554 3032 14610 3088
rect 14646 2760 14702 2816
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 14186 1536 14242 1592
rect 15658 7792 15714 7848
rect 15658 6160 15714 6216
rect 15474 4120 15530 4176
rect 16762 12960 16818 13016
rect 16578 10512 16634 10568
rect 16486 8880 16542 8936
rect 17130 16632 17186 16688
rect 16118 5244 16120 5264
rect 16120 5244 16172 5264
rect 16172 5244 16174 5264
rect 16118 5208 16174 5244
rect 16210 1964 16266 2000
rect 16210 1944 16212 1964
rect 16212 1944 16264 1964
rect 16264 1944 16266 1964
rect 18694 20712 18750 20768
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18602 20440 18658 20496
rect 17590 17856 17646 17912
rect 17866 17856 17922 17912
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18050 19252 18052 19272
rect 18052 19252 18104 19272
rect 18104 19252 18106 19272
rect 18050 19216 18106 19252
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18142 17992 18198 18048
rect 18234 17584 18290 17640
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 17590 13776 17646 13832
rect 17498 11600 17554 11656
rect 17498 11192 17554 11248
rect 17038 3984 17094 4040
rect 17682 12824 17738 12880
rect 17866 12280 17922 12336
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18326 15544 18382 15600
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18970 20304 19026 20360
rect 18970 19896 19026 19952
rect 19338 21664 19394 21720
rect 18694 18400 18750 18456
rect 18694 17720 18750 17776
rect 18694 17176 18750 17232
rect 18602 14884 18658 14920
rect 18602 14864 18604 14884
rect 18604 14864 18656 14884
rect 18656 14864 18658 14884
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18418 13776 18474 13832
rect 18326 13232 18382 13288
rect 18510 13268 18512 13288
rect 18512 13268 18564 13288
rect 18564 13268 18566 13288
rect 18510 13232 18566 13268
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18510 12688 18566 12744
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18326 11756 18382 11792
rect 18326 11736 18328 11756
rect 18328 11736 18380 11756
rect 18380 11736 18382 11756
rect 17958 11328 18014 11384
rect 18418 11192 18474 11248
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 17866 10648 17922 10704
rect 18510 9968 18566 10024
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18326 9424 18382 9480
rect 18234 8880 18290 8936
rect 18602 9016 18658 9072
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 17958 8064 18014 8120
rect 17590 1944 17646 2000
rect 15290 584 15346 640
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18142 5752 18198 5808
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 17958 4800 18014 4856
rect 18694 6160 18750 6216
rect 17958 4528 18014 4584
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 17958 4276 18014 4312
rect 17958 4256 17960 4276
rect 17960 4256 18012 4276
rect 18012 4256 18014 4276
rect 18050 3576 18106 3632
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 19890 21256 19946 21312
rect 19890 19352 19946 19408
rect 19246 17448 19302 17504
rect 18970 10920 19026 10976
rect 18878 10784 18934 10840
rect 18970 9152 19026 9208
rect 18418 2932 18420 2952
rect 18420 2932 18472 2952
rect 18472 2932 18474 2952
rect 18418 2896 18474 2932
rect 18142 2488 18198 2544
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 19154 9424 19210 9480
rect 19062 3440 19118 3496
rect 20626 18808 20682 18864
rect 21270 19760 21326 19816
rect 20442 17040 20498 17096
rect 20442 14184 20498 14240
rect 20626 14592 20682 14648
rect 20994 16088 21050 16144
rect 21178 16496 21234 16552
rect 21086 15136 21142 15192
rect 20534 13776 20590 13832
rect 20626 13232 20682 13288
rect 20442 10376 20498 10432
rect 20166 9152 20222 9208
rect 21362 9988 21418 10024
rect 21362 9968 21364 9988
rect 21364 9968 21416 9988
rect 21416 9968 21418 9988
rect 20994 9424 21050 9480
rect 20258 6704 20314 6760
rect 20534 4120 20590 4176
rect 19154 2352 19210 2408
rect 18878 992 18934 1048
rect 20810 7148 20812 7168
rect 20812 7148 20864 7168
rect 20864 7148 20866 7168
rect 20810 7112 20866 7148
rect 20718 3984 20774 4040
rect 20626 3848 20682 3904
rect 20902 3032 20958 3088
rect 20718 2896 20774 2952
rect 17774 176 17830 232
<< metal3 >>
rect 19057 22674 19123 22677
rect 22200 22674 23000 22704
rect 19057 22672 23000 22674
rect 19057 22616 19062 22672
rect 19118 22616 23000 22672
rect 19057 22614 23000 22616
rect 19057 22611 19123 22614
rect 22200 22584 23000 22614
rect 18873 22266 18939 22269
rect 22200 22266 23000 22296
rect 18873 22264 23000 22266
rect 18873 22208 18878 22264
rect 18934 22208 23000 22264
rect 18873 22206 23000 22208
rect 18873 22203 18939 22206
rect 22200 22176 23000 22206
rect 19333 21722 19399 21725
rect 22200 21722 23000 21752
rect 19333 21720 23000 21722
rect 19333 21664 19338 21720
rect 19394 21664 23000 21720
rect 19333 21662 23000 21664
rect 19333 21659 19399 21662
rect 22200 21632 23000 21662
rect 19885 21314 19951 21317
rect 22200 21314 23000 21344
rect 19885 21312 23000 21314
rect 19885 21256 19890 21312
rect 19946 21256 23000 21312
rect 19885 21254 23000 21256
rect 19885 21251 19951 21254
rect 22200 21224 23000 21254
rect 18689 20770 18755 20773
rect 22200 20770 23000 20800
rect 18689 20768 23000 20770
rect 18689 20712 18694 20768
rect 18750 20712 23000 20768
rect 18689 20710 23000 20712
rect 18689 20707 18755 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 22200 20680 23000 20710
rect 18270 20639 18590 20640
rect 16389 20498 16455 20501
rect 18597 20498 18663 20501
rect 16389 20496 18663 20498
rect 16389 20440 16394 20496
rect 16450 20440 18602 20496
rect 18658 20440 18663 20496
rect 16389 20438 18663 20440
rect 16389 20435 16455 20438
rect 18597 20435 18663 20438
rect 18965 20362 19031 20365
rect 22200 20362 23000 20392
rect 18965 20360 23000 20362
rect 18965 20304 18970 20360
rect 19026 20304 23000 20360
rect 18965 20302 23000 20304
rect 18965 20299 19031 20302
rect 22200 20272 23000 20302
rect 10777 20226 10843 20229
rect 14457 20226 14523 20229
rect 10777 20224 14523 20226
rect 10777 20168 10782 20224
rect 10838 20168 14462 20224
rect 14518 20168 14523 20224
rect 10777 20166 14523 20168
rect 10777 20163 10843 20166
rect 14457 20163 14523 20166
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 13537 19954 13603 19957
rect 18965 19954 19031 19957
rect 13537 19952 19031 19954
rect 13537 19896 13542 19952
rect 13598 19896 18970 19952
rect 19026 19896 19031 19952
rect 13537 19894 19031 19896
rect 13537 19891 13603 19894
rect 18965 19891 19031 19894
rect 11145 19818 11211 19821
rect 12157 19818 12223 19821
rect 11145 19816 12223 19818
rect 11145 19760 11150 19816
rect 11206 19760 12162 19816
rect 12218 19760 12223 19816
rect 11145 19758 12223 19760
rect 11145 19755 11211 19758
rect 12157 19755 12223 19758
rect 21265 19818 21331 19821
rect 22200 19818 23000 19848
rect 21265 19816 23000 19818
rect 21265 19760 21270 19816
rect 21326 19760 23000 19816
rect 21265 19758 23000 19760
rect 21265 19755 21331 19758
rect 22200 19728 23000 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 19885 19410 19951 19413
rect 22200 19410 23000 19440
rect 19885 19408 23000 19410
rect 19885 19352 19890 19408
rect 19946 19352 23000 19408
rect 19885 19350 23000 19352
rect 19885 19347 19951 19350
rect 22200 19320 23000 19350
rect 10133 19274 10199 19277
rect 14181 19274 14247 19277
rect 18045 19274 18111 19277
rect 10133 19272 18111 19274
rect 10133 19216 10138 19272
rect 10194 19216 14186 19272
rect 14242 19216 18050 19272
rect 18106 19216 18111 19272
rect 10133 19214 18111 19216
rect 10133 19211 10199 19214
rect 14181 19211 14247 19214
rect 18045 19211 18111 19214
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 11881 18866 11947 18869
rect 12433 18866 12499 18869
rect 20621 18866 20687 18869
rect 22200 18866 23000 18896
rect 11881 18864 12534 18866
rect 11881 18808 11886 18864
rect 11942 18808 12438 18864
rect 12494 18808 12534 18864
rect 11881 18806 12534 18808
rect 20621 18864 23000 18866
rect 20621 18808 20626 18864
rect 20682 18808 23000 18864
rect 20621 18806 23000 18808
rect 11881 18803 11947 18806
rect 12433 18803 12499 18806
rect 20621 18803 20687 18806
rect 22200 18776 23000 18806
rect 12801 18730 12867 18733
rect 16297 18730 16363 18733
rect 12801 18728 16363 18730
rect 12801 18672 12806 18728
rect 12862 18672 16302 18728
rect 16358 18672 16363 18728
rect 12801 18670 16363 18672
rect 12801 18667 12867 18670
rect 16297 18667 16363 18670
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 18689 18458 18755 18461
rect 22200 18458 23000 18488
rect 18689 18456 23000 18458
rect 18689 18400 18694 18456
rect 18750 18400 23000 18456
rect 18689 18398 23000 18400
rect 18689 18395 18755 18398
rect 22200 18368 23000 18398
rect 18137 18050 18203 18053
rect 22200 18050 23000 18080
rect 18137 18048 23000 18050
rect 18137 17992 18142 18048
rect 18198 17992 23000 18048
rect 18137 17990 23000 17992
rect 18137 17987 18203 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22200 17960 23000 17990
rect 14805 17919 15125 17920
rect 15745 17914 15811 17917
rect 17585 17914 17651 17917
rect 17861 17914 17927 17917
rect 15745 17912 17927 17914
rect 15745 17856 15750 17912
rect 15806 17856 17590 17912
rect 17646 17856 17866 17912
rect 17922 17856 17927 17912
rect 15745 17854 17927 17856
rect 15745 17851 15811 17854
rect 17585 17851 17651 17854
rect 17861 17851 17927 17854
rect 14825 17778 14891 17781
rect 18689 17778 18755 17781
rect 14825 17776 18755 17778
rect 14825 17720 14830 17776
rect 14886 17720 18694 17776
rect 18750 17720 18755 17776
rect 14825 17718 18755 17720
rect 14825 17715 14891 17718
rect 18689 17715 18755 17718
rect 9857 17642 9923 17645
rect 13486 17642 13492 17644
rect 9857 17640 13492 17642
rect 9857 17584 9862 17640
rect 9918 17584 13492 17640
rect 9857 17582 13492 17584
rect 9857 17579 9923 17582
rect 13486 17580 13492 17582
rect 13556 17642 13562 17644
rect 13629 17642 13695 17645
rect 13556 17640 13695 17642
rect 13556 17584 13634 17640
rect 13690 17584 13695 17640
rect 13556 17582 13695 17584
rect 13556 17580 13562 17582
rect 13629 17579 13695 17582
rect 15745 17642 15811 17645
rect 18229 17642 18295 17645
rect 15745 17640 18295 17642
rect 15745 17584 15750 17640
rect 15806 17584 18234 17640
rect 18290 17584 18295 17640
rect 15745 17582 18295 17584
rect 15745 17579 15811 17582
rect 18229 17579 18295 17582
rect 19241 17506 19307 17509
rect 22200 17506 23000 17536
rect 19241 17504 23000 17506
rect 19241 17448 19246 17504
rect 19302 17448 23000 17504
rect 19241 17446 23000 17448
rect 19241 17443 19307 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 22200 17416 23000 17446
rect 18270 17375 18590 17376
rect 0 17234 800 17264
rect 3417 17234 3483 17237
rect 0 17232 3483 17234
rect 0 17176 3422 17232
rect 3478 17176 3483 17232
rect 0 17174 3483 17176
rect 0 17144 800 17174
rect 3417 17171 3483 17174
rect 11697 17234 11763 17237
rect 18689 17234 18755 17237
rect 11697 17232 18755 17234
rect 11697 17176 11702 17232
rect 11758 17176 18694 17232
rect 18750 17176 18755 17232
rect 11697 17174 18755 17176
rect 11697 17171 11763 17174
rect 18689 17171 18755 17174
rect 20437 17098 20503 17101
rect 22200 17098 23000 17128
rect 20437 17096 23000 17098
rect 20437 17040 20442 17096
rect 20498 17040 23000 17096
rect 20437 17038 23000 17040
rect 20437 17035 20503 17038
rect 22200 17008 23000 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 10317 16690 10383 16693
rect 17125 16690 17191 16693
rect 10317 16688 17191 16690
rect 10317 16632 10322 16688
rect 10378 16632 17130 16688
rect 17186 16632 17191 16688
rect 10317 16630 17191 16632
rect 10317 16627 10383 16630
rect 17125 16627 17191 16630
rect 21173 16554 21239 16557
rect 22200 16554 23000 16584
rect 21173 16552 23000 16554
rect 21173 16496 21178 16552
rect 21234 16496 23000 16552
rect 21173 16494 23000 16496
rect 21173 16491 21239 16494
rect 22200 16464 23000 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 11053 16146 11119 16149
rect 11513 16146 11579 16149
rect 11053 16144 11579 16146
rect 11053 16088 11058 16144
rect 11114 16088 11518 16144
rect 11574 16088 11579 16144
rect 11053 16086 11579 16088
rect 11053 16083 11119 16086
rect 11513 16083 11579 16086
rect 20989 16146 21055 16149
rect 22200 16146 23000 16176
rect 20989 16144 23000 16146
rect 20989 16088 20994 16144
rect 21050 16088 23000 16144
rect 20989 16086 23000 16088
rect 20989 16083 21055 16086
rect 22200 16056 23000 16086
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 8385 15738 8451 15741
rect 10593 15740 10659 15741
rect 10542 15738 10548 15740
rect 8385 15736 10548 15738
rect 10612 15738 10659 15740
rect 12433 15738 12499 15741
rect 10612 15736 12499 15738
rect 8385 15680 8390 15736
rect 8446 15680 10548 15736
rect 10654 15680 12438 15736
rect 12494 15680 12499 15736
rect 8385 15678 10548 15680
rect 8385 15675 8451 15678
rect 10542 15676 10548 15678
rect 10612 15678 12499 15680
rect 10612 15676 10659 15678
rect 10593 15675 10659 15676
rect 12433 15675 12499 15678
rect 18321 15602 18387 15605
rect 22200 15602 23000 15632
rect 18321 15600 23000 15602
rect 18321 15544 18326 15600
rect 18382 15544 23000 15600
rect 18321 15542 23000 15544
rect 18321 15539 18387 15542
rect 22200 15512 23000 15542
rect 16021 15466 16087 15469
rect 11102 15464 16087 15466
rect 11102 15408 16026 15464
rect 16082 15408 16087 15464
rect 11102 15406 16087 15408
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 8937 15194 9003 15197
rect 9949 15194 10015 15197
rect 10358 15194 10364 15196
rect 8937 15192 10364 15194
rect 8937 15136 8942 15192
rect 8998 15136 9954 15192
rect 10010 15136 10364 15192
rect 8937 15134 10364 15136
rect 8937 15131 9003 15134
rect 9949 15131 10015 15134
rect 10358 15132 10364 15134
rect 10428 15194 10434 15196
rect 11102 15194 11162 15406
rect 16021 15403 16087 15406
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 10428 15134 11162 15194
rect 21081 15194 21147 15197
rect 22200 15194 23000 15224
rect 21081 15192 23000 15194
rect 21081 15136 21086 15192
rect 21142 15136 23000 15192
rect 21081 15134 23000 15136
rect 10428 15132 10434 15134
rect 21081 15131 21147 15134
rect 22200 15104 23000 15134
rect 13445 15058 13511 15061
rect 14365 15058 14431 15061
rect 13445 15056 14431 15058
rect 13445 15000 13450 15056
rect 13506 15000 14370 15056
rect 14426 15000 14431 15056
rect 13445 14998 14431 15000
rect 13445 14995 13511 14998
rect 14365 14995 14431 14998
rect 10133 14922 10199 14925
rect 12433 14922 12499 14925
rect 10133 14920 12499 14922
rect 10133 14864 10138 14920
rect 10194 14864 12438 14920
rect 12494 14864 12499 14920
rect 10133 14862 12499 14864
rect 10133 14859 10199 14862
rect 12433 14859 12499 14862
rect 15469 14922 15535 14925
rect 18597 14922 18663 14925
rect 15469 14920 18663 14922
rect 15469 14864 15474 14920
rect 15530 14864 18602 14920
rect 18658 14864 18663 14920
rect 15469 14862 18663 14864
rect 15469 14859 15535 14862
rect 18597 14859 18663 14862
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 20621 14650 20687 14653
rect 22200 14650 23000 14680
rect 20621 14648 23000 14650
rect 20621 14592 20626 14648
rect 20682 14592 23000 14648
rect 20621 14590 23000 14592
rect 20621 14587 20687 14590
rect 22200 14560 23000 14590
rect 11881 14514 11947 14517
rect 12198 14514 12204 14516
rect 11881 14512 12204 14514
rect 11881 14456 11886 14512
rect 11942 14456 12204 14512
rect 11881 14454 12204 14456
rect 11881 14451 11947 14454
rect 12198 14452 12204 14454
rect 12268 14452 12274 14516
rect 12617 14514 12683 14517
rect 16665 14514 16731 14517
rect 12617 14512 16731 14514
rect 12617 14456 12622 14512
rect 12678 14456 16670 14512
rect 16726 14456 16731 14512
rect 12617 14454 16731 14456
rect 12617 14451 12683 14454
rect 16665 14451 16731 14454
rect 20437 14242 20503 14245
rect 22200 14242 23000 14272
rect 20437 14240 23000 14242
rect 20437 14184 20442 14240
rect 20498 14184 23000 14240
rect 20437 14182 23000 14184
rect 20437 14179 20503 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 22200 14152 23000 14182
rect 18270 14111 18590 14112
rect 10777 13970 10843 13973
rect 12893 13970 12959 13973
rect 13169 13970 13235 13973
rect 10777 13968 13235 13970
rect 10777 13912 10782 13968
rect 10838 13912 12898 13968
rect 12954 13912 13174 13968
rect 13230 13912 13235 13968
rect 10777 13910 13235 13912
rect 10777 13907 10843 13910
rect 12893 13907 12959 13910
rect 13169 13907 13235 13910
rect 15193 13834 15259 13837
rect 14598 13832 15259 13834
rect 14598 13776 15198 13832
rect 15254 13776 15259 13832
rect 14598 13774 15259 13776
rect 14598 13698 14658 13774
rect 15193 13771 15259 13774
rect 16113 13834 16179 13837
rect 17585 13834 17651 13837
rect 18413 13834 18479 13837
rect 16113 13832 18479 13834
rect 16113 13776 16118 13832
rect 16174 13776 17590 13832
rect 17646 13776 18418 13832
rect 18474 13776 18479 13832
rect 16113 13774 18479 13776
rect 16113 13771 16179 13774
rect 17585 13771 17651 13774
rect 18413 13771 18479 13774
rect 20529 13834 20595 13837
rect 22200 13834 23000 13864
rect 20529 13832 23000 13834
rect 20529 13776 20534 13832
rect 20590 13776 23000 13832
rect 20529 13774 23000 13776
rect 20529 13771 20595 13774
rect 22200 13744 23000 13774
rect 9584 13638 14658 13698
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 9584 13565 9644 13638
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 9581 13560 9647 13565
rect 9581 13504 9586 13560
rect 9642 13504 9647 13560
rect 9581 13499 9647 13504
rect 12157 13426 12223 13429
rect 12157 13424 18154 13426
rect 12157 13368 12162 13424
rect 12218 13368 18154 13424
rect 12157 13366 18154 13368
rect 12157 13363 12223 13366
rect 9765 13290 9831 13293
rect 15469 13290 15535 13293
rect 18094 13292 18154 13366
rect 9765 13288 15535 13290
rect 9765 13232 9770 13288
rect 9826 13232 15474 13288
rect 15530 13232 15535 13288
rect 9765 13230 15535 13232
rect 9765 13227 9831 13230
rect 15469 13227 15535 13230
rect 18086 13228 18092 13292
rect 18156 13290 18162 13292
rect 18321 13290 18387 13293
rect 18156 13288 18387 13290
rect 18156 13232 18326 13288
rect 18382 13232 18387 13288
rect 18156 13230 18387 13232
rect 18156 13228 18162 13230
rect 18321 13227 18387 13230
rect 18505 13290 18571 13293
rect 18822 13290 18828 13292
rect 18505 13288 18828 13290
rect 18505 13232 18510 13288
rect 18566 13232 18828 13288
rect 18505 13230 18828 13232
rect 18505 13227 18571 13230
rect 18822 13228 18828 13230
rect 18892 13228 18898 13292
rect 20621 13290 20687 13293
rect 22200 13290 23000 13320
rect 20621 13288 23000 13290
rect 20621 13232 20626 13288
rect 20682 13232 23000 13288
rect 20621 13230 23000 13232
rect 20621 13227 20687 13230
rect 22200 13200 23000 13230
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 15745 13018 15811 13021
rect 16757 13018 16823 13021
rect 15745 13016 16823 13018
rect 15745 12960 15750 13016
rect 15806 12960 16762 13016
rect 16818 12960 16823 13016
rect 15745 12958 16823 12960
rect 15745 12955 15811 12958
rect 16757 12955 16823 12958
rect 10869 12882 10935 12885
rect 12065 12882 12131 12885
rect 10869 12880 12131 12882
rect 10869 12824 10874 12880
rect 10930 12824 12070 12880
rect 12126 12824 12131 12880
rect 10869 12822 12131 12824
rect 10869 12819 10935 12822
rect 12065 12819 12131 12822
rect 12341 12882 12407 12885
rect 12801 12882 12867 12885
rect 12341 12880 12867 12882
rect 12341 12824 12346 12880
rect 12402 12824 12806 12880
rect 12862 12824 12867 12880
rect 12341 12822 12867 12824
rect 12341 12819 12407 12822
rect 12801 12819 12867 12822
rect 17677 12882 17743 12885
rect 22200 12882 23000 12912
rect 17677 12880 23000 12882
rect 17677 12824 17682 12880
rect 17738 12824 23000 12880
rect 17677 12822 23000 12824
rect 17677 12819 17743 12822
rect 22200 12792 23000 12822
rect 9949 12746 10015 12749
rect 11789 12746 11855 12749
rect 18505 12746 18571 12749
rect 9949 12744 18571 12746
rect 9949 12688 9954 12744
rect 10010 12688 11794 12744
rect 11850 12688 18510 12744
rect 18566 12688 18571 12744
rect 9949 12686 18571 12688
rect 9949 12683 10015 12686
rect 11789 12683 11855 12686
rect 18505 12683 18571 12686
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 8845 12474 8911 12477
rect 8664 12472 8911 12474
rect 8664 12416 8850 12472
rect 8906 12416 8911 12472
rect 8664 12414 8911 12416
rect 8664 12205 8724 12414
rect 8845 12411 8911 12414
rect 12249 12474 12315 12477
rect 14641 12476 14707 12477
rect 13486 12474 13492 12476
rect 12249 12472 13492 12474
rect 12249 12416 12254 12472
rect 12310 12416 13492 12472
rect 12249 12414 13492 12416
rect 12249 12411 12315 12414
rect 13486 12412 13492 12414
rect 13556 12412 13562 12476
rect 14590 12474 14596 12476
rect 14550 12414 14596 12474
rect 14660 12472 14707 12476
rect 14702 12416 14707 12472
rect 14590 12412 14596 12414
rect 14660 12412 14707 12416
rect 14641 12411 14707 12412
rect 10593 12340 10659 12341
rect 10542 12276 10548 12340
rect 10612 12338 10659 12340
rect 17861 12338 17927 12341
rect 22200 12338 23000 12368
rect 10612 12336 10704 12338
rect 10654 12280 10704 12336
rect 10612 12278 10704 12280
rect 17861 12336 23000 12338
rect 17861 12280 17866 12336
rect 17922 12280 23000 12336
rect 17861 12278 23000 12280
rect 10612 12276 10659 12278
rect 10593 12275 10659 12276
rect 17861 12275 17927 12278
rect 22200 12248 23000 12278
rect 8661 12200 8727 12205
rect 8661 12144 8666 12200
rect 8722 12144 8727 12200
rect 8661 12139 8727 12144
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 22200 11930 23000 11960
rect 18830 11870 23000 11930
rect 14181 11794 14247 11797
rect 18321 11794 18387 11797
rect 14181 11792 18387 11794
rect 14181 11736 14186 11792
rect 14242 11736 18326 11792
rect 18382 11736 18387 11792
rect 14181 11734 18387 11736
rect 14181 11731 14247 11734
rect 18321 11731 18387 11734
rect 17493 11658 17559 11661
rect 18830 11658 18890 11870
rect 22200 11840 23000 11870
rect 17493 11656 18890 11658
rect 17493 11600 17498 11656
rect 17554 11600 18890 11656
rect 17493 11598 18890 11600
rect 17493 11595 17559 11598
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 17953 11386 18019 11389
rect 22200 11386 23000 11416
rect 17953 11384 23000 11386
rect 17953 11328 17958 11384
rect 18014 11328 23000 11384
rect 17953 11326 23000 11328
rect 17953 11323 18019 11326
rect 22200 11296 23000 11326
rect 17493 11250 17559 11253
rect 18413 11250 18479 11253
rect 17493 11248 18479 11250
rect 17493 11192 17498 11248
rect 17554 11192 18418 11248
rect 18474 11192 18479 11248
rect 17493 11190 18479 11192
rect 17493 11187 17559 11190
rect 18413 11187 18479 11190
rect 10317 10980 10383 10981
rect 10317 10978 10364 10980
rect 10272 10976 10364 10978
rect 10272 10920 10322 10976
rect 10272 10918 10364 10920
rect 10317 10916 10364 10918
rect 10428 10916 10434 10980
rect 18965 10978 19031 10981
rect 22200 10978 23000 11008
rect 18965 10976 23000 10978
rect 18965 10920 18970 10976
rect 19026 10920 23000 10976
rect 18965 10918 23000 10920
rect 10317 10915 10383 10916
rect 18965 10915 19031 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 22200 10888 23000 10918
rect 18270 10847 18590 10848
rect 18873 10844 18939 10845
rect 18822 10780 18828 10844
rect 18892 10842 18939 10844
rect 18892 10840 18984 10842
rect 18934 10784 18984 10840
rect 18892 10782 18984 10784
rect 18892 10780 18939 10782
rect 18873 10779 18939 10780
rect 17861 10706 17927 10709
rect 18086 10706 18092 10708
rect 17861 10704 18092 10706
rect 17861 10648 17866 10704
rect 17922 10648 18092 10704
rect 17861 10646 18092 10648
rect 17861 10643 17927 10646
rect 18086 10644 18092 10646
rect 18156 10644 18162 10708
rect 11237 10570 11303 10573
rect 16573 10570 16639 10573
rect 11237 10568 16639 10570
rect 11237 10512 11242 10568
rect 11298 10512 16578 10568
rect 16634 10512 16639 10568
rect 11237 10510 16639 10512
rect 11237 10507 11303 10510
rect 16573 10507 16639 10510
rect 20437 10434 20503 10437
rect 22200 10434 23000 10464
rect 20437 10432 23000 10434
rect 20437 10376 20442 10432
rect 20498 10376 23000 10432
rect 20437 10374 23000 10376
rect 20437 10371 20503 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 22200 10344 23000 10374
rect 14805 10303 15125 10304
rect 11605 10162 11671 10165
rect 12525 10162 12591 10165
rect 11605 10160 12591 10162
rect 11605 10104 11610 10160
rect 11666 10104 12530 10160
rect 12586 10104 12591 10160
rect 11605 10102 12591 10104
rect 11605 10099 11671 10102
rect 12525 10099 12591 10102
rect 13169 10162 13235 10165
rect 14733 10162 14799 10165
rect 13169 10160 14799 10162
rect 13169 10104 13174 10160
rect 13230 10104 14738 10160
rect 14794 10104 14799 10160
rect 13169 10102 14799 10104
rect 13169 10099 13235 10102
rect 14733 10099 14799 10102
rect 10501 10026 10567 10029
rect 12893 10026 12959 10029
rect 18505 10026 18571 10029
rect 10501 10024 18571 10026
rect 10501 9968 10506 10024
rect 10562 9968 12898 10024
rect 12954 9968 18510 10024
rect 18566 9968 18571 10024
rect 10501 9966 18571 9968
rect 10501 9963 10567 9966
rect 12893 9963 12959 9966
rect 18505 9963 18571 9966
rect 21357 10026 21423 10029
rect 22200 10026 23000 10056
rect 21357 10024 23000 10026
rect 21357 9968 21362 10024
rect 21418 9968 23000 10024
rect 21357 9966 23000 9968
rect 21357 9963 21423 9966
rect 22200 9936 23000 9966
rect 14089 9890 14155 9893
rect 14549 9890 14615 9893
rect 14089 9888 14615 9890
rect 14089 9832 14094 9888
rect 14150 9832 14554 9888
rect 14610 9832 14615 9888
rect 14089 9830 14615 9832
rect 14089 9827 14155 9830
rect 14549 9827 14615 9830
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 14590 9692 14596 9756
rect 14660 9754 14666 9756
rect 14825 9754 14891 9757
rect 14660 9752 14891 9754
rect 14660 9696 14830 9752
rect 14886 9696 14891 9752
rect 14660 9694 14891 9696
rect 14660 9692 14666 9694
rect 14825 9691 14891 9694
rect 14825 9618 14891 9621
rect 15285 9618 15351 9621
rect 14825 9616 15351 9618
rect 14825 9560 14830 9616
rect 14886 9560 15290 9616
rect 15346 9560 15351 9616
rect 14825 9558 15351 9560
rect 14825 9555 14891 9558
rect 15285 9555 15351 9558
rect 11605 9482 11671 9485
rect 18321 9482 18387 9485
rect 11605 9480 18387 9482
rect 11605 9424 11610 9480
rect 11666 9424 18326 9480
rect 18382 9424 18387 9480
rect 11605 9422 18387 9424
rect 11605 9419 11671 9422
rect 18321 9419 18387 9422
rect 19149 9482 19215 9485
rect 20989 9482 21055 9485
rect 22200 9482 23000 9512
rect 19149 9480 23000 9482
rect 19149 9424 19154 9480
rect 19210 9424 20994 9480
rect 21050 9424 23000 9480
rect 19149 9422 23000 9424
rect 19149 9419 19215 9422
rect 20989 9419 21055 9422
rect 22200 9392 23000 9422
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 18965 9210 19031 9213
rect 20161 9210 20227 9213
rect 18965 9208 20227 9210
rect 18965 9152 18970 9208
rect 19026 9152 20166 9208
rect 20222 9152 20227 9208
rect 18965 9150 20227 9152
rect 18965 9147 19031 9150
rect 20161 9147 20227 9150
rect 18597 9074 18663 9077
rect 22200 9074 23000 9104
rect 18597 9072 23000 9074
rect 18597 9016 18602 9072
rect 18658 9016 23000 9072
rect 18597 9014 23000 9016
rect 18597 9011 18663 9014
rect 22200 8984 23000 9014
rect 10041 8938 10107 8941
rect 13261 8938 13327 8941
rect 16481 8938 16547 8941
rect 10041 8936 16547 8938
rect 10041 8880 10046 8936
rect 10102 8880 13266 8936
rect 13322 8880 16486 8936
rect 16542 8880 16547 8936
rect 10041 8878 16547 8880
rect 10041 8875 10107 8878
rect 13261 8875 13327 8878
rect 16481 8875 16547 8878
rect 18229 8938 18295 8941
rect 18229 8936 18890 8938
rect 18229 8880 18234 8936
rect 18290 8880 18890 8936
rect 18229 8878 18890 8880
rect 18229 8875 18295 8878
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 18830 8666 18890 8878
rect 22200 8666 23000 8696
rect 18830 8606 23000 8666
rect 22200 8576 23000 8606
rect 12198 8196 12204 8260
rect 12268 8258 12274 8260
rect 12341 8258 12407 8261
rect 12268 8256 12407 8258
rect 12268 8200 12346 8256
rect 12402 8200 12407 8256
rect 12268 8198 12407 8200
rect 12268 8196 12274 8198
rect 12341 8195 12407 8198
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 17953 8122 18019 8125
rect 22200 8122 23000 8152
rect 17953 8120 23000 8122
rect 17953 8064 17958 8120
rect 18014 8064 23000 8120
rect 17953 8062 23000 8064
rect 17953 8059 18019 8062
rect 22200 8032 23000 8062
rect 15653 7850 15719 7853
rect 15653 7848 18752 7850
rect 15653 7792 15658 7848
rect 15714 7792 18752 7848
rect 15653 7790 18752 7792
rect 15653 7787 15719 7790
rect 18692 7714 18752 7790
rect 22200 7714 23000 7744
rect 18692 7654 23000 7714
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 22200 7624 23000 7654
rect 18270 7583 18590 7584
rect 10133 7444 10199 7445
rect 10133 7442 10180 7444
rect 10088 7440 10180 7442
rect 10088 7384 10138 7440
rect 10088 7382 10180 7384
rect 10133 7380 10180 7382
rect 10244 7380 10250 7444
rect 10133 7379 10199 7380
rect 20805 7170 20871 7173
rect 22200 7170 23000 7200
rect 20805 7168 23000 7170
rect 20805 7112 20810 7168
rect 20866 7112 23000 7168
rect 20805 7110 23000 7112
rect 20805 7107 20871 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 22200 7080 23000 7110
rect 14805 7039 15125 7040
rect 10041 7032 10107 7037
rect 10041 6976 10046 7032
rect 10102 6976 10107 7032
rect 10041 6971 10107 6976
rect 9673 6898 9739 6901
rect 10044 6898 10104 6971
rect 9673 6896 10104 6898
rect 9673 6840 9678 6896
rect 9734 6840 10104 6896
rect 9673 6838 10104 6840
rect 9673 6835 9739 6838
rect 8661 6762 8727 6765
rect 9305 6762 9371 6765
rect 8661 6760 9371 6762
rect 8661 6704 8666 6760
rect 8722 6704 9310 6760
rect 9366 6704 9371 6760
rect 8661 6702 9371 6704
rect 8661 6699 8727 6702
rect 9305 6699 9371 6702
rect 20253 6762 20319 6765
rect 22200 6762 23000 6792
rect 20253 6760 23000 6762
rect 20253 6704 20258 6760
rect 20314 6704 23000 6760
rect 20253 6702 23000 6704
rect 20253 6699 20319 6702
rect 22200 6672 23000 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 10869 6218 10935 6221
rect 15653 6218 15719 6221
rect 10869 6216 15719 6218
rect 10869 6160 10874 6216
rect 10930 6160 15658 6216
rect 15714 6160 15719 6216
rect 10869 6158 15719 6160
rect 10869 6155 10935 6158
rect 15653 6155 15719 6158
rect 18689 6218 18755 6221
rect 22200 6218 23000 6248
rect 18689 6216 23000 6218
rect 18689 6160 18694 6216
rect 18750 6160 23000 6216
rect 18689 6158 23000 6160
rect 18689 6155 18755 6158
rect 22200 6128 23000 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 0 5810 800 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 800 5750
rect 4061 5747 4127 5750
rect 11881 5810 11947 5813
rect 14825 5810 14891 5813
rect 11881 5808 14891 5810
rect 11881 5752 11886 5808
rect 11942 5752 14830 5808
rect 14886 5752 14891 5808
rect 11881 5750 14891 5752
rect 11881 5747 11947 5750
rect 14825 5747 14891 5750
rect 18137 5810 18203 5813
rect 22200 5810 23000 5840
rect 18137 5808 23000 5810
rect 18137 5752 18142 5808
rect 18198 5752 23000 5808
rect 18137 5750 23000 5752
rect 18137 5747 18203 5750
rect 22200 5720 23000 5750
rect 12341 5674 12407 5677
rect 13905 5674 13971 5677
rect 12341 5672 13971 5674
rect 12341 5616 12346 5672
rect 12402 5616 13910 5672
rect 13966 5616 13971 5672
rect 12341 5614 13971 5616
rect 12341 5611 12407 5614
rect 13905 5611 13971 5614
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 16113 5266 16179 5269
rect 22200 5266 23000 5296
rect 16113 5264 23000 5266
rect 16113 5208 16118 5264
rect 16174 5208 23000 5264
rect 16113 5206 23000 5208
rect 16113 5203 16179 5206
rect 22200 5176 23000 5206
rect 10961 5130 11027 5133
rect 12341 5130 12407 5133
rect 10961 5128 12407 5130
rect 10961 5072 10966 5128
rect 11022 5072 12346 5128
rect 12402 5072 12407 5128
rect 10961 5070 12407 5072
rect 10961 5067 11027 5070
rect 12341 5067 12407 5070
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 17953 4858 18019 4861
rect 22200 4858 23000 4888
rect 17953 4856 23000 4858
rect 17953 4800 17958 4856
rect 18014 4800 23000 4856
rect 17953 4798 23000 4800
rect 17953 4795 18019 4798
rect 22200 4768 23000 4798
rect 17953 4586 18019 4589
rect 17953 4584 18890 4586
rect 17953 4528 17958 4584
rect 18014 4528 18890 4584
rect 17953 4526 18890 4528
rect 17953 4523 18019 4526
rect 18830 4450 18890 4526
rect 22200 4450 23000 4480
rect 18830 4390 23000 4450
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 22200 4360 23000 4390
rect 18270 4319 18590 4320
rect 17953 4314 18019 4317
rect 15334 4312 18019 4314
rect 15334 4256 17958 4312
rect 18014 4256 18019 4312
rect 15334 4254 18019 4256
rect 10041 4178 10107 4181
rect 15334 4178 15394 4254
rect 17953 4251 18019 4254
rect 10041 4176 15394 4178
rect 10041 4120 10046 4176
rect 10102 4120 15394 4176
rect 10041 4118 15394 4120
rect 15469 4178 15535 4181
rect 20529 4178 20595 4181
rect 15469 4176 20595 4178
rect 15469 4120 15474 4176
rect 15530 4120 20534 4176
rect 20590 4120 20595 4176
rect 15469 4118 20595 4120
rect 10041 4115 10107 4118
rect 15469 4115 15535 4118
rect 20529 4115 20595 4118
rect 8845 4042 8911 4045
rect 10501 4042 10567 4045
rect 8845 4040 10567 4042
rect 8845 3984 8850 4040
rect 8906 3984 10506 4040
rect 10562 3984 10567 4040
rect 8845 3982 10567 3984
rect 8845 3979 8911 3982
rect 10501 3979 10567 3982
rect 12433 4042 12499 4045
rect 17033 4042 17099 4045
rect 20713 4042 20779 4045
rect 12433 4040 20779 4042
rect 12433 3984 12438 4040
rect 12494 3984 17038 4040
rect 17094 3984 20718 4040
rect 20774 3984 20779 4040
rect 12433 3982 20779 3984
rect 12433 3979 12499 3982
rect 17033 3979 17099 3982
rect 20713 3979 20779 3982
rect 20621 3906 20687 3909
rect 22200 3906 23000 3936
rect 20621 3904 23000 3906
rect 20621 3848 20626 3904
rect 20682 3848 23000 3904
rect 20621 3846 23000 3848
rect 20621 3843 20687 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22200 3816 23000 3846
rect 14805 3775 15125 3776
rect 9397 3770 9463 3773
rect 9397 3768 14658 3770
rect 9397 3712 9402 3768
rect 9458 3712 14658 3768
rect 9397 3710 14658 3712
rect 9397 3707 9463 3710
rect 11973 3634 12039 3637
rect 13721 3634 13787 3637
rect 11973 3632 13787 3634
rect 11973 3576 11978 3632
rect 12034 3576 13726 3632
rect 13782 3576 13787 3632
rect 11973 3574 13787 3576
rect 14598 3634 14658 3710
rect 18045 3634 18111 3637
rect 14598 3632 18111 3634
rect 14598 3576 18050 3632
rect 18106 3576 18111 3632
rect 14598 3574 18111 3576
rect 11973 3571 12039 3574
rect 13721 3571 13787 3574
rect 18045 3571 18111 3574
rect 841 3498 907 3501
rect 13905 3498 13971 3501
rect 841 3496 13971 3498
rect 841 3440 846 3496
rect 902 3440 13910 3496
rect 13966 3440 13971 3496
rect 841 3438 13971 3440
rect 841 3435 907 3438
rect 13905 3435 13971 3438
rect 19057 3498 19123 3501
rect 22200 3498 23000 3528
rect 19057 3496 23000 3498
rect 19057 3440 19062 3496
rect 19118 3440 23000 3496
rect 19057 3438 23000 3440
rect 19057 3435 19123 3438
rect 22200 3408 23000 3438
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 10501 3090 10567 3093
rect 14549 3090 14615 3093
rect 20897 3090 20963 3093
rect 10501 3088 20963 3090
rect 10501 3032 10506 3088
rect 10562 3032 14554 3088
rect 14610 3032 20902 3088
rect 20958 3032 20963 3088
rect 10501 3030 20963 3032
rect 10501 3027 10567 3030
rect 14549 3027 14615 3030
rect 20897 3027 20963 3030
rect 9857 2954 9923 2957
rect 10961 2954 11027 2957
rect 18413 2954 18479 2957
rect 9857 2952 10794 2954
rect 9857 2896 9862 2952
rect 9918 2896 10794 2952
rect 9857 2894 10794 2896
rect 9857 2891 9923 2894
rect 10734 2818 10794 2894
rect 10961 2952 18479 2954
rect 10961 2896 10966 2952
rect 11022 2896 18418 2952
rect 18474 2896 18479 2952
rect 10961 2894 18479 2896
rect 10961 2891 11027 2894
rect 18413 2891 18479 2894
rect 20713 2954 20779 2957
rect 22200 2954 23000 2984
rect 20713 2952 23000 2954
rect 20713 2896 20718 2952
rect 20774 2896 23000 2952
rect 20713 2894 23000 2896
rect 20713 2891 20779 2894
rect 22200 2864 23000 2894
rect 14641 2818 14707 2821
rect 10734 2816 14707 2818
rect 10734 2760 14646 2816
rect 14702 2760 14707 2816
rect 10734 2758 14707 2760
rect 14641 2755 14707 2758
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 18137 2546 18203 2549
rect 22200 2546 23000 2576
rect 18137 2544 23000 2546
rect 18137 2488 18142 2544
rect 18198 2488 23000 2544
rect 18137 2486 23000 2488
rect 18137 2483 18203 2486
rect 22200 2456 23000 2486
rect 10133 2412 10199 2413
rect 10133 2410 10180 2412
rect 10052 2408 10180 2410
rect 10244 2410 10250 2412
rect 19149 2410 19215 2413
rect 10244 2408 19215 2410
rect 10052 2352 10138 2408
rect 10244 2352 19154 2408
rect 19210 2352 19215 2408
rect 10052 2350 10180 2352
rect 10133 2348 10180 2350
rect 10244 2350 19215 2352
rect 10244 2348 10250 2350
rect 10133 2347 10199 2348
rect 19149 2347 19215 2350
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 16205 2002 16271 2005
rect 17585 2002 17651 2005
rect 22200 2002 23000 2032
rect 16205 2000 23000 2002
rect 16205 1944 16210 2000
rect 16266 1944 17590 2000
rect 17646 1944 23000 2000
rect 16205 1942 23000 1944
rect 16205 1939 16271 1942
rect 17585 1939 17651 1942
rect 22200 1912 23000 1942
rect 14181 1594 14247 1597
rect 22200 1594 23000 1624
rect 14181 1592 23000 1594
rect 14181 1536 14186 1592
rect 14242 1536 23000 1592
rect 14181 1534 23000 1536
rect 14181 1531 14247 1534
rect 22200 1504 23000 1534
rect 18873 1050 18939 1053
rect 22200 1050 23000 1080
rect 18873 1048 23000 1050
rect 18873 992 18878 1048
rect 18934 992 23000 1048
rect 18873 990 23000 992
rect 18873 987 18939 990
rect 22200 960 23000 990
rect 15285 642 15351 645
rect 22200 642 23000 672
rect 15285 640 23000 642
rect 15285 584 15290 640
rect 15346 584 23000 640
rect 15285 582 23000 584
rect 15285 579 15351 582
rect 22200 552 23000 582
rect 17769 234 17835 237
rect 22200 234 23000 264
rect 17769 232 23000 234
rect 17769 176 17774 232
rect 17830 176 23000 232
rect 17769 174 23000 176
rect 17769 171 17835 174
rect 22200 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 13492 17580 13556 17644
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 10548 15736 10612 15740
rect 10548 15680 10598 15736
rect 10598 15680 10612 15736
rect 10548 15676 10612 15680
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 10364 15132 10428 15196
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 12204 14452 12268 14516
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 18092 13228 18156 13292
rect 18828 13228 18892 13292
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 13492 12412 13556 12476
rect 14596 12472 14660 12476
rect 14596 12416 14646 12472
rect 14646 12416 14660 12472
rect 14596 12412 14660 12416
rect 10548 12336 10612 12340
rect 10548 12280 10598 12336
rect 10598 12280 10612 12336
rect 10548 12276 10612 12280
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 10364 10976 10428 10980
rect 10364 10920 10378 10976
rect 10378 10920 10428 10976
rect 10364 10916 10428 10920
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 18828 10840 18892 10844
rect 18828 10784 18878 10840
rect 18878 10784 18892 10840
rect 18828 10780 18892 10784
rect 18092 10644 18156 10708
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 14596 9692 14660 9756
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 12204 8196 12268 8260
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 10180 7440 10244 7444
rect 10180 7384 10194 7440
rect 10194 7384 10244 7440
rect 10180 7380 10244 7384
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 10180 2408 10244 2412
rect 10180 2352 10194 2408
rect 10194 2352 10244 2408
rect 10180 2348 10244 2352
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 13491 17644 13557 17645
rect 13491 17580 13492 17644
rect 13556 17580 13557 17644
rect 13491 17579 13557 17580
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 10547 15740 10613 15741
rect 10547 15676 10548 15740
rect 10612 15676 10613 15740
rect 10547 15675 10613 15676
rect 10363 15196 10429 15197
rect 10363 15132 10364 15196
rect 10428 15132 10429 15196
rect 10363 15131 10429 15132
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 10366 10981 10426 15131
rect 10550 12341 10610 15675
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 12203 14516 12269 14517
rect 12203 14452 12204 14516
rect 12268 14452 12269 14516
rect 12203 14451 12269 14452
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 10547 12340 10613 12341
rect 10547 12276 10548 12340
rect 10612 12276 10613 12340
rect 10547 12275 10613 12276
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 10363 10980 10429 10981
rect 10363 10916 10364 10980
rect 10428 10916 10429 10980
rect 10363 10915 10429 10916
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 12206 8261 12266 14451
rect 13494 12477 13554 17579
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18091 13292 18157 13293
rect 18091 13228 18092 13292
rect 18156 13228 18157 13292
rect 18091 13227 18157 13228
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 13491 12476 13557 12477
rect 13491 12412 13492 12476
rect 13556 12412 13557 12476
rect 13491 12411 13557 12412
rect 14595 12476 14661 12477
rect 14595 12412 14596 12476
rect 14660 12412 14661 12476
rect 14595 12411 14661 12412
rect 14598 9757 14658 12411
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 18094 10709 18154 13227
rect 18270 13088 18591 14112
rect 18827 13292 18893 13293
rect 18827 13228 18828 13292
rect 18892 13228 18893 13292
rect 18827 13227 18893 13228
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18091 10708 18157 10709
rect 18091 10644 18092 10708
rect 18156 10644 18157 10708
rect 18091 10643 18157 10644
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14595 9756 14661 9757
rect 14595 9692 14596 9756
rect 14660 9692 14661 9756
rect 14595 9691 14661 9692
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 12203 8260 12269 8261
rect 12203 8196 12204 8260
rect 12268 8196 12269 8260
rect 12203 8195 12269 8196
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 10179 7444 10245 7445
rect 10179 7380 10180 7444
rect 10244 7380 10245 7444
rect 10179 7379 10245 7380
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 10182 2413 10242 7379
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 10179 2412 10245 2413
rect 10179 2348 10180 2412
rect 10244 2348 10245 2412
rect 10179 2347 10245 2348
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 9824 18591 10848
rect 18830 10845 18890 13227
rect 18827 10844 18893 10845
rect 18827 10780 18828 10844
rect 18892 10780 18893 10844
rect 18827 10779 18893 10780
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__decap_12  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608910539
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1608910539
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608910539
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608910539
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_82 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8648 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_74
timestamp 1608910539
transform 1 0 7912 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_83
timestamp 1608910539
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79
timestamp 1608910539
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75
timestamp 1608910539
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1608910539
transform 1 0 8556 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1608910539
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87
timestamp 1608910539
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1608910539
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1608910539
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp 1608910539
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_89
timestamp 1608910539
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1608910539
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1608910539
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1608910539
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_97
timestamp 1608910539
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1608910539
transform 1 0 10028 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1608910539
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 10212 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_103
timestamp 1608910539
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1608910539
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1608910539
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107
timestamp 1608910539
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11132 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_123
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1608910539
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1608910539
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_115
timestamp 1608910539
transform 1 0 11684 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608910539
transform 1 0 11960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608910539
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12512 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1608910539
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_130
timestamp 1608910539
transform 1 0 13064 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1608910539
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_139
timestamp 1608910539
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1608910539
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13432 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13340 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14444 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608910539
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1608910539
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_159
timestamp 1608910539
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1608910539
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 15548 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15916 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16100 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608910539
transform 1 0 14628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1608910539
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1608910539
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1608910539
transform 1 0 17756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_170
timestamp 1608910539
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16928 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1608910539
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1608910539
transform 1 0 19228 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191
timestamp 1608910539
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19044 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608910539
transform 1 0 18860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_204
timestamp 1608910539
transform 1 0 19872 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1608910539
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20148 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608910539
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608910539
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_213
timestamp 1608910539
transform 1 0 20700 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1608910539
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608910539
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1608910539
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608910539
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1608910539
transform 1 0 21252 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_220
timestamp 1608910539
transform 1 0 21344 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608910539
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608910539
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1608910539
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608910539
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_80
timestamp 1608910539
transform 1 0 8464 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1608910539
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_103
timestamp 1608910539
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_99
timestamp 1608910539
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_95
timestamp 1608910539
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1608910539
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1608910539
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1608910539
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_118
timestamp 1608910539
transform 1 0 11960 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_114
timestamp 1608910539
transform 1 0 11592 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10764 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12052 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_140
timestamp 1608910539
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_135
timestamp 1608910539
transform 1 0 13524 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1608910539
transform 1 0 16284 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_157
timestamp 1608910539
transform 1 0 15548 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1608910539
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15732 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _040_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_185
timestamp 1608910539
transform 1 0 18124 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18308 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16652 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_203
timestamp 1608910539
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19964 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1608910539
transform 1 0 21252 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_211
timestamp 1608910539
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608910539
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608910539
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608910539
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608910539
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608910539
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608910539
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1608910539
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_74
timestamp 1608910539
transform 1 0 7912 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1608910539
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_90
timestamp 1608910539
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_86
timestamp 1608910539
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1608910539
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1608910539
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9568 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10580 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1608910539
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608910539
transform 1 0 12512 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_128
timestamp 1608910539
transform 1 0 12880 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13248 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1608910539
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_154
timestamp 1608910539
transform 1 0 15272 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_148
timestamp 1608910539
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15548 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608910539
transform 1 0 14904 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1608910539
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1608910539
transform 1 0 17480 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1608910539
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608910539
transform 1 0 17112 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608910539
transform 1 0 16560 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_206
timestamp 1608910539
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1608910539
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1608910539
transform 1 0 20240 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18584 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1608910539
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_217
timestamp 1608910539
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608910539
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608910539
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1608910539
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1608910539
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1608910539
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1608910539
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1608910539
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_86
timestamp 1608910539
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1608910539
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_4_125
timestamp 1608910539
transform 1 0 12604 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_120
timestamp 1608910539
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_109
timestamp 1608910539
transform 1 0 11132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11316 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1608910539
transform 1 0 12328 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1608910539
transform 1 0 14352 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12880 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1608910539
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1608910539
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1608910539
transform 1 0 16284 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608910539
transform 1 0 14720 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_183
timestamp 1608910539
transform 1 0 17940 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_179
timestamp 1608910539
transform 1 0 17572 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_174
timestamp 1608910539
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608910539
transform 1 0 18032 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608910539
transform 1 0 17296 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_199
timestamp 1608910539
transform 1 0 19412 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1608910539
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18584 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1608910539
transform 1 0 19596 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1608910539
transform 1 0 21252 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1608910539
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608910539
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608910539
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1608910539
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608910539
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608910539
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1608910539
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_81
timestamp 1608910539
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_78
timestamp 1608910539
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_74
timestamp 1608910539
transform 1 0 7912 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_97
timestamp 1608910539
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1608910539
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_89
timestamp 1608910539
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1608910539
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1608910539
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10212 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1608910539
transform 1 0 12604 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp 1608910539
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_108
timestamp 1608910539
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11224 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_143
timestamp 1608910539
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_138
timestamp 1608910539
transform 1 0 13800 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12972 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14444 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_161
timestamp 1608910539
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 16100 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_179
timestamp 1608910539
transform 1 0 17572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_200
timestamp 1608910539
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 19688 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1608910539
transform 1 0 21528 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1608910539
transform 1 0 21160 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608910539
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608910539
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1608910539
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608910539
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608910539
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608910539
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1608910539
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp 1608910539
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_56
timestamp 1608910539
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1608910539
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_72
timestamp 1608910539
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_68
timestamp 1608910539
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1608910539
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_78
timestamp 1608910539
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7912 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_90
timestamp 1608910539
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1608910539
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_86
timestamp 1608910539
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608910539
transform 1 0 9568 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_99
timestamp 1608910539
transform 1 0 10212 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_95
timestamp 1608910539
transform 1 0 9844 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_98
timestamp 1608910539
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10304 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10304 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_109
timestamp 1608910539
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11316 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_125
timestamp 1608910539
transform 1 0 12604 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1608910539
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_121
timestamp 1608910539
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_116
timestamp 1608910539
transform 1 0 11776 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12052 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12420 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_142
timestamp 1608910539
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_131
timestamp 1608910539
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_139
timestamp 1608910539
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 14076 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13340 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1608910539
transform 1 0 12880 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_150
timestamp 1608910539
transform 1 0 14904 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_146
timestamp 1608910539
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp 1608910539
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15272 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_163
timestamp 1608910539
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1608910539
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16284 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 16284 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_186
timestamp 1608910539
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1608910539
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_174
timestamp 1608910539
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_174
timestamp 1608910539
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 17296 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608910539
transform 1 0 17296 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_190
timestamp 1608910539
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1608910539
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_192
timestamp 1608910539
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608910539
transform 1 0 18952 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_208
timestamp 1608910539
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_201
timestamp 1608910539
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 19412 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19780 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18768 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1608910539
transform 1 0 21252 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1608910539
transform 1 0 21252 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1608910539
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 20424 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608910539
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608910539
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608910539
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_56
timestamp 1608910539
transform 1 0 6256 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1608910539
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1608910539
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1608910539
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_64
timestamp 1608910539
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1608910539
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1608910539
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10672 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_122
timestamp 1608910539
transform 1 0 12328 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_118
timestamp 1608910539
transform 1 0 11960 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_113
timestamp 1608910539
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11684 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12420 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_139
timestamp 1608910539
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1608910539
transform 1 0 14076 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_160
timestamp 1608910539
transform 1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_156
timestamp 1608910539
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp 1608910539
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 15640 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16100 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_172
timestamp 1608910539
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 17112 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1608910539
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 1608910539
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 19136 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1608910539
transform 1 0 21528 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_218
timestamp 1608910539
transform 1 0 21160 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1608910539
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608910539
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1608910539
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1608910539
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1608910539
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608910539
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1608910539
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_77
timestamp 1608910539
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_73
timestamp 1608910539
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_70
timestamp 1608910539
transform 1 0 7544 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 8372 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_95
timestamp 1608910539
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10028 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_125
timestamp 1608910539
transform 1 0 12604 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp 1608910539
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1608910539
transform 1 0 11500 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_143
timestamp 1608910539
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1608910539
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_129
timestamp 1608910539
transform 1 0 12972 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13432 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1608910539
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_147
timestamp 1608910539
transform 1 0 14628 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 14904 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1608910539
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_170
timestamp 1608910539
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1608910539
transform 1 0 16928 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_198
timestamp 1608910539
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1608910539
transform 1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1608910539
transform 1 0 19504 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_220
timestamp 1608910539
transform 1 0 21344 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_209
timestamp 1608910539
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1608910539
transform 1 0 20516 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1608910539
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608910539
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1608910539
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1608910539
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1608910539
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_78
timestamp 1608910539
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_68
timestamp 1608910539
transform 1 0 7360 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1608910539
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608910539
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8832 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_117
timestamp 1608910539
transform 1 0 11868 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_106
timestamp 1608910539
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11040 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12236 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1608910539
transform 1 0 14076 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_137
timestamp 1608910539
transform 1 0 13708 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1608910539
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_180
timestamp 1608910539
transform 1 0 17664 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_175
timestamp 1608910539
transform 1 0 17204 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_170
timestamp 1608910539
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 16928 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 17848 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1608910539
transform 1 0 19044 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1608910539
transform 1 0 18676 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19136 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_222
timestamp 1608910539
transform 1 0 21528 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_218
timestamp 1608910539
transform 1 0 21160 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1608910539
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1608910539
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1608910539
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1608910539
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1608910539
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608910539
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1608910539
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1608910539
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_74
timestamp 1608910539
transform 1 0 7912 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_88
timestamp 1608910539
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1608910539
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9384 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1608910539
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1608910539
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_106
timestamp 1608910539
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11040 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_143
timestamp 1608910539
transform 1 0 14260 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1608910539
transform 1 0 13892 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14352 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_160
timestamp 1608910539
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16008 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_187
timestamp 1608910539
transform 1 0 18308 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_180
timestamp 1608910539
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_176
timestamp 1608910539
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_171
timestamp 1608910539
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 17020 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1608910539
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18676 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 19688 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_222
timestamp 1608910539
transform 1 0 21528 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_218
timestamp 1608910539
transform 1 0 21160 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1608910539
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608910539
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1608910539
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1608910539
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1608910539
transform 1 0 8464 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1608910539
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_99
timestamp 1608910539
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_93
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1608910539
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_86
timestamp 1608910539
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10396 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608910539
transform 1 0 9936 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_121
timestamp 1608910539
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1608910539
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 12420 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 11408 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_137
timestamp 1608910539
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_126
timestamp 1608910539
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 12880 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13892 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1608910539
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1608910539
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_148
timestamp 1608910539
transform 1 0 14720 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_172
timestamp 1608910539
transform 1 0 16928 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_167
timestamp 1608910539
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 16652 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 17112 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_201
timestamp 1608910539
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_190
timestamp 1608910539
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18768 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19780 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1608910539
transform 1 0 21528 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1608910539
transform 1 0 21160 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1608910539
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1608910539
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1608910539
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1608910539
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1608910539
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1608910539
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1608910539
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1608910539
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1608910539
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608910539
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1608910539
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1608910539
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1608910539
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_82
timestamp 1608910539
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_74
timestamp 1608910539
transform 1 0 7912 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1608910539
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_86
timestamp 1608910539
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_86
timestamp 1608910539
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_98
timestamp 1608910539
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_104
timestamp 1608910539
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10304 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9200 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_116
timestamp 1608910539
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_125
timestamp 1608910539
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1608910539
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_115
timestamp 1608910539
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 11868 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10856 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 11960 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_14_145
timestamp 1608910539
transform 1 0 14444 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_134
timestamp 1608910539
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_145
timestamp 1608910539
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_141
timestamp 1608910539
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_130
timestamp 1608910539
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 12788 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13248 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1608910539
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1608910539
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 14628 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608910539
transform 1 0 14720 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1608910539
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_161
timestamp 1608910539
transform 1 0 15916 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16284 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1608910539
transform 1 0 15640 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16284 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_183
timestamp 1608910539
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_171
timestamp 1608910539
transform 1 0 16836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_184
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1608910539
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18124 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1608910539
transform 1 0 17112 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18308 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_14_199
timestamp 1608910539
transform 1 0 19412 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1608910539
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_207
timestamp 1608910539
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_203
timestamp 1608910539
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1608910539
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19688 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608910539
transform 1 0 19136 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1608910539
transform 1 0 21068 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1608910539
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_218
timestamp 1608910539
transform 1 0 21160 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1608910539
transform 1 0 20332 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1608910539
transform 1 0 21436 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_222
timestamp 1608910539
transform 1 0 21528 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 21252 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1608910539
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1608910539
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1608910539
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608910539
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1608910539
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_74
timestamp 1608910539
transform 1 0 7912 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_103
timestamp 1608910539
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1608910539
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 1608910539
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 9016 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9752 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_123
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1608910539
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_114
timestamp 1608910539
transform 1 0 11592 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_135
timestamp 1608910539
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13708 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12696 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1608910539
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_146
timestamp 1608910539
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1608910539
transform 1 0 15732 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 14720 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608910539
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_168
timestamp 1608910539
transform 1 0 16560 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16928 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_197
timestamp 1608910539
transform 1 0 19228 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_193
timestamp 1608910539
transform 1 0 18860 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 19320 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_220
timestamp 1608910539
transform 1 0 21344 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_214
timestamp 1608910539
transform 1 0 20792 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1608910539
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608910539
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1608910539
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1608910539
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1608910539
transform 1 0 8464 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1608910539
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_102
timestamp 1608910539
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608910539
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_86
timestamp 1608910539
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_111
timestamp 1608910539
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_106
timestamp 1608910539
transform 1 0 10856 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11500 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1608910539
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 13156 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_16_157
timestamp 1608910539
transform 1 0 15548 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1608910539
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15916 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_177
timestamp 1608910539
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 17572 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1608910539
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_195
timestamp 1608910539
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_222
timestamp 1608910539
transform 1 0 21528 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1608910539
transform 1 0 21160 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1608910539
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608910539
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1608910539
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1608910539
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1608910539
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608910539
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1608910539
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_80
timestamp 1608910539
transform 1 0 8464 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_74
timestamp 1608910539
transform 1 0 7912 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8556 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_97
timestamp 1608910539
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10212 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1608910539
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_115
timestamp 1608910539
transform 1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1608910539
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_126
timestamp 1608910539
transform 1 0 12696 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12972 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_163
timestamp 1608910539
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14628 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1608910539
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_171
timestamp 1608910539
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_167
timestamp 1608910539
transform 1 0 16468 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16928 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_208
timestamp 1608910539
transform 1 0 20240 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_190
timestamp 1608910539
transform 1 0 18584 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18768 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_220
timestamp 1608910539
transform 1 0 21344 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1608910539
transform 1 0 20516 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1608910539
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608910539
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1608910539
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1608910539
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_81
timestamp 1608910539
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1608910539
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_74
timestamp 1608910539
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_68
timestamp 1608910539
transform 1 0 7360 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_102
timestamp 1608910539
transform 1 0 10488 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1608910539
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1608910539
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608910539
transform 1 0 9108 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_121
timestamp 1608910539
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12420 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10764 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_140
timestamp 1608910539
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_132
timestamp 1608910539
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13432 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1608910539
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_181
timestamp 1608910539
transform 1 0 17756 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1608910539
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1608910539
transform 1 0 18032 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 16928 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1608910539
transform 1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 19136 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1608910539
transform 1 0 21252 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1608910539
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608910539
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608910539
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1608910539
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1608910539
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1608910539
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1608910539
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1608910539
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_56
timestamp 1608910539
transform 1 0 6256 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1608910539
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_62
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608910539
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1608910539
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1608910539
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1608910539
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_70
timestamp 1608910539
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1608910539
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_78
timestamp 1608910539
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_74
timestamp 1608910539
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_74
timestamp 1608910539
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8096 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1608910539
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_96
timestamp 1608910539
transform 1 0 9936 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_92
timestamp 1608910539
transform 1 0 9568 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10028 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8832 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9752 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1608910539
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_106
timestamp 1608910539
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1608910539
transform 1 0 11040 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11408 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_121
timestamp 1608910539
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1608910539
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_117
timestamp 1608910539
transform 1 0 11868 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1608910539
transform 1 0 12420 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_140
timestamp 1608910539
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_132
timestamp 1608910539
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_140
timestamp 1608910539
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_129
timestamp 1608910539
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13432 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1608910539
transform 1 0 13156 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 14168 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1608910539
transform 1 0 14168 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_154
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1608910539
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_151
timestamp 1608910539
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15180 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15364 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_164
timestamp 1608910539
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_159
timestamp 1608910539
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15916 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16376 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_182
timestamp 1608910539
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1608910539
transform 1 0 18308 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1608910539
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1608910539
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16928 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18032 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1608910539
transform 1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_207
timestamp 1608910539
transform 1 0 20148 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 19136 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18676 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1608910539
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1608910539
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1608910539
transform 1 0 21252 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608910539
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1608910539
transform 1 0 20424 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20884 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1608910539
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1608910539
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1608910539
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1608910539
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1608910539
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_64
timestamp 1608910539
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_68
timestamp 1608910539
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7544 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_72
timestamp 1608910539
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_76
timestamp 1608910539
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_80
timestamp 1608910539
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1608910539
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp 1608910539
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_88
timestamp 1608910539
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_84
timestamp 1608910539
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 9752 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10212 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1608910539
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_115
timestamp 1608910539
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608910539
transform 1 0 11868 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1608910539
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608910539
transform 1 0 14076 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1608910539
transform 1 0 16376 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1608910539
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_150
timestamp 1608910539
transform 1 0 14904 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1608910539
transform 1 0 15180 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1608910539
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_177
timestamp 1608910539
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 16560 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_193
timestamp 1608910539
transform 1 0 18860 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 19228 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1608910539
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_213
timestamp 1608910539
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20884 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1608910539
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608910539
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1608910539
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1608910539
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_76
timestamp 1608910539
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_72
timestamp 1608910539
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_68
timestamp 1608910539
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_64
timestamp 1608910539
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8280 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1608910539
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1608910539
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_120
timestamp 1608910539
transform 1 0 12144 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1608910539
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11316 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12512 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_133
timestamp 1608910539
transform 1 0 13340 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13524 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1608910539
transform 1 0 16100 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1608910539
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1608910539
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18124 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 16468 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_201
timestamp 1608910539
transform 1 0 19596 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1608910539
transform 1 0 19780 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_219
timestamp 1608910539
transform 1 0 21252 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1608910539
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608910539
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1608910539
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1608910539
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1608910539
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1608910539
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_62
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1608910539
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_51
timestamp 1608910539
transform 1 0 5796 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1608910539
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_74
timestamp 1608910539
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_70
timestamp 1608910539
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_65
timestamp 1608910539
transform 1 0 7084 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6900 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8464 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_102
timestamp 1608910539
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_97
timestamp 1608910539
transform 1 0 10028 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_89
timestamp 1608910539
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 10672 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 9476 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1608910539
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1608910539
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1608910539
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_106
timestamp 1608910539
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 11408 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_142
timestamp 1608910539
transform 1 0 14168 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_129
timestamp 1608910539
transform 1 0 12972 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13340 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_163
timestamp 1608910539
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_146
timestamp 1608910539
transform 1 0 14536 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 16284 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 14628 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_187
timestamp 1608910539
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1608910539
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_174
timestamp 1608910539
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 17296 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608910539
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_205
timestamp 1608910539
transform 1 0 19964 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1608910539
transform 1 0 20148 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18492 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1608910539
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_216
timestamp 1608910539
transform 1 0 20976 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608910539
transform 1 0 21160 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1608910539
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1608910539
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_61
timestamp 1608910539
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_57
timestamp 1608910539
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_53
timestamp 1608910539
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_50
timestamp 1608910539
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_44
timestamp 1608910539
transform 1 0 5152 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6532 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_76
timestamp 1608910539
transform 1 0 8096 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_65
timestamp 1608910539
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8372 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7268 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_96
timestamp 1608910539
transform 1 0 9936 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1608910539
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10212 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_119
timestamp 1608910539
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_108
timestamp 1608910539
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1608910539
transform 1 0 12236 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1608910539
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_130
timestamp 1608910539
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13248 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608910539
transform 1 0 14260 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_158
timestamp 1608910539
transform 1 0 15640 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_154
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1608910539
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_146
timestamp 1608910539
transform 1 0 14536 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 15916 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608910539
transform 1 0 15364 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608910539
transform 1 0 14720 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_175
timestamp 1608910539
transform 1 0 17204 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1608910539
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 17480 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1608910539
transform 1 0 16928 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_205
timestamp 1608910539
transform 1 0 19964 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1608910539
transform 1 0 18952 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19136 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608910539
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1608910539
transform 1 0 21252 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1608910539
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608910539
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1608910539
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1608910539
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1608910539
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1608910539
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1608910539
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_51
timestamp 1608910539
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1608910539
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 8464 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_96
timestamp 1608910539
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10120 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1608910539
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_114
timestamp 1608910539
transform 1 0 11592 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1608910539
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13432 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_161
timestamp 1608910539
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_150
timestamp 1608910539
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16100 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1608910539
transform 1 0 15088 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_184
timestamp 1608910539
transform 1 0 18032 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1608910539
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1608910539
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608910539
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17112 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608910539
transform 1 0 18124 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_200
timestamp 1608910539
transform 1 0 19504 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_189
timestamp 1608910539
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19872 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18676 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1608910539
transform 1 0 21252 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_213
timestamp 1608910539
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608910539
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1608910539
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1608910539
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1608910539
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1608910539
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1608910539
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_44
timestamp 1608910539
transform 1 0 5152 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_51
timestamp 1608910539
transform 1 0 5796 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_53
timestamp 1608910539
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_50
timestamp 1608910539
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6164 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1608910539
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_61
timestamp 1608910539
transform 1 0 6716 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1608910539
transform 1 0 6348 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6532 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608910539
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_80
timestamp 1608910539
transform 1 0 8464 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_83
timestamp 1608910539
transform 1 0 8740 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_65
timestamp 1608910539
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6900 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7268 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6992 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_89
timestamp 1608910539
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1608910539
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1608910539
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_87
timestamp 1608910539
transform 1 0 9108 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1608910539
transform 1 0 9476 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_100
timestamp 1608910539
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_103
timestamp 1608910539
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1608910539
transform 1 0 10120 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 9936 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 10304 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 10488 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1608910539
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_108
timestamp 1608910539
transform 1 0 11040 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_121
timestamp 1608910539
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608910539
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11316 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10764 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_144
timestamp 1608910539
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_126
timestamp 1608910539
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_139
timestamp 1608910539
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14076 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12880 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1608910539
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_155
timestamp 1608910539
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1608910539
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1608910539
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15548 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1608910539
transform 1 0 14536 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1608910539
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1608910539
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16560 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16652 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_184
timestamp 1608910539
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1608910539
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_187
timestamp 1608910539
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_182
timestamp 1608910539
transform 1 0 17848 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_178
timestamp 1608910539
transform 1 0 17480 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608910539
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608910539
transform 1 0 17940 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18308 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_27_203
timestamp 1608910539
transform 1 0 19780 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_203
timestamp 1608910539
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_198
timestamp 1608910539
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19964 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18492 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20056 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608910539
transform 1 0 19504 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_220
timestamp 1608910539
transform 1 0 21344 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_212
timestamp 1608910539
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1608910539
transform 1 0 21252 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_211
timestamp 1608910539
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608910539
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20792 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608910539
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1608910539
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1608910539
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608910539
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1608910539
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1608910539
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608910539
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_60
timestamp 1608910539
transform 1 0 6624 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_56
timestamp 1608910539
transform 1 0 6256 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1608910539
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_67
timestamp 1608910539
transform 1 0 7268 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1608910539
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7636 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1608910539
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1608910539
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_87
timestamp 1608910539
transform 1 0 9108 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608910539
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10672 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_118
timestamp 1608910539
transform 1 0 11960 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_113
timestamp 1608910539
transform 1 0 11500 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1608910539
transform 1 0 11776 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12144 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_142
timestamp 1608910539
transform 1 0 14168 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_131
timestamp 1608910539
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_126
timestamp 1608910539
transform 1 0 12696 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1608910539
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13340 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_160
timestamp 1608910539
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1608910539
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_146
timestamp 1608910539
transform 1 0 14536 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608910539
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15272 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16008 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1608910539
transform 1 0 14628 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_178
timestamp 1608910539
transform 1 0 17480 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 17664 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_207
timestamp 1608910539
transform 1 0 20148 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_196
timestamp 1608910539
transform 1 0 19136 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19320 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1608910539
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1608910539
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608910539
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608910539
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20884 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1608910539
transform 1 0 20332 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1608910539
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1608910539
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608910539
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1608910539
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1608910539
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1608910539
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1608910539
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1608910539
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608910539
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_78
timestamp 1608910539
transform 1 0 8280 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_67
timestamp 1608910539
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7452 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 8648 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_29_103
timestamp 1608910539
transform 1 0 10580 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_98
timestamp 1608910539
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1608910539
transform 1 0 10304 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1608910539
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_116
timestamp 1608910539
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_108
timestamp 1608910539
transform 1 0 11040 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1608910539
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608910539
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11224 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_141
timestamp 1608910539
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_136
timestamp 1608910539
transform 1 0 13616 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp 1608910539
transform 1 0 13248 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 14260 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1608910539
transform 1 0 13708 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1608910539
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_159
timestamp 1608910539
transform 1 0 15732 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1608910539
transform 1 0 16008 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1608910539
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_177
timestamp 1608910539
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1608910539
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608910539
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16560 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18032 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_200
timestamp 1608910539
transform 1 0 19504 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19688 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_222
timestamp 1608910539
transform 1 0 21528 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_218
timestamp 1608910539
transform 1 0 21160 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_211
timestamp 1608910539
transform 1 0 20516 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608910539
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608910539
transform 1 0 20792 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1608910539
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1608910539
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608910539
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1608910539
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1608910539
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608910539
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1608910539
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1608910539
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1608910539
transform 1 0 8648 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_78
timestamp 1608910539
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_68
timestamp 1608910539
transform 1 0 7360 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 8096 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 8464 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1608910539
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_86
timestamp 1608910539
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1608910539
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608910539
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1608910539
transform 1 0 12144 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_109
timestamp 1608910539
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1608910539
transform 1 0 12328 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11316 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_141
timestamp 1608910539
transform 1 0 14076 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_137
timestamp 1608910539
transform 1 0 13708 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_131
timestamp 1608910539
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608910539
transform 1 0 13340 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1608910539
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1608910539
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608910539
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15456 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_184
timestamp 1608910539
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_178
timestamp 1608910539
transform 1 0 17480 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_172
timestamp 1608910539
transform 1 0 16928 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1608910539
transform 1 0 17664 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1608910539
transform 1 0 17112 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608910539
transform 1 0 18216 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_205
timestamp 1608910539
transform 1 0 19964 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_201
timestamp 1608910539
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1608910539
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18768 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608910539
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1608910539
transform 1 0 21252 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1608910539
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608910539
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608910539
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608910539
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1608910539
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1608910539
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608910539
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1608910539
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1608910539
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1608910539
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1608910539
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1608910539
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608910539
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_83
timestamp 1608910539
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_79
timestamp 1608910539
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_74
timestamp 1608910539
transform 1 0 7912 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608910539
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_95
timestamp 1608910539
transform 1 0 9844 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1608910539
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_87
timestamp 1608910539
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 8924 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10212 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1608910539
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_115
timestamp 1608910539
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608910539
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1608910539
transform 1 0 11868 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1608910539
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14076 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_157
timestamp 1608910539
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15732 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1608910539
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1608910539
transform 1 0 17480 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_168
timestamp 1608910539
transform 1 0 16560 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608910539
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16928 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_203
timestamp 1608910539
transform 1 0 19780 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_199
timestamp 1608910539
transform 1 0 19412 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_190
timestamp 1608910539
transform 1 0 18584 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 19872 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 18860 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_220
timestamp 1608910539
transform 1 0 21344 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_216
timestamp 1608910539
transform 1 0 20976 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608910539
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1608910539
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1608910539
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608910539
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1608910539
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1608910539
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608910539
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1608910539
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1608910539
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1608910539
transform 1 0 8464 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1608910539
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_95
timestamp 1608910539
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1608910539
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_86
timestamp 1608910539
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608910539
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10028 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1608910539
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_106
timestamp 1608910539
transform 1 0 10856 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11132 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1608910539
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_139
timestamp 1608910539
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_129
timestamp 1608910539
transform 1 0 12972 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13064 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608910539
transform 1 0 14076 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_163
timestamp 1608910539
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1608910539
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608910539
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1608910539
transform 1 0 16284 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608910539
transform 1 0 14628 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_186
timestamp 1608910539
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_180
timestamp 1608910539
transform 1 0 17664 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_175
timestamp 1608910539
transform 1 0 17204 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_169
timestamp 1608910539
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1608910539
transform 1 0 16836 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608910539
transform 1 0 17848 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1608910539
transform 1 0 17388 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_206
timestamp 1608910539
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_200
timestamp 1608910539
transform 1 0 19504 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_196
timestamp 1608910539
transform 1 0 19136 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_190
timestamp 1608910539
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 19320 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1608910539
transform 1 0 18400 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608910539
transform 1 0 18768 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608910539
transform 1 0 19688 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608910539
transform 1 0 20240 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1608910539
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1608910539
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608910539
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608910539
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20884 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1608910539
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1608910539
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608910539
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1608910539
transform 1 0 4048 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1608910539
transform 1 0 3588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608910539
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_56
timestamp 1608910539
transform 1 0 6256 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1608910539
transform 1 0 5152 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608910539
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_75
timestamp 1608910539
transform 1 0 8004 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_63
timestamp 1608910539
transform 1 0 6900 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_87
timestamp 1608910539
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1608910539
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_91
timestamp 1608910539
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_94
timestamp 1608910539
transform 1 0 9752 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608910539
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_97
timestamp 1608910539
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1608910539
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1608910539
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_101
timestamp 1608910539
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1608910539
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_122
timestamp 1608910539
transform 1 0 12328 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_117
timestamp 1608910539
transform 1 0 11868 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_111
timestamp 1608910539
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_105
timestamp 1608910539
transform 1 0 10764 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1608910539
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1608910539
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608910539
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608910539
transform 1 0 11500 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608910539
transform 1 0 10948 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_143
timestamp 1608910539
transform 1 0 14260 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_137
timestamp 1608910539
transform 1 0 13708 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_131
timestamp 1608910539
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_127
timestamp 1608910539
transform 1 0 12788 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1608910539
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1608910539
transform 1 0 13340 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1608910539
transform 1 0 13892 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1608910539
transform 1 0 14444 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1608910539
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_160
timestamp 1608910539
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_153
timestamp 1608910539
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_149
timestamp 1608910539
transform 1 0 14812 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 14996 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608910539
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1608910539
transform 1 0 15456 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1608910539
transform 1 0 16008 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_187
timestamp 1608910539
transform 1 0 18308 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_184
timestamp 1608910539
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_178
timestamp 1608910539
transform 1 0 17480 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_172
timestamp 1608910539
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608910539
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1608910539
transform 1 0 16560 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1608910539
transform 1 0 17112 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1608910539
transform 1 0 17664 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_206
timestamp 1608910539
transform 1 0 20056 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_200
timestamp 1608910539
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_194
timestamp 1608910539
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608910539
transform 1 0 18584 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608910539
transform 1 0 19136 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608910539
transform 1 0 19688 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_220
timestamp 1608910539
transform 1 0 21344 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1608910539
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_210
timestamp 1608910539
transform 1 0 20424 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1608910539
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608910539
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608910539
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608910539
transform 1 0 20516 0 1 20128
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 800 6 bottom_left_grid_pin_1_
port 0 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 ccff_tail
port 2 nsew signal tristate
rlabel metal3 s 22200 3816 23000 3936 6 chanx_right_in[0]
port 3 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[10]
port 4 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[11]
port 5 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[12]
port 6 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[13]
port 7 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[14]
port 8 nsew signal input
rlabel metal3 s 22200 10888 23000 11008 6 chanx_right_in[15]
port 9 nsew signal input
rlabel metal3 s 22200 11296 23000 11416 6 chanx_right_in[16]
port 10 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[17]
port 11 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[18]
port 12 nsew signal input
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_in[19]
port 13 nsew signal input
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[1]
port 14 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[2]
port 15 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[3]
port 16 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[4]
port 17 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[5]
port 18 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[6]
port 19 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[7]
port 20 nsew signal input
rlabel metal3 s 22200 7624 23000 7744 6 chanx_right_in[8]
port 21 nsew signal input
rlabel metal3 s 22200 8032 23000 8152 6 chanx_right_in[9]
port 22 nsew signal input
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_out[0]
port 23 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[10]
port 24 nsew signal tristate
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[11]
port 25 nsew signal tristate
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[12]
port 26 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[13]
port 27 nsew signal tristate
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[14]
port 28 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[15]
port 29 nsew signal tristate
rlabel metal3 s 22200 20680 23000 20800 6 chanx_right_out[16]
port 30 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[17]
port 31 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[18]
port 32 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[19]
port 33 nsew signal tristate
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[1]
port 34 nsew signal tristate
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[2]
port 35 nsew signal tristate
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[3]
port 36 nsew signal tristate
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[4]
port 37 nsew signal tristate
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[5]
port 38 nsew signal tristate
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[6]
port 39 nsew signal tristate
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[7]
port 40 nsew signal tristate
rlabel metal3 s 22200 17008 23000 17128 6 chanx_right_out[8]
port 41 nsew signal tristate
rlabel metal3 s 22200 17416 23000 17536 6 chanx_right_out[9]
port 42 nsew signal tristate
rlabel metal2 s 846 0 902 800 6 chany_bottom_in[0]
port 43 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[10]
port 44 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_in[11]
port 45 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 chany_bottom_in[12]
port 46 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[13]
port 47 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[14]
port 48 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[15]
port 49 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[16]
port 50 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[17]
port 51 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[18]
port 52 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[19]
port 53 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_in[1]
port 54 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 chany_bottom_in[2]
port 55 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 chany_bottom_in[3]
port 56 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 chany_bottom_in[4]
port 57 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 chany_bottom_in[5]
port 58 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_in[6]
port 59 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 chany_bottom_in[7]
port 60 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 chany_bottom_in[8]
port 61 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 chany_bottom_in[9]
port 62 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_out[0]
port 63 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[10]
port 64 nsew signal tristate
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[11]
port 65 nsew signal tristate
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_out[12]
port 66 nsew signal tristate
rlabel metal2 s 19338 0 19394 800 6 chany_bottom_out[13]
port 67 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_out[14]
port 68 nsew signal tristate
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[15]
port 69 nsew signal tristate
rlabel metal2 s 20994 0 21050 800 6 chany_bottom_out[16]
port 70 nsew signal tristate
rlabel metal2 s 21546 0 21602 800 6 chany_bottom_out[17]
port 71 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 chany_bottom_out[18]
port 72 nsew signal tristate
rlabel metal2 s 22650 0 22706 800 6 chany_bottom_out[19]
port 73 nsew signal tristate
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_out[1]
port 74 nsew signal tristate
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_out[2]
port 75 nsew signal tristate
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[3]
port 76 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_out[4]
port 77 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 chany_bottom_out[5]
port 78 nsew signal tristate
rlabel metal2 s 15382 0 15438 800 6 chany_bottom_out[6]
port 79 nsew signal tristate
rlabel metal2 s 15934 0 15990 800 6 chany_bottom_out[7]
port 80 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[8]
port 81 nsew signal tristate
rlabel metal2 s 17038 0 17094 800 6 chany_bottom_out[9]
port 82 nsew signal tristate
rlabel metal2 s 846 22200 902 23000 6 chany_top_in[0]
port 83 nsew signal input
rlabel metal2 s 6458 22200 6514 23000 6 chany_top_in[10]
port 84 nsew signal input
rlabel metal2 s 7010 22200 7066 23000 6 chany_top_in[11]
port 85 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[12]
port 86 nsew signal input
rlabel metal2 s 8114 22200 8170 23000 6 chany_top_in[13]
port 87 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[14]
port 88 nsew signal input
rlabel metal2 s 9218 22200 9274 23000 6 chany_top_in[15]
port 89 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[16]
port 90 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[17]
port 91 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_in[18]
port 92 nsew signal input
rlabel metal2 s 11426 22200 11482 23000 6 chany_top_in[19]
port 93 nsew signal input
rlabel metal2 s 1398 22200 1454 23000 6 chany_top_in[1]
port 94 nsew signal input
rlabel metal2 s 1950 22200 2006 23000 6 chany_top_in[2]
port 95 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 chany_top_in[3]
port 96 nsew signal input
rlabel metal2 s 3054 22200 3110 23000 6 chany_top_in[4]
port 97 nsew signal input
rlabel metal2 s 3606 22200 3662 23000 6 chany_top_in[5]
port 98 nsew signal input
rlabel metal2 s 4158 22200 4214 23000 6 chany_top_in[6]
port 99 nsew signal input
rlabel metal2 s 4710 22200 4766 23000 6 chany_top_in[7]
port 100 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[8]
port 101 nsew signal input
rlabel metal2 s 5814 22200 5870 23000 6 chany_top_in[9]
port 102 nsew signal input
rlabel metal2 s 12070 22200 12126 23000 6 chany_top_out[0]
port 103 nsew signal tristate
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 104 nsew signal tristate
rlabel metal2 s 18234 22200 18290 23000 6 chany_top_out[11]
port 105 nsew signal tristate
rlabel metal2 s 18786 22200 18842 23000 6 chany_top_out[12]
port 106 nsew signal tristate
rlabel metal2 s 19338 22200 19394 23000 6 chany_top_out[13]
port 107 nsew signal tristate
rlabel metal2 s 19890 22200 19946 23000 6 chany_top_out[14]
port 108 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[15]
port 109 nsew signal tristate
rlabel metal2 s 20994 22200 21050 23000 6 chany_top_out[16]
port 110 nsew signal tristate
rlabel metal2 s 21546 22200 21602 23000 6 chany_top_out[17]
port 111 nsew signal tristate
rlabel metal2 s 22098 22200 22154 23000 6 chany_top_out[18]
port 112 nsew signal tristate
rlabel metal2 s 22650 22200 22706 23000 6 chany_top_out[19]
port 113 nsew signal tristate
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_out[1]
port 114 nsew signal tristate
rlabel metal2 s 13174 22200 13230 23000 6 chany_top_out[2]
port 115 nsew signal tristate
rlabel metal2 s 13726 22200 13782 23000 6 chany_top_out[3]
port 116 nsew signal tristate
rlabel metal2 s 14278 22200 14334 23000 6 chany_top_out[4]
port 117 nsew signal tristate
rlabel metal2 s 14830 22200 14886 23000 6 chany_top_out[5]
port 118 nsew signal tristate
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[6]
port 119 nsew signal tristate
rlabel metal2 s 15934 22200 15990 23000 6 chany_top_out[7]
port 120 nsew signal tristate
rlabel metal2 s 16486 22200 16542 23000 6 chany_top_out[8]
port 121 nsew signal tristate
rlabel metal2 s 17038 22200 17094 23000 6 chany_top_out[9]
port 122 nsew signal tristate
rlabel metal3 s 22200 22584 23000 22704 6 prog_clk_0_E_in
port 123 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 124 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 125 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 126 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_37_
port 127 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_38_
port 128 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_39_
port 129 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_40_
port 130 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_41_
port 131 nsew signal input
rlabel metal2 s 294 22200 350 23000 6 top_left_grid_pin_1_
port 132 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 133 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 134 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 135 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 136 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 137 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
