magic
tech sky130A
magscale 1 2
timestamp 1605109083
<< locali >>
rect 21649 5083 21683 5321
rect 19809 2907 19843 3009
rect 23305 2975 23339 3145
<< viali >>
rect 23489 24361 23523 24395
rect 10241 23817 10275 23851
rect 13001 23817 13035 23851
rect 17785 23817 17819 23851
rect 24777 23817 24811 23851
rect 10057 23613 10091 23647
rect 12817 23613 12851 23647
rect 13369 23613 13403 23647
rect 18061 23613 18095 23647
rect 24593 23613 24627 23647
rect 25145 23613 25179 23647
rect 18306 23545 18340 23579
rect 10701 23477 10735 23511
rect 19441 23477 19475 23511
rect 25145 23273 25179 23307
rect 12081 23205 12115 23239
rect 23949 23205 23983 23239
rect 11805 23137 11839 23171
rect 23673 23137 23707 23171
rect 24961 23137 24995 23171
rect 18153 22933 18187 22967
rect 24777 22729 24811 22763
rect 24593 22525 24627 22559
rect 25145 22525 25179 22559
rect 25513 22457 25547 22491
rect 11805 22389 11839 22423
rect 23857 22389 23891 22423
rect 10057 22049 10091 22083
rect 17049 22049 17083 22083
rect 10333 21981 10367 22015
rect 17233 21913 17267 21947
rect 17049 21641 17083 21675
rect 24777 21641 24811 21675
rect 13737 21505 13771 21539
rect 13461 21437 13495 21471
rect 14197 21437 14231 21471
rect 24593 21437 24627 21471
rect 25145 21437 25179 21471
rect 10057 21301 10091 21335
rect 24777 21097 24811 21131
rect 16221 21029 16255 21063
rect 15945 20961 15979 20995
rect 24593 20961 24627 20995
rect 25145 20553 25179 20587
rect 23949 20417 23983 20451
rect 23673 20349 23707 20383
rect 24961 20349 24995 20383
rect 25513 20349 25547 20383
rect 15945 20213 15979 20247
rect 23489 20213 23523 20247
rect 24593 20213 24627 20247
rect 24777 20009 24811 20043
rect 21465 19941 21499 19975
rect 21189 19873 21223 19907
rect 24593 19873 24627 19907
rect 23673 19261 23707 19295
rect 23949 19261 23983 19295
rect 24961 19261 24995 19295
rect 25513 19261 25547 19295
rect 21189 19125 21223 19159
rect 23489 19125 23523 19159
rect 24593 19125 24627 19159
rect 25145 19125 25179 19159
rect 11161 18785 11195 18819
rect 16037 18785 16071 18819
rect 16313 18785 16347 18819
rect 11345 18649 11379 18683
rect 13185 18173 13219 18207
rect 13921 18173 13955 18207
rect 13461 18105 13495 18139
rect 11161 18037 11195 18071
rect 16037 18037 16071 18071
rect 24777 17833 24811 17867
rect 10517 17765 10551 17799
rect 10241 17697 10275 17731
rect 24593 17697 24627 17731
rect 24777 17289 24811 17323
rect 16037 17221 16071 17255
rect 12449 17085 12483 17119
rect 13185 17085 13219 17119
rect 15853 17085 15887 17119
rect 16405 17085 16439 17119
rect 24593 17085 24627 17119
rect 25145 17085 25179 17119
rect 12725 17017 12759 17051
rect 10241 16949 10275 16983
rect 24409 16949 24443 16983
rect 24777 16745 24811 16779
rect 15577 16677 15611 16711
rect 15301 16609 15335 16643
rect 24593 16609 24627 16643
rect 24777 16201 24811 16235
rect 24501 16133 24535 16167
rect 18337 16065 18371 16099
rect 18061 15997 18095 16031
rect 24593 15997 24627 16031
rect 25145 15997 25179 16031
rect 15301 15861 15335 15895
rect 18797 15861 18831 15895
rect 25053 15657 25087 15691
rect 23857 15589 23891 15623
rect 23581 15521 23615 15555
rect 24869 15521 24903 15555
rect 25513 15113 25547 15147
rect 24225 14977 24259 15011
rect 23489 14909 23523 14943
rect 24041 14909 24075 14943
rect 25329 14909 25363 14943
rect 25881 14909 25915 14943
rect 23857 14773 23891 14807
rect 24869 14773 24903 14807
rect 23397 14501 23431 14535
rect 23121 14433 23155 14467
rect 24593 14433 24627 14467
rect 20913 14365 20947 14399
rect 24777 14229 24811 14263
rect 24777 14025 24811 14059
rect 25145 14025 25179 14059
rect 23121 13821 23155 13855
rect 24593 13821 24627 13855
rect 19349 13685 19383 13719
rect 21281 13685 21315 13719
rect 22293 13685 22327 13719
rect 24409 13685 24443 13719
rect 20913 13481 20947 13515
rect 21281 13481 21315 13515
rect 23121 13481 23155 13515
rect 24777 13481 24811 13515
rect 16313 13345 16347 13379
rect 21373 13345 21407 13379
rect 23029 13345 23063 13379
rect 24593 13345 24627 13379
rect 18153 13277 18187 13311
rect 18889 13277 18923 13311
rect 21465 13277 21499 13311
rect 23213 13277 23247 13311
rect 17785 13141 17819 13175
rect 20085 13141 20119 13175
rect 22661 13141 22695 13175
rect 23857 13141 23891 13175
rect 16313 12937 16347 12971
rect 21097 12937 21131 12971
rect 22385 12937 22419 12971
rect 23397 12937 23431 12971
rect 24593 12937 24627 12971
rect 25789 12937 25823 12971
rect 18429 12869 18463 12903
rect 18981 12801 19015 12835
rect 19809 12801 19843 12835
rect 20545 12801 20579 12835
rect 24133 12801 24167 12835
rect 18337 12733 18371 12767
rect 18797 12733 18831 12767
rect 20361 12733 20395 12767
rect 23857 12733 23891 12767
rect 25145 12733 25179 12767
rect 17877 12665 17911 12699
rect 19533 12665 19567 12699
rect 20453 12665 20487 12699
rect 21465 12665 21499 12699
rect 18889 12597 18923 12631
rect 19993 12597 20027 12631
rect 21741 12597 21775 12631
rect 22477 12597 22511 12631
rect 22937 12597 22971 12631
rect 25329 12597 25363 12631
rect 18521 12393 18555 12427
rect 19257 12393 19291 12427
rect 22293 12393 22327 12427
rect 24133 12393 24167 12427
rect 17417 12325 17451 12359
rect 17141 12257 17175 12291
rect 19625 12257 19659 12291
rect 21169 12257 21203 12291
rect 24041 12257 24075 12291
rect 25237 12257 25271 12291
rect 16129 12189 16163 12223
rect 19717 12189 19751 12223
rect 19809 12189 19843 12223
rect 20913 12189 20947 12223
rect 24225 12189 24259 12223
rect 19165 12121 19199 12155
rect 20269 12053 20303 12087
rect 22845 12053 22879 12087
rect 23489 12053 23523 12087
rect 23673 12053 23707 12087
rect 24685 12053 24719 12087
rect 25421 12053 25455 12087
rect 18981 11849 19015 11883
rect 20821 11849 20855 11883
rect 21373 11849 21407 11883
rect 23489 11849 23523 11883
rect 25697 11849 25731 11883
rect 18429 11713 18463 11747
rect 22477 11713 22511 11747
rect 22661 11713 22695 11747
rect 16405 11645 16439 11679
rect 19441 11645 19475 11679
rect 21925 11645 21959 11679
rect 22385 11645 22419 11679
rect 23673 11645 23707 11679
rect 16681 11577 16715 11611
rect 17233 11577 17267 11611
rect 19686 11577 19720 11611
rect 23918 11577 23952 11611
rect 17509 11509 17543 11543
rect 19349 11509 19383 11543
rect 22017 11509 22051 11543
rect 23121 11509 23155 11543
rect 25053 11509 25087 11543
rect 16681 11305 16715 11339
rect 19717 11305 19751 11339
rect 20269 11305 20303 11339
rect 22753 11305 22787 11339
rect 23765 11305 23799 11339
rect 17049 11237 17083 11271
rect 24124 11237 24158 11271
rect 13921 11169 13955 11203
rect 15301 11169 15335 11203
rect 18337 11169 18371 11203
rect 18593 11169 18627 11203
rect 20637 11169 20671 11203
rect 21281 11169 21315 11203
rect 21640 11169 21674 11203
rect 14197 11101 14231 11135
rect 15485 11101 15519 11135
rect 17141 11101 17175 11135
rect 17325 11101 17359 11135
rect 21373 11101 21407 11135
rect 23857 11101 23891 11135
rect 16589 11033 16623 11067
rect 25237 11033 25271 11067
rect 18153 10965 18187 10999
rect 23397 10965 23431 10999
rect 14197 10761 14231 10795
rect 16773 10761 16807 10795
rect 17141 10761 17175 10795
rect 17785 10761 17819 10795
rect 20085 10761 20119 10795
rect 20637 10761 20671 10795
rect 21465 10761 21499 10795
rect 21925 10761 21959 10795
rect 23489 10761 23523 10795
rect 21833 10625 21867 10659
rect 22477 10625 22511 10659
rect 14565 10557 14599 10591
rect 14749 10557 14783 10591
rect 18061 10557 18095 10591
rect 18317 10557 18351 10591
rect 20821 10557 20855 10591
rect 22293 10557 22327 10591
rect 23673 10557 23707 10591
rect 14994 10489 15028 10523
rect 23121 10489 23155 10523
rect 23918 10489 23952 10523
rect 13737 10421 13771 10455
rect 16129 10421 16163 10455
rect 17509 10421 17543 10455
rect 19441 10421 19475 10455
rect 21005 10421 21039 10455
rect 22385 10421 22419 10455
rect 25053 10421 25087 10455
rect 25605 10421 25639 10455
rect 25973 10421 26007 10455
rect 13645 10217 13679 10251
rect 15485 10217 15519 10251
rect 17509 10217 17543 10251
rect 18429 10217 18463 10251
rect 18613 10217 18647 10251
rect 20269 10217 20303 10251
rect 20913 10217 20947 10251
rect 21281 10217 21315 10251
rect 22385 10217 22419 10251
rect 22937 10217 22971 10251
rect 23397 10217 23431 10251
rect 24041 10217 24075 10251
rect 24501 10217 24535 10251
rect 16374 10149 16408 10183
rect 23305 10149 23339 10183
rect 14013 10081 14047 10115
rect 14105 10081 14139 10115
rect 18981 10081 19015 10115
rect 24869 10081 24903 10115
rect 24961 10081 24995 10115
rect 14197 10013 14231 10047
rect 16129 10013 16163 10047
rect 19073 10013 19107 10047
rect 19165 10013 19199 10047
rect 21373 10013 21407 10047
rect 21557 10013 21591 10047
rect 23581 10013 23615 10047
rect 25053 10013 25087 10047
rect 22661 9945 22695 9979
rect 24317 9945 24351 9979
rect 13093 9877 13127 9911
rect 13553 9877 13587 9911
rect 14841 9877 14875 9911
rect 15945 9877 15979 9911
rect 18153 9877 18187 9911
rect 20729 9877 20763 9911
rect 21925 9877 21959 9911
rect 13369 9673 13403 9707
rect 20913 9673 20947 9707
rect 23029 9673 23063 9707
rect 23397 9673 23431 9707
rect 25605 9673 25639 9707
rect 25973 9673 26007 9707
rect 17877 9605 17911 9639
rect 19901 9605 19935 9639
rect 21373 9605 21407 9639
rect 16681 9537 16715 9571
rect 17141 9537 17175 9571
rect 20545 9537 20579 9571
rect 22201 9537 22235 9571
rect 13461 9469 13495 9503
rect 13717 9469 13751 9503
rect 15945 9469 15979 9503
rect 16497 9469 16531 9503
rect 18521 9469 18555 9503
rect 21557 9469 21591 9503
rect 23673 9469 23707 9503
rect 23929 9469 23963 9503
rect 13001 9401 13035 9435
rect 16589 9401 16623 9435
rect 18788 9401 18822 9435
rect 22109 9401 22143 9435
rect 12449 9333 12483 9367
rect 14841 9333 14875 9367
rect 15669 9333 15703 9367
rect 16129 9333 16163 9367
rect 18337 9333 18371 9367
rect 21189 9333 21223 9367
rect 21649 9333 21683 9367
rect 22017 9333 22051 9367
rect 25053 9333 25087 9367
rect 10517 9129 10551 9163
rect 13461 9129 13495 9163
rect 14013 9129 14047 9163
rect 14381 9129 14415 9163
rect 15301 9129 15335 9163
rect 16681 9129 16715 9163
rect 18613 9129 18647 9163
rect 19257 9129 19291 9163
rect 20729 9129 20763 9163
rect 23029 9129 23063 9163
rect 24869 9129 24903 9163
rect 21180 9061 21214 9095
rect 10885 8993 10919 9027
rect 12337 8993 12371 9027
rect 15669 8993 15703 9027
rect 17489 8993 17523 9027
rect 20913 8993 20947 9027
rect 23756 8993 23790 9027
rect 10425 8925 10459 8959
rect 10977 8925 11011 8959
rect 11069 8925 11103 8959
rect 12081 8925 12115 8959
rect 15117 8925 15151 8959
rect 15761 8925 15795 8959
rect 15945 8925 15979 8959
rect 17233 8925 17267 8959
rect 19809 8925 19843 8959
rect 23489 8925 23523 8959
rect 20269 8857 20303 8891
rect 11529 8789 11563 8823
rect 16405 8789 16439 8823
rect 17049 8789 17083 8823
rect 19717 8789 19751 8823
rect 22293 8789 22327 8823
rect 23397 8789 23431 8823
rect 10793 8585 10827 8619
rect 13277 8585 13311 8619
rect 13461 8585 13495 8619
rect 16865 8585 16899 8619
rect 19165 8585 19199 8619
rect 21281 8585 21315 8619
rect 21833 8585 21867 8619
rect 23121 8585 23155 8619
rect 24777 8585 24811 8619
rect 9965 8517 9999 8551
rect 12081 8517 12115 8551
rect 14841 8517 14875 8551
rect 18061 8517 18095 8551
rect 22201 8517 22235 8551
rect 22661 8517 22695 8551
rect 23673 8517 23707 8551
rect 10609 8449 10643 8483
rect 11437 8449 11471 8483
rect 14013 8449 14047 8483
rect 14565 8449 14599 8483
rect 18705 8449 18739 8483
rect 19533 8449 19567 8483
rect 24317 8449 24351 8483
rect 25421 8449 25455 8483
rect 11161 8381 11195 8415
rect 13829 8381 13863 8415
rect 13921 8381 13955 8415
rect 15209 8381 15243 8415
rect 15485 8381 15519 8415
rect 15752 8381 15786 8415
rect 17509 8381 17543 8415
rect 19809 8381 19843 8415
rect 19901 8381 19935 8415
rect 22477 8381 22511 8415
rect 23489 8381 23523 8415
rect 24041 8381 24075 8415
rect 25237 8381 25271 8415
rect 25973 8381 26007 8415
rect 10333 8313 10367 8347
rect 11253 8313 11287 8347
rect 12449 8313 12483 8347
rect 13001 8313 13035 8347
rect 17877 8313 17911 8347
rect 20146 8313 20180 8347
rect 15025 8245 15059 8279
rect 18429 8245 18463 8279
rect 18521 8245 18555 8279
rect 19625 8245 19659 8279
rect 24133 8245 24167 8279
rect 25145 8245 25179 8279
rect 9781 8041 9815 8075
rect 12173 8041 12207 8075
rect 13277 8041 13311 8075
rect 16681 8041 16715 8075
rect 17233 8041 17267 8075
rect 19165 8041 19199 8075
rect 21097 8041 21131 8075
rect 23029 8041 23063 8075
rect 23121 8041 23155 8075
rect 24133 8041 24167 8075
rect 10609 7973 10643 8007
rect 11060 7973 11094 8007
rect 13645 7973 13679 8007
rect 18521 7973 18555 8007
rect 20361 7973 20395 8007
rect 21557 7973 21591 8007
rect 23765 7973 23799 8007
rect 24685 7973 24719 8007
rect 15117 7905 15151 7939
rect 15568 7905 15602 7939
rect 18429 7905 18463 7939
rect 19717 7905 19751 7939
rect 21465 7905 21499 7939
rect 24593 7905 24627 7939
rect 10793 7837 10827 7871
rect 13737 7837 13771 7871
rect 13829 7837 13863 7871
rect 15301 7837 15335 7871
rect 18613 7837 18647 7871
rect 21741 7837 21775 7871
rect 23213 7837 23247 7871
rect 24777 7837 24811 7871
rect 12817 7769 12851 7803
rect 22569 7769 22603 7803
rect 13185 7701 13219 7735
rect 14749 7701 14783 7735
rect 14933 7701 14967 7735
rect 17601 7701 17635 7735
rect 18061 7701 18095 7735
rect 19441 7701 19475 7735
rect 19901 7701 19935 7735
rect 20729 7701 20763 7735
rect 22109 7701 22143 7735
rect 22661 7701 22695 7735
rect 24225 7701 24259 7735
rect 25237 7701 25271 7735
rect 11253 7497 11287 7531
rect 13093 7497 13127 7531
rect 15761 7497 15795 7531
rect 21373 7497 21407 7531
rect 22661 7497 22695 7531
rect 23029 7497 23063 7531
rect 23673 7497 23707 7531
rect 24685 7497 24719 7531
rect 20913 7429 20947 7463
rect 23489 7429 23523 7463
rect 13277 7361 13311 7395
rect 16405 7361 16439 7395
rect 16773 7361 16807 7395
rect 21281 7361 21315 7395
rect 21925 7361 21959 7395
rect 24133 7361 24167 7395
rect 24225 7361 24259 7395
rect 26341 7361 26375 7395
rect 9873 7293 9907 7327
rect 13544 7293 13578 7327
rect 15301 7293 15335 7327
rect 18889 7293 18923 7327
rect 21741 7293 21775 7327
rect 24041 7293 24075 7327
rect 25237 7293 25271 7327
rect 25973 7293 26007 7327
rect 9781 7225 9815 7259
rect 10118 7225 10152 7259
rect 12817 7225 12851 7259
rect 16129 7225 16163 7259
rect 18337 7225 18371 7259
rect 19156 7225 19190 7259
rect 21833 7225 21867 7259
rect 25513 7225 25547 7259
rect 9321 7157 9355 7191
rect 14657 7157 14691 7191
rect 15577 7157 15611 7191
rect 16221 7157 16255 7191
rect 17325 7157 17359 7191
rect 17785 7157 17819 7191
rect 18613 7157 18647 7191
rect 20269 7157 20303 7191
rect 25053 7157 25087 7191
rect 13185 6953 13219 6987
rect 13737 6953 13771 6987
rect 15577 6953 15611 6987
rect 19165 6953 19199 6987
rect 22937 6953 22971 6987
rect 23489 6953 23523 6987
rect 24961 6953 24995 6987
rect 14933 6885 14967 6919
rect 17601 6885 17635 6919
rect 19625 6885 19659 6919
rect 23848 6885 23882 6919
rect 8585 6817 8619 6851
rect 10057 6817 10091 6851
rect 10885 6817 10919 6851
rect 12061 6817 12095 6851
rect 16037 6817 16071 6851
rect 17141 6817 17175 6851
rect 17693 6817 17727 6851
rect 21169 6817 21203 6851
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 11805 6749 11839 6783
rect 16129 6749 16163 6783
rect 16313 6749 16347 6783
rect 17785 6749 17819 6783
rect 19717 6749 19751 6783
rect 19809 6749 19843 6783
rect 20913 6749 20947 6783
rect 23581 6749 23615 6783
rect 9689 6681 9723 6715
rect 15669 6681 15703 6715
rect 17233 6681 17267 6715
rect 19257 6681 19291 6715
rect 9045 6613 9079 6647
rect 11161 6613 11195 6647
rect 14105 6613 14139 6647
rect 14657 6613 14691 6647
rect 18337 6613 18371 6647
rect 18797 6613 18831 6647
rect 20361 6613 20395 6647
rect 20637 6613 20671 6647
rect 22293 6613 22327 6647
rect 8953 6409 8987 6443
rect 10425 6409 10459 6443
rect 11529 6409 11563 6443
rect 11897 6409 11931 6443
rect 12449 6409 12483 6443
rect 15209 6409 15243 6443
rect 16681 6409 16715 6443
rect 18889 6409 18923 6443
rect 19349 6409 19383 6443
rect 23121 6409 23155 6443
rect 25053 6409 25087 6443
rect 15117 6341 15151 6375
rect 13001 6273 13035 6307
rect 15761 6273 15795 6307
rect 19809 6273 19843 6307
rect 19901 6273 19935 6307
rect 20913 6273 20947 6307
rect 23673 6273 23707 6307
rect 9045 6205 9079 6239
rect 16221 6205 16255 6239
rect 16865 6205 16899 6239
rect 18245 6205 18279 6239
rect 19717 6205 19751 6239
rect 21005 6205 21039 6239
rect 21272 6205 21306 6239
rect 9290 6137 9324 6171
rect 12817 6137 12851 6171
rect 15577 6137 15611 6171
rect 23489 6137 23523 6171
rect 23940 6137 23974 6171
rect 11069 6069 11103 6103
rect 12265 6069 12299 6103
rect 12909 6069 12943 6103
rect 13461 6069 13495 6103
rect 14197 6069 14231 6103
rect 14657 6069 14691 6103
rect 15669 6069 15703 6103
rect 17049 6069 17083 6103
rect 17509 6069 17543 6103
rect 17785 6069 17819 6103
rect 18429 6069 18463 6103
rect 19257 6069 19291 6103
rect 20453 6069 20487 6103
rect 22385 6069 22419 6103
rect 25605 6069 25639 6103
rect 8585 5865 8619 5899
rect 9137 5865 9171 5899
rect 9873 5865 9907 5899
rect 10241 5865 10275 5899
rect 11897 5865 11931 5899
rect 13001 5865 13035 5899
rect 18797 5865 18831 5899
rect 19165 5865 19199 5899
rect 20361 5865 20395 5899
rect 20637 5865 20671 5899
rect 20913 5865 20947 5899
rect 21281 5865 21315 5899
rect 23673 5865 23707 5899
rect 24041 5865 24075 5899
rect 12541 5797 12575 5831
rect 17040 5797 17074 5831
rect 23581 5797 23615 5831
rect 10517 5729 10551 5763
rect 10784 5729 10818 5763
rect 13369 5729 13403 5763
rect 15669 5729 15703 5763
rect 19625 5729 19659 5763
rect 19717 5729 19751 5763
rect 22569 5729 22603 5763
rect 25237 5729 25271 5763
rect 13461 5661 13495 5695
rect 13553 5661 13587 5695
rect 15577 5661 15611 5695
rect 16589 5661 16623 5695
rect 16773 5661 16807 5695
rect 19809 5661 19843 5695
rect 21373 5661 21407 5695
rect 21465 5661 21499 5695
rect 23213 5661 23247 5695
rect 24133 5661 24167 5695
rect 24225 5661 24259 5695
rect 12909 5593 12943 5627
rect 15117 5593 15151 5627
rect 19257 5593 19291 5627
rect 22753 5593 22787 5627
rect 24685 5593 24719 5627
rect 25053 5593 25087 5627
rect 15853 5525 15887 5559
rect 18153 5525 18187 5559
rect 22109 5525 22143 5559
rect 22477 5525 22511 5559
rect 25421 5525 25455 5559
rect 10701 5321 10735 5355
rect 12265 5321 12299 5355
rect 17141 5321 17175 5355
rect 18889 5321 18923 5355
rect 19349 5321 19383 5355
rect 21465 5321 21499 5355
rect 21649 5321 21683 5355
rect 22017 5321 22051 5355
rect 23121 5321 23155 5355
rect 23489 5321 23523 5355
rect 25605 5321 25639 5355
rect 17417 5253 17451 5287
rect 21097 5253 21131 5287
rect 11345 5185 11379 5219
rect 11897 5185 11931 5219
rect 19901 5185 19935 5219
rect 8217 5117 8251 5151
rect 8677 5117 8711 5151
rect 12633 5117 12667 5151
rect 12900 5117 12934 5151
rect 15117 5117 15151 5151
rect 18245 5117 18279 5151
rect 20913 5117 20947 5151
rect 22661 5185 22695 5219
rect 21833 5117 21867 5151
rect 22385 5117 22419 5151
rect 22477 5117 22511 5151
rect 23673 5117 23707 5151
rect 8585 5049 8619 5083
rect 8944 5049 8978 5083
rect 14657 5049 14691 5083
rect 15362 5049 15396 5083
rect 19717 5049 19751 5083
rect 20453 5049 20487 5083
rect 21649 5049 21683 5083
rect 23940 5049 23974 5083
rect 10057 4981 10091 5015
rect 10977 4981 11011 5015
rect 14013 4981 14047 5015
rect 15025 4981 15059 5015
rect 16497 4981 16531 5015
rect 17785 4981 17819 5015
rect 18429 4981 18463 5015
rect 19165 4981 19199 5015
rect 19809 4981 19843 5015
rect 20821 4981 20855 5015
rect 25053 4981 25087 5015
rect 25973 4981 26007 5015
rect 9413 4777 9447 4811
rect 9689 4777 9723 4811
rect 11621 4777 11655 4811
rect 12449 4777 12483 4811
rect 14013 4777 14047 4811
rect 16681 4777 16715 4811
rect 17785 4777 17819 4811
rect 19073 4777 19107 4811
rect 20729 4777 20763 4811
rect 23397 4777 23431 4811
rect 23949 4777 23983 4811
rect 24317 4777 24351 4811
rect 24501 4777 24535 4811
rect 24961 4777 24995 4811
rect 12173 4709 12207 4743
rect 12900 4709 12934 4743
rect 17693 4709 17727 4743
rect 22262 4709 22296 4743
rect 24869 4709 24903 4743
rect 10057 4641 10091 4675
rect 15568 4641 15602 4675
rect 18153 4641 18187 4675
rect 19717 4641 19751 4675
rect 20913 4641 20947 4675
rect 22017 4641 22051 4675
rect 8585 4573 8619 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 11437 4573 11471 4607
rect 12633 4573 12667 4607
rect 14657 4573 14691 4607
rect 15117 4573 15151 4607
rect 15301 4573 15335 4607
rect 18245 4573 18279 4607
rect 18429 4573 18463 4607
rect 19441 4573 19475 4607
rect 25145 4573 25179 4607
rect 21097 4505 21131 4539
rect 8217 4437 8251 4471
rect 9045 4437 9079 4471
rect 10701 4437 10735 4471
rect 17325 4437 17359 4471
rect 19901 4437 19935 4471
rect 20269 4437 20303 4471
rect 21833 4437 21867 4471
rect 25605 4437 25639 4471
rect 11069 4233 11103 4267
rect 15945 4233 15979 4267
rect 17141 4233 17175 4267
rect 19533 4233 19567 4267
rect 21005 4233 21039 4267
rect 23121 4233 23155 4267
rect 25881 4233 25915 4267
rect 8769 4097 8803 4131
rect 9505 4097 9539 4131
rect 12173 4097 12207 4131
rect 13093 4097 13127 4131
rect 14933 4097 14967 4131
rect 15485 4097 15519 4131
rect 16497 4097 16531 4131
rect 17417 4097 17451 4131
rect 18521 4097 18555 4131
rect 18613 4097 18647 4131
rect 20085 4097 20119 4131
rect 20269 4097 20303 4131
rect 22385 4097 22419 4131
rect 22753 4097 22787 4131
rect 8033 4029 8067 4063
rect 8493 4029 8527 4063
rect 9689 4029 9723 4063
rect 12909 4029 12943 4063
rect 13921 4029 13955 4063
rect 14841 4029 14875 4063
rect 16405 4029 16439 4063
rect 19993 4029 20027 4063
rect 23949 4029 23983 4063
rect 24216 4029 24250 4063
rect 9934 3961 9968 3995
rect 11897 3961 11931 3995
rect 13001 3961 13035 3995
rect 14749 3961 14783 3995
rect 16313 3961 16347 3995
rect 19165 3961 19199 3995
rect 22201 3961 22235 3995
rect 7665 3893 7699 3927
rect 8125 3893 8159 3927
rect 8585 3893 8619 3927
rect 9229 3893 9263 3927
rect 12541 3893 12575 3927
rect 14197 3893 14231 3927
rect 14381 3893 14415 3927
rect 15761 3893 15795 3927
rect 17785 3893 17819 3927
rect 18061 3893 18095 3927
rect 18429 3893 18463 3927
rect 19625 3893 19659 3927
rect 21557 3893 21591 3927
rect 21741 3893 21775 3927
rect 22109 3893 22143 3927
rect 25329 3893 25363 3927
rect 26249 3893 26283 3927
rect 7021 3689 7055 3723
rect 8033 3689 8067 3723
rect 9965 3689 9999 3723
rect 10977 3689 11011 3723
rect 13921 3689 13955 3723
rect 15117 3689 15151 3723
rect 15945 3689 15979 3723
rect 20177 3689 20211 3723
rect 21097 3689 21131 3723
rect 22937 3689 22971 3723
rect 24041 3689 24075 3723
rect 24501 3689 24535 3723
rect 25053 3689 25087 3723
rect 25789 3689 25823 3723
rect 7573 3621 7607 3655
rect 11774 3621 11808 3655
rect 13461 3621 13495 3655
rect 19533 3621 19567 3655
rect 20545 3621 20579 3655
rect 23673 3621 23707 3655
rect 25421 3621 25455 3655
rect 8401 3553 8435 3587
rect 10333 3553 10367 3587
rect 14013 3553 14047 3587
rect 15301 3553 15335 3587
rect 16753 3553 16787 3587
rect 19073 3553 19107 3587
rect 19625 3553 19659 3587
rect 21557 3553 21591 3587
rect 21824 3553 21858 3587
rect 24409 3553 24443 3587
rect 8493 3485 8527 3519
rect 8677 3485 8711 3519
rect 9137 3485 9171 3519
rect 10425 3485 10459 3519
rect 10609 3485 10643 3519
rect 11529 3485 11563 3519
rect 16497 3485 16531 3519
rect 19809 3485 19843 3519
rect 24685 3485 24719 3519
rect 14657 3417 14691 3451
rect 19165 3417 19199 3451
rect 7941 3349 7975 3383
rect 9505 3349 9539 3383
rect 11437 3349 11471 3383
rect 12909 3349 12943 3383
rect 14197 3349 14231 3383
rect 15485 3349 15519 3383
rect 16313 3349 16347 3383
rect 17877 3349 17911 3383
rect 18429 3349 18463 3383
rect 7481 3145 7515 3179
rect 7849 3145 7883 3179
rect 9045 3145 9079 3179
rect 10885 3145 10919 3179
rect 11529 3145 11563 3179
rect 12633 3145 12667 3179
rect 13737 3145 13771 3179
rect 16129 3145 16163 3179
rect 20085 3145 20119 3179
rect 21925 3145 21959 3179
rect 22477 3145 22511 3179
rect 23305 3145 23339 3179
rect 23673 3145 23707 3179
rect 24685 3145 24719 3179
rect 25145 3145 25179 3179
rect 26157 3145 26191 3179
rect 7941 3077 7975 3111
rect 19441 3077 19475 3111
rect 8585 3009 8619 3043
rect 9505 3009 9539 3043
rect 13093 3009 13127 3043
rect 13277 3009 13311 3043
rect 17785 3009 17819 3043
rect 19809 3009 19843 3043
rect 23121 3009 23155 3043
rect 6929 2941 6963 2975
rect 9321 2941 9355 2975
rect 9772 2941 9806 2975
rect 12173 2941 12207 2975
rect 14197 2941 14231 2975
rect 16589 2941 16623 2975
rect 16681 2941 16715 2975
rect 17233 2941 17267 2975
rect 18061 2941 18095 2975
rect 18317 2941 18351 2975
rect 25881 3077 25915 3111
rect 24225 3009 24259 3043
rect 20545 2941 20579 2975
rect 23305 2941 23339 2975
rect 24041 2941 24075 2975
rect 8401 2873 8435 2907
rect 11897 2873 11931 2907
rect 13001 2873 13035 2907
rect 14105 2873 14139 2907
rect 14442 2873 14476 2907
rect 19809 2873 19843 2907
rect 20453 2873 20487 2907
rect 20812 2873 20846 2907
rect 23489 2873 23523 2907
rect 24133 2873 24167 2907
rect 6653 2805 6687 2839
rect 8309 2805 8343 2839
rect 15577 2805 15611 2839
rect 16865 2805 16899 2839
rect 25421 2805 25455 2839
rect 7113 2601 7147 2635
rect 8125 2601 8159 2635
rect 9597 2601 9631 2635
rect 10517 2601 10551 2635
rect 10977 2601 11011 2635
rect 11437 2601 11471 2635
rect 12081 2601 12115 2635
rect 15301 2601 15335 2635
rect 16865 2601 16899 2635
rect 19717 2601 19751 2635
rect 21189 2601 21223 2635
rect 21649 2601 21683 2635
rect 22293 2601 22327 2635
rect 22661 2601 22695 2635
rect 23857 2601 23891 2635
rect 24409 2601 24443 2635
rect 25145 2601 25179 2635
rect 12449 2533 12483 2567
rect 12900 2533 12934 2567
rect 15730 2533 15764 2567
rect 17417 2533 17451 2567
rect 21005 2533 21039 2567
rect 23489 2533 23523 2567
rect 24501 2533 24535 2567
rect 7665 2465 7699 2499
rect 8493 2465 8527 2499
rect 9873 2465 9907 2499
rect 11345 2465 11379 2499
rect 12633 2465 12667 2499
rect 14565 2465 14599 2499
rect 15485 2465 15519 2499
rect 18593 2465 18627 2499
rect 20637 2465 20671 2499
rect 21557 2465 21591 2499
rect 22845 2465 22879 2499
rect 25605 2465 25639 2499
rect 8033 2397 8067 2431
rect 8585 2397 8619 2431
rect 8769 2397 8803 2431
rect 11621 2397 11655 2431
rect 18061 2397 18095 2431
rect 18337 2397 18371 2431
rect 21833 2397 21867 2431
rect 24593 2397 24627 2431
rect 25421 2397 25455 2431
rect 6745 2329 6779 2363
rect 9229 2329 9263 2363
rect 24041 2329 24075 2363
rect 10057 2261 10091 2295
rect 10793 2261 10827 2295
rect 14013 2261 14047 2295
rect 23029 2261 23063 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 12986 24828 12992 24880
rect 13044 24868 13050 24880
rect 24762 24868 24768 24880
rect 13044 24840 24768 24868
rect 13044 24828 13050 24840
rect 24762 24828 24768 24840
rect 24820 24828 24826 24880
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 23477 24395 23535 24401
rect 23477 24361 23489 24395
rect 23523 24392 23535 24395
rect 24210 24392 24216 24404
rect 23523 24364 24216 24392
rect 23523 24361 23535 24364
rect 23477 24355 23535 24361
rect 24210 24352 24216 24364
rect 24268 24352 24274 24404
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 10134 23808 10140 23860
rect 10192 23848 10198 23860
rect 10229 23851 10287 23857
rect 10229 23848 10241 23851
rect 10192 23820 10241 23848
rect 10192 23808 10198 23820
rect 10229 23817 10241 23820
rect 10275 23817 10287 23851
rect 12986 23848 12992 23860
rect 12947 23820 12992 23848
rect 10229 23811 10287 23817
rect 12986 23808 12992 23820
rect 13044 23808 13050 23860
rect 17494 23808 17500 23860
rect 17552 23848 17558 23860
rect 17773 23851 17831 23857
rect 17773 23848 17785 23851
rect 17552 23820 17785 23848
rect 17552 23808 17558 23820
rect 17773 23817 17785 23820
rect 17819 23817 17831 23851
rect 17773 23811 17831 23817
rect 10045 23647 10103 23653
rect 10045 23613 10057 23647
rect 10091 23644 10103 23647
rect 10091 23616 10732 23644
rect 10091 23613 10103 23616
rect 10045 23607 10103 23613
rect 10704 23520 10732 23616
rect 12342 23604 12348 23656
rect 12400 23644 12406 23656
rect 12805 23647 12863 23653
rect 12805 23644 12817 23647
rect 12400 23616 12817 23644
rect 12400 23604 12406 23616
rect 12805 23613 12817 23616
rect 12851 23644 12863 23647
rect 13357 23647 13415 23653
rect 13357 23644 13369 23647
rect 12851 23616 13369 23644
rect 12851 23613 12863 23616
rect 12805 23607 12863 23613
rect 13357 23613 13369 23616
rect 13403 23613 13415 23647
rect 13357 23607 13415 23613
rect 17788 23576 17816 23811
rect 24670 23808 24676 23860
rect 24728 23848 24734 23860
rect 24765 23851 24823 23857
rect 24765 23848 24777 23851
rect 24728 23820 24777 23848
rect 24728 23808 24734 23820
rect 24765 23817 24777 23820
rect 24811 23817 24823 23851
rect 24765 23811 24823 23817
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23644 18107 23647
rect 18138 23644 18144 23656
rect 18095 23616 18144 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 18138 23604 18144 23616
rect 18196 23604 18202 23656
rect 23934 23604 23940 23656
rect 23992 23644 23998 23656
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 23992 23616 24593 23644
rect 23992 23604 23998 23616
rect 24581 23613 24593 23616
rect 24627 23644 24639 23647
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 24627 23616 25145 23644
rect 24627 23613 24639 23616
rect 24581 23607 24639 23613
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 18294 23579 18352 23585
rect 18294 23576 18306 23579
rect 17788 23548 18306 23576
rect 18294 23545 18306 23548
rect 18340 23545 18352 23579
rect 18294 23539 18352 23545
rect 3510 23468 3516 23520
rect 3568 23508 3574 23520
rect 4062 23508 4068 23520
rect 3568 23480 4068 23508
rect 3568 23468 3574 23480
rect 4062 23468 4068 23480
rect 4120 23468 4126 23520
rect 10686 23508 10692 23520
rect 10647 23480 10692 23508
rect 10686 23468 10692 23480
rect 10744 23468 10750 23520
rect 19426 23508 19432 23520
rect 19387 23480 19432 23508
rect 19426 23468 19432 23480
rect 19484 23468 19490 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 24854 23264 24860 23316
rect 24912 23304 24918 23316
rect 25133 23307 25191 23313
rect 25133 23304 25145 23307
rect 24912 23276 25145 23304
rect 24912 23264 24918 23276
rect 25133 23273 25145 23276
rect 25179 23273 25191 23307
rect 25133 23267 25191 23273
rect 12069 23239 12127 23245
rect 12069 23205 12081 23239
rect 12115 23236 12127 23239
rect 12342 23236 12348 23248
rect 12115 23208 12348 23236
rect 12115 23205 12127 23208
rect 12069 23199 12127 23205
rect 12342 23196 12348 23208
rect 12400 23196 12406 23248
rect 23934 23236 23940 23248
rect 23895 23208 23940 23236
rect 23934 23196 23940 23208
rect 23992 23196 23998 23248
rect 11790 23168 11796 23180
rect 11751 23140 11796 23168
rect 11790 23128 11796 23140
rect 11848 23128 11854 23180
rect 23661 23171 23719 23177
rect 23661 23137 23673 23171
rect 23707 23168 23719 23171
rect 23842 23168 23848 23180
rect 23707 23140 23848 23168
rect 23707 23137 23719 23140
rect 23661 23131 23719 23137
rect 23842 23128 23848 23140
rect 23900 23128 23906 23180
rect 24946 23168 24952 23180
rect 24907 23140 24952 23168
rect 24946 23128 24952 23140
rect 25004 23128 25010 23180
rect 18141 22967 18199 22973
rect 18141 22933 18153 22967
rect 18187 22964 18199 22967
rect 18230 22964 18236 22976
rect 18187 22936 18236 22964
rect 18187 22933 18199 22936
rect 18141 22927 18199 22933
rect 18230 22924 18236 22936
rect 18288 22924 18294 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 24210 22720 24216 22772
rect 24268 22760 24274 22772
rect 24765 22763 24823 22769
rect 24765 22760 24777 22763
rect 24268 22732 24777 22760
rect 24268 22720 24274 22732
rect 24765 22729 24777 22732
rect 24811 22729 24823 22763
rect 24765 22723 24823 22729
rect 24026 22584 24032 22636
rect 24084 22624 24090 22636
rect 24210 22624 24216 22636
rect 24084 22596 24216 22624
rect 24084 22584 24090 22596
rect 24210 22584 24216 22596
rect 24268 22584 24274 22636
rect 24578 22556 24584 22568
rect 24539 22528 24584 22556
rect 24578 22516 24584 22528
rect 24636 22556 24642 22568
rect 25133 22559 25191 22565
rect 25133 22556 25145 22559
rect 24636 22528 25145 22556
rect 24636 22516 24642 22528
rect 25133 22525 25145 22528
rect 25179 22525 25191 22559
rect 25133 22519 25191 22525
rect 24946 22448 24952 22500
rect 25004 22488 25010 22500
rect 25501 22491 25559 22497
rect 25501 22488 25513 22491
rect 25004 22460 25513 22488
rect 25004 22448 25010 22460
rect 25501 22457 25513 22460
rect 25547 22457 25559 22491
rect 25501 22451 25559 22457
rect 11790 22420 11796 22432
rect 11751 22392 11796 22420
rect 11790 22380 11796 22392
rect 11848 22380 11854 22432
rect 23842 22420 23848 22432
rect 23803 22392 23848 22420
rect 23842 22380 23848 22392
rect 23900 22380 23906 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 10042 22080 10048 22092
rect 10003 22052 10048 22080
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 17034 22080 17040 22092
rect 16995 22052 17040 22080
rect 17034 22040 17040 22052
rect 17092 22040 17098 22092
rect 10318 22012 10324 22024
rect 10279 21984 10324 22012
rect 10318 21972 10324 21984
rect 10376 21972 10382 22024
rect 17218 21944 17224 21956
rect 17179 21916 17224 21944
rect 17218 21904 17224 21916
rect 17276 21904 17282 21956
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 17034 21672 17040 21684
rect 16995 21644 17040 21672
rect 17034 21632 17040 21644
rect 17092 21632 17098 21684
rect 24670 21632 24676 21684
rect 24728 21672 24734 21684
rect 24765 21675 24823 21681
rect 24765 21672 24777 21675
rect 24728 21644 24777 21672
rect 24728 21632 24734 21644
rect 24765 21641 24777 21644
rect 24811 21641 24823 21675
rect 24765 21635 24823 21641
rect 13722 21536 13728 21548
rect 13683 21508 13728 21536
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 12986 21428 12992 21480
rect 13044 21468 13050 21480
rect 13449 21471 13507 21477
rect 13449 21468 13461 21471
rect 13044 21440 13461 21468
rect 13044 21428 13050 21440
rect 13449 21437 13461 21440
rect 13495 21468 13507 21471
rect 14185 21471 14243 21477
rect 14185 21468 14197 21471
rect 13495 21440 14197 21468
rect 13495 21437 13507 21440
rect 13449 21431 13507 21437
rect 14185 21437 14197 21440
rect 14231 21437 14243 21471
rect 14185 21431 14243 21437
rect 23934 21428 23940 21480
rect 23992 21468 23998 21480
rect 24581 21471 24639 21477
rect 24581 21468 24593 21471
rect 23992 21440 24593 21468
rect 23992 21428 23998 21440
rect 24581 21437 24593 21440
rect 24627 21468 24639 21471
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24627 21440 25145 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 9674 21292 9680 21344
rect 9732 21332 9738 21344
rect 10042 21332 10048 21344
rect 9732 21304 10048 21332
rect 9732 21292 9738 21304
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 16206 21292 16212 21344
rect 16264 21332 16270 21344
rect 17034 21332 17040 21344
rect 16264 21304 17040 21332
rect 16264 21292 16270 21304
rect 17034 21292 17040 21304
rect 17092 21292 17098 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 24762 21128 24768 21140
rect 24723 21100 24768 21128
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 16206 21060 16212 21072
rect 16167 21032 16212 21060
rect 16206 21020 16212 21032
rect 16264 21020 16270 21072
rect 15838 20952 15844 21004
rect 15896 20992 15902 21004
rect 15933 20995 15991 21001
rect 15933 20992 15945 20995
rect 15896 20964 15945 20992
rect 15896 20952 15902 20964
rect 15933 20961 15945 20964
rect 15979 20961 15991 20995
rect 15933 20955 15991 20961
rect 24581 20995 24639 21001
rect 24581 20961 24593 20995
rect 24627 20992 24639 20995
rect 24670 20992 24676 21004
rect 24627 20964 24676 20992
rect 24627 20961 24639 20964
rect 24581 20955 24639 20961
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 25130 20584 25136 20596
rect 25091 20556 25136 20584
rect 25130 20544 25136 20556
rect 25188 20544 25194 20596
rect 23934 20448 23940 20460
rect 23895 20420 23940 20448
rect 23934 20408 23940 20420
rect 23992 20408 23998 20460
rect 23661 20383 23719 20389
rect 23661 20380 23673 20383
rect 23492 20352 23673 20380
rect 23492 20256 23520 20352
rect 23661 20349 23673 20352
rect 23707 20349 23719 20383
rect 23661 20343 23719 20349
rect 24854 20340 24860 20392
rect 24912 20380 24918 20392
rect 24949 20383 25007 20389
rect 24949 20380 24961 20383
rect 24912 20352 24961 20380
rect 24912 20340 24918 20352
rect 24949 20349 24961 20352
rect 24995 20380 25007 20383
rect 25501 20383 25559 20389
rect 25501 20380 25513 20383
rect 24995 20352 25513 20380
rect 24995 20349 25007 20352
rect 24949 20343 25007 20349
rect 25501 20349 25513 20352
rect 25547 20349 25559 20383
rect 25501 20343 25559 20349
rect 15838 20204 15844 20256
rect 15896 20244 15902 20256
rect 15933 20247 15991 20253
rect 15933 20244 15945 20247
rect 15896 20216 15945 20244
rect 15896 20204 15902 20216
rect 15933 20213 15945 20216
rect 15979 20213 15991 20247
rect 23474 20244 23480 20256
rect 23435 20216 23480 20244
rect 15933 20207 15991 20213
rect 23474 20204 23480 20216
rect 23532 20204 23538 20256
rect 24578 20244 24584 20256
rect 24539 20216 24584 20244
rect 24578 20204 24584 20216
rect 24636 20204 24642 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 24026 20000 24032 20052
rect 24084 20040 24090 20052
rect 24765 20043 24823 20049
rect 24765 20040 24777 20043
rect 24084 20012 24777 20040
rect 24084 20000 24090 20012
rect 24765 20009 24777 20012
rect 24811 20009 24823 20043
rect 24765 20003 24823 20009
rect 21450 19972 21456 19984
rect 21411 19944 21456 19972
rect 21450 19932 21456 19944
rect 21508 19932 21514 19984
rect 20898 19864 20904 19916
rect 20956 19904 20962 19916
rect 21177 19907 21235 19913
rect 21177 19904 21189 19907
rect 20956 19876 21189 19904
rect 20956 19864 20962 19876
rect 21177 19873 21189 19876
rect 21223 19873 21235 19907
rect 21177 19867 21235 19873
rect 24026 19864 24032 19916
rect 24084 19904 24090 19916
rect 24581 19907 24639 19913
rect 24581 19904 24593 19907
rect 24084 19876 24593 19904
rect 24084 19864 24090 19876
rect 24581 19873 24593 19876
rect 24627 19873 24639 19907
rect 24581 19867 24639 19873
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 24854 19360 24860 19372
rect 24780 19332 24860 19360
rect 23661 19295 23719 19301
rect 23661 19292 23673 19295
rect 23492 19264 23673 19292
rect 23492 19168 23520 19264
rect 23661 19261 23673 19264
rect 23707 19261 23719 19295
rect 23661 19255 23719 19261
rect 23937 19295 23995 19301
rect 23937 19261 23949 19295
rect 23983 19292 23995 19295
rect 24780 19292 24808 19332
rect 24854 19320 24860 19332
rect 24912 19320 24918 19372
rect 24946 19292 24952 19304
rect 23983 19264 24808 19292
rect 24907 19264 24952 19292
rect 23983 19261 23995 19264
rect 23937 19255 23995 19261
rect 24946 19252 24952 19264
rect 25004 19292 25010 19304
rect 25501 19295 25559 19301
rect 25501 19292 25513 19295
rect 25004 19264 25513 19292
rect 25004 19252 25010 19264
rect 25501 19261 25513 19264
rect 25547 19261 25559 19295
rect 25501 19255 25559 19261
rect 20898 19116 20904 19168
rect 20956 19156 20962 19168
rect 21177 19159 21235 19165
rect 21177 19156 21189 19159
rect 20956 19128 21189 19156
rect 20956 19116 20962 19128
rect 21177 19125 21189 19128
rect 21223 19125 21235 19159
rect 23474 19156 23480 19168
rect 23435 19128 23480 19156
rect 21177 19119 21235 19125
rect 23474 19116 23480 19128
rect 23532 19116 23538 19168
rect 24578 19156 24584 19168
rect 24539 19128 24584 19156
rect 24578 19116 24584 19128
rect 24636 19116 24642 19168
rect 24854 19116 24860 19168
rect 24912 19156 24918 19168
rect 25133 19159 25191 19165
rect 25133 19156 25145 19159
rect 24912 19128 25145 19156
rect 24912 19116 24918 19128
rect 25133 19125 25145 19128
rect 25179 19125 25191 19159
rect 25133 19119 25191 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11149 18819 11207 18825
rect 11149 18816 11161 18819
rect 11112 18788 11161 18816
rect 11112 18776 11118 18788
rect 11149 18785 11161 18788
rect 11195 18785 11207 18819
rect 16022 18816 16028 18828
rect 15983 18788 16028 18816
rect 11149 18779 11207 18785
rect 16022 18776 16028 18788
rect 16080 18776 16086 18828
rect 16298 18816 16304 18828
rect 16259 18788 16304 18816
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 11330 18680 11336 18692
rect 11291 18652 11336 18680
rect 11330 18640 11336 18652
rect 11388 18640 11394 18692
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 13173 18207 13231 18213
rect 13173 18173 13185 18207
rect 13219 18204 13231 18207
rect 13262 18204 13268 18216
rect 13219 18176 13268 18204
rect 13219 18173 13231 18176
rect 13173 18167 13231 18173
rect 13262 18164 13268 18176
rect 13320 18204 13326 18216
rect 13909 18207 13967 18213
rect 13909 18204 13921 18207
rect 13320 18176 13921 18204
rect 13320 18164 13326 18176
rect 13909 18173 13921 18176
rect 13955 18173 13967 18207
rect 13909 18167 13967 18173
rect 13446 18136 13452 18148
rect 13407 18108 13452 18136
rect 13446 18096 13452 18108
rect 13504 18096 13510 18148
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11149 18071 11207 18077
rect 11149 18068 11161 18071
rect 11112 18040 11161 18068
rect 11112 18028 11118 18040
rect 11149 18037 11161 18040
rect 11195 18037 11207 18071
rect 11149 18031 11207 18037
rect 15286 18028 15292 18080
rect 15344 18068 15350 18080
rect 16022 18068 16028 18080
rect 15344 18040 16028 18068
rect 15344 18028 15350 18040
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 24670 17824 24676 17876
rect 24728 17864 24734 17876
rect 24765 17867 24823 17873
rect 24765 17864 24777 17867
rect 24728 17836 24777 17864
rect 24728 17824 24734 17836
rect 24765 17833 24777 17836
rect 24811 17833 24823 17867
rect 24765 17827 24823 17833
rect 10505 17799 10563 17805
rect 10505 17765 10517 17799
rect 10551 17796 10563 17799
rect 10962 17796 10968 17808
rect 10551 17768 10968 17796
rect 10551 17765 10563 17768
rect 10505 17759 10563 17765
rect 10962 17756 10968 17768
rect 11020 17756 11026 17808
rect 10134 17688 10140 17740
rect 10192 17728 10198 17740
rect 10229 17731 10287 17737
rect 10229 17728 10241 17731
rect 10192 17700 10241 17728
rect 10192 17688 10198 17700
rect 10229 17697 10241 17700
rect 10275 17697 10287 17731
rect 10229 17691 10287 17697
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 25130 17728 25136 17740
rect 24627 17700 25136 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 25130 17688 25136 17700
rect 25188 17688 25194 17740
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 24762 17320 24768 17332
rect 24723 17292 24768 17320
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 16022 17252 16028 17264
rect 15983 17224 16028 17252
rect 16022 17212 16028 17224
rect 16080 17212 16086 17264
rect 12342 17076 12348 17128
rect 12400 17116 12406 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12400 17088 12449 17116
rect 12400 17076 12406 17088
rect 12437 17085 12449 17088
rect 12483 17116 12495 17119
rect 13173 17119 13231 17125
rect 13173 17116 13185 17119
rect 12483 17088 13185 17116
rect 12483 17085 12495 17088
rect 12437 17079 12495 17085
rect 13173 17085 13185 17088
rect 13219 17085 13231 17119
rect 13173 17079 13231 17085
rect 15562 17076 15568 17128
rect 15620 17116 15626 17128
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 15620 17088 15853 17116
rect 15620 17076 15626 17088
rect 15841 17085 15853 17088
rect 15887 17116 15899 17119
rect 16393 17119 16451 17125
rect 16393 17116 16405 17119
rect 15887 17088 16405 17116
rect 15887 17085 15899 17088
rect 15841 17079 15899 17085
rect 16393 17085 16405 17088
rect 16439 17085 16451 17119
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 16393 17079 16451 17085
rect 24412 17088 24593 17116
rect 12710 17048 12716 17060
rect 12671 17020 12716 17048
rect 12710 17008 12716 17020
rect 12768 17008 12774 17060
rect 24412 16992 24440 17088
rect 24581 17085 24593 17088
rect 24627 17085 24639 17119
rect 25130 17116 25136 17128
rect 25091 17088 25136 17116
rect 24581 17079 24639 17085
rect 25130 17076 25136 17088
rect 25188 17076 25194 17128
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 10192 16952 10241 16980
rect 10192 16940 10198 16952
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 24394 16980 24400 16992
rect 24355 16952 24400 16980
rect 10229 16943 10287 16949
rect 24394 16940 24400 16952
rect 24452 16940 24458 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 24026 16736 24032 16788
rect 24084 16776 24090 16788
rect 24765 16779 24823 16785
rect 24765 16776 24777 16779
rect 24084 16748 24777 16776
rect 24084 16736 24090 16748
rect 24765 16745 24777 16748
rect 24811 16745 24823 16779
rect 24765 16739 24823 16745
rect 15562 16708 15568 16720
rect 15523 16680 15568 16708
rect 15562 16668 15568 16680
rect 15620 16668 15626 16720
rect 15289 16643 15347 16649
rect 15289 16609 15301 16643
rect 15335 16640 15347 16643
rect 15378 16640 15384 16652
rect 15335 16612 15384 16640
rect 15335 16609 15347 16612
rect 15289 16603 15347 16609
rect 15378 16600 15384 16612
rect 15436 16600 15442 16652
rect 24581 16643 24639 16649
rect 24581 16609 24593 16643
rect 24627 16640 24639 16643
rect 24670 16640 24676 16652
rect 24627 16612 24676 16640
rect 24627 16609 24639 16612
rect 24581 16603 24639 16609
rect 24670 16600 24676 16612
rect 24728 16600 24734 16652
rect 24210 16396 24216 16448
rect 24268 16436 24274 16448
rect 24946 16436 24952 16448
rect 24268 16408 24952 16436
rect 24268 16396 24274 16408
rect 24946 16396 24952 16408
rect 25004 16396 25010 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 24762 16232 24768 16244
rect 24723 16204 24768 16232
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 24489 16167 24547 16173
rect 24489 16133 24501 16167
rect 24535 16164 24547 16167
rect 24670 16164 24676 16176
rect 24535 16136 24676 16164
rect 24535 16133 24547 16136
rect 24489 16127 24547 16133
rect 24670 16124 24676 16136
rect 24728 16124 24734 16176
rect 18322 16096 18328 16108
rect 18283 16068 18328 16096
rect 18322 16056 18328 16068
rect 18380 16056 18386 16108
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18095 16000 18736 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18708 15904 18736 16000
rect 24210 15988 24216 16040
rect 24268 16028 24274 16040
rect 24581 16031 24639 16037
rect 24581 16028 24593 16031
rect 24268 16000 24593 16028
rect 24268 15988 24274 16000
rect 24581 15997 24593 16000
rect 24627 16028 24639 16031
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24627 16000 25145 16028
rect 24627 15997 24639 16000
rect 24581 15991 24639 15997
rect 25133 15997 25145 16000
rect 25179 15997 25191 16031
rect 25133 15991 25191 15997
rect 15194 15852 15200 15904
rect 15252 15892 15258 15904
rect 15289 15895 15347 15901
rect 15289 15892 15301 15895
rect 15252 15864 15301 15892
rect 15252 15852 15258 15864
rect 15289 15861 15301 15864
rect 15335 15892 15347 15895
rect 15378 15892 15384 15904
rect 15335 15864 15384 15892
rect 15335 15861 15347 15864
rect 15289 15855 15347 15861
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 18690 15852 18696 15904
rect 18748 15892 18754 15904
rect 18785 15895 18843 15901
rect 18785 15892 18797 15895
rect 18748 15864 18797 15892
rect 18748 15852 18754 15864
rect 18785 15861 18797 15864
rect 18831 15861 18843 15895
rect 18785 15855 18843 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 25038 15688 25044 15700
rect 24999 15660 25044 15688
rect 25038 15648 25044 15660
rect 25096 15648 25102 15700
rect 23845 15623 23903 15629
rect 23845 15589 23857 15623
rect 23891 15620 23903 15623
rect 24670 15620 24676 15632
rect 23891 15592 24676 15620
rect 23891 15589 23903 15592
rect 23845 15583 23903 15589
rect 24670 15580 24676 15592
rect 24728 15580 24734 15632
rect 23474 15512 23480 15564
rect 23532 15552 23538 15564
rect 23569 15555 23627 15561
rect 23569 15552 23581 15555
rect 23532 15524 23581 15552
rect 23532 15512 23538 15524
rect 23569 15521 23581 15524
rect 23615 15521 23627 15555
rect 24854 15552 24860 15564
rect 24815 15524 24860 15552
rect 23569 15515 23627 15521
rect 24854 15512 24860 15524
rect 24912 15512 24918 15564
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 25498 15144 25504 15156
rect 25459 15116 25504 15144
rect 25498 15104 25504 15116
rect 25556 15104 25562 15156
rect 24210 15008 24216 15020
rect 24171 14980 24216 15008
rect 24210 14968 24216 14980
rect 24268 14968 24274 15020
rect 23474 14940 23480 14952
rect 23435 14912 23480 14940
rect 23474 14900 23480 14912
rect 23532 14900 23538 14952
rect 24029 14943 24087 14949
rect 24029 14940 24041 14943
rect 23860 14912 24041 14940
rect 23658 14764 23664 14816
rect 23716 14804 23722 14816
rect 23860 14813 23888 14912
rect 24029 14909 24041 14912
rect 24075 14909 24087 14943
rect 24029 14903 24087 14909
rect 25317 14943 25375 14949
rect 25317 14909 25329 14943
rect 25363 14940 25375 14943
rect 25406 14940 25412 14952
rect 25363 14912 25412 14940
rect 25363 14909 25375 14912
rect 25317 14903 25375 14909
rect 25406 14900 25412 14912
rect 25464 14940 25470 14952
rect 25869 14943 25927 14949
rect 25869 14940 25881 14943
rect 25464 14912 25881 14940
rect 25464 14900 25470 14912
rect 25869 14909 25881 14912
rect 25915 14909 25927 14943
rect 25869 14903 25927 14909
rect 23845 14807 23903 14813
rect 23845 14804 23857 14807
rect 23716 14776 23857 14804
rect 23716 14764 23722 14776
rect 23845 14773 23857 14776
rect 23891 14773 23903 14807
rect 24854 14804 24860 14816
rect 24815 14776 24860 14804
rect 23845 14767 23903 14773
rect 24854 14764 24860 14776
rect 24912 14764 24918 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 23382 14532 23388 14544
rect 23343 14504 23388 14532
rect 23382 14492 23388 14504
rect 23440 14492 23446 14544
rect 23106 14464 23112 14476
rect 23067 14436 23112 14464
rect 23106 14424 23112 14436
rect 23164 14424 23170 14476
rect 24581 14467 24639 14473
rect 24581 14433 24593 14467
rect 24627 14464 24639 14467
rect 24762 14464 24768 14476
rect 24627 14436 24768 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 24762 14424 24768 14436
rect 24820 14424 24826 14476
rect 20901 14399 20959 14405
rect 20901 14365 20913 14399
rect 20947 14396 20959 14399
rect 21266 14396 21272 14408
rect 20947 14368 21272 14396
rect 20947 14365 20959 14368
rect 20901 14359 20959 14365
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 24762 14260 24768 14272
rect 24723 14232 24768 14260
rect 24762 14220 24768 14232
rect 24820 14220 24826 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 24118 14016 24124 14068
rect 24176 14056 24182 14068
rect 24765 14059 24823 14065
rect 24765 14056 24777 14059
rect 24176 14028 24777 14056
rect 24176 14016 24182 14028
rect 24765 14025 24777 14028
rect 24811 14025 24823 14059
rect 24765 14019 24823 14025
rect 24854 14016 24860 14068
rect 24912 14056 24918 14068
rect 25133 14059 25191 14065
rect 25133 14056 25145 14059
rect 24912 14028 25145 14056
rect 24912 14016 24918 14028
rect 25133 14025 25145 14028
rect 25179 14025 25191 14059
rect 25133 14019 25191 14025
rect 21818 13812 21824 13864
rect 21876 13852 21882 13864
rect 23106 13852 23112 13864
rect 21876 13824 23112 13852
rect 21876 13812 21882 13824
rect 23106 13812 23112 13824
rect 23164 13812 23170 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 24412 13824 24593 13852
rect 19337 13719 19395 13725
rect 19337 13685 19349 13719
rect 19383 13716 19395 13719
rect 20438 13716 20444 13728
rect 19383 13688 20444 13716
rect 19383 13685 19395 13688
rect 19337 13679 19395 13685
rect 20438 13676 20444 13688
rect 20496 13676 20502 13728
rect 21269 13719 21327 13725
rect 21269 13685 21281 13719
rect 21315 13716 21327 13719
rect 21726 13716 21732 13728
rect 21315 13688 21732 13716
rect 21315 13685 21327 13688
rect 21269 13679 21327 13685
rect 21726 13676 21732 13688
rect 21784 13676 21790 13728
rect 22278 13716 22284 13728
rect 22239 13688 22284 13716
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 24118 13676 24124 13728
rect 24176 13716 24182 13728
rect 24412 13725 24440 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 24397 13719 24455 13725
rect 24397 13716 24409 13719
rect 24176 13688 24409 13716
rect 24176 13676 24182 13688
rect 24397 13685 24409 13688
rect 24443 13685 24455 13719
rect 24397 13679 24455 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 20898 13512 20904 13524
rect 20859 13484 20904 13512
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 21266 13512 21272 13524
rect 21227 13484 21272 13512
rect 21266 13472 21272 13484
rect 21324 13472 21330 13524
rect 23109 13515 23167 13521
rect 23109 13481 23121 13515
rect 23155 13512 23167 13515
rect 23382 13512 23388 13524
rect 23155 13484 23388 13512
rect 23155 13481 23167 13484
rect 23109 13475 23167 13481
rect 23382 13472 23388 13484
rect 23440 13472 23446 13524
rect 23566 13472 23572 13524
rect 23624 13512 23630 13524
rect 24765 13515 24823 13521
rect 24765 13512 24777 13515
rect 23624 13484 24777 13512
rect 23624 13472 23630 13484
rect 24765 13481 24777 13484
rect 24811 13481 24823 13515
rect 24765 13475 24823 13481
rect 16298 13376 16304 13388
rect 16259 13348 16304 13376
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 21361 13379 21419 13385
rect 21361 13345 21373 13379
rect 21407 13376 21419 13379
rect 21542 13376 21548 13388
rect 21407 13348 21548 13376
rect 21407 13345 21419 13348
rect 21361 13339 21419 13345
rect 21542 13336 21548 13348
rect 21600 13336 21606 13388
rect 22922 13336 22928 13388
rect 22980 13376 22986 13388
rect 23017 13379 23075 13385
rect 23017 13376 23029 13379
rect 22980 13348 23029 13376
rect 22980 13336 22986 13348
rect 23017 13345 23029 13348
rect 23063 13345 23075 13379
rect 23017 13339 23075 13345
rect 24026 13336 24032 13388
rect 24084 13376 24090 13388
rect 24581 13379 24639 13385
rect 24581 13376 24593 13379
rect 24084 13348 24593 13376
rect 24084 13336 24090 13348
rect 24581 13345 24593 13348
rect 24627 13345 24639 13379
rect 24581 13339 24639 13345
rect 18138 13308 18144 13320
rect 18099 13280 18144 13308
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 18782 13268 18788 13320
rect 18840 13308 18846 13320
rect 18877 13311 18935 13317
rect 18877 13308 18889 13311
rect 18840 13280 18889 13308
rect 18840 13268 18846 13280
rect 18877 13277 18889 13280
rect 18923 13277 18935 13311
rect 18877 13271 18935 13277
rect 21453 13311 21511 13317
rect 21453 13277 21465 13311
rect 21499 13308 21511 13311
rect 21634 13308 21640 13320
rect 21499 13280 21640 13308
rect 21499 13277 21511 13280
rect 21453 13271 21511 13277
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 23198 13308 23204 13320
rect 23159 13280 23204 13308
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 17770 13172 17776 13184
rect 17731 13144 17776 13172
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 20073 13175 20131 13181
rect 20073 13141 20085 13175
rect 20119 13172 20131 13175
rect 20530 13172 20536 13184
rect 20119 13144 20536 13172
rect 20119 13141 20131 13144
rect 20073 13135 20131 13141
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 22646 13172 22652 13184
rect 22607 13144 22652 13172
rect 22646 13132 22652 13144
rect 22704 13132 22710 13184
rect 23842 13172 23848 13184
rect 23803 13144 23848 13172
rect 23842 13132 23848 13144
rect 23900 13132 23906 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 16298 12968 16304 12980
rect 16259 12940 16304 12968
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 21085 12971 21143 12977
rect 21085 12937 21097 12971
rect 21131 12968 21143 12971
rect 21266 12968 21272 12980
rect 21131 12940 21272 12968
rect 21131 12937 21143 12940
rect 21085 12931 21143 12937
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 22373 12971 22431 12977
rect 22373 12937 22385 12971
rect 22419 12968 22431 12971
rect 23198 12968 23204 12980
rect 22419 12940 23204 12968
rect 22419 12937 22431 12940
rect 22373 12931 22431 12937
rect 23198 12928 23204 12940
rect 23256 12928 23262 12980
rect 23382 12968 23388 12980
rect 23343 12940 23388 12968
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 24026 12928 24032 12980
rect 24084 12968 24090 12980
rect 24581 12971 24639 12977
rect 24581 12968 24593 12971
rect 24084 12940 24593 12968
rect 24084 12928 24090 12940
rect 24581 12937 24593 12940
rect 24627 12937 24639 12971
rect 25774 12968 25780 12980
rect 25735 12940 25780 12968
rect 24581 12931 24639 12937
rect 25774 12928 25780 12940
rect 25832 12928 25838 12980
rect 18414 12900 18420 12912
rect 18375 12872 18420 12900
rect 18414 12860 18420 12872
rect 18472 12860 18478 12912
rect 18966 12832 18972 12844
rect 18927 12804 18972 12832
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 19518 12792 19524 12844
rect 19576 12832 19582 12844
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 19576 12804 19809 12832
rect 19576 12792 19582 12804
rect 19797 12801 19809 12804
rect 19843 12832 19855 12835
rect 20530 12832 20536 12844
rect 19843 12804 20392 12832
rect 20491 12804 20536 12832
rect 19843 12801 19855 12804
rect 19797 12795 19855 12801
rect 18325 12767 18383 12773
rect 18325 12733 18337 12767
rect 18371 12764 18383 12767
rect 18782 12764 18788 12776
rect 18371 12736 18788 12764
rect 18371 12733 18383 12736
rect 18325 12727 18383 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 20364 12773 20392 12804
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 24118 12832 24124 12844
rect 24079 12804 24124 12832
rect 24118 12792 24124 12804
rect 24176 12792 24182 12844
rect 20349 12767 20407 12773
rect 20349 12733 20361 12767
rect 20395 12733 20407 12767
rect 23842 12764 23848 12776
rect 23803 12736 23848 12764
rect 20349 12727 20407 12733
rect 23842 12724 23848 12736
rect 23900 12724 23906 12776
rect 25133 12767 25191 12773
rect 25133 12733 25145 12767
rect 25179 12764 25191 12767
rect 25774 12764 25780 12776
rect 25179 12736 25780 12764
rect 25179 12733 25191 12736
rect 25133 12727 25191 12733
rect 25774 12724 25780 12736
rect 25832 12724 25838 12776
rect 17865 12699 17923 12705
rect 17865 12665 17877 12699
rect 17911 12696 17923 12699
rect 17911 12668 18644 12696
rect 17911 12665 17923 12668
rect 17865 12659 17923 12665
rect 18616 12640 18644 12668
rect 19334 12656 19340 12708
rect 19392 12696 19398 12708
rect 19521 12699 19579 12705
rect 19521 12696 19533 12699
rect 19392 12668 19533 12696
rect 19392 12656 19398 12668
rect 19521 12665 19533 12668
rect 19567 12696 19579 12699
rect 20441 12699 20499 12705
rect 20441 12696 20453 12699
rect 19567 12668 20453 12696
rect 19567 12665 19579 12668
rect 19521 12659 19579 12665
rect 20441 12665 20453 12668
rect 20487 12665 20499 12699
rect 20441 12659 20499 12665
rect 21453 12699 21511 12705
rect 21453 12665 21465 12699
rect 21499 12696 21511 12699
rect 21634 12696 21640 12708
rect 21499 12668 21640 12696
rect 21499 12665 21511 12668
rect 21453 12659 21511 12665
rect 21634 12656 21640 12668
rect 21692 12656 21698 12708
rect 18598 12588 18604 12640
rect 18656 12628 18662 12640
rect 18877 12631 18935 12637
rect 18877 12628 18889 12631
rect 18656 12600 18889 12628
rect 18656 12588 18662 12600
rect 18877 12597 18889 12600
rect 18923 12597 18935 12631
rect 19978 12628 19984 12640
rect 19939 12600 19984 12628
rect 18877 12591 18935 12597
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 21266 12588 21272 12640
rect 21324 12628 21330 12640
rect 21542 12628 21548 12640
rect 21324 12600 21548 12628
rect 21324 12588 21330 12600
rect 21542 12588 21548 12600
rect 21600 12628 21606 12640
rect 21729 12631 21787 12637
rect 21729 12628 21741 12631
rect 21600 12600 21741 12628
rect 21600 12588 21606 12600
rect 21729 12597 21741 12600
rect 21775 12597 21787 12631
rect 21729 12591 21787 12597
rect 22465 12631 22523 12637
rect 22465 12597 22477 12631
rect 22511 12628 22523 12631
rect 22738 12628 22744 12640
rect 22511 12600 22744 12628
rect 22511 12597 22523 12600
rect 22465 12591 22523 12597
rect 22738 12588 22744 12600
rect 22796 12588 22802 12640
rect 22922 12628 22928 12640
rect 22883 12600 22928 12628
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 25314 12628 25320 12640
rect 25275 12600 25320 12628
rect 25314 12588 25320 12600
rect 25372 12588 25378 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 18509 12427 18567 12433
rect 18509 12393 18521 12427
rect 18555 12424 18567 12427
rect 18966 12424 18972 12436
rect 18555 12396 18972 12424
rect 18555 12393 18567 12396
rect 18509 12387 18567 12393
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 19242 12424 19248 12436
rect 19203 12396 19248 12424
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21910 12424 21916 12436
rect 20772 12396 21916 12424
rect 20772 12384 20778 12396
rect 21910 12384 21916 12396
rect 21968 12424 21974 12436
rect 22281 12427 22339 12433
rect 22281 12424 22293 12427
rect 21968 12396 22293 12424
rect 21968 12384 21974 12396
rect 22281 12393 22293 12396
rect 22327 12393 22339 12427
rect 22281 12387 22339 12393
rect 23750 12384 23756 12436
rect 23808 12424 23814 12436
rect 24121 12427 24179 12433
rect 24121 12424 24133 12427
rect 23808 12396 24133 12424
rect 23808 12384 23814 12396
rect 24121 12393 24133 12396
rect 24167 12424 24179 12427
rect 24302 12424 24308 12436
rect 24167 12396 24308 12424
rect 24167 12393 24179 12396
rect 24121 12387 24179 12393
rect 24302 12384 24308 12396
rect 24360 12384 24366 12436
rect 17402 12356 17408 12368
rect 17363 12328 17408 12356
rect 17402 12316 17408 12328
rect 17460 12316 17466 12368
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12288 17187 12291
rect 17494 12288 17500 12300
rect 17175 12260 17500 12288
rect 17175 12257 17187 12260
rect 17129 12251 17187 12257
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19613 12291 19671 12297
rect 19613 12288 19625 12291
rect 19392 12260 19625 12288
rect 19392 12248 19398 12260
rect 19613 12257 19625 12260
rect 19659 12257 19671 12291
rect 21157 12291 21215 12297
rect 21157 12288 21169 12291
rect 19613 12251 19671 12257
rect 20824 12260 21169 12288
rect 16117 12223 16175 12229
rect 16117 12189 16129 12223
rect 16163 12220 16175 12223
rect 17034 12220 17040 12232
rect 16163 12192 17040 12220
rect 16163 12189 16175 12192
rect 16117 12183 16175 12189
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 19702 12220 19708 12232
rect 19663 12192 19708 12220
rect 19702 12180 19708 12192
rect 19760 12180 19766 12232
rect 19797 12223 19855 12229
rect 19797 12189 19809 12223
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 19153 12155 19211 12161
rect 19153 12121 19165 12155
rect 19199 12152 19211 12155
rect 19812 12152 19840 12183
rect 20824 12164 20852 12260
rect 21157 12257 21169 12260
rect 21203 12257 21215 12291
rect 24026 12288 24032 12300
rect 23987 12260 24032 12288
rect 21157 12251 21215 12257
rect 24026 12248 24032 12260
rect 24084 12248 24090 12300
rect 25225 12291 25283 12297
rect 25225 12257 25237 12291
rect 25271 12288 25283 12291
rect 25682 12288 25688 12300
rect 25271 12260 25688 12288
rect 25271 12257 25283 12260
rect 25225 12251 25283 12257
rect 25682 12248 25688 12260
rect 25740 12248 25746 12300
rect 20901 12223 20959 12229
rect 20901 12189 20913 12223
rect 20947 12189 20959 12223
rect 20901 12183 20959 12189
rect 20806 12152 20812 12164
rect 19199 12124 20812 12152
rect 19199 12121 19211 12124
rect 19153 12115 19211 12121
rect 20806 12112 20812 12124
rect 20864 12112 20870 12164
rect 20254 12084 20260 12096
rect 20215 12056 20260 12084
rect 20254 12044 20260 12056
rect 20312 12084 20318 12096
rect 20916 12084 20944 12183
rect 24210 12180 24216 12232
rect 24268 12220 24274 12232
rect 24268 12192 24313 12220
rect 24268 12180 24274 12192
rect 20312 12056 20944 12084
rect 20312 12044 20318 12056
rect 22462 12044 22468 12096
rect 22520 12084 22526 12096
rect 22646 12084 22652 12096
rect 22520 12056 22652 12084
rect 22520 12044 22526 12056
rect 22646 12044 22652 12056
rect 22704 12084 22710 12096
rect 22833 12087 22891 12093
rect 22833 12084 22845 12087
rect 22704 12056 22845 12084
rect 22704 12044 22710 12056
rect 22833 12053 22845 12056
rect 22879 12053 22891 12087
rect 22833 12047 22891 12053
rect 23198 12044 23204 12096
rect 23256 12084 23262 12096
rect 23474 12084 23480 12096
rect 23256 12056 23480 12084
rect 23256 12044 23262 12056
rect 23474 12044 23480 12056
rect 23532 12044 23538 12096
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 23661 12087 23719 12093
rect 23661 12084 23673 12087
rect 23624 12056 23673 12084
rect 23624 12044 23630 12056
rect 23661 12053 23673 12056
rect 23707 12053 23719 12087
rect 23661 12047 23719 12053
rect 24118 12044 24124 12096
rect 24176 12084 24182 12096
rect 24673 12087 24731 12093
rect 24673 12084 24685 12087
rect 24176 12056 24685 12084
rect 24176 12044 24182 12056
rect 24673 12053 24685 12056
rect 24719 12053 24731 12087
rect 24673 12047 24731 12053
rect 24854 12044 24860 12096
rect 24912 12084 24918 12096
rect 25409 12087 25467 12093
rect 25409 12084 25421 12087
rect 24912 12056 25421 12084
rect 24912 12044 24918 12056
rect 25409 12053 25421 12056
rect 25455 12053 25467 12087
rect 25409 12047 25467 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 18969 11883 19027 11889
rect 18969 11849 18981 11883
rect 19015 11880 19027 11883
rect 19702 11880 19708 11892
rect 19015 11852 19708 11880
rect 19015 11849 19027 11852
rect 18969 11843 19027 11849
rect 19702 11840 19708 11852
rect 19760 11840 19766 11892
rect 20806 11880 20812 11892
rect 20767 11852 20812 11880
rect 20806 11840 20812 11852
rect 20864 11880 20870 11892
rect 21361 11883 21419 11889
rect 21361 11880 21373 11883
rect 20864 11852 21373 11880
rect 20864 11840 20870 11852
rect 21361 11849 21373 11852
rect 21407 11849 21419 11883
rect 21361 11843 21419 11849
rect 22922 11840 22928 11892
rect 22980 11880 22986 11892
rect 23477 11883 23535 11889
rect 23477 11880 23489 11883
rect 22980 11852 23489 11880
rect 22980 11840 22986 11852
rect 23477 11849 23489 11852
rect 23523 11880 23535 11883
rect 23934 11880 23940 11892
rect 23523 11852 23940 11880
rect 23523 11849 23535 11852
rect 23477 11843 23535 11849
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 25682 11880 25688 11892
rect 25643 11852 25688 11880
rect 25682 11840 25688 11852
rect 25740 11840 25746 11892
rect 18414 11744 18420 11756
rect 18375 11716 18420 11744
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 22462 11744 22468 11756
rect 22423 11716 22468 11744
rect 22462 11704 22468 11716
rect 22520 11704 22526 11756
rect 22649 11747 22707 11753
rect 22649 11713 22661 11747
rect 22695 11744 22707 11747
rect 23106 11744 23112 11756
rect 22695 11716 23112 11744
rect 22695 11713 22707 11716
rect 22649 11707 22707 11713
rect 23106 11704 23112 11716
rect 23164 11704 23170 11756
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11676 16451 11679
rect 16439 11648 17264 11676
rect 16439 11645 16451 11648
rect 16393 11639 16451 11645
rect 16669 11611 16727 11617
rect 16669 11577 16681 11611
rect 16715 11608 16727 11611
rect 16758 11608 16764 11620
rect 16715 11580 16764 11608
rect 16715 11577 16727 11580
rect 16669 11571 16727 11577
rect 16758 11568 16764 11580
rect 16816 11568 16822 11620
rect 17236 11617 17264 11648
rect 18230 11636 18236 11688
rect 18288 11676 18294 11688
rect 19429 11679 19487 11685
rect 19429 11676 19441 11679
rect 18288 11648 19441 11676
rect 18288 11636 18294 11648
rect 19429 11645 19441 11648
rect 19475 11676 19487 11679
rect 20254 11676 20260 11688
rect 19475 11648 20260 11676
rect 19475 11645 19487 11648
rect 19429 11639 19487 11645
rect 20254 11636 20260 11648
rect 20312 11636 20318 11688
rect 21913 11679 21971 11685
rect 21913 11645 21925 11679
rect 21959 11676 21971 11679
rect 22278 11676 22284 11688
rect 21959 11648 22284 11676
rect 21959 11645 21971 11648
rect 21913 11639 21971 11645
rect 22278 11636 22284 11648
rect 22336 11676 22342 11688
rect 22373 11679 22431 11685
rect 22373 11676 22385 11679
rect 22336 11648 22385 11676
rect 22336 11636 22342 11648
rect 22373 11645 22385 11648
rect 22419 11645 22431 11679
rect 22373 11639 22431 11645
rect 23661 11679 23719 11685
rect 23661 11645 23673 11679
rect 23707 11676 23719 11679
rect 23707 11648 24072 11676
rect 23707 11645 23719 11648
rect 23661 11639 23719 11645
rect 24044 11620 24072 11648
rect 17221 11611 17279 11617
rect 17221 11577 17233 11611
rect 17267 11608 17279 11611
rect 17402 11608 17408 11620
rect 17267 11580 17408 11608
rect 17267 11577 17279 11580
rect 17221 11571 17279 11577
rect 17402 11568 17408 11580
rect 17460 11568 17466 11620
rect 18966 11568 18972 11620
rect 19024 11608 19030 11620
rect 19518 11608 19524 11620
rect 19024 11580 19524 11608
rect 19024 11568 19030 11580
rect 19518 11568 19524 11580
rect 19576 11608 19582 11620
rect 19674 11611 19732 11617
rect 19674 11608 19686 11611
rect 19576 11580 19686 11608
rect 19576 11568 19582 11580
rect 19674 11577 19686 11580
rect 19720 11577 19732 11611
rect 19674 11571 19732 11577
rect 22738 11568 22744 11620
rect 22796 11608 22802 11620
rect 23474 11608 23480 11620
rect 22796 11580 23480 11608
rect 22796 11568 22802 11580
rect 23474 11568 23480 11580
rect 23532 11608 23538 11620
rect 23906 11611 23964 11617
rect 23906 11608 23918 11611
rect 23532 11580 23918 11608
rect 23532 11568 23538 11580
rect 23906 11577 23918 11580
rect 23952 11577 23964 11611
rect 23906 11571 23964 11577
rect 24026 11568 24032 11620
rect 24084 11568 24090 11620
rect 17494 11540 17500 11552
rect 17455 11512 17500 11540
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 19334 11540 19340 11552
rect 19295 11512 19340 11540
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 20714 11500 20720 11552
rect 20772 11540 20778 11552
rect 22005 11543 22063 11549
rect 22005 11540 22017 11543
rect 20772 11512 22017 11540
rect 20772 11500 20778 11512
rect 22005 11509 22017 11512
rect 22051 11509 22063 11543
rect 23106 11540 23112 11552
rect 23067 11512 23112 11540
rect 22005 11503 22063 11509
rect 23106 11500 23112 11512
rect 23164 11500 23170 11552
rect 25038 11540 25044 11552
rect 24999 11512 25044 11540
rect 25038 11500 25044 11512
rect 25096 11500 25102 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 16669 11339 16727 11345
rect 16669 11305 16681 11339
rect 16715 11336 16727 11339
rect 17494 11336 17500 11348
rect 16715 11308 17500 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 17494 11296 17500 11308
rect 17552 11296 17558 11348
rect 19518 11296 19524 11348
rect 19576 11336 19582 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 19576 11308 19717 11336
rect 19576 11296 19582 11308
rect 19705 11305 19717 11308
rect 19751 11336 19763 11339
rect 20257 11339 20315 11345
rect 20257 11336 20269 11339
rect 19751 11308 20269 11336
rect 19751 11305 19763 11308
rect 19705 11299 19763 11305
rect 20257 11305 20269 11308
rect 20303 11305 20315 11339
rect 22738 11336 22744 11348
rect 22699 11308 22744 11336
rect 20257 11299 20315 11305
rect 22738 11296 22744 11308
rect 22796 11296 22802 11348
rect 23750 11336 23756 11348
rect 23711 11308 23756 11336
rect 23750 11296 23756 11308
rect 23808 11296 23814 11348
rect 23842 11296 23848 11348
rect 23900 11336 23906 11348
rect 24026 11336 24032 11348
rect 23900 11308 24032 11336
rect 23900 11296 23906 11308
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 17034 11268 17040 11280
rect 16995 11240 17040 11268
rect 17034 11228 17040 11240
rect 17092 11228 17098 11280
rect 22002 11268 22008 11280
rect 21468 11240 22008 11268
rect 21468 11212 21496 11240
rect 22002 11228 22008 11240
rect 22060 11228 22066 11280
rect 23106 11228 23112 11280
rect 23164 11268 23170 11280
rect 23474 11268 23480 11280
rect 23164 11240 23480 11268
rect 23164 11228 23170 11240
rect 23474 11228 23480 11240
rect 23532 11268 23538 11280
rect 24112 11271 24170 11277
rect 24112 11268 24124 11271
rect 23532 11240 24124 11268
rect 23532 11228 23538 11240
rect 24112 11237 24124 11240
rect 24158 11268 24170 11271
rect 25038 11268 25044 11280
rect 24158 11240 25044 11268
rect 24158 11237 24170 11240
rect 24112 11231 24170 11237
rect 25038 11228 25044 11240
rect 25096 11228 25102 11280
rect 13906 11200 13912 11212
rect 13867 11172 13912 11200
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 15378 11200 15384 11212
rect 15335 11172 15384 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 18230 11160 18236 11212
rect 18288 11200 18294 11212
rect 18325 11203 18383 11209
rect 18325 11200 18337 11203
rect 18288 11172 18337 11200
rect 18288 11160 18294 11172
rect 18325 11169 18337 11172
rect 18371 11169 18383 11203
rect 18325 11163 18383 11169
rect 18414 11160 18420 11212
rect 18472 11200 18478 11212
rect 18581 11203 18639 11209
rect 18581 11200 18593 11203
rect 18472 11172 18593 11200
rect 18472 11160 18478 11172
rect 18581 11169 18593 11172
rect 18627 11169 18639 11203
rect 18581 11163 18639 11169
rect 20254 11160 20260 11212
rect 20312 11200 20318 11212
rect 20625 11203 20683 11209
rect 20625 11200 20637 11203
rect 20312 11172 20637 11200
rect 20312 11160 20318 11172
rect 20625 11169 20637 11172
rect 20671 11169 20683 11203
rect 20625 11163 20683 11169
rect 21269 11203 21327 11209
rect 21269 11169 21281 11203
rect 21315 11200 21327 11203
rect 21450 11200 21456 11212
rect 21315 11172 21456 11200
rect 21315 11169 21327 11172
rect 21269 11163 21327 11169
rect 14185 11135 14243 11141
rect 14185 11101 14197 11135
rect 14231 11132 14243 11135
rect 14274 11132 14280 11144
rect 14231 11104 14280 11132
rect 14231 11101 14243 11104
rect 14185 11095 14243 11101
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 15470 11132 15476 11144
rect 15431 11104 15476 11132
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 17129 11135 17187 11141
rect 17129 11101 17141 11135
rect 17175 11101 17187 11135
rect 17310 11132 17316 11144
rect 17271 11104 17316 11132
rect 17129 11095 17187 11101
rect 16574 11064 16580 11076
rect 16535 11036 16580 11064
rect 16574 11024 16580 11036
rect 16632 11064 16638 11076
rect 17144 11064 17172 11095
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 20640 11132 20668 11163
rect 21450 11160 21456 11172
rect 21508 11160 21514 11212
rect 21628 11203 21686 11209
rect 21628 11169 21640 11203
rect 21674 11200 21686 11203
rect 21910 11200 21916 11212
rect 21674 11172 21916 11200
rect 21674 11169 21686 11172
rect 21628 11163 21686 11169
rect 21910 11160 21916 11172
rect 21968 11160 21974 11212
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 20640 11104 21373 11132
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 23750 11092 23756 11144
rect 23808 11132 23814 11144
rect 23845 11135 23903 11141
rect 23845 11132 23857 11135
rect 23808 11104 23857 11132
rect 23808 11092 23814 11104
rect 23845 11101 23857 11104
rect 23891 11101 23903 11135
rect 23845 11095 23903 11101
rect 25225 11067 25283 11073
rect 25225 11064 25237 11067
rect 16632 11036 17172 11064
rect 24780 11036 25237 11064
rect 16632 11024 16638 11036
rect 18138 10996 18144 11008
rect 18099 10968 18144 10996
rect 18138 10956 18144 10968
rect 18196 10956 18202 11008
rect 23385 10999 23443 11005
rect 23385 10965 23397 10999
rect 23431 10996 23443 10999
rect 23842 10996 23848 11008
rect 23431 10968 23848 10996
rect 23431 10965 23443 10968
rect 23385 10959 23443 10965
rect 23842 10956 23848 10968
rect 23900 10996 23906 11008
rect 24210 10996 24216 11008
rect 23900 10968 24216 10996
rect 23900 10956 23906 10968
rect 24210 10956 24216 10968
rect 24268 10996 24274 11008
rect 24780 10996 24808 11036
rect 25225 11033 25237 11036
rect 25271 11033 25283 11067
rect 25225 11027 25283 11033
rect 24268 10968 24808 10996
rect 24268 10956 24274 10968
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14185 10795 14243 10801
rect 14185 10792 14197 10795
rect 13964 10764 14197 10792
rect 13964 10752 13970 10764
rect 14185 10761 14197 10764
rect 14231 10761 14243 10795
rect 14185 10755 14243 10761
rect 16761 10795 16819 10801
rect 16761 10761 16773 10795
rect 16807 10792 16819 10795
rect 17034 10792 17040 10804
rect 16807 10764 17040 10792
rect 16807 10761 16819 10764
rect 16761 10755 16819 10761
rect 17034 10752 17040 10764
rect 17092 10752 17098 10804
rect 17129 10795 17187 10801
rect 17129 10761 17141 10795
rect 17175 10792 17187 10795
rect 17310 10792 17316 10804
rect 17175 10764 17316 10792
rect 17175 10761 17187 10764
rect 17129 10755 17187 10761
rect 17310 10752 17316 10764
rect 17368 10792 17374 10804
rect 17773 10795 17831 10801
rect 17773 10792 17785 10795
rect 17368 10764 17785 10792
rect 17368 10752 17374 10764
rect 17773 10761 17785 10764
rect 17819 10761 17831 10795
rect 17773 10755 17831 10761
rect 20073 10795 20131 10801
rect 20073 10761 20085 10795
rect 20119 10792 20131 10795
rect 20254 10792 20260 10804
rect 20119 10764 20260 10792
rect 20119 10761 20131 10764
rect 20073 10755 20131 10761
rect 17788 10656 17816 10755
rect 20254 10752 20260 10764
rect 20312 10792 20318 10804
rect 20625 10795 20683 10801
rect 20625 10792 20637 10795
rect 20312 10764 20637 10792
rect 20312 10752 20318 10764
rect 20625 10761 20637 10764
rect 20671 10761 20683 10795
rect 20625 10755 20683 10761
rect 21453 10795 21511 10801
rect 21453 10761 21465 10795
rect 21499 10792 21511 10795
rect 21542 10792 21548 10804
rect 21499 10764 21548 10792
rect 21499 10761 21511 10764
rect 21453 10755 21511 10761
rect 17788 10628 18184 10656
rect 14182 10548 14188 10600
rect 14240 10588 14246 10600
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 14240 10560 14565 10588
rect 14240 10548 14246 10560
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 14734 10588 14740 10600
rect 14695 10560 14740 10588
rect 14553 10551 14611 10557
rect 14568 10520 14596 10551
rect 14734 10548 14740 10560
rect 14792 10548 14798 10600
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10557 18107 10591
rect 18156 10588 18184 10628
rect 18305 10591 18363 10597
rect 18305 10588 18317 10591
rect 18156 10560 18317 10588
rect 18049 10551 18107 10557
rect 18305 10557 18317 10560
rect 18351 10557 18363 10591
rect 18305 10551 18363 10557
rect 20809 10591 20867 10597
rect 20809 10557 20821 10591
rect 20855 10588 20867 10591
rect 21468 10588 21496 10755
rect 21542 10752 21548 10764
rect 21600 10752 21606 10804
rect 21818 10752 21824 10804
rect 21876 10792 21882 10804
rect 21913 10795 21971 10801
rect 21913 10792 21925 10795
rect 21876 10764 21925 10792
rect 21876 10752 21882 10764
rect 21913 10761 21925 10764
rect 21959 10761 21971 10795
rect 23474 10792 23480 10804
rect 23435 10764 23480 10792
rect 21913 10755 21971 10761
rect 23474 10752 23480 10764
rect 23532 10752 23538 10804
rect 21821 10659 21879 10665
rect 21821 10625 21833 10659
rect 21867 10656 21879 10659
rect 21910 10656 21916 10668
rect 21867 10628 21916 10656
rect 21867 10625 21879 10628
rect 21821 10619 21879 10625
rect 21910 10616 21916 10628
rect 21968 10616 21974 10668
rect 22462 10656 22468 10668
rect 22423 10628 22468 10656
rect 22462 10616 22468 10628
rect 22520 10616 22526 10668
rect 20855 10560 21496 10588
rect 20855 10557 20867 10560
rect 20809 10551 20867 10557
rect 14982 10523 15040 10529
rect 14982 10520 14994 10523
rect 14568 10492 14994 10520
rect 14982 10489 14994 10492
rect 15028 10489 15040 10523
rect 18064 10520 18092 10551
rect 22094 10548 22100 10600
rect 22152 10588 22158 10600
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 22152 10560 22293 10588
rect 22152 10548 22158 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 23661 10591 23719 10597
rect 23661 10557 23673 10591
rect 23707 10588 23719 10591
rect 23750 10588 23756 10600
rect 23707 10560 23756 10588
rect 23707 10557 23719 10560
rect 23661 10551 23719 10557
rect 23750 10548 23756 10560
rect 23808 10588 23814 10600
rect 23808 10560 25360 10588
rect 23808 10548 23814 10560
rect 18138 10520 18144 10532
rect 18064 10492 18144 10520
rect 14982 10483 15040 10489
rect 18138 10480 18144 10492
rect 18196 10480 18202 10532
rect 23109 10523 23167 10529
rect 23109 10489 23121 10523
rect 23155 10520 23167 10523
rect 23842 10520 23848 10532
rect 23155 10492 23848 10520
rect 23155 10489 23167 10492
rect 23109 10483 23167 10489
rect 23842 10480 23848 10492
rect 23900 10529 23906 10532
rect 23900 10523 23964 10529
rect 23900 10489 23918 10523
rect 23952 10489 23964 10523
rect 23900 10483 23964 10489
rect 23900 10480 23906 10483
rect 25332 10464 25360 10560
rect 13722 10452 13728 10464
rect 13683 10424 13728 10452
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 16114 10452 16120 10464
rect 16075 10424 16120 10452
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 17497 10455 17555 10461
rect 17497 10421 17509 10455
rect 17543 10452 17555 10455
rect 18414 10452 18420 10464
rect 17543 10424 18420 10452
rect 17543 10421 17555 10424
rect 17497 10415 17555 10421
rect 18414 10412 18420 10424
rect 18472 10452 18478 10464
rect 19429 10455 19487 10461
rect 19429 10452 19441 10455
rect 18472 10424 19441 10452
rect 18472 10412 18478 10424
rect 19429 10421 19441 10424
rect 19475 10421 19487 10455
rect 20990 10452 20996 10464
rect 20951 10424 20996 10452
rect 19429 10415 19487 10421
rect 20990 10412 20996 10424
rect 21048 10412 21054 10464
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 22373 10455 22431 10461
rect 22373 10452 22385 10455
rect 22152 10424 22385 10452
rect 22152 10412 22158 10424
rect 22373 10421 22385 10424
rect 22419 10421 22431 10455
rect 22373 10415 22431 10421
rect 24026 10412 24032 10464
rect 24084 10452 24090 10464
rect 25041 10455 25099 10461
rect 25041 10452 25053 10455
rect 24084 10424 25053 10452
rect 24084 10412 24090 10424
rect 25041 10421 25053 10424
rect 25087 10421 25099 10455
rect 25041 10415 25099 10421
rect 25314 10412 25320 10464
rect 25372 10452 25378 10464
rect 25593 10455 25651 10461
rect 25593 10452 25605 10455
rect 25372 10424 25605 10452
rect 25372 10412 25378 10424
rect 25593 10421 25605 10424
rect 25639 10452 25651 10455
rect 25961 10455 26019 10461
rect 25961 10452 25973 10455
rect 25639 10424 25973 10452
rect 25639 10421 25651 10424
rect 25593 10415 25651 10421
rect 25961 10421 25973 10424
rect 26007 10421 26019 10455
rect 25961 10415 26019 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 13630 10248 13636 10260
rect 13591 10220 13636 10248
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 15473 10251 15531 10257
rect 15473 10248 15485 10251
rect 15436 10220 15485 10248
rect 15436 10208 15442 10220
rect 15473 10217 15485 10220
rect 15519 10217 15531 10251
rect 15473 10211 15531 10217
rect 17310 10208 17316 10260
rect 17368 10248 17374 10260
rect 17497 10251 17555 10257
rect 17497 10248 17509 10251
rect 17368 10220 17509 10248
rect 17368 10208 17374 10220
rect 17497 10217 17509 10220
rect 17543 10217 17555 10251
rect 18414 10248 18420 10260
rect 18375 10220 18420 10248
rect 17497 10211 17555 10217
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18598 10248 18604 10260
rect 18559 10220 18604 10248
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 20254 10248 20260 10260
rect 20215 10220 20260 10248
rect 20254 10208 20260 10220
rect 20312 10208 20318 10260
rect 20901 10251 20959 10257
rect 20901 10217 20913 10251
rect 20947 10217 20959 10251
rect 20901 10211 20959 10217
rect 16114 10140 16120 10192
rect 16172 10180 16178 10192
rect 16362 10183 16420 10189
rect 16362 10180 16374 10183
rect 16172 10152 16374 10180
rect 16172 10140 16178 10152
rect 16362 10149 16374 10152
rect 16408 10149 16420 10183
rect 18432 10180 18460 10208
rect 20916 10180 20944 10211
rect 21174 10208 21180 10260
rect 21232 10248 21238 10260
rect 21269 10251 21327 10257
rect 21269 10248 21281 10251
rect 21232 10220 21281 10248
rect 21232 10208 21238 10220
rect 21269 10217 21281 10220
rect 21315 10217 21327 10251
rect 21269 10211 21327 10217
rect 22373 10251 22431 10257
rect 22373 10217 22385 10251
rect 22419 10248 22431 10251
rect 22462 10248 22468 10260
rect 22419 10220 22468 10248
rect 22419 10217 22431 10220
rect 22373 10211 22431 10217
rect 22462 10208 22468 10220
rect 22520 10208 22526 10260
rect 22922 10248 22928 10260
rect 22883 10220 22928 10248
rect 22922 10208 22928 10220
rect 22980 10208 22986 10260
rect 23382 10248 23388 10260
rect 23343 10220 23388 10248
rect 23382 10208 23388 10220
rect 23440 10208 23446 10260
rect 24026 10248 24032 10260
rect 23987 10220 24032 10248
rect 24026 10208 24032 10220
rect 24084 10208 24090 10260
rect 24486 10248 24492 10260
rect 24447 10220 24492 10248
rect 24486 10208 24492 10220
rect 24544 10208 24550 10260
rect 21358 10180 21364 10192
rect 18432 10152 19196 10180
rect 20916 10152 21364 10180
rect 16362 10143 16420 10149
rect 13354 10072 13360 10124
rect 13412 10112 13418 10124
rect 13722 10112 13728 10124
rect 13412 10084 13728 10112
rect 13412 10072 13418 10084
rect 13722 10072 13728 10084
rect 13780 10112 13786 10124
rect 14001 10115 14059 10121
rect 14001 10112 14013 10115
rect 13780 10084 14013 10112
rect 13780 10072 13786 10084
rect 14001 10081 14013 10084
rect 14047 10081 14059 10115
rect 14001 10075 14059 10081
rect 14090 10072 14096 10124
rect 14148 10112 14154 10124
rect 14148 10084 14193 10112
rect 14148 10072 14154 10084
rect 18322 10072 18328 10124
rect 18380 10112 18386 10124
rect 18969 10115 19027 10121
rect 18969 10112 18981 10115
rect 18380 10084 18981 10112
rect 18380 10072 18386 10084
rect 18969 10081 18981 10084
rect 19015 10081 19027 10115
rect 18969 10075 19027 10081
rect 14182 10044 14188 10056
rect 14143 10016 14188 10044
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 16117 10047 16175 10053
rect 16117 10044 16129 10047
rect 15948 10016 16129 10044
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 13081 9911 13139 9917
rect 13081 9908 13093 9911
rect 12860 9880 13093 9908
rect 12860 9868 12866 9880
rect 13081 9877 13093 9880
rect 13127 9877 13139 9911
rect 13538 9908 13544 9920
rect 13499 9880 13544 9908
rect 13081 9871 13139 9877
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 14829 9911 14887 9917
rect 14829 9908 14841 9911
rect 14792 9880 14841 9908
rect 14792 9868 14798 9880
rect 14829 9877 14841 9880
rect 14875 9908 14887 9911
rect 15378 9908 15384 9920
rect 14875 9880 15384 9908
rect 14875 9877 14887 9880
rect 14829 9871 14887 9877
rect 15378 9868 15384 9880
rect 15436 9908 15442 9920
rect 15948 9917 15976 10016
rect 16117 10013 16129 10016
rect 16163 10013 16175 10047
rect 16117 10007 16175 10013
rect 17954 10004 17960 10056
rect 18012 10044 18018 10056
rect 19058 10044 19064 10056
rect 18012 10016 19064 10044
rect 18012 10004 18018 10016
rect 19058 10004 19064 10016
rect 19116 10004 19122 10056
rect 19168 10053 19196 10152
rect 21358 10140 21364 10152
rect 21416 10140 21422 10192
rect 21726 10140 21732 10192
rect 21784 10180 21790 10192
rect 23014 10180 23020 10192
rect 21784 10152 23020 10180
rect 21784 10140 21790 10152
rect 23014 10140 23020 10152
rect 23072 10180 23078 10192
rect 23293 10183 23351 10189
rect 23293 10180 23305 10183
rect 23072 10152 23305 10180
rect 23072 10140 23078 10152
rect 23293 10149 23305 10152
rect 23339 10149 23351 10183
rect 23293 10143 23351 10149
rect 24854 10112 24860 10124
rect 24815 10084 24860 10112
rect 24854 10072 24860 10084
rect 24912 10072 24918 10124
rect 24949 10115 25007 10121
rect 24949 10081 24961 10115
rect 24995 10112 25007 10115
rect 25774 10112 25780 10124
rect 24995 10084 25780 10112
rect 24995 10081 25007 10084
rect 24949 10075 25007 10081
rect 25774 10072 25780 10084
rect 25832 10072 25838 10124
rect 19153 10047 19211 10053
rect 19153 10013 19165 10047
rect 19199 10013 19211 10047
rect 21361 10047 21419 10053
rect 21361 10044 21373 10047
rect 19153 10007 19211 10013
rect 20732 10016 21373 10044
rect 20732 9920 20760 10016
rect 21361 10013 21373 10016
rect 21407 10013 21419 10047
rect 21542 10044 21548 10056
rect 21503 10016 21548 10044
rect 21361 10007 21419 10013
rect 21542 10004 21548 10016
rect 21600 10004 21606 10056
rect 23474 10004 23480 10056
rect 23532 10044 23538 10056
rect 23569 10047 23627 10053
rect 23569 10044 23581 10047
rect 23532 10016 23581 10044
rect 23532 10004 23538 10016
rect 23569 10013 23581 10016
rect 23615 10044 23627 10047
rect 24026 10044 24032 10056
rect 23615 10016 24032 10044
rect 23615 10013 23627 10016
rect 23569 10007 23627 10013
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 25041 10047 25099 10053
rect 25041 10013 25053 10047
rect 25087 10013 25099 10047
rect 25041 10007 25099 10013
rect 22094 9936 22100 9988
rect 22152 9976 22158 9988
rect 22649 9979 22707 9985
rect 22649 9976 22661 9979
rect 22152 9948 22661 9976
rect 22152 9936 22158 9948
rect 22649 9945 22661 9948
rect 22695 9945 22707 9979
rect 24302 9976 24308 9988
rect 24263 9948 24308 9976
rect 22649 9939 22707 9945
rect 24302 9936 24308 9948
rect 24360 9976 24366 9988
rect 25056 9976 25084 10007
rect 24360 9948 25084 9976
rect 24360 9936 24366 9948
rect 15933 9911 15991 9917
rect 15933 9908 15945 9911
rect 15436 9880 15945 9908
rect 15436 9868 15442 9880
rect 15933 9877 15945 9880
rect 15979 9877 15991 9911
rect 18138 9908 18144 9920
rect 18099 9880 18144 9908
rect 15933 9871 15991 9877
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 20714 9908 20720 9920
rect 20675 9880 20720 9908
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 21910 9908 21916 9920
rect 21871 9880 21916 9908
rect 21910 9868 21916 9880
rect 21968 9868 21974 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 13354 9704 13360 9716
rect 13315 9676 13360 9704
rect 13354 9664 13360 9676
rect 13412 9664 13418 9716
rect 20254 9664 20260 9716
rect 20312 9704 20318 9716
rect 20901 9707 20959 9713
rect 20312 9676 20760 9704
rect 20312 9664 20318 9676
rect 17865 9639 17923 9645
rect 17865 9605 17877 9639
rect 17911 9636 17923 9639
rect 17954 9636 17960 9648
rect 17911 9608 17960 9636
rect 17911 9605 17923 9608
rect 17865 9599 17923 9605
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 19886 9636 19892 9648
rect 19847 9608 19892 9636
rect 19886 9596 19892 9608
rect 19944 9596 19950 9648
rect 20732 9636 20760 9676
rect 20901 9673 20913 9707
rect 20947 9704 20959 9707
rect 21174 9704 21180 9716
rect 20947 9676 21180 9704
rect 20947 9673 20959 9676
rect 20901 9667 20959 9673
rect 21174 9664 21180 9676
rect 21232 9664 21238 9716
rect 23014 9704 23020 9716
rect 22975 9676 23020 9704
rect 23014 9664 23020 9676
rect 23072 9664 23078 9716
rect 23385 9707 23443 9713
rect 23385 9673 23397 9707
rect 23431 9704 23443 9707
rect 23474 9704 23480 9716
rect 23431 9676 23480 9704
rect 23431 9673 23443 9676
rect 23385 9667 23443 9673
rect 23474 9664 23480 9676
rect 23532 9664 23538 9716
rect 24854 9664 24860 9716
rect 24912 9704 24918 9716
rect 25593 9707 25651 9713
rect 25593 9704 25605 9707
rect 24912 9676 25605 9704
rect 24912 9664 24918 9676
rect 25593 9673 25605 9676
rect 25639 9673 25651 9707
rect 25593 9667 25651 9673
rect 25774 9664 25780 9716
rect 25832 9704 25838 9716
rect 25961 9707 26019 9713
rect 25961 9704 25973 9707
rect 25832 9676 25973 9704
rect 25832 9664 25838 9676
rect 25961 9673 25973 9676
rect 26007 9673 26019 9707
rect 25961 9667 26019 9673
rect 20990 9636 20996 9648
rect 20732 9608 20996 9636
rect 20990 9596 20996 9608
rect 21048 9636 21054 9648
rect 21361 9639 21419 9645
rect 21361 9636 21373 9639
rect 21048 9608 21373 9636
rect 21048 9596 21054 9608
rect 21361 9605 21373 9608
rect 21407 9605 21419 9639
rect 21361 9599 21419 9605
rect 16114 9528 16120 9580
rect 16172 9568 16178 9580
rect 16666 9568 16672 9580
rect 16172 9540 16672 9568
rect 16172 9528 16178 9540
rect 16666 9528 16672 9540
rect 16724 9568 16730 9580
rect 17129 9571 17187 9577
rect 17129 9568 17141 9571
rect 16724 9540 17141 9568
rect 16724 9528 16730 9540
rect 17129 9537 17141 9540
rect 17175 9537 17187 9571
rect 17129 9531 17187 9537
rect 20533 9571 20591 9577
rect 20533 9537 20545 9571
rect 20579 9568 20591 9571
rect 22189 9571 22247 9577
rect 22189 9568 22201 9571
rect 20579 9540 22201 9568
rect 20579 9537 20591 9540
rect 20533 9531 20591 9537
rect 21744 9512 21772 9540
rect 22189 9537 22201 9540
rect 22235 9537 22247 9571
rect 23492 9568 23520 9664
rect 23492 9540 23796 9568
rect 22189 9531 22247 9537
rect 12802 9460 12808 9512
rect 12860 9500 12866 9512
rect 13449 9503 13507 9509
rect 13449 9500 13461 9503
rect 12860 9472 13461 9500
rect 12860 9460 12866 9472
rect 13449 9469 13461 9472
rect 13495 9469 13507 9503
rect 13449 9463 13507 9469
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 13705 9503 13763 9509
rect 13705 9500 13717 9503
rect 13596 9472 13717 9500
rect 13596 9460 13602 9472
rect 13705 9469 13717 9472
rect 13751 9469 13763 9503
rect 13705 9463 13763 9469
rect 14734 9460 14740 9512
rect 14792 9500 14798 9512
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 14792 9472 15945 9500
rect 14792 9460 14798 9472
rect 15933 9469 15945 9472
rect 15979 9500 15991 9503
rect 16485 9503 16543 9509
rect 16485 9500 16497 9503
rect 15979 9472 16497 9500
rect 15979 9469 15991 9472
rect 15933 9463 15991 9469
rect 16485 9469 16497 9472
rect 16531 9469 16543 9503
rect 16485 9463 16543 9469
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 18196 9472 18521 9500
rect 18196 9460 18202 9472
rect 18509 9469 18521 9472
rect 18555 9500 18567 9503
rect 19518 9500 19524 9512
rect 18555 9472 19524 9500
rect 18555 9469 18567 9472
rect 18509 9463 18567 9469
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 21450 9460 21456 9512
rect 21508 9500 21514 9512
rect 21545 9503 21603 9509
rect 21545 9500 21557 9503
rect 21508 9472 21557 9500
rect 21508 9460 21514 9472
rect 21545 9469 21557 9472
rect 21591 9469 21603 9503
rect 21545 9463 21603 9469
rect 21726 9460 21732 9512
rect 21784 9460 21790 9512
rect 23474 9460 23480 9512
rect 23532 9500 23538 9512
rect 23661 9503 23719 9509
rect 23661 9500 23673 9503
rect 23532 9472 23673 9500
rect 23532 9460 23538 9472
rect 23661 9469 23673 9472
rect 23707 9469 23719 9503
rect 23768 9500 23796 9540
rect 23917 9503 23975 9509
rect 23917 9500 23929 9503
rect 23768 9472 23929 9500
rect 23661 9463 23719 9469
rect 23917 9469 23929 9472
rect 23963 9469 23975 9503
rect 23917 9463 23975 9469
rect 12989 9435 13047 9441
rect 12989 9401 13001 9435
rect 13035 9432 13047 9435
rect 14182 9432 14188 9444
rect 13035 9404 14188 9432
rect 13035 9401 13047 9404
rect 12989 9395 13047 9401
rect 14182 9392 14188 9404
rect 14240 9432 14246 9444
rect 18782 9441 18788 9444
rect 16577 9435 16635 9441
rect 16577 9432 16589 9435
rect 14240 9404 14872 9432
rect 14240 9392 14246 9404
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 13078 9364 13084 9376
rect 12483 9336 13084 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 14844 9373 14872 9404
rect 16040 9404 16589 9432
rect 16040 9376 16068 9404
rect 16577 9401 16589 9404
rect 16623 9401 16635 9435
rect 18776 9432 18788 9441
rect 18743 9404 18788 9432
rect 16577 9395 16635 9401
rect 18776 9395 18788 9404
rect 18782 9392 18788 9395
rect 18840 9392 18846 9444
rect 22097 9435 22155 9441
rect 22097 9432 22109 9435
rect 21192 9404 22109 9432
rect 14829 9367 14887 9373
rect 14829 9333 14841 9367
rect 14875 9333 14887 9367
rect 14829 9327 14887 9333
rect 15657 9367 15715 9373
rect 15657 9333 15669 9367
rect 15703 9364 15715 9367
rect 16022 9364 16028 9376
rect 15703 9336 16028 9364
rect 15703 9333 15715 9336
rect 15657 9327 15715 9333
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 16117 9367 16175 9373
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 16390 9364 16396 9376
rect 16163 9336 16396 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 18322 9364 18328 9376
rect 18283 9336 18328 9364
rect 18322 9324 18328 9336
rect 18380 9324 18386 9376
rect 20898 9324 20904 9376
rect 20956 9364 20962 9376
rect 21192 9373 21220 9404
rect 22097 9401 22109 9404
rect 22143 9401 22155 9435
rect 22097 9395 22155 9401
rect 21177 9367 21235 9373
rect 21177 9364 21189 9367
rect 20956 9336 21189 9364
rect 20956 9324 20962 9336
rect 21177 9333 21189 9336
rect 21223 9333 21235 9367
rect 21177 9327 21235 9333
rect 21266 9324 21272 9376
rect 21324 9364 21330 9376
rect 21637 9367 21695 9373
rect 21637 9364 21649 9367
rect 21324 9336 21649 9364
rect 21324 9324 21330 9336
rect 21637 9333 21649 9336
rect 21683 9333 21695 9367
rect 21637 9327 21695 9333
rect 21910 9324 21916 9376
rect 21968 9364 21974 9376
rect 22005 9367 22063 9373
rect 22005 9364 22017 9367
rect 21968 9336 22017 9364
rect 21968 9324 21974 9336
rect 22005 9333 22017 9336
rect 22051 9333 22063 9367
rect 25038 9364 25044 9376
rect 24999 9336 25044 9364
rect 22005 9327 22063 9333
rect 25038 9324 25044 9336
rect 25096 9324 25102 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 10505 9163 10563 9169
rect 10505 9129 10517 9163
rect 10551 9160 10563 9163
rect 10686 9160 10692 9172
rect 10551 9132 10692 9160
rect 10551 9129 10563 9132
rect 10505 9123 10563 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 13449 9163 13507 9169
rect 13449 9129 13461 9163
rect 13495 9160 13507 9163
rect 13538 9160 13544 9172
rect 13495 9132 13544 9160
rect 13495 9129 13507 9132
rect 13449 9123 13507 9129
rect 13538 9120 13544 9132
rect 13596 9160 13602 9172
rect 13998 9160 14004 9172
rect 13596 9132 14004 9160
rect 13596 9120 13602 9132
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14090 9120 14096 9172
rect 14148 9160 14154 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 14148 9132 14381 9160
rect 14148 9120 14154 9132
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 15286 9160 15292 9172
rect 15247 9132 15292 9160
rect 14369 9123 14427 9129
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 16666 9160 16672 9172
rect 16627 9132 16672 9160
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 18601 9163 18659 9169
rect 18601 9129 18613 9163
rect 18647 9160 18659 9163
rect 18782 9160 18788 9172
rect 18647 9132 18788 9160
rect 18647 9129 18659 9132
rect 18601 9123 18659 9129
rect 18782 9120 18788 9132
rect 18840 9160 18846 9172
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 18840 9132 19257 9160
rect 18840 9120 18846 9132
rect 19245 9129 19257 9132
rect 19291 9160 19303 9163
rect 20717 9163 20775 9169
rect 20717 9160 20729 9163
rect 19291 9132 20729 9160
rect 19291 9129 19303 9132
rect 19245 9123 19303 9129
rect 20717 9129 20729 9132
rect 20763 9160 20775 9163
rect 21542 9160 21548 9172
rect 20763 9132 21548 9160
rect 20763 9129 20775 9132
rect 20717 9123 20775 9129
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 23017 9163 23075 9169
rect 23017 9129 23029 9163
rect 23063 9160 23075 9163
rect 23382 9160 23388 9172
rect 23063 9132 23388 9160
rect 23063 9129 23075 9132
rect 23017 9123 23075 9129
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 24854 9160 24860 9172
rect 24815 9132 24860 9160
rect 24854 9120 24860 9132
rect 24912 9120 24918 9172
rect 21168 9095 21226 9101
rect 21168 9061 21180 9095
rect 21214 9092 21226 9095
rect 21266 9092 21272 9104
rect 21214 9064 21272 9092
rect 21214 9061 21226 9064
rect 21168 9055 21226 9061
rect 21266 9052 21272 9064
rect 21324 9092 21330 9104
rect 21818 9092 21824 9104
rect 21324 9064 21824 9092
rect 21324 9052 21330 9064
rect 21818 9052 21824 9064
rect 21876 9052 21882 9104
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10744 8996 10885 9024
rect 10744 8984 10750 8996
rect 10873 8993 10885 8996
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 12325 9027 12383 9033
rect 12325 9024 12337 9027
rect 12216 8996 12337 9024
rect 12216 8984 12222 8996
rect 12325 8993 12337 8996
rect 12371 8993 12383 9027
rect 12325 8987 12383 8993
rect 14826 8984 14832 9036
rect 14884 9024 14890 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 14884 8996 15669 9024
rect 14884 8984 14890 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 16850 8984 16856 9036
rect 16908 9024 16914 9036
rect 17477 9027 17535 9033
rect 17477 9024 17489 9027
rect 16908 8996 17489 9024
rect 16908 8984 16914 8996
rect 17477 8993 17489 8996
rect 17523 8993 17535 9027
rect 17477 8987 17535 8993
rect 20901 9027 20959 9033
rect 20901 8993 20913 9027
rect 20947 9024 20959 9027
rect 20990 9024 20996 9036
rect 20947 8996 20996 9024
rect 20947 8993 20959 8996
rect 20901 8987 20959 8993
rect 20990 8984 20996 8996
rect 21048 9024 21054 9036
rect 23744 9027 23802 9033
rect 21048 8996 23520 9024
rect 21048 8984 21054 8996
rect 23492 8968 23520 8996
rect 23744 8993 23756 9027
rect 23790 9024 23802 9027
rect 25038 9024 25044 9036
rect 23790 8996 25044 9024
rect 23790 8993 23802 8996
rect 23744 8987 23802 8993
rect 25038 8984 25044 8996
rect 25096 8984 25102 9036
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8956 10471 8959
rect 10778 8956 10784 8968
rect 10459 8928 10784 8956
rect 10459 8925 10471 8928
rect 10413 8919 10471 8925
rect 10778 8916 10784 8928
rect 10836 8956 10842 8968
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10836 8928 10977 8956
rect 10836 8916 10842 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 12069 8959 12127 8965
rect 11112 8928 11157 8956
rect 11112 8916 11118 8928
rect 12069 8925 12081 8959
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 15105 8959 15163 8965
rect 15105 8925 15117 8959
rect 15151 8956 15163 8959
rect 15746 8956 15752 8968
rect 15151 8928 15752 8956
rect 15151 8925 15163 8928
rect 15105 8919 15163 8925
rect 11514 8820 11520 8832
rect 11475 8792 11520 8820
rect 11514 8780 11520 8792
rect 11572 8780 11578 8832
rect 12084 8820 12112 8919
rect 15746 8916 15752 8928
rect 15804 8916 15810 8968
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8956 15991 8959
rect 17221 8959 17279 8965
rect 17221 8956 17233 8959
rect 15979 8928 16436 8956
rect 15979 8925 15991 8928
rect 15933 8919 15991 8925
rect 12802 8820 12808 8832
rect 12084 8792 12808 8820
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 16408 8829 16436 8928
rect 17052 8928 17233 8956
rect 17052 8832 17080 8928
rect 17221 8925 17233 8928
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8956 19855 8959
rect 20622 8956 20628 8968
rect 19843 8928 20628 8956
rect 19843 8925 19855 8928
rect 19797 8919 19855 8925
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 23474 8956 23480 8968
rect 23387 8928 23480 8956
rect 23474 8916 23480 8928
rect 23532 8916 23538 8968
rect 19518 8848 19524 8900
rect 19576 8888 19582 8900
rect 20257 8891 20315 8897
rect 20257 8888 20269 8891
rect 19576 8860 20269 8888
rect 19576 8848 19582 8860
rect 20257 8857 20269 8860
rect 20303 8857 20315 8891
rect 20257 8851 20315 8857
rect 16393 8823 16451 8829
rect 16393 8789 16405 8823
rect 16439 8820 16451 8823
rect 16482 8820 16488 8832
rect 16439 8792 16488 8820
rect 16439 8789 16451 8792
rect 16393 8783 16451 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 17034 8820 17040 8832
rect 16995 8792 17040 8820
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 19705 8823 19763 8829
rect 19705 8789 19717 8823
rect 19751 8820 19763 8823
rect 19794 8820 19800 8832
rect 19751 8792 19800 8820
rect 19751 8789 19763 8792
rect 19705 8783 19763 8789
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 22278 8820 22284 8832
rect 22239 8792 22284 8820
rect 22278 8780 22284 8792
rect 22336 8780 22342 8832
rect 23385 8823 23443 8829
rect 23385 8789 23397 8823
rect 23431 8820 23443 8823
rect 23492 8820 23520 8916
rect 24854 8820 24860 8832
rect 23431 8792 24860 8820
rect 23431 8789 23443 8792
rect 23385 8783 23443 8789
rect 24854 8780 24860 8792
rect 24912 8820 24918 8832
rect 25314 8820 25320 8832
rect 24912 8792 25320 8820
rect 24912 8780 24918 8792
rect 25314 8780 25320 8792
rect 25372 8780 25378 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 10778 8616 10784 8628
rect 10739 8588 10784 8616
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 13265 8619 13323 8625
rect 13265 8616 13277 8619
rect 13228 8588 13277 8616
rect 13228 8576 13234 8588
rect 13265 8585 13277 8588
rect 13311 8585 13323 8619
rect 13265 8579 13323 8585
rect 13449 8619 13507 8625
rect 13449 8585 13461 8619
rect 13495 8616 13507 8619
rect 14090 8616 14096 8628
rect 13495 8588 14096 8616
rect 13495 8585 13507 8588
rect 13449 8579 13507 8585
rect 9953 8551 10011 8557
rect 9953 8517 9965 8551
rect 9999 8548 10011 8551
rect 11054 8548 11060 8560
rect 9999 8520 11060 8548
rect 9999 8517 10011 8520
rect 9953 8511 10011 8517
rect 11054 8508 11060 8520
rect 11112 8548 11118 8560
rect 12069 8551 12127 8557
rect 12069 8548 12081 8551
rect 11112 8520 12081 8548
rect 11112 8508 11118 8520
rect 12069 8517 12081 8520
rect 12115 8548 12127 8551
rect 12158 8548 12164 8560
rect 12115 8520 12164 8548
rect 12115 8517 12127 8520
rect 12069 8511 12127 8517
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 10594 8480 10600 8492
rect 10555 8452 10600 8480
rect 10594 8440 10600 8452
rect 10652 8480 10658 8492
rect 11425 8483 11483 8489
rect 10652 8452 11192 8480
rect 10652 8440 10658 8452
rect 11164 8421 11192 8452
rect 11425 8449 11437 8483
rect 11471 8480 11483 8483
rect 11514 8480 11520 8492
rect 11471 8452 11520 8480
rect 11471 8449 11483 8452
rect 11425 8443 11483 8449
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 12526 8412 12532 8424
rect 11149 8375 11207 8381
rect 11256 8384 12532 8412
rect 11256 8353 11284 8384
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 13280 8412 13308 8579
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 16850 8616 16856 8628
rect 16811 8588 16856 8616
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 19150 8616 19156 8628
rect 19111 8588 19156 8616
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 19794 8576 19800 8628
rect 19852 8616 19858 8628
rect 21266 8616 21272 8628
rect 19852 8588 20852 8616
rect 21227 8588 21272 8616
rect 19852 8576 19858 8588
rect 13354 8508 13360 8560
rect 13412 8548 13418 8560
rect 14826 8548 14832 8560
rect 13412 8520 14136 8548
rect 14787 8520 14832 8548
rect 13412 8508 13418 8520
rect 13998 8480 14004 8492
rect 13959 8452 14004 8480
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 13817 8415 13875 8421
rect 13817 8412 13829 8415
rect 13280 8384 13829 8412
rect 13817 8381 13829 8384
rect 13863 8381 13875 8415
rect 13817 8375 13875 8381
rect 13909 8415 13967 8421
rect 13909 8381 13921 8415
rect 13955 8412 13967 8415
rect 14108 8412 14136 8520
rect 14826 8508 14832 8520
rect 14884 8508 14890 8560
rect 17862 8508 17868 8560
rect 17920 8548 17926 8560
rect 18049 8551 18107 8557
rect 18049 8548 18061 8551
rect 17920 8520 18061 8548
rect 17920 8508 17926 8520
rect 18049 8517 18061 8520
rect 18095 8517 18107 8551
rect 18049 8511 18107 8517
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8480 14611 8483
rect 14599 8452 15608 8480
rect 14599 8449 14611 8452
rect 14553 8443 14611 8449
rect 15102 8412 15108 8424
rect 13955 8384 15108 8412
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 15197 8415 15255 8421
rect 15197 8381 15209 8415
rect 15243 8381 15255 8415
rect 15197 8375 15255 8381
rect 10321 8347 10379 8353
rect 10321 8313 10333 8347
rect 10367 8344 10379 8347
rect 11241 8347 11299 8353
rect 11241 8344 11253 8347
rect 10367 8316 11253 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 11241 8313 11253 8316
rect 11287 8313 11299 8347
rect 11241 8307 11299 8313
rect 12434 8304 12440 8356
rect 12492 8344 12498 8356
rect 12989 8347 13047 8353
rect 12492 8316 12537 8344
rect 12492 8304 12498 8316
rect 12989 8313 13001 8347
rect 13035 8344 13047 8347
rect 13354 8344 13360 8356
rect 13035 8316 13360 8344
rect 13035 8313 13047 8316
rect 12989 8307 13047 8313
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 13446 8304 13452 8356
rect 13504 8344 13510 8356
rect 15212 8344 15240 8375
rect 15286 8372 15292 8424
rect 15344 8412 15350 8424
rect 15473 8415 15531 8421
rect 15473 8412 15485 8415
rect 15344 8384 15485 8412
rect 15344 8372 15350 8384
rect 15473 8381 15485 8384
rect 15519 8381 15531 8415
rect 15580 8412 15608 8452
rect 18506 8440 18512 8492
rect 18564 8480 18570 8492
rect 18693 8483 18751 8489
rect 18693 8480 18705 8483
rect 18564 8452 18705 8480
rect 18564 8440 18570 8452
rect 18693 8449 18705 8452
rect 18739 8480 18751 8483
rect 19168 8480 19196 8576
rect 20824 8548 20852 8588
rect 21266 8576 21272 8588
rect 21324 8616 21330 8628
rect 21821 8619 21879 8625
rect 21821 8616 21833 8619
rect 21324 8588 21833 8616
rect 21324 8576 21330 8588
rect 21821 8585 21833 8588
rect 21867 8585 21879 8619
rect 21821 8579 21879 8585
rect 23109 8619 23167 8625
rect 23109 8585 23121 8619
rect 23155 8616 23167 8619
rect 23198 8616 23204 8628
rect 23155 8588 23204 8616
rect 23155 8585 23167 8588
rect 23109 8579 23167 8585
rect 21450 8548 21456 8560
rect 20824 8520 21456 8548
rect 21450 8508 21456 8520
rect 21508 8548 21514 8560
rect 22189 8551 22247 8557
rect 22189 8548 22201 8551
rect 21508 8520 22201 8548
rect 21508 8508 21514 8520
rect 22189 8517 22201 8520
rect 22235 8517 22247 8551
rect 22646 8548 22652 8560
rect 22607 8520 22652 8548
rect 22189 8511 22247 8517
rect 22646 8508 22652 8520
rect 22704 8508 22710 8560
rect 18739 8452 19196 8480
rect 19521 8483 19579 8489
rect 18739 8449 18751 8452
rect 18693 8443 18751 8449
rect 19521 8449 19533 8483
rect 19567 8480 19579 8483
rect 19567 8452 20024 8480
rect 19567 8449 19579 8452
rect 19521 8443 19579 8449
rect 15740 8415 15798 8421
rect 15740 8412 15752 8415
rect 15580 8384 15752 8412
rect 15473 8375 15531 8381
rect 15740 8381 15752 8384
rect 15786 8412 15798 8415
rect 16482 8412 16488 8424
rect 15786 8384 16488 8412
rect 15786 8381 15798 8384
rect 15740 8375 15798 8381
rect 16482 8372 16488 8384
rect 16540 8372 16546 8424
rect 17497 8415 17555 8421
rect 17497 8381 17509 8415
rect 17543 8412 17555 8415
rect 19794 8412 19800 8424
rect 17543 8384 18552 8412
rect 19755 8384 19800 8412
rect 17543 8381 17555 8384
rect 17497 8375 17555 8381
rect 16390 8344 16396 8356
rect 13504 8316 15056 8344
rect 13504 8304 13510 8316
rect 15028 8285 15056 8316
rect 15120 8316 16396 8344
rect 15120 8288 15148 8316
rect 16390 8304 16396 8316
rect 16448 8304 16454 8356
rect 17865 8347 17923 8353
rect 17865 8313 17877 8347
rect 17911 8344 17923 8347
rect 17911 8316 18460 8344
rect 17911 8313 17923 8316
rect 17865 8307 17923 8313
rect 18432 8288 18460 8316
rect 15013 8279 15071 8285
rect 15013 8245 15025 8279
rect 15059 8245 15071 8279
rect 15013 8239 15071 8245
rect 15102 8236 15108 8288
rect 15160 8236 15166 8288
rect 18414 8276 18420 8288
rect 18375 8248 18420 8276
rect 18414 8236 18420 8248
rect 18472 8236 18478 8288
rect 18524 8285 18552 8384
rect 19794 8372 19800 8384
rect 19852 8372 19858 8424
rect 19889 8415 19947 8421
rect 19889 8381 19901 8415
rect 19935 8381 19947 8415
rect 19889 8375 19947 8381
rect 19904 8344 19932 8375
rect 19996 8356 20024 8452
rect 22465 8415 22523 8421
rect 22465 8381 22477 8415
rect 22511 8412 22523 8415
rect 23124 8412 23152 8579
rect 23198 8576 23204 8588
rect 23256 8576 23262 8628
rect 24765 8619 24823 8625
rect 24765 8585 24777 8619
rect 24811 8616 24823 8619
rect 25038 8616 25044 8628
rect 24811 8588 25044 8616
rect 24811 8585 24823 8588
rect 24765 8579 24823 8585
rect 23474 8508 23480 8560
rect 23532 8548 23538 8560
rect 23661 8551 23719 8557
rect 23661 8548 23673 8551
rect 23532 8520 23673 8548
rect 23532 8508 23538 8520
rect 23661 8517 23673 8520
rect 23707 8517 23719 8551
rect 23661 8511 23719 8517
rect 24118 8440 24124 8492
rect 24176 8480 24182 8492
rect 24305 8483 24363 8489
rect 24305 8480 24317 8483
rect 24176 8452 24317 8480
rect 24176 8440 24182 8452
rect 24305 8449 24317 8452
rect 24351 8480 24363 8483
rect 24780 8480 24808 8579
rect 25038 8576 25044 8588
rect 25096 8576 25102 8628
rect 25406 8480 25412 8492
rect 24351 8452 24808 8480
rect 25367 8452 25412 8480
rect 24351 8449 24363 8452
rect 24305 8443 24363 8449
rect 25406 8440 25412 8452
rect 25464 8440 25470 8492
rect 22511 8384 23152 8412
rect 23477 8415 23535 8421
rect 22511 8381 22523 8384
rect 22465 8375 22523 8381
rect 23477 8381 23489 8415
rect 23523 8412 23535 8415
rect 23934 8412 23940 8424
rect 23523 8384 23940 8412
rect 23523 8381 23535 8384
rect 23477 8375 23535 8381
rect 23934 8372 23940 8384
rect 23992 8412 23998 8424
rect 24029 8415 24087 8421
rect 24029 8412 24041 8415
rect 23992 8384 24041 8412
rect 23992 8372 23998 8384
rect 24029 8381 24041 8384
rect 24075 8381 24087 8415
rect 25222 8412 25228 8424
rect 25183 8384 25228 8412
rect 24029 8375 24087 8381
rect 25222 8372 25228 8384
rect 25280 8412 25286 8424
rect 25961 8415 26019 8421
rect 25961 8412 25973 8415
rect 25280 8384 25973 8412
rect 25280 8372 25286 8384
rect 25961 8381 25973 8384
rect 26007 8381 26019 8415
rect 25961 8375 26019 8381
rect 19628 8316 19932 8344
rect 18509 8279 18567 8285
rect 18509 8245 18521 8279
rect 18555 8276 18567 8279
rect 18598 8276 18604 8288
rect 18555 8248 18604 8276
rect 18555 8245 18567 8248
rect 18509 8239 18567 8245
rect 18598 8236 18604 8248
rect 18656 8236 18662 8288
rect 19518 8236 19524 8288
rect 19576 8276 19582 8288
rect 19628 8285 19656 8316
rect 19978 8304 19984 8356
rect 20036 8344 20042 8356
rect 20134 8347 20192 8353
rect 20134 8344 20146 8347
rect 20036 8316 20146 8344
rect 20036 8304 20042 8316
rect 20134 8313 20146 8316
rect 20180 8313 20192 8347
rect 20134 8307 20192 8313
rect 19613 8279 19671 8285
rect 19613 8276 19625 8279
rect 19576 8248 19625 8276
rect 19576 8236 19582 8248
rect 19613 8245 19625 8248
rect 19659 8245 19671 8279
rect 19613 8239 19671 8245
rect 24121 8279 24179 8285
rect 24121 8245 24133 8279
rect 24167 8276 24179 8279
rect 24210 8276 24216 8288
rect 24167 8248 24216 8276
rect 24167 8245 24179 8248
rect 24121 8239 24179 8245
rect 24210 8236 24216 8248
rect 24268 8236 24274 8288
rect 24854 8236 24860 8288
rect 24912 8276 24918 8288
rect 25133 8279 25191 8285
rect 25133 8276 25145 8279
rect 24912 8248 25145 8276
rect 24912 8236 24918 8248
rect 25133 8245 25145 8248
rect 25179 8276 25191 8279
rect 25682 8276 25688 8288
rect 25179 8248 25688 8276
rect 25179 8245 25191 8248
rect 25133 8239 25191 8245
rect 25682 8236 25688 8248
rect 25740 8236 25746 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 9769 8075 9827 8081
rect 9769 8041 9781 8075
rect 9815 8072 9827 8075
rect 10778 8072 10784 8084
rect 9815 8044 10784 8072
rect 9815 8041 9827 8044
rect 9769 8035 9827 8041
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 12158 8072 12164 8084
rect 12119 8044 12164 8072
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 13262 8072 13268 8084
rect 13223 8044 13268 8072
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 16574 8032 16580 8084
rect 16632 8072 16638 8084
rect 16669 8075 16727 8081
rect 16669 8072 16681 8075
rect 16632 8044 16681 8072
rect 16632 8032 16638 8044
rect 16669 8041 16681 8044
rect 16715 8041 16727 8075
rect 16669 8035 16727 8041
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 17221 8075 17279 8081
rect 17221 8072 17233 8075
rect 16908 8044 17233 8072
rect 16908 8032 16914 8044
rect 17221 8041 17233 8044
rect 17267 8041 17279 8075
rect 17221 8035 17279 8041
rect 19153 8075 19211 8081
rect 19153 8041 19165 8075
rect 19199 8072 19211 8075
rect 19242 8072 19248 8084
rect 19199 8044 19248 8072
rect 19199 8041 19211 8044
rect 19153 8035 19211 8041
rect 19242 8032 19248 8044
rect 19300 8072 19306 8084
rect 19426 8072 19432 8084
rect 19300 8044 19432 8072
rect 19300 8032 19306 8044
rect 19426 8032 19432 8044
rect 19484 8032 19490 8084
rect 21085 8075 21143 8081
rect 21085 8041 21097 8075
rect 21131 8072 21143 8075
rect 22002 8072 22008 8084
rect 21131 8044 22008 8072
rect 21131 8041 21143 8044
rect 21085 8035 21143 8041
rect 22002 8032 22008 8044
rect 22060 8032 22066 8084
rect 22554 8032 22560 8084
rect 22612 8072 22618 8084
rect 23014 8072 23020 8084
rect 22612 8044 23020 8072
rect 22612 8032 22618 8044
rect 23014 8032 23020 8044
rect 23072 8032 23078 8084
rect 23109 8075 23167 8081
rect 23109 8041 23121 8075
rect 23155 8072 23167 8075
rect 23382 8072 23388 8084
rect 23155 8044 23388 8072
rect 23155 8041 23167 8044
rect 23109 8035 23167 8041
rect 23382 8032 23388 8044
rect 23440 8032 23446 8084
rect 24118 8072 24124 8084
rect 24079 8044 24124 8072
rect 24118 8032 24124 8044
rect 24176 8032 24182 8084
rect 10597 8007 10655 8013
rect 10597 7973 10609 8007
rect 10643 8004 10655 8007
rect 10686 8004 10692 8016
rect 10643 7976 10692 8004
rect 10643 7973 10655 7976
rect 10597 7967 10655 7973
rect 10686 7964 10692 7976
rect 10744 7964 10750 8016
rect 11048 8007 11106 8013
rect 11048 7973 11060 8007
rect 11094 8004 11106 8007
rect 11514 8004 11520 8016
rect 11094 7976 11520 8004
rect 11094 7973 11106 7976
rect 11048 7967 11106 7973
rect 11514 7964 11520 7976
rect 11572 7964 11578 8016
rect 13078 7964 13084 8016
rect 13136 8004 13142 8016
rect 13633 8007 13691 8013
rect 13633 8004 13645 8007
rect 13136 7976 13645 8004
rect 13136 7964 13142 7976
rect 13633 7973 13645 7976
rect 13679 7973 13691 8007
rect 13633 7967 13691 7973
rect 18509 8007 18567 8013
rect 18509 7973 18521 8007
rect 18555 8004 18567 8007
rect 18598 8004 18604 8016
rect 18555 7976 18604 8004
rect 18555 7973 18567 7976
rect 18509 7967 18567 7973
rect 18598 7964 18604 7976
rect 18656 7964 18662 8016
rect 20349 8007 20407 8013
rect 20349 7973 20361 8007
rect 20395 8004 20407 8007
rect 21545 8007 21603 8013
rect 21545 8004 21557 8007
rect 20395 7976 21557 8004
rect 20395 7973 20407 7976
rect 20349 7967 20407 7973
rect 21545 7973 21557 7976
rect 21591 8004 21603 8007
rect 21634 8004 21640 8016
rect 21591 7976 21640 8004
rect 21591 7973 21603 7976
rect 21545 7967 21603 7973
rect 21634 7964 21640 7976
rect 21692 7964 21698 8016
rect 23753 8007 23811 8013
rect 23753 7973 23765 8007
rect 23799 8004 23811 8007
rect 24210 8004 24216 8016
rect 23799 7976 24216 8004
rect 23799 7973 23811 7976
rect 23753 7967 23811 7973
rect 24210 7964 24216 7976
rect 24268 7964 24274 8016
rect 24673 8007 24731 8013
rect 24673 7973 24685 8007
rect 24719 8004 24731 8007
rect 24762 8004 24768 8016
rect 24719 7976 24768 8004
rect 24719 7973 24731 7976
rect 24673 7967 24731 7973
rect 24762 7964 24768 7976
rect 24820 7964 24826 8016
rect 15102 7936 15108 7948
rect 14752 7908 15108 7936
rect 10778 7868 10784 7880
rect 10739 7840 10784 7868
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 13722 7868 13728 7880
rect 13683 7840 13728 7868
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 13817 7871 13875 7877
rect 13817 7837 13829 7871
rect 13863 7837 13875 7871
rect 13817 7831 13875 7837
rect 12802 7800 12808 7812
rect 12715 7772 12808 7800
rect 12802 7760 12808 7772
rect 12860 7800 12866 7812
rect 13446 7800 13452 7812
rect 12860 7772 13452 7800
rect 12860 7760 12866 7772
rect 13446 7760 13452 7772
rect 13504 7760 13510 7812
rect 13538 7760 13544 7812
rect 13596 7800 13602 7812
rect 13832 7800 13860 7831
rect 13596 7772 13860 7800
rect 13596 7760 13602 7772
rect 13170 7732 13176 7744
rect 13131 7704 13176 7732
rect 13170 7692 13176 7704
rect 13228 7692 13234 7744
rect 14642 7692 14648 7744
rect 14700 7732 14706 7744
rect 14752 7741 14780 7908
rect 15102 7896 15108 7908
rect 15160 7896 15166 7948
rect 15556 7939 15614 7945
rect 15556 7905 15568 7939
rect 15602 7936 15614 7939
rect 16390 7936 16396 7948
rect 15602 7908 16396 7936
rect 15602 7905 15614 7908
rect 15556 7899 15614 7905
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 18414 7936 18420 7948
rect 18375 7908 18420 7936
rect 18414 7896 18420 7908
rect 18472 7896 18478 7948
rect 19705 7939 19763 7945
rect 19705 7905 19717 7939
rect 19751 7936 19763 7939
rect 21453 7939 21511 7945
rect 19751 7908 20392 7936
rect 19751 7905 19763 7908
rect 19705 7899 19763 7905
rect 20364 7880 20392 7908
rect 21453 7905 21465 7939
rect 21499 7936 21511 7939
rect 21499 7908 22324 7936
rect 21499 7905 21511 7908
rect 21453 7899 21511 7905
rect 15286 7868 15292 7880
rect 14936 7840 15292 7868
rect 14737 7735 14795 7741
rect 14737 7732 14749 7735
rect 14700 7704 14749 7732
rect 14700 7692 14706 7704
rect 14737 7701 14749 7704
rect 14783 7701 14795 7735
rect 14737 7695 14795 7701
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 14936 7741 14964 7840
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 17678 7828 17684 7880
rect 17736 7868 17742 7880
rect 18601 7871 18659 7877
rect 18601 7868 18613 7871
rect 17736 7840 18613 7868
rect 17736 7828 17742 7840
rect 18601 7837 18613 7840
rect 18647 7837 18659 7871
rect 18601 7831 18659 7837
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 21726 7868 21732 7880
rect 21687 7840 21732 7868
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 19610 7760 19616 7812
rect 19668 7800 19674 7812
rect 20898 7800 20904 7812
rect 19668 7772 20904 7800
rect 19668 7760 19674 7772
rect 20898 7760 20904 7772
rect 20956 7760 20962 7812
rect 22296 7800 22324 7908
rect 23474 7896 23480 7948
rect 23532 7936 23538 7948
rect 24581 7939 24639 7945
rect 24581 7936 24593 7939
rect 23532 7908 24593 7936
rect 23532 7896 23538 7908
rect 24581 7905 24593 7908
rect 24627 7905 24639 7939
rect 24581 7899 24639 7905
rect 22370 7828 22376 7880
rect 22428 7868 22434 7880
rect 23201 7871 23259 7877
rect 23201 7868 23213 7871
rect 22428 7840 23213 7868
rect 22428 7828 22434 7840
rect 23201 7837 23213 7840
rect 23247 7837 23259 7871
rect 23201 7831 23259 7837
rect 24210 7828 24216 7880
rect 24268 7868 24274 7880
rect 24765 7871 24823 7877
rect 24765 7868 24777 7871
rect 24268 7840 24777 7868
rect 24268 7828 24274 7840
rect 24765 7837 24777 7840
rect 24811 7837 24823 7871
rect 24765 7831 24823 7837
rect 22557 7803 22615 7809
rect 22557 7800 22569 7803
rect 22296 7772 22569 7800
rect 22557 7769 22569 7772
rect 22603 7800 22615 7803
rect 23290 7800 23296 7812
rect 22603 7772 23296 7800
rect 22603 7769 22615 7772
rect 22557 7763 22615 7769
rect 23290 7760 23296 7772
rect 23348 7760 23354 7812
rect 14921 7735 14979 7741
rect 14921 7732 14933 7735
rect 14884 7704 14933 7732
rect 14884 7692 14890 7704
rect 14921 7701 14933 7704
rect 14967 7732 14979 7735
rect 17034 7732 17040 7744
rect 14967 7704 17040 7732
rect 14967 7701 14979 7704
rect 14921 7695 14979 7701
rect 17034 7692 17040 7704
rect 17092 7732 17098 7744
rect 17589 7735 17647 7741
rect 17589 7732 17601 7735
rect 17092 7704 17601 7732
rect 17092 7692 17098 7704
rect 17589 7701 17601 7704
rect 17635 7701 17647 7735
rect 17589 7695 17647 7701
rect 17954 7692 17960 7744
rect 18012 7732 18018 7744
rect 18049 7735 18107 7741
rect 18049 7732 18061 7735
rect 18012 7704 18061 7732
rect 18012 7692 18018 7704
rect 18049 7701 18061 7704
rect 18095 7701 18107 7735
rect 19426 7732 19432 7744
rect 19387 7704 19432 7732
rect 18049 7695 18107 7701
rect 19426 7692 19432 7704
rect 19484 7692 19490 7744
rect 19889 7735 19947 7741
rect 19889 7701 19901 7735
rect 19935 7732 19947 7735
rect 20162 7732 20168 7744
rect 19935 7704 20168 7732
rect 19935 7701 19947 7704
rect 19889 7695 19947 7701
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 20714 7732 20720 7744
rect 20675 7704 20720 7732
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 22094 7692 22100 7744
rect 22152 7732 22158 7744
rect 22646 7732 22652 7744
rect 22152 7704 22197 7732
rect 22607 7704 22652 7732
rect 22152 7692 22158 7704
rect 22646 7692 22652 7704
rect 22704 7692 22710 7744
rect 24118 7692 24124 7744
rect 24176 7732 24182 7744
rect 24213 7735 24271 7741
rect 24213 7732 24225 7735
rect 24176 7704 24225 7732
rect 24176 7692 24182 7704
rect 24213 7701 24225 7704
rect 24259 7732 24271 7735
rect 25225 7735 25283 7741
rect 25225 7732 25237 7735
rect 24259 7704 25237 7732
rect 24259 7701 24271 7704
rect 24213 7695 24271 7701
rect 25225 7701 25237 7704
rect 25271 7701 25283 7735
rect 25225 7695 25283 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 11241 7531 11299 7537
rect 11241 7528 11253 7531
rect 11020 7500 11253 7528
rect 11020 7488 11026 7500
rect 11241 7497 11253 7500
rect 11287 7528 11299 7531
rect 11514 7528 11520 7540
rect 11287 7500 11520 7528
rect 11287 7497 11299 7500
rect 11241 7491 11299 7497
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 13078 7528 13084 7540
rect 13039 7500 13084 7528
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 14826 7528 14832 7540
rect 13228 7500 14832 7528
rect 13228 7488 13234 7500
rect 13280 7401 13308 7500
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 15746 7528 15752 7540
rect 15707 7500 15752 7528
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 21358 7528 21364 7540
rect 21319 7500 21364 7528
rect 21358 7488 21364 7500
rect 21416 7488 21422 7540
rect 22370 7488 22376 7540
rect 22428 7528 22434 7540
rect 22649 7531 22707 7537
rect 22649 7528 22661 7531
rect 22428 7500 22661 7528
rect 22428 7488 22434 7500
rect 22649 7497 22661 7500
rect 22695 7497 22707 7531
rect 23014 7528 23020 7540
rect 22975 7500 23020 7528
rect 22649 7491 22707 7497
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 23658 7528 23664 7540
rect 23619 7500 23664 7528
rect 23658 7488 23664 7500
rect 23716 7488 23722 7540
rect 23842 7488 23848 7540
rect 23900 7528 23906 7540
rect 24210 7528 24216 7540
rect 23900 7500 24216 7528
rect 23900 7488 23906 7500
rect 24210 7488 24216 7500
rect 24268 7528 24274 7540
rect 24673 7531 24731 7537
rect 24673 7528 24685 7531
rect 24268 7500 24685 7528
rect 24268 7488 24274 7500
rect 24673 7497 24685 7500
rect 24719 7497 24731 7531
rect 24673 7491 24731 7497
rect 26234 7488 26240 7540
rect 26292 7528 26298 7540
rect 26878 7528 26884 7540
rect 26292 7500 26884 7528
rect 26292 7488 26298 7500
rect 26878 7488 26884 7500
rect 26936 7488 26942 7540
rect 20901 7463 20959 7469
rect 20901 7429 20913 7463
rect 20947 7460 20959 7463
rect 21450 7460 21456 7472
rect 20947 7432 21456 7460
rect 20947 7429 20959 7432
rect 20901 7423 20959 7429
rect 21450 7420 21456 7432
rect 21508 7460 21514 7472
rect 21726 7460 21732 7472
rect 21508 7432 21732 7460
rect 21508 7420 21514 7432
rect 21726 7420 21732 7432
rect 21784 7420 21790 7472
rect 23477 7463 23535 7469
rect 23477 7429 23489 7463
rect 23523 7460 23535 7463
rect 23523 7432 24256 7460
rect 23523 7429 23535 7432
rect 23477 7423 23535 7429
rect 24228 7404 24256 7432
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7361 13323 7395
rect 16390 7392 16396 7404
rect 16303 7364 16396 7392
rect 13265 7355 13323 7361
rect 16390 7352 16396 7364
rect 16448 7392 16454 7404
rect 16761 7395 16819 7401
rect 16761 7392 16773 7395
rect 16448 7364 16773 7392
rect 16448 7352 16454 7364
rect 16761 7361 16773 7364
rect 16807 7361 16819 7395
rect 21266 7392 21272 7404
rect 21179 7364 21272 7392
rect 16761 7355 16819 7361
rect 21266 7352 21272 7364
rect 21324 7392 21330 7404
rect 21913 7395 21971 7401
rect 21913 7392 21925 7395
rect 21324 7364 21925 7392
rect 21324 7352 21330 7364
rect 21913 7361 21925 7364
rect 21959 7361 21971 7395
rect 24118 7392 24124 7404
rect 24079 7364 24124 7392
rect 21913 7355 21971 7361
rect 24118 7352 24124 7364
rect 24176 7352 24182 7404
rect 24210 7352 24216 7404
rect 24268 7392 24274 7404
rect 26329 7395 26387 7401
rect 26329 7392 26341 7395
rect 24268 7364 24361 7392
rect 24688 7364 26341 7392
rect 24268 7352 24274 7364
rect 13538 7333 13544 7336
rect 9861 7327 9919 7333
rect 9861 7324 9873 7327
rect 9324 7296 9873 7324
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 9324 7197 9352 7296
rect 9861 7293 9873 7296
rect 9907 7293 9919 7327
rect 13532 7324 13544 7333
rect 9861 7287 9919 7293
rect 13372 7296 13544 7324
rect 9769 7259 9827 7265
rect 9769 7225 9781 7259
rect 9815 7256 9827 7259
rect 10042 7256 10048 7268
rect 9815 7228 10048 7256
rect 9815 7225 9827 7228
rect 9769 7219 9827 7225
rect 10042 7216 10048 7228
rect 10100 7265 10106 7268
rect 10100 7259 10164 7265
rect 10100 7225 10118 7259
rect 10152 7225 10164 7259
rect 10100 7219 10164 7225
rect 12805 7259 12863 7265
rect 12805 7225 12817 7259
rect 12851 7256 12863 7259
rect 13372 7256 13400 7296
rect 13532 7287 13544 7296
rect 13538 7284 13544 7287
rect 13596 7284 13602 7336
rect 15286 7324 15292 7336
rect 15199 7296 15292 7324
rect 15286 7284 15292 7296
rect 15344 7324 15350 7336
rect 15344 7296 16252 7324
rect 15344 7284 15350 7296
rect 16117 7259 16175 7265
rect 16117 7256 16129 7259
rect 12851 7228 13400 7256
rect 15580 7228 16129 7256
rect 12851 7225 12863 7228
rect 12805 7219 12863 7225
rect 10100 7216 10106 7219
rect 15580 7200 15608 7228
rect 16117 7225 16129 7228
rect 16163 7225 16175 7259
rect 16117 7219 16175 7225
rect 9309 7191 9367 7197
rect 9309 7188 9321 7191
rect 9088 7160 9321 7188
rect 9088 7148 9094 7160
rect 9309 7157 9321 7160
rect 9355 7157 9367 7191
rect 14642 7188 14648 7200
rect 14603 7160 14648 7188
rect 9309 7151 9367 7157
rect 14642 7148 14648 7160
rect 14700 7148 14706 7200
rect 15562 7188 15568 7200
rect 15523 7160 15568 7188
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 16224 7197 16252 7296
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 18877 7327 18935 7333
rect 18877 7324 18889 7327
rect 18104 7296 18889 7324
rect 18104 7284 18110 7296
rect 18877 7293 18889 7296
rect 18923 7324 18935 7327
rect 19426 7324 19432 7336
rect 18923 7296 19432 7324
rect 18923 7293 18935 7296
rect 18877 7287 18935 7293
rect 19426 7284 19432 7296
rect 19484 7284 19490 7336
rect 20714 7284 20720 7336
rect 20772 7324 20778 7336
rect 21729 7327 21787 7333
rect 21729 7324 21741 7327
rect 20772 7296 21741 7324
rect 20772 7284 20778 7296
rect 21729 7293 21741 7296
rect 21775 7293 21787 7327
rect 21729 7287 21787 7293
rect 23658 7284 23664 7336
rect 23716 7324 23722 7336
rect 24029 7327 24087 7333
rect 24029 7324 24041 7327
rect 23716 7296 24041 7324
rect 23716 7284 23722 7296
rect 24029 7293 24041 7296
rect 24075 7324 24087 7327
rect 24688 7324 24716 7364
rect 26329 7361 26341 7364
rect 26375 7361 26387 7395
rect 26329 7355 26387 7361
rect 25222 7324 25228 7336
rect 24075 7296 24716 7324
rect 25183 7296 25228 7324
rect 24075 7293 24087 7296
rect 24029 7287 24087 7293
rect 25222 7284 25228 7296
rect 25280 7324 25286 7336
rect 25961 7327 26019 7333
rect 25961 7324 25973 7327
rect 25280 7296 25973 7324
rect 25280 7284 25286 7296
rect 25961 7293 25973 7296
rect 26007 7293 26019 7327
rect 25961 7287 26019 7293
rect 18325 7259 18383 7265
rect 18325 7225 18337 7259
rect 18371 7256 18383 7259
rect 18414 7256 18420 7268
rect 18371 7228 18420 7256
rect 18371 7225 18383 7228
rect 18325 7219 18383 7225
rect 18414 7216 18420 7228
rect 18472 7256 18478 7268
rect 19144 7259 19202 7265
rect 18472 7228 19104 7256
rect 18472 7216 18478 7228
rect 16209 7191 16267 7197
rect 16209 7157 16221 7191
rect 16255 7188 16267 7191
rect 16298 7188 16304 7200
rect 16255 7160 16304 7188
rect 16255 7157 16267 7160
rect 16209 7151 16267 7157
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 17313 7191 17371 7197
rect 17313 7157 17325 7191
rect 17359 7188 17371 7191
rect 17586 7188 17592 7200
rect 17359 7160 17592 7188
rect 17359 7157 17371 7160
rect 17313 7151 17371 7157
rect 17586 7148 17592 7160
rect 17644 7148 17650 7200
rect 17678 7148 17684 7200
rect 17736 7188 17742 7200
rect 17773 7191 17831 7197
rect 17773 7188 17785 7191
rect 17736 7160 17785 7188
rect 17736 7148 17742 7160
rect 17773 7157 17785 7160
rect 17819 7157 17831 7191
rect 18598 7188 18604 7200
rect 18559 7160 18604 7188
rect 17773 7151 17831 7157
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 19076 7188 19104 7228
rect 19144 7225 19156 7259
rect 19190 7256 19202 7259
rect 19242 7256 19248 7268
rect 19190 7228 19248 7256
rect 19190 7225 19202 7228
rect 19144 7219 19202 7225
rect 19242 7216 19248 7228
rect 19300 7216 19306 7268
rect 20530 7216 20536 7268
rect 20588 7256 20594 7268
rect 21821 7259 21879 7265
rect 21821 7256 21833 7259
rect 20588 7228 21833 7256
rect 20588 7216 20594 7228
rect 21821 7225 21833 7228
rect 21867 7256 21879 7259
rect 22094 7256 22100 7268
rect 21867 7228 22100 7256
rect 21867 7225 21879 7228
rect 21821 7219 21879 7225
rect 22094 7216 22100 7228
rect 22152 7216 22158 7268
rect 25498 7256 25504 7268
rect 25459 7228 25504 7256
rect 25498 7216 25504 7228
rect 25556 7216 25562 7268
rect 19426 7188 19432 7200
rect 19076 7160 19432 7188
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 20254 7188 20260 7200
rect 20215 7160 20260 7188
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 24762 7148 24768 7200
rect 24820 7188 24826 7200
rect 25041 7191 25099 7197
rect 25041 7188 25053 7191
rect 24820 7160 25053 7188
rect 24820 7148 24826 7160
rect 25041 7157 25053 7160
rect 25087 7157 25099 7191
rect 25041 7151 25099 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 13173 6987 13231 6993
rect 13173 6953 13185 6987
rect 13219 6984 13231 6987
rect 13538 6984 13544 6996
rect 13219 6956 13544 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 13538 6944 13544 6956
rect 13596 6984 13602 6996
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 13596 6956 13737 6984
rect 13596 6944 13602 6956
rect 13725 6953 13737 6956
rect 13771 6953 13783 6987
rect 13725 6947 13783 6953
rect 14642 6944 14648 6996
rect 14700 6984 14706 6996
rect 15565 6987 15623 6993
rect 15565 6984 15577 6987
rect 14700 6956 15577 6984
rect 14700 6944 14706 6956
rect 15565 6953 15577 6956
rect 15611 6984 15623 6987
rect 16390 6984 16396 6996
rect 15611 6956 16396 6984
rect 15611 6953 15623 6956
rect 15565 6947 15623 6953
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 19153 6987 19211 6993
rect 19153 6953 19165 6987
rect 19199 6984 19211 6987
rect 19242 6984 19248 6996
rect 19199 6956 19248 6984
rect 19199 6953 19211 6956
rect 19153 6947 19211 6953
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 20162 6944 20168 6996
rect 20220 6984 20226 6996
rect 22830 6984 22836 6996
rect 20220 6956 22836 6984
rect 20220 6944 20226 6956
rect 22830 6944 22836 6956
rect 22888 6944 22894 6996
rect 22925 6987 22983 6993
rect 22925 6953 22937 6987
rect 22971 6984 22983 6987
rect 23382 6984 23388 6996
rect 22971 6956 23388 6984
rect 22971 6953 22983 6956
rect 22925 6947 22983 6953
rect 23382 6944 23388 6956
rect 23440 6944 23446 6996
rect 23474 6944 23480 6996
rect 23532 6984 23538 6996
rect 23532 6956 23577 6984
rect 23532 6944 23538 6956
rect 24210 6944 24216 6996
rect 24268 6984 24274 6996
rect 24949 6987 25007 6993
rect 24949 6984 24961 6987
rect 24268 6956 24961 6984
rect 24268 6944 24274 6956
rect 24949 6953 24961 6956
rect 24995 6953 25007 6987
rect 24949 6947 25007 6953
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 14921 6919 14979 6925
rect 14921 6916 14933 6919
rect 14792 6888 14933 6916
rect 14792 6876 14798 6888
rect 14921 6885 14933 6888
rect 14967 6885 14979 6919
rect 17586 6916 17592 6928
rect 17547 6888 17592 6916
rect 14921 6879 14979 6885
rect 17586 6876 17592 6888
rect 17644 6876 17650 6928
rect 8573 6851 8631 6857
rect 8573 6817 8585 6851
rect 8619 6848 8631 6851
rect 9858 6848 9864 6860
rect 8619 6820 9864 6848
rect 8619 6817 8631 6820
rect 8573 6811 8631 6817
rect 9858 6808 9864 6820
rect 9916 6848 9922 6860
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 9916 6820 10057 6848
rect 9916 6808 9922 6820
rect 10045 6817 10057 6820
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 10873 6851 10931 6857
rect 10873 6817 10885 6851
rect 10919 6848 10931 6851
rect 10962 6848 10968 6860
rect 10919 6820 10968 6848
rect 10919 6817 10931 6820
rect 10873 6811 10931 6817
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 12049 6851 12107 6857
rect 12049 6848 12061 6851
rect 11940 6820 12061 6848
rect 11940 6808 11946 6820
rect 12049 6817 12061 6820
rect 12095 6817 12107 6851
rect 12049 6811 12107 6817
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 16206 6848 16212 6860
rect 16071 6820 16212 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 16206 6808 16212 6820
rect 16264 6808 16270 6860
rect 17129 6851 17187 6857
rect 17129 6817 17141 6851
rect 17175 6848 17187 6851
rect 17681 6851 17739 6857
rect 17681 6848 17693 6851
rect 17175 6820 17693 6848
rect 17175 6817 17187 6820
rect 17129 6811 17187 6817
rect 17681 6817 17693 6820
rect 17727 6848 17739 6851
rect 17862 6848 17868 6860
rect 17727 6820 17868 6848
rect 17727 6817 17739 6820
rect 17681 6811 17739 6817
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 19260 6848 19288 6944
rect 19610 6916 19616 6928
rect 19523 6888 19616 6916
rect 19610 6876 19616 6888
rect 19668 6916 19674 6928
rect 20438 6916 20444 6928
rect 19668 6888 20444 6916
rect 19668 6876 19674 6888
rect 20438 6876 20444 6888
rect 20496 6876 20502 6928
rect 23842 6925 23848 6928
rect 23836 6916 23848 6925
rect 23803 6888 23848 6916
rect 23836 6879 23848 6888
rect 23842 6876 23848 6879
rect 23900 6876 23906 6928
rect 19260 6820 19840 6848
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 9674 6712 9680 6724
rect 9635 6684 9680 6712
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 10042 6672 10048 6724
rect 10100 6712 10106 6724
rect 10244 6712 10272 6743
rect 10778 6740 10784 6792
rect 10836 6780 10842 6792
rect 11793 6783 11851 6789
rect 11793 6780 11805 6783
rect 10836 6752 11805 6780
rect 10836 6740 10842 6752
rect 10100 6684 10272 6712
rect 10100 6672 10106 6684
rect 11164 6656 11192 6752
rect 11793 6749 11805 6752
rect 11839 6749 11851 6783
rect 16114 6780 16120 6792
rect 16075 6752 16120 6780
rect 11793 6743 11851 6749
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16301 6783 16359 6789
rect 16301 6749 16313 6783
rect 16347 6780 16359 6783
rect 16850 6780 16856 6792
rect 16347 6752 16856 6780
rect 16347 6749 16359 6752
rect 16301 6743 16359 6749
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 17770 6780 17776 6792
rect 17731 6752 17776 6780
rect 17770 6740 17776 6752
rect 17828 6740 17834 6792
rect 19518 6740 19524 6792
rect 19576 6780 19582 6792
rect 19812 6789 19840 6820
rect 20806 6808 20812 6860
rect 20864 6848 20870 6860
rect 21157 6851 21215 6857
rect 21157 6848 21169 6851
rect 20864 6820 21169 6848
rect 20864 6808 20870 6820
rect 21157 6817 21169 6820
rect 21203 6817 21215 6851
rect 21157 6811 21215 6817
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 19576 6752 19717 6780
rect 19576 6740 19582 6752
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 19797 6783 19855 6789
rect 19797 6749 19809 6783
rect 19843 6749 19855 6783
rect 20898 6780 20904 6792
rect 20859 6752 20904 6780
rect 19797 6743 19855 6749
rect 20898 6740 20904 6752
rect 20956 6740 20962 6792
rect 23566 6780 23572 6792
rect 21928 6752 23572 6780
rect 15654 6712 15660 6724
rect 15615 6684 15660 6712
rect 15654 6672 15660 6684
rect 15712 6672 15718 6724
rect 17218 6712 17224 6724
rect 17179 6684 17224 6712
rect 17218 6672 17224 6684
rect 17276 6672 17282 6724
rect 19245 6715 19303 6721
rect 19245 6681 19257 6715
rect 19291 6712 19303 6715
rect 19291 6684 20668 6712
rect 19291 6681 19303 6684
rect 19245 6675 19303 6681
rect 20640 6656 20668 6684
rect 9030 6644 9036 6656
rect 8991 6616 9036 6644
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 11146 6644 11152 6656
rect 11107 6616 11152 6644
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 14090 6644 14096 6656
rect 14051 6616 14096 6644
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14645 6647 14703 6653
rect 14645 6613 14657 6647
rect 14691 6644 14703 6647
rect 14734 6644 14740 6656
rect 14691 6616 14740 6644
rect 14691 6613 14703 6616
rect 14645 6607 14703 6613
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 18325 6647 18383 6653
rect 18325 6644 18337 6647
rect 18104 6616 18337 6644
rect 18104 6604 18110 6616
rect 18325 6613 18337 6616
rect 18371 6613 18383 6647
rect 18782 6644 18788 6656
rect 18743 6616 18788 6644
rect 18325 6607 18383 6613
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 20346 6644 20352 6656
rect 20307 6616 20352 6644
rect 20346 6604 20352 6616
rect 20404 6604 20410 6656
rect 20622 6644 20628 6656
rect 20583 6616 20628 6644
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 20898 6604 20904 6656
rect 20956 6644 20962 6656
rect 21928 6644 21956 6752
rect 23566 6740 23572 6752
rect 23624 6740 23630 6792
rect 22278 6644 22284 6656
rect 20956 6616 21956 6644
rect 22239 6616 22284 6644
rect 20956 6604 20962 6616
rect 22278 6604 22284 6616
rect 22336 6604 22342 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 8941 6443 8999 6449
rect 8941 6409 8953 6443
rect 8987 6440 8999 6443
rect 10042 6440 10048 6452
rect 8987 6412 10048 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 10042 6400 10048 6412
rect 10100 6440 10106 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 10100 6412 10425 6440
rect 10100 6400 10106 6412
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 10413 6403 10471 6409
rect 11517 6443 11575 6449
rect 11517 6409 11529 6443
rect 11563 6440 11575 6443
rect 11882 6440 11888 6452
rect 11563 6412 11888 6440
rect 11563 6409 11575 6412
rect 11517 6403 11575 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12437 6443 12495 6449
rect 12437 6409 12449 6443
rect 12483 6440 12495 6443
rect 13722 6440 13728 6452
rect 12483 6412 13728 6440
rect 12483 6409 12495 6412
rect 12437 6403 12495 6409
rect 13722 6400 13728 6412
rect 13780 6440 13786 6452
rect 14090 6440 14096 6452
rect 13780 6412 14096 6440
rect 13780 6400 13786 6412
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 15197 6443 15255 6449
rect 15197 6409 15209 6443
rect 15243 6440 15255 6443
rect 15838 6440 15844 6452
rect 15243 6412 15844 6440
rect 15243 6409 15255 6412
rect 15197 6403 15255 6409
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 16669 6443 16727 6449
rect 16669 6409 16681 6443
rect 16715 6440 16727 6443
rect 16850 6440 16856 6452
rect 16715 6412 16856 6440
rect 16715 6409 16727 6412
rect 16669 6403 16727 6409
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 18874 6440 18880 6452
rect 18835 6412 18880 6440
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 19337 6443 19395 6449
rect 19337 6409 19349 6443
rect 19383 6440 19395 6443
rect 20530 6440 20536 6452
rect 19383 6412 20536 6440
rect 19383 6409 19395 6412
rect 19337 6403 19395 6409
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 23109 6443 23167 6449
rect 23109 6409 23121 6443
rect 23155 6440 23167 6443
rect 23842 6440 23848 6452
rect 23155 6412 23848 6440
rect 23155 6409 23167 6412
rect 23109 6403 23167 6409
rect 23842 6400 23848 6412
rect 23900 6440 23906 6452
rect 25041 6443 25099 6449
rect 25041 6440 25053 6443
rect 23900 6412 25053 6440
rect 23900 6400 23906 6412
rect 25041 6409 25053 6412
rect 25087 6409 25099 6443
rect 25041 6403 25099 6409
rect 11900 6304 11928 6400
rect 15105 6375 15163 6381
rect 15105 6341 15117 6375
rect 15151 6372 15163 6375
rect 16114 6372 16120 6384
rect 15151 6344 16120 6372
rect 15151 6341 15163 6344
rect 15105 6335 15163 6341
rect 16114 6332 16120 6344
rect 16172 6332 16178 6384
rect 19058 6332 19064 6384
rect 19116 6372 19122 6384
rect 19116 6344 19932 6372
rect 19116 6332 19122 6344
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 11900 6276 13001 6304
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 15746 6304 15752 6316
rect 15707 6276 15752 6304
rect 12989 6267 13047 6273
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 18782 6264 18788 6316
rect 18840 6304 18846 6316
rect 19334 6304 19340 6316
rect 18840 6276 19340 6304
rect 18840 6264 18846 6276
rect 19334 6264 19340 6276
rect 19392 6304 19398 6316
rect 19904 6313 19932 6344
rect 19797 6307 19855 6313
rect 19797 6304 19809 6307
rect 19392 6276 19809 6304
rect 19392 6264 19398 6276
rect 19797 6273 19809 6276
rect 19843 6273 19855 6307
rect 19797 6267 19855 6273
rect 19889 6307 19947 6313
rect 19889 6273 19901 6307
rect 19935 6304 19947 6307
rect 20254 6304 20260 6316
rect 19935 6276 20260 6304
rect 19935 6273 19947 6276
rect 19889 6267 19947 6273
rect 20254 6264 20260 6276
rect 20312 6304 20318 6316
rect 20530 6304 20536 6316
rect 20312 6276 20536 6304
rect 20312 6264 20318 6276
rect 20530 6264 20536 6276
rect 20588 6304 20594 6316
rect 20806 6304 20812 6316
rect 20588 6276 20812 6304
rect 20588 6264 20594 6276
rect 20806 6264 20812 6276
rect 20864 6264 20870 6316
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6304 20959 6307
rect 20947 6276 21128 6304
rect 20947 6273 20959 6276
rect 20901 6267 20959 6273
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 9030 6236 9036 6248
rect 8720 6208 9036 6236
rect 8720 6196 8726 6208
rect 9030 6196 9036 6208
rect 9088 6196 9094 6248
rect 16206 6236 16212 6248
rect 16167 6208 16212 6236
rect 16206 6196 16212 6208
rect 16264 6196 16270 6248
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6236 16911 6239
rect 18233 6239 18291 6245
rect 16899 6208 17540 6236
rect 16899 6205 16911 6208
rect 16853 6199 16911 6205
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 9278 6171 9336 6177
rect 9278 6168 9290 6171
rect 9180 6140 9290 6168
rect 9180 6128 9186 6140
rect 9278 6137 9290 6140
rect 9324 6137 9336 6171
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 9278 6131 9336 6137
rect 12268 6140 12817 6168
rect 12268 6112 12296 6140
rect 12805 6137 12817 6140
rect 12851 6137 12863 6171
rect 15565 6171 15623 6177
rect 15565 6168 15577 6171
rect 12805 6131 12863 6137
rect 14660 6140 15577 6168
rect 14660 6112 14688 6140
rect 15565 6137 15577 6140
rect 15611 6137 15623 6171
rect 15565 6131 15623 6137
rect 17512 6112 17540 6208
rect 18233 6205 18245 6239
rect 18279 6236 18291 6239
rect 18874 6236 18880 6248
rect 18279 6208 18880 6236
rect 18279 6205 18291 6208
rect 18233 6199 18291 6205
rect 18874 6196 18880 6208
rect 18932 6196 18938 6248
rect 19705 6239 19763 6245
rect 19705 6205 19717 6239
rect 19751 6236 19763 6239
rect 20622 6236 20628 6248
rect 19751 6208 20628 6236
rect 19751 6205 19763 6208
rect 19705 6199 19763 6205
rect 20622 6196 20628 6208
rect 20680 6196 20686 6248
rect 20993 6239 21051 6245
rect 20993 6205 21005 6239
rect 21039 6205 21051 6239
rect 21100 6236 21128 6276
rect 23566 6264 23572 6316
rect 23624 6304 23630 6316
rect 23661 6307 23719 6313
rect 23661 6304 23673 6307
rect 23624 6276 23673 6304
rect 23624 6264 23630 6276
rect 23661 6273 23673 6276
rect 23707 6273 23719 6307
rect 23661 6267 23719 6273
rect 21266 6245 21272 6248
rect 21260 6236 21272 6245
rect 21100 6208 21272 6236
rect 20993 6199 21051 6205
rect 21260 6199 21272 6208
rect 21324 6236 21330 6248
rect 22278 6236 22284 6248
rect 21324 6208 22284 6236
rect 20898 6128 20904 6180
rect 20956 6168 20962 6180
rect 21008 6168 21036 6199
rect 21266 6196 21272 6199
rect 21324 6196 21330 6208
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 21358 6168 21364 6180
rect 20956 6140 21364 6168
rect 20956 6128 20962 6140
rect 21358 6128 21364 6140
rect 21416 6128 21422 6180
rect 22646 6128 22652 6180
rect 22704 6168 22710 6180
rect 23477 6171 23535 6177
rect 23477 6168 23489 6171
rect 22704 6140 23489 6168
rect 22704 6128 22710 6140
rect 23477 6137 23489 6140
rect 23523 6168 23535 6171
rect 23928 6171 23986 6177
rect 23928 6168 23940 6171
rect 23523 6140 23940 6168
rect 23523 6137 23535 6140
rect 23477 6131 23535 6137
rect 23928 6137 23940 6140
rect 23974 6168 23986 6171
rect 24578 6168 24584 6180
rect 23974 6140 24584 6168
rect 23974 6137 23986 6140
rect 23928 6131 23986 6137
rect 24578 6128 24584 6140
rect 24636 6128 24642 6180
rect 10686 6060 10692 6112
rect 10744 6100 10750 6112
rect 11057 6103 11115 6109
rect 11057 6100 11069 6103
rect 10744 6072 11069 6100
rect 10744 6060 10750 6072
rect 11057 6069 11069 6072
rect 11103 6100 11115 6103
rect 11146 6100 11152 6112
rect 11103 6072 11152 6100
rect 11103 6069 11115 6072
rect 11057 6063 11115 6069
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 12250 6100 12256 6112
rect 12211 6072 12256 6100
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12894 6100 12900 6112
rect 12855 6072 12900 6100
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13446 6100 13452 6112
rect 13407 6072 13452 6100
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 14182 6100 14188 6112
rect 14143 6072 14188 6100
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 14642 6100 14648 6112
rect 14603 6072 14648 6100
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 15657 6103 15715 6109
rect 15657 6069 15669 6103
rect 15703 6100 15715 6103
rect 15930 6100 15936 6112
rect 15703 6072 15936 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 17034 6100 17040 6112
rect 16995 6072 17040 6100
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 17494 6100 17500 6112
rect 17455 6072 17500 6100
rect 17494 6060 17500 6072
rect 17552 6060 17558 6112
rect 17770 6100 17776 6112
rect 17731 6072 17776 6100
rect 17770 6060 17776 6072
rect 17828 6060 17834 6112
rect 18417 6103 18475 6109
rect 18417 6069 18429 6103
rect 18463 6100 18475 6103
rect 18966 6100 18972 6112
rect 18463 6072 18972 6100
rect 18463 6069 18475 6072
rect 18417 6063 18475 6069
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 19245 6103 19303 6109
rect 19245 6069 19257 6103
rect 19291 6100 19303 6103
rect 19518 6100 19524 6112
rect 19291 6072 19524 6100
rect 19291 6069 19303 6072
rect 19245 6063 19303 6069
rect 19518 6060 19524 6072
rect 19576 6060 19582 6112
rect 20438 6100 20444 6112
rect 20351 6072 20444 6100
rect 20438 6060 20444 6072
rect 20496 6100 20502 6112
rect 22186 6100 22192 6112
rect 20496 6072 22192 6100
rect 20496 6060 20502 6072
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 22370 6100 22376 6112
rect 22331 6072 22376 6100
rect 22370 6060 22376 6072
rect 22428 6060 22434 6112
rect 25038 6060 25044 6112
rect 25096 6100 25102 6112
rect 25593 6103 25651 6109
rect 25593 6100 25605 6103
rect 25096 6072 25605 6100
rect 25096 6060 25102 6072
rect 25593 6069 25605 6072
rect 25639 6069 25651 6103
rect 25593 6063 25651 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 8570 5896 8576 5908
rect 8531 5868 8576 5896
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 9122 5896 9128 5908
rect 9083 5868 9128 5896
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 9858 5896 9864 5908
rect 9819 5868 9864 5896
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10134 5856 10140 5908
rect 10192 5896 10198 5908
rect 10229 5899 10287 5905
rect 10229 5896 10241 5899
rect 10192 5868 10241 5896
rect 10192 5856 10198 5868
rect 10229 5865 10241 5868
rect 10275 5865 10287 5899
rect 11882 5896 11888 5908
rect 11843 5868 11888 5896
rect 10229 5859 10287 5865
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 12986 5896 12992 5908
rect 12947 5868 12992 5896
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 18322 5896 18328 5908
rect 13320 5868 18328 5896
rect 13320 5856 13326 5868
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 18785 5899 18843 5905
rect 18785 5865 18797 5899
rect 18831 5896 18843 5899
rect 19058 5896 19064 5908
rect 18831 5868 19064 5896
rect 18831 5865 18843 5868
rect 18785 5859 18843 5865
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 19153 5899 19211 5905
rect 19153 5865 19165 5899
rect 19199 5896 19211 5899
rect 19242 5896 19248 5908
rect 19199 5868 19248 5896
rect 19199 5865 19211 5868
rect 19153 5859 19211 5865
rect 19242 5856 19248 5868
rect 19300 5856 19306 5908
rect 19426 5856 19432 5908
rect 19484 5896 19490 5908
rect 20346 5896 20352 5908
rect 19484 5868 19748 5896
rect 20307 5868 20352 5896
rect 19484 5856 19490 5868
rect 12526 5828 12532 5840
rect 12439 5800 12532 5828
rect 12526 5788 12532 5800
rect 12584 5828 12590 5840
rect 12894 5828 12900 5840
rect 12584 5800 12900 5828
rect 12584 5788 12590 5800
rect 12894 5788 12900 5800
rect 12952 5788 12958 5840
rect 17028 5831 17086 5837
rect 17028 5797 17040 5831
rect 17074 5828 17086 5831
rect 17218 5828 17224 5840
rect 17074 5800 17224 5828
rect 17074 5797 17086 5800
rect 17028 5791 17086 5797
rect 17218 5788 17224 5800
rect 17276 5788 17282 5840
rect 10505 5763 10563 5769
rect 10505 5729 10517 5763
rect 10551 5760 10563 5763
rect 10594 5760 10600 5772
rect 10551 5732 10600 5760
rect 10551 5729 10563 5732
rect 10505 5723 10563 5729
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 10778 5769 10784 5772
rect 10772 5723 10784 5769
rect 10836 5760 10842 5772
rect 10836 5732 10872 5760
rect 10778 5720 10784 5723
rect 10836 5720 10842 5732
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 13357 5763 13415 5769
rect 13357 5760 13369 5763
rect 12400 5732 13369 5760
rect 12400 5720 12406 5732
rect 13357 5729 13369 5732
rect 13403 5729 13415 5763
rect 15654 5760 15660 5772
rect 15615 5732 15660 5760
rect 13357 5723 13415 5729
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 13449 5695 13507 5701
rect 13449 5692 13461 5695
rect 12492 5664 13461 5692
rect 12492 5652 12498 5664
rect 13449 5661 13461 5664
rect 13495 5661 13507 5695
rect 13449 5655 13507 5661
rect 13538 5652 13544 5704
rect 13596 5692 13602 5704
rect 15565 5695 15623 5701
rect 15565 5692 15577 5695
rect 13596 5664 13641 5692
rect 13740 5664 15577 5692
rect 13596 5652 13602 5664
rect 12894 5624 12900 5636
rect 12807 5596 12900 5624
rect 12894 5584 12900 5596
rect 12952 5624 12958 5636
rect 13740 5624 13768 5664
rect 15565 5661 15577 5664
rect 15611 5692 15623 5695
rect 15746 5692 15752 5704
rect 15611 5664 15752 5692
rect 15611 5661 15623 5664
rect 15565 5655 15623 5661
rect 15746 5652 15752 5664
rect 15804 5692 15810 5704
rect 16390 5692 16396 5704
rect 15804 5664 16396 5692
rect 15804 5652 15810 5664
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 16577 5695 16635 5701
rect 16577 5661 16589 5695
rect 16623 5692 16635 5695
rect 16666 5692 16672 5704
rect 16623 5664 16672 5692
rect 16623 5661 16635 5664
rect 16577 5655 16635 5661
rect 16666 5652 16672 5664
rect 16724 5692 16730 5704
rect 16761 5695 16819 5701
rect 16761 5692 16773 5695
rect 16724 5664 16773 5692
rect 16724 5652 16730 5664
rect 16761 5661 16773 5664
rect 16807 5661 16819 5695
rect 19260 5692 19288 5856
rect 19426 5720 19432 5772
rect 19484 5760 19490 5772
rect 19720 5769 19748 5868
rect 20346 5856 20352 5868
rect 20404 5856 20410 5908
rect 20530 5856 20536 5908
rect 20588 5896 20594 5908
rect 20625 5899 20683 5905
rect 20625 5896 20637 5899
rect 20588 5868 20637 5896
rect 20588 5856 20594 5868
rect 20625 5865 20637 5868
rect 20671 5865 20683 5899
rect 20625 5859 20683 5865
rect 20714 5856 20720 5908
rect 20772 5896 20778 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 20772 5868 20913 5896
rect 20772 5856 20778 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 21174 5856 21180 5908
rect 21232 5896 21238 5908
rect 21269 5899 21327 5905
rect 21269 5896 21281 5899
rect 21232 5868 21281 5896
rect 21232 5856 21238 5868
rect 21269 5865 21281 5868
rect 21315 5865 21327 5899
rect 23658 5896 23664 5908
rect 23619 5868 23664 5896
rect 21269 5859 21327 5865
rect 23658 5856 23664 5868
rect 23716 5856 23722 5908
rect 23750 5856 23756 5908
rect 23808 5896 23814 5908
rect 24029 5899 24087 5905
rect 24029 5896 24041 5899
rect 23808 5868 24041 5896
rect 23808 5856 23814 5868
rect 24029 5865 24041 5868
rect 24075 5865 24087 5899
rect 24029 5859 24087 5865
rect 23569 5831 23627 5837
rect 23569 5797 23581 5831
rect 23615 5828 23627 5831
rect 23842 5828 23848 5840
rect 23615 5800 23848 5828
rect 23615 5797 23627 5800
rect 23569 5791 23627 5797
rect 23842 5788 23848 5800
rect 23900 5828 23906 5840
rect 23900 5800 24164 5828
rect 23900 5788 23906 5800
rect 19613 5763 19671 5769
rect 19613 5760 19625 5763
rect 19484 5732 19625 5760
rect 19484 5720 19490 5732
rect 19613 5729 19625 5732
rect 19659 5729 19671 5763
rect 19613 5723 19671 5729
rect 19705 5763 19763 5769
rect 19705 5729 19717 5763
rect 19751 5760 19763 5763
rect 20162 5760 20168 5772
rect 19751 5732 20168 5760
rect 19751 5729 19763 5732
rect 19705 5723 19763 5729
rect 20162 5720 20168 5732
rect 20220 5720 20226 5772
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 22557 5763 22615 5769
rect 20772 5732 21496 5760
rect 20772 5720 20778 5732
rect 19797 5695 19855 5701
rect 19797 5692 19809 5695
rect 19260 5664 19809 5692
rect 16761 5655 16819 5661
rect 19797 5661 19809 5664
rect 19843 5692 19855 5695
rect 19886 5692 19892 5704
rect 19843 5664 19892 5692
rect 19843 5661 19855 5664
rect 19797 5655 19855 5661
rect 19886 5652 19892 5664
rect 19944 5652 19950 5704
rect 21468 5701 21496 5732
rect 22557 5729 22569 5763
rect 22603 5760 22615 5763
rect 23106 5760 23112 5772
rect 22603 5732 23112 5760
rect 22603 5729 22615 5732
rect 22557 5723 22615 5729
rect 23106 5720 23112 5732
rect 23164 5720 23170 5772
rect 23290 5720 23296 5772
rect 23348 5760 23354 5772
rect 23658 5760 23664 5772
rect 23348 5732 23664 5760
rect 23348 5720 23354 5732
rect 23658 5720 23664 5732
rect 23716 5720 23722 5772
rect 24136 5760 24164 5800
rect 24136 5732 24256 5760
rect 21361 5695 21419 5701
rect 21361 5661 21373 5695
rect 21407 5661 21419 5695
rect 21361 5655 21419 5661
rect 21453 5695 21511 5701
rect 21453 5661 21465 5695
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 12952 5596 13768 5624
rect 15105 5627 15163 5633
rect 12952 5584 12958 5596
rect 15105 5593 15117 5627
rect 15151 5624 15163 5627
rect 15930 5624 15936 5636
rect 15151 5596 15936 5624
rect 15151 5593 15163 5596
rect 15105 5587 15163 5593
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 19245 5627 19303 5633
rect 19245 5593 19257 5627
rect 19291 5624 19303 5627
rect 21082 5624 21088 5636
rect 19291 5596 21088 5624
rect 19291 5593 19303 5596
rect 19245 5587 19303 5593
rect 21082 5584 21088 5596
rect 21140 5624 21146 5636
rect 21376 5624 21404 5655
rect 22002 5652 22008 5704
rect 22060 5692 22066 5704
rect 24228 5701 24256 5732
rect 24670 5720 24676 5772
rect 24728 5760 24734 5772
rect 25225 5763 25283 5769
rect 25225 5760 25237 5763
rect 24728 5732 25237 5760
rect 24728 5720 24734 5732
rect 25225 5729 25237 5732
rect 25271 5760 25283 5763
rect 25590 5760 25596 5772
rect 25271 5732 25596 5760
rect 25271 5729 25283 5732
rect 25225 5723 25283 5729
rect 25590 5720 25596 5732
rect 25648 5720 25654 5772
rect 23201 5695 23259 5701
rect 23201 5692 23213 5695
rect 22060 5664 23213 5692
rect 22060 5652 22066 5664
rect 23201 5661 23213 5664
rect 23247 5692 23259 5695
rect 24121 5695 24179 5701
rect 24121 5692 24133 5695
rect 23247 5664 24133 5692
rect 23247 5661 23259 5664
rect 23201 5655 23259 5661
rect 24121 5661 24133 5664
rect 24167 5661 24179 5695
rect 24121 5655 24179 5661
rect 24213 5695 24271 5701
rect 24213 5661 24225 5695
rect 24259 5661 24271 5695
rect 24213 5655 24271 5661
rect 21140 5596 21404 5624
rect 21140 5584 21146 5596
rect 21910 5584 21916 5636
rect 21968 5624 21974 5636
rect 22741 5627 22799 5633
rect 22741 5624 22753 5627
rect 21968 5596 22753 5624
rect 21968 5584 21974 5596
rect 22741 5593 22753 5596
rect 22787 5593 22799 5627
rect 22741 5587 22799 5593
rect 23566 5584 23572 5636
rect 23624 5624 23630 5636
rect 24673 5627 24731 5633
rect 24673 5624 24685 5627
rect 23624 5596 24685 5624
rect 23624 5584 23630 5596
rect 24673 5593 24685 5596
rect 24719 5624 24731 5627
rect 25038 5624 25044 5636
rect 24719 5596 25044 5624
rect 24719 5593 24731 5596
rect 24673 5587 24731 5593
rect 25038 5584 25044 5596
rect 25096 5584 25102 5636
rect 15838 5556 15844 5568
rect 15799 5528 15844 5556
rect 15838 5516 15844 5528
rect 15896 5516 15902 5568
rect 16574 5516 16580 5568
rect 16632 5556 16638 5568
rect 17770 5556 17776 5568
rect 16632 5528 17776 5556
rect 16632 5516 16638 5528
rect 17770 5516 17776 5528
rect 17828 5556 17834 5568
rect 18141 5559 18199 5565
rect 18141 5556 18153 5559
rect 17828 5528 18153 5556
rect 17828 5516 17834 5528
rect 18141 5525 18153 5528
rect 18187 5525 18199 5559
rect 18141 5519 18199 5525
rect 22094 5516 22100 5568
rect 22152 5556 22158 5568
rect 22465 5559 22523 5565
rect 22152 5528 22197 5556
rect 22152 5516 22158 5528
rect 22465 5525 22477 5559
rect 22511 5556 22523 5559
rect 22646 5556 22652 5568
rect 22511 5528 22652 5556
rect 22511 5525 22523 5528
rect 22465 5519 22523 5525
rect 22646 5516 22652 5528
rect 22704 5516 22710 5568
rect 25406 5556 25412 5568
rect 25367 5528 25412 5556
rect 25406 5516 25412 5528
rect 25464 5516 25470 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 10689 5355 10747 5361
rect 10689 5321 10701 5355
rect 10735 5352 10747 5355
rect 10778 5352 10784 5364
rect 10735 5324 10784 5352
rect 10735 5321 10747 5324
rect 10689 5315 10747 5321
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 12253 5355 12311 5361
rect 12253 5352 12265 5355
rect 11348 5324 12265 5352
rect 11348 5225 11376 5324
rect 12253 5321 12265 5324
rect 12299 5352 12311 5355
rect 12342 5352 12348 5364
rect 12299 5324 12348 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 17129 5355 17187 5361
rect 17129 5321 17141 5355
rect 17175 5352 17187 5355
rect 17218 5352 17224 5364
rect 17175 5324 17224 5352
rect 17175 5321 17187 5324
rect 17129 5315 17187 5321
rect 17218 5312 17224 5324
rect 17276 5352 17282 5364
rect 18506 5352 18512 5364
rect 17276 5324 18512 5352
rect 17276 5312 17282 5324
rect 18506 5312 18512 5324
rect 18564 5312 18570 5364
rect 18877 5355 18935 5361
rect 18877 5321 18889 5355
rect 18923 5352 18935 5355
rect 19150 5352 19156 5364
rect 18923 5324 19156 5352
rect 18923 5321 18935 5324
rect 18877 5315 18935 5321
rect 16666 5244 16672 5296
rect 16724 5284 16730 5296
rect 17405 5287 17463 5293
rect 17405 5284 17417 5287
rect 16724 5256 17417 5284
rect 16724 5244 16730 5256
rect 17405 5253 17417 5256
rect 17451 5253 17463 5287
rect 17405 5247 17463 5253
rect 11333 5219 11391 5225
rect 11333 5185 11345 5219
rect 11379 5185 11391 5219
rect 11333 5179 11391 5185
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5216 11943 5219
rect 12342 5216 12348 5228
rect 11931 5188 12348 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 12342 5176 12348 5188
rect 12400 5176 12406 5228
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8662 5148 8668 5160
rect 8251 5120 8668 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 12894 5157 12900 5160
rect 12621 5151 12679 5157
rect 12621 5117 12633 5151
rect 12667 5117 12679 5151
rect 12888 5148 12900 5157
rect 12855 5120 12900 5148
rect 12621 5111 12679 5117
rect 12888 5111 12900 5120
rect 8573 5083 8631 5089
rect 8573 5049 8585 5083
rect 8619 5080 8631 5083
rect 8932 5083 8990 5089
rect 8932 5080 8944 5083
rect 8619 5052 8944 5080
rect 8619 5049 8631 5052
rect 8573 5043 8631 5049
rect 8932 5049 8944 5052
rect 8978 5080 8990 5083
rect 9490 5080 9496 5092
rect 8978 5052 9496 5080
rect 8978 5049 8990 5052
rect 8932 5043 8990 5049
rect 9490 5040 9496 5052
rect 9548 5040 9554 5092
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 12636 5080 12664 5111
rect 12894 5108 12900 5111
rect 12952 5108 12958 5160
rect 14734 5108 14740 5160
rect 14792 5148 14798 5160
rect 15102 5148 15108 5160
rect 14792 5120 15108 5148
rect 14792 5108 14798 5120
rect 15102 5108 15108 5120
rect 15160 5108 15166 5160
rect 16482 5108 16488 5160
rect 16540 5108 16546 5160
rect 18233 5151 18291 5157
rect 18233 5117 18245 5151
rect 18279 5148 18291 5151
rect 18892 5148 18920 5315
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 19334 5352 19340 5364
rect 19295 5324 19340 5352
rect 19334 5312 19340 5324
rect 19392 5312 19398 5364
rect 21174 5312 21180 5364
rect 21232 5352 21238 5364
rect 21453 5355 21511 5361
rect 21453 5352 21465 5355
rect 21232 5324 21465 5352
rect 21232 5312 21238 5324
rect 21453 5321 21465 5324
rect 21499 5321 21511 5355
rect 21453 5315 21511 5321
rect 21637 5355 21695 5361
rect 21637 5321 21649 5355
rect 21683 5352 21695 5355
rect 22002 5352 22008 5364
rect 21683 5324 21864 5352
rect 21963 5324 22008 5352
rect 21683 5321 21695 5324
rect 21637 5315 21695 5321
rect 21085 5287 21143 5293
rect 21085 5253 21097 5287
rect 21131 5284 21143 5287
rect 21726 5284 21732 5296
rect 21131 5256 21732 5284
rect 21131 5253 21143 5256
rect 21085 5247 21143 5253
rect 21726 5244 21732 5256
rect 21784 5244 21790 5296
rect 21836 5284 21864 5324
rect 22002 5312 22008 5324
rect 22060 5312 22066 5364
rect 23106 5352 23112 5364
rect 23067 5324 23112 5352
rect 23106 5312 23112 5324
rect 23164 5312 23170 5364
rect 23477 5355 23535 5361
rect 23477 5321 23489 5355
rect 23523 5352 23535 5355
rect 23658 5352 23664 5364
rect 23523 5324 23664 5352
rect 23523 5321 23535 5324
rect 23477 5315 23535 5321
rect 23658 5312 23664 5324
rect 23716 5312 23722 5364
rect 25590 5352 25596 5364
rect 25551 5324 25596 5352
rect 25590 5312 25596 5324
rect 25648 5312 25654 5364
rect 22094 5284 22100 5296
rect 21836 5256 22100 5284
rect 22094 5244 22100 5256
rect 22152 5284 22158 5296
rect 22152 5256 22508 5284
rect 22152 5244 22158 5256
rect 19886 5216 19892 5228
rect 19847 5188 19892 5216
rect 19886 5176 19892 5188
rect 19944 5176 19950 5228
rect 20898 5148 20904 5160
rect 18279 5120 18920 5148
rect 20859 5120 20904 5148
rect 18279 5117 18291 5120
rect 18233 5111 18291 5117
rect 20898 5108 20904 5120
rect 20956 5108 20962 5160
rect 21818 5148 21824 5160
rect 21779 5120 21824 5148
rect 21818 5108 21824 5120
rect 21876 5148 21882 5160
rect 22480 5157 22508 5256
rect 22646 5216 22652 5228
rect 22607 5188 22652 5216
rect 22646 5176 22652 5188
rect 22704 5176 22710 5228
rect 22373 5151 22431 5157
rect 22373 5148 22385 5151
rect 21876 5120 22385 5148
rect 21876 5108 21882 5120
rect 22373 5117 22385 5120
rect 22419 5117 22431 5151
rect 22373 5111 22431 5117
rect 22465 5151 22523 5157
rect 22465 5117 22477 5151
rect 22511 5148 22523 5151
rect 23382 5148 23388 5160
rect 22511 5120 23388 5148
rect 22511 5117 22523 5120
rect 22465 5111 22523 5117
rect 23382 5108 23388 5120
rect 23440 5108 23446 5160
rect 23658 5148 23664 5160
rect 23619 5120 23664 5148
rect 23658 5108 23664 5120
rect 23716 5108 23722 5160
rect 25038 5148 25044 5160
rect 23768 5120 25044 5148
rect 13446 5080 13452 5092
rect 12400 5052 13452 5080
rect 12400 5040 12406 5052
rect 13446 5040 13452 5052
rect 13504 5040 13510 5092
rect 14645 5083 14703 5089
rect 14645 5049 14657 5083
rect 14691 5080 14703 5083
rect 15350 5083 15408 5089
rect 15350 5080 15362 5083
rect 14691 5052 15362 5080
rect 14691 5049 14703 5052
rect 14645 5043 14703 5049
rect 15350 5049 15362 5052
rect 15396 5080 15408 5083
rect 16500 5080 16528 5108
rect 15396 5052 16528 5080
rect 15396 5049 15408 5052
rect 15350 5043 15408 5049
rect 18598 5040 18604 5092
rect 18656 5080 18662 5092
rect 19705 5083 19763 5089
rect 18656 5052 19380 5080
rect 18656 5040 18662 5052
rect 9122 4972 9128 5024
rect 9180 5012 9186 5024
rect 10045 5015 10103 5021
rect 10045 5012 10057 5015
rect 9180 4984 10057 5012
rect 9180 4972 9186 4984
rect 10045 4981 10057 4984
rect 10091 4981 10103 5015
rect 10045 4975 10103 4981
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 10965 5015 11023 5021
rect 10965 5012 10977 5015
rect 10744 4984 10977 5012
rect 10744 4972 10750 4984
rect 10965 4981 10977 4984
rect 11011 4981 11023 5015
rect 10965 4975 11023 4981
rect 12986 4972 12992 5024
rect 13044 5012 13050 5024
rect 14001 5015 14059 5021
rect 14001 5012 14013 5015
rect 13044 4984 14013 5012
rect 13044 4972 13050 4984
rect 14001 4981 14013 4984
rect 14047 4981 14059 5015
rect 15010 5012 15016 5024
rect 14971 4984 15016 5012
rect 14001 4975 14059 4981
rect 15010 4972 15016 4984
rect 15068 4972 15074 5024
rect 16482 5012 16488 5024
rect 16443 4984 16488 5012
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17770 4972 17776 4984
rect 17828 5012 17834 5024
rect 18046 5012 18052 5024
rect 17828 4984 18052 5012
rect 17828 4972 17834 4984
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 18414 5012 18420 5024
rect 18375 4984 18420 5012
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 19150 5012 19156 5024
rect 19111 4984 19156 5012
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 19352 5012 19380 5052
rect 19705 5049 19717 5083
rect 19751 5080 19763 5083
rect 20070 5080 20076 5092
rect 19751 5052 20076 5080
rect 19751 5049 19763 5052
rect 19705 5043 19763 5049
rect 20070 5040 20076 5052
rect 20128 5040 20134 5092
rect 20162 5040 20168 5092
rect 20220 5080 20226 5092
rect 20441 5083 20499 5089
rect 20441 5080 20453 5083
rect 20220 5052 20453 5080
rect 20220 5040 20226 5052
rect 20441 5049 20453 5052
rect 20487 5080 20499 5083
rect 21637 5083 21695 5089
rect 21637 5080 21649 5083
rect 20487 5052 21649 5080
rect 20487 5049 20499 5052
rect 20441 5043 20499 5049
rect 21637 5049 21649 5052
rect 21683 5049 21695 5083
rect 21637 5043 21695 5049
rect 23106 5040 23112 5092
rect 23164 5080 23170 5092
rect 23768 5080 23796 5120
rect 25038 5108 25044 5120
rect 25096 5108 25102 5160
rect 23934 5089 23940 5092
rect 23928 5080 23940 5089
rect 23164 5052 23796 5080
rect 23895 5052 23940 5080
rect 23164 5040 23170 5052
rect 23928 5043 23940 5052
rect 23934 5040 23940 5043
rect 23992 5040 23998 5092
rect 24670 5040 24676 5092
rect 24728 5080 24734 5092
rect 24728 5052 25084 5080
rect 24728 5040 24734 5052
rect 19797 5015 19855 5021
rect 19797 5012 19809 5015
rect 19352 4984 19809 5012
rect 19797 4981 19809 4984
rect 19843 5012 19855 5015
rect 20806 5012 20812 5024
rect 19843 4984 20812 5012
rect 19843 4981 19855 4984
rect 19797 4975 19855 4981
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 25056 5021 25084 5052
rect 25041 5015 25099 5021
rect 25041 4981 25053 5015
rect 25087 5012 25099 5015
rect 25130 5012 25136 5024
rect 25087 4984 25136 5012
rect 25087 4981 25099 4984
rect 25041 4975 25099 4981
rect 25130 4972 25136 4984
rect 25188 4972 25194 5024
rect 25590 4972 25596 5024
rect 25648 5012 25654 5024
rect 25961 5015 26019 5021
rect 25961 5012 25973 5015
rect 25648 4984 25973 5012
rect 25648 4972 25654 4984
rect 25961 4981 25973 4984
rect 26007 4981 26019 5015
rect 25961 4975 26019 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 9122 4768 9128 4820
rect 9180 4808 9186 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9180 4780 9413 4808
rect 9180 4768 9186 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 10134 4808 10140 4820
rect 9723 4780 10140 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 9416 4740 9444 4771
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 11606 4808 11612 4820
rect 11567 4780 11612 4808
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 13538 4808 13544 4820
rect 12492 4780 13544 4808
rect 12492 4768 12498 4780
rect 13538 4768 13544 4780
rect 13596 4808 13602 4820
rect 14001 4811 14059 4817
rect 14001 4808 14013 4811
rect 13596 4780 14013 4808
rect 13596 4768 13602 4780
rect 14001 4777 14013 4780
rect 14047 4777 14059 4811
rect 14001 4771 14059 4777
rect 16390 4768 16396 4820
rect 16448 4808 16454 4820
rect 16669 4811 16727 4817
rect 16669 4808 16681 4811
rect 16448 4780 16681 4808
rect 16448 4768 16454 4780
rect 16669 4777 16681 4780
rect 16715 4777 16727 4811
rect 16669 4771 16727 4777
rect 17586 4768 17592 4820
rect 17644 4808 17650 4820
rect 17773 4811 17831 4817
rect 17773 4808 17785 4811
rect 17644 4780 17785 4808
rect 17644 4768 17650 4780
rect 17773 4777 17785 4780
rect 17819 4777 17831 4811
rect 17773 4771 17831 4777
rect 19061 4811 19119 4817
rect 19061 4777 19073 4811
rect 19107 4808 19119 4811
rect 19242 4808 19248 4820
rect 19107 4780 19248 4808
rect 19107 4777 19119 4780
rect 19061 4771 19119 4777
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 20714 4808 20720 4820
rect 20675 4780 20720 4808
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 22462 4768 22468 4820
rect 22520 4808 22526 4820
rect 23385 4811 23443 4817
rect 23385 4808 23397 4811
rect 22520 4780 23397 4808
rect 22520 4768 22526 4780
rect 23385 4777 23397 4780
rect 23431 4808 23443 4811
rect 23934 4808 23940 4820
rect 23431 4780 23940 4808
rect 23431 4777 23443 4780
rect 23385 4771 23443 4777
rect 23934 4768 23940 4780
rect 23992 4768 23998 4820
rect 24210 4768 24216 4820
rect 24268 4808 24274 4820
rect 24305 4811 24363 4817
rect 24305 4808 24317 4811
rect 24268 4780 24317 4808
rect 24268 4768 24274 4780
rect 24305 4777 24317 4780
rect 24351 4777 24363 4811
rect 24305 4771 24363 4777
rect 24489 4811 24547 4817
rect 24489 4777 24501 4811
rect 24535 4808 24547 4811
rect 24762 4808 24768 4820
rect 24535 4780 24768 4808
rect 24535 4777 24547 4780
rect 24489 4771 24547 4777
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 24949 4811 25007 4817
rect 24949 4777 24961 4811
rect 24995 4808 25007 4811
rect 25222 4808 25228 4820
rect 24995 4780 25228 4808
rect 24995 4777 25007 4780
rect 24949 4771 25007 4777
rect 25222 4768 25228 4780
rect 25280 4768 25286 4820
rect 12161 4743 12219 4749
rect 9416 4712 10272 4740
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 9732 4644 10057 4672
rect 9732 4632 9738 4644
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 10045 4635 10103 4641
rect 8570 4604 8576 4616
rect 8531 4576 8576 4604
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 10244 4613 10272 4712
rect 12161 4709 12173 4743
rect 12207 4740 12219 4743
rect 12888 4743 12946 4749
rect 12888 4740 12900 4743
rect 12207 4712 12900 4740
rect 12207 4709 12219 4712
rect 12161 4703 12219 4709
rect 12888 4709 12900 4712
rect 12934 4740 12946 4743
rect 12986 4740 12992 4752
rect 12934 4712 12992 4740
rect 12934 4709 12946 4712
rect 12888 4703 12946 4709
rect 12986 4700 12992 4712
rect 13044 4700 13050 4752
rect 17681 4743 17739 4749
rect 17681 4709 17693 4743
rect 17727 4740 17739 4743
rect 17862 4740 17868 4752
rect 17727 4712 17868 4740
rect 17727 4709 17739 4712
rect 17681 4703 17739 4709
rect 17862 4700 17868 4712
rect 17920 4700 17926 4752
rect 21450 4700 21456 4752
rect 21508 4740 21514 4752
rect 22250 4743 22308 4749
rect 22250 4740 22262 4743
rect 21508 4712 22262 4740
rect 21508 4700 21514 4712
rect 22250 4709 22262 4712
rect 22296 4740 22308 4743
rect 23014 4740 23020 4752
rect 22296 4712 23020 4740
rect 22296 4709 22308 4712
rect 22250 4703 22308 4709
rect 23014 4700 23020 4712
rect 23072 4700 23078 4752
rect 24857 4743 24915 4749
rect 24857 4709 24869 4743
rect 24903 4740 24915 4743
rect 25038 4740 25044 4752
rect 24903 4712 25044 4740
rect 24903 4709 24915 4712
rect 24857 4703 24915 4709
rect 25038 4700 25044 4712
rect 25096 4700 25102 4752
rect 15562 4681 15568 4684
rect 15556 4672 15568 4681
rect 15523 4644 15568 4672
rect 15556 4635 15568 4644
rect 15562 4632 15568 4635
rect 15620 4632 15626 4684
rect 17402 4632 17408 4684
rect 17460 4672 17466 4684
rect 18141 4675 18199 4681
rect 18141 4672 18153 4675
rect 17460 4644 18153 4672
rect 17460 4632 17466 4644
rect 18141 4641 18153 4644
rect 18187 4641 18199 4675
rect 18141 4635 18199 4641
rect 19518 4632 19524 4684
rect 19576 4672 19582 4684
rect 19705 4675 19763 4681
rect 19705 4672 19717 4675
rect 19576 4644 19717 4672
rect 19576 4632 19582 4644
rect 19705 4641 19717 4644
rect 19751 4672 19763 4675
rect 19978 4672 19984 4684
rect 19751 4644 19984 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 20990 4672 20996 4684
rect 20947 4644 20996 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 21542 4632 21548 4684
rect 21600 4672 21606 4684
rect 22005 4675 22063 4681
rect 22005 4672 22017 4675
rect 21600 4644 22017 4672
rect 21600 4632 21606 4644
rect 22005 4641 22017 4644
rect 22051 4672 22063 4675
rect 23658 4672 23664 4684
rect 22051 4644 23664 4672
rect 22051 4641 22063 4644
rect 22005 4635 22063 4641
rect 23658 4632 23664 4644
rect 23716 4632 23722 4684
rect 10137 4607 10195 4613
rect 10137 4573 10149 4607
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 9766 4496 9772 4548
rect 9824 4536 9830 4548
rect 10152 4536 10180 4567
rect 10686 4564 10692 4616
rect 10744 4604 10750 4616
rect 11425 4607 11483 4613
rect 11425 4604 11437 4607
rect 10744 4576 11437 4604
rect 10744 4564 10750 4576
rect 11425 4573 11437 4576
rect 11471 4604 11483 4607
rect 12342 4604 12348 4616
rect 11471 4576 12348 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 12342 4564 12348 4576
rect 12400 4604 12406 4616
rect 12526 4604 12532 4616
rect 12400 4576 12532 4604
rect 12400 4564 12406 4576
rect 12526 4564 12532 4576
rect 12584 4604 12590 4616
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 12584 4576 12633 4604
rect 12584 4564 12590 4576
rect 12621 4573 12633 4576
rect 12667 4573 12679 4607
rect 12621 4567 12679 4573
rect 14645 4607 14703 4613
rect 14645 4573 14657 4607
rect 14691 4604 14703 4607
rect 15102 4604 15108 4616
rect 14691 4576 15108 4604
rect 14691 4573 14703 4576
rect 14645 4567 14703 4573
rect 15102 4564 15108 4576
rect 15160 4604 15166 4616
rect 15289 4607 15347 4613
rect 15289 4604 15301 4607
rect 15160 4576 15301 4604
rect 15160 4564 15166 4576
rect 15289 4573 15301 4576
rect 15335 4573 15347 4607
rect 15289 4567 15347 4573
rect 10962 4536 10968 4548
rect 9824 4508 10968 4536
rect 9824 4496 9830 4508
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 8202 4468 8208 4480
rect 8163 4440 8208 4468
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 9030 4468 9036 4480
rect 8720 4440 9036 4468
rect 8720 4428 8726 4440
rect 9030 4428 9036 4440
rect 9088 4428 9094 4480
rect 10686 4468 10692 4480
rect 10647 4440 10692 4468
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 15304 4468 15332 4567
rect 17954 4564 17960 4616
rect 18012 4604 18018 4616
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 18012 4576 18245 4604
rect 18012 4564 18018 4576
rect 18233 4573 18245 4576
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 18417 4607 18475 4613
rect 18417 4573 18429 4607
rect 18463 4604 18475 4607
rect 18506 4604 18512 4616
rect 18463 4576 18512 4604
rect 18463 4573 18475 4576
rect 18417 4567 18475 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 19426 4604 19432 4616
rect 19339 4576 19432 4604
rect 19426 4564 19432 4576
rect 19484 4604 19490 4616
rect 20070 4604 20076 4616
rect 19484 4576 20076 4604
rect 19484 4564 19490 4576
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 25130 4604 25136 4616
rect 25091 4576 25136 4604
rect 25130 4564 25136 4576
rect 25188 4564 25194 4616
rect 19978 4496 19984 4548
rect 20036 4536 20042 4548
rect 21085 4539 21143 4545
rect 21085 4536 21097 4539
rect 20036 4508 21097 4536
rect 20036 4496 20042 4508
rect 21085 4505 21097 4508
rect 21131 4505 21143 4539
rect 21085 4499 21143 4505
rect 16206 4468 16212 4480
rect 15304 4440 16212 4468
rect 16206 4428 16212 4440
rect 16264 4468 16270 4480
rect 16666 4468 16672 4480
rect 16264 4440 16672 4468
rect 16264 4428 16270 4440
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 17313 4471 17371 4477
rect 17313 4437 17325 4471
rect 17359 4468 17371 4471
rect 17862 4468 17868 4480
rect 17359 4440 17868 4468
rect 17359 4437 17371 4440
rect 17313 4431 17371 4437
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 19886 4468 19892 4480
rect 19847 4440 19892 4468
rect 19886 4428 19892 4440
rect 19944 4428 19950 4480
rect 20254 4468 20260 4480
rect 20215 4440 20260 4468
rect 20254 4428 20260 4440
rect 20312 4428 20318 4480
rect 21821 4471 21879 4477
rect 21821 4437 21833 4471
rect 21867 4468 21879 4471
rect 22002 4468 22008 4480
rect 21867 4440 22008 4468
rect 21867 4437 21879 4440
rect 21821 4431 21879 4437
rect 22002 4428 22008 4440
rect 22060 4428 22066 4480
rect 23658 4428 23664 4480
rect 23716 4468 23722 4480
rect 25590 4468 25596 4480
rect 23716 4440 25596 4468
rect 23716 4428 23722 4440
rect 25590 4428 25596 4440
rect 25648 4428 25654 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 10778 4264 10784 4276
rect 8864 4236 10784 4264
rect 8202 4156 8208 4208
rect 8260 4196 8266 4208
rect 8864 4196 8892 4236
rect 10778 4224 10784 4236
rect 10836 4264 10842 4276
rect 11057 4267 11115 4273
rect 11057 4264 11069 4267
rect 10836 4236 11069 4264
rect 10836 4224 10842 4236
rect 11057 4233 11069 4236
rect 11103 4233 11115 4267
rect 15930 4264 15936 4276
rect 15891 4236 15936 4264
rect 11057 4227 11115 4233
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 17129 4267 17187 4273
rect 17129 4233 17141 4267
rect 17175 4264 17187 4267
rect 17218 4264 17224 4276
rect 17175 4236 17224 4264
rect 17175 4233 17187 4236
rect 17129 4227 17187 4233
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 19518 4264 19524 4276
rect 19479 4236 19524 4264
rect 19518 4224 19524 4236
rect 19576 4224 19582 4276
rect 20990 4264 20996 4276
rect 20951 4236 20996 4264
rect 20990 4224 20996 4236
rect 21048 4224 21054 4276
rect 23014 4224 23020 4276
rect 23072 4264 23078 4276
rect 23109 4267 23167 4273
rect 23109 4264 23121 4267
rect 23072 4236 23121 4264
rect 23072 4224 23078 4236
rect 23109 4233 23121 4236
rect 23155 4233 23167 4267
rect 23109 4227 23167 4233
rect 25222 4224 25228 4276
rect 25280 4264 25286 4276
rect 25869 4267 25927 4273
rect 25869 4264 25881 4267
rect 25280 4236 25881 4264
rect 25280 4224 25286 4236
rect 25869 4233 25881 4236
rect 25915 4233 25927 4267
rect 25869 4227 25927 4233
rect 23382 4196 23388 4208
rect 8260 4168 8892 4196
rect 20088 4168 23388 4196
rect 8260 4156 8266 4168
rect 8772 4137 8800 4168
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4097 8815 4131
rect 9490 4128 9496 4140
rect 9451 4100 9496 4128
rect 8757 4091 8815 4097
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 12066 4088 12072 4140
rect 12124 4128 12130 4140
rect 12161 4131 12219 4137
rect 12161 4128 12173 4131
rect 12124 4100 12173 4128
rect 12124 4088 12130 4100
rect 12161 4097 12173 4100
rect 12207 4097 12219 4131
rect 12161 4091 12219 4097
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 8067 4032 8493 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8481 4029 8493 4032
rect 8527 4060 8539 4063
rect 8570 4060 8576 4072
rect 8527 4032 8576 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 9030 4020 9036 4072
rect 9088 4060 9094 4072
rect 9582 4060 9588 4072
rect 9088 4032 9588 4060
rect 9088 4020 9094 4032
rect 9582 4020 9588 4032
rect 9640 4060 9646 4072
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9640 4032 9689 4060
rect 9640 4020 9646 4032
rect 9677 4029 9689 4032
rect 9723 4060 9735 4063
rect 10686 4060 10692 4072
rect 9723 4032 10692 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 12176 4060 12204 4091
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 13081 4131 13139 4137
rect 13081 4128 13093 4131
rect 13044 4100 13093 4128
rect 13044 4088 13050 4100
rect 13081 4097 13093 4100
rect 13127 4097 13139 4131
rect 14918 4128 14924 4140
rect 14879 4100 14924 4128
rect 13081 4091 13139 4097
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 15473 4131 15531 4137
rect 15473 4097 15485 4131
rect 15519 4128 15531 4131
rect 15562 4128 15568 4140
rect 15519 4100 15568 4128
rect 15519 4097 15531 4100
rect 15473 4091 15531 4097
rect 15562 4088 15568 4100
rect 15620 4128 15626 4140
rect 16482 4128 16488 4140
rect 15620 4100 16488 4128
rect 15620 4088 15626 4100
rect 16482 4088 16488 4100
rect 16540 4088 16546 4140
rect 17402 4128 17408 4140
rect 17363 4100 17408 4128
rect 17402 4088 17408 4100
rect 17460 4088 17466 4140
rect 18046 4088 18052 4140
rect 18104 4128 18110 4140
rect 18509 4131 18567 4137
rect 18509 4128 18521 4131
rect 18104 4100 18521 4128
rect 18104 4088 18110 4100
rect 18509 4097 18521 4100
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 18598 4088 18604 4140
rect 18656 4128 18662 4140
rect 20088 4137 20116 4168
rect 23382 4156 23388 4168
rect 23440 4156 23446 4208
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 18656 4100 18701 4128
rect 19904 4100 20085 4128
rect 18656 4088 18662 4100
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12176 4032 12909 4060
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 13909 4063 13967 4069
rect 13909 4029 13921 4063
rect 13955 4060 13967 4063
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 13955 4032 14841 4060
rect 13955 4029 13967 4032
rect 13909 4023 13967 4029
rect 14829 4029 14841 4032
rect 14875 4060 14887 4063
rect 15930 4060 15936 4072
rect 14875 4032 15936 4060
rect 14875 4029 14887 4032
rect 14829 4023 14887 4029
rect 15930 4020 15936 4032
rect 15988 4060 15994 4072
rect 16393 4063 16451 4069
rect 16393 4060 16405 4063
rect 15988 4032 16405 4060
rect 15988 4020 15994 4032
rect 16393 4029 16405 4032
rect 16439 4029 16451 4063
rect 16393 4023 16451 4029
rect 18138 4020 18144 4072
rect 18196 4060 18202 4072
rect 18690 4060 18696 4072
rect 18196 4032 18696 4060
rect 18196 4020 18202 4032
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 7668 3964 8616 3992
rect 7668 3936 7696 3964
rect 7650 3924 7656 3936
rect 7611 3896 7656 3924
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 8588 3933 8616 3964
rect 9490 3952 9496 4004
rect 9548 3992 9554 4004
rect 9922 3995 9980 4001
rect 9922 3992 9934 3995
rect 9548 3964 9934 3992
rect 9548 3952 9554 3964
rect 9922 3961 9934 3964
rect 9968 3961 9980 3995
rect 9922 3955 9980 3961
rect 11885 3995 11943 4001
rect 11885 3961 11897 3995
rect 11931 3992 11943 3995
rect 12066 3992 12072 4004
rect 11931 3964 12072 3992
rect 11931 3961 11943 3964
rect 11885 3955 11943 3961
rect 12066 3952 12072 3964
rect 12124 3992 12130 4004
rect 12989 3995 13047 4001
rect 12989 3992 13001 3995
rect 12124 3964 13001 3992
rect 12124 3952 12130 3964
rect 12989 3961 13001 3964
rect 13035 3992 13047 3995
rect 13078 3992 13084 4004
rect 13035 3964 13084 3992
rect 13035 3961 13047 3964
rect 12989 3955 13047 3961
rect 13078 3952 13084 3964
rect 13136 3952 13142 4004
rect 14737 3995 14795 4001
rect 14737 3992 14749 3995
rect 14200 3964 14749 3992
rect 14200 3936 14228 3964
rect 14737 3961 14749 3964
rect 14783 3961 14795 3995
rect 16301 3995 16359 4001
rect 16301 3992 16313 3995
rect 14737 3955 14795 3961
rect 15764 3964 16313 3992
rect 8573 3927 8631 3933
rect 8573 3893 8585 3927
rect 8619 3893 8631 3927
rect 8573 3887 8631 3893
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 9217 3927 9275 3933
rect 9217 3924 9229 3927
rect 8812 3896 9229 3924
rect 8812 3884 8818 3896
rect 9217 3893 9229 3896
rect 9263 3924 9275 3927
rect 9766 3924 9772 3936
rect 9263 3896 9772 3924
rect 9263 3893 9275 3896
rect 9217 3887 9275 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12529 3927 12587 3933
rect 12529 3924 12541 3927
rect 12492 3896 12541 3924
rect 12492 3884 12498 3896
rect 12529 3893 12541 3896
rect 12575 3893 12587 3927
rect 14182 3924 14188 3936
rect 14143 3896 14188 3924
rect 12529 3887 12587 3893
rect 14182 3884 14188 3896
rect 14240 3884 14246 3936
rect 14366 3924 14372 3936
rect 14327 3896 14372 3924
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 15654 3884 15660 3936
rect 15712 3924 15718 3936
rect 15764 3933 15792 3964
rect 16301 3961 16313 3964
rect 16347 3961 16359 3995
rect 16301 3955 16359 3961
rect 17862 3952 17868 4004
rect 17920 3992 17926 4004
rect 19150 3992 19156 4004
rect 17920 3964 18460 3992
rect 19063 3964 19156 3992
rect 17920 3952 17926 3964
rect 18432 3936 18460 3964
rect 19150 3952 19156 3964
rect 19208 3992 19214 4004
rect 19904 3992 19932 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20254 4128 20260 4140
rect 20215 4100 20260 4128
rect 20073 4091 20131 4097
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 22370 4128 22376 4140
rect 22331 4100 22376 4128
rect 22370 4088 22376 4100
rect 22428 4128 22434 4140
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 22428 4100 22753 4128
rect 22428 4088 22434 4100
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 22741 4091 22799 4097
rect 19981 4063 20039 4069
rect 19981 4029 19993 4063
rect 20027 4060 20039 4063
rect 20162 4060 20168 4072
rect 20027 4032 20168 4060
rect 20027 4029 20039 4032
rect 19981 4023 20039 4029
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 23290 4020 23296 4072
rect 23348 4060 23354 4072
rect 23934 4060 23940 4072
rect 23348 4032 23940 4060
rect 23348 4020 23354 4032
rect 23934 4020 23940 4032
rect 23992 4020 23998 4072
rect 24210 4069 24216 4072
rect 24204 4060 24216 4069
rect 24171 4032 24216 4060
rect 24204 4023 24216 4032
rect 24210 4020 24216 4023
rect 24268 4020 24274 4072
rect 22189 3995 22247 4001
rect 22189 3992 22201 3995
rect 19208 3964 19932 3992
rect 21560 3964 22201 3992
rect 19208 3952 19214 3964
rect 15749 3927 15807 3933
rect 15749 3924 15761 3927
rect 15712 3896 15761 3924
rect 15712 3884 15718 3896
rect 15749 3893 15761 3896
rect 15795 3893 15807 3927
rect 15749 3887 15807 3893
rect 17586 3884 17592 3936
rect 17644 3924 17650 3936
rect 17773 3927 17831 3933
rect 17773 3924 17785 3927
rect 17644 3896 17785 3924
rect 17644 3884 17650 3896
rect 17773 3893 17785 3896
rect 17819 3924 17831 3927
rect 17954 3924 17960 3936
rect 17819 3896 17960 3924
rect 17819 3893 17831 3896
rect 17773 3887 17831 3893
rect 17954 3884 17960 3896
rect 18012 3884 18018 3936
rect 18049 3927 18107 3933
rect 18049 3893 18061 3927
rect 18095 3924 18107 3927
rect 18138 3924 18144 3936
rect 18095 3896 18144 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 18414 3924 18420 3936
rect 18375 3896 18420 3924
rect 18414 3884 18420 3896
rect 18472 3884 18478 3936
rect 19518 3884 19524 3936
rect 19576 3924 19582 3936
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 19576 3896 19625 3924
rect 19576 3884 19582 3896
rect 19613 3893 19625 3896
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 21450 3884 21456 3936
rect 21508 3924 21514 3936
rect 21560 3933 21588 3964
rect 22189 3961 22201 3964
rect 22235 3961 22247 3995
rect 22189 3955 22247 3961
rect 21545 3927 21603 3933
rect 21545 3924 21557 3927
rect 21508 3896 21557 3924
rect 21508 3884 21514 3896
rect 21545 3893 21557 3896
rect 21591 3893 21603 3927
rect 21545 3887 21603 3893
rect 21634 3884 21640 3936
rect 21692 3924 21698 3936
rect 21729 3927 21787 3933
rect 21729 3924 21741 3927
rect 21692 3896 21741 3924
rect 21692 3884 21698 3896
rect 21729 3893 21741 3896
rect 21775 3893 21787 3927
rect 21729 3887 21787 3893
rect 22002 3884 22008 3936
rect 22060 3924 22066 3936
rect 22094 3924 22100 3936
rect 22060 3896 22100 3924
rect 22060 3884 22066 3896
rect 22094 3884 22100 3896
rect 22152 3924 22158 3936
rect 25314 3924 25320 3936
rect 22152 3896 22245 3924
rect 25275 3896 25320 3924
rect 22152 3884 22158 3896
rect 25314 3884 25320 3896
rect 25372 3884 25378 3936
rect 26234 3924 26240 3936
rect 26195 3896 26240 3924
rect 26234 3884 26240 3896
rect 26292 3884 26298 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 7006 3720 7012 3732
rect 6967 3692 7012 3720
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7650 3680 7656 3732
rect 7708 3720 7714 3732
rect 8021 3723 8079 3729
rect 8021 3720 8033 3723
rect 7708 3692 8033 3720
rect 7708 3680 7714 3692
rect 8021 3689 8033 3692
rect 8067 3689 8079 3723
rect 9950 3720 9956 3732
rect 9911 3692 9956 3720
rect 8021 3683 8079 3689
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 10965 3723 11023 3729
rect 10965 3720 10977 3723
rect 10744 3692 10977 3720
rect 10744 3680 10750 3692
rect 10965 3689 10977 3692
rect 11011 3720 11023 3723
rect 11011 3692 11468 3720
rect 11011 3689 11023 3692
rect 10965 3683 11023 3689
rect 7561 3655 7619 3661
rect 7561 3621 7573 3655
rect 7607 3652 7619 3655
rect 8478 3652 8484 3664
rect 7607 3624 8484 3652
rect 7607 3621 7619 3624
rect 7561 3615 7619 3621
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 8386 3584 8392 3596
rect 8347 3556 8392 3584
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 8754 3584 8760 3596
rect 8496 3556 8760 3584
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 8496 3525 8524 3556
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 9306 3544 9312 3596
rect 9364 3584 9370 3596
rect 10321 3587 10379 3593
rect 10321 3584 10333 3587
rect 9364 3556 10333 3584
rect 9364 3544 9370 3556
rect 10321 3553 10333 3556
rect 10367 3553 10379 3587
rect 10962 3584 10968 3596
rect 10321 3547 10379 3553
rect 10428 3556 10968 3584
rect 10428 3525 10456 3556
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 8481 3519 8539 3525
rect 8481 3516 8493 3519
rect 7524 3488 8493 3516
rect 7524 3476 7530 3488
rect 8481 3485 8493 3488
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 8665 3519 8723 3525
rect 8665 3485 8677 3519
rect 8711 3485 8723 3519
rect 8665 3479 8723 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3516 9183 3519
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 9171 3488 10425 3516
rect 9171 3485 9183 3488
rect 9125 3479 9183 3485
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3516 10655 3519
rect 11054 3516 11060 3528
rect 10643 3488 11060 3516
rect 10643 3485 10655 3488
rect 10597 3479 10655 3485
rect 8680 3448 8708 3479
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 11440 3516 11468 3692
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 13909 3723 13967 3729
rect 13909 3720 13921 3723
rect 13136 3692 13921 3720
rect 13136 3680 13142 3692
rect 13909 3689 13921 3692
rect 13955 3720 13967 3723
rect 14366 3720 14372 3732
rect 13955 3692 14372 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 15105 3723 15163 3729
rect 15105 3689 15117 3723
rect 15151 3720 15163 3723
rect 15562 3720 15568 3732
rect 15151 3692 15568 3720
rect 15151 3689 15163 3692
rect 15105 3683 15163 3689
rect 15562 3680 15568 3692
rect 15620 3680 15626 3732
rect 15930 3720 15936 3732
rect 15891 3692 15936 3720
rect 15930 3680 15936 3692
rect 15988 3680 15994 3732
rect 20162 3720 20168 3732
rect 20123 3692 20168 3720
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 21082 3720 21088 3732
rect 21043 3692 21088 3720
rect 21082 3680 21088 3692
rect 21140 3680 21146 3732
rect 22925 3723 22983 3729
rect 22925 3689 22937 3723
rect 22971 3720 22983 3723
rect 23014 3720 23020 3732
rect 22971 3692 23020 3720
rect 22971 3689 22983 3692
rect 22925 3683 22983 3689
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 23474 3680 23480 3732
rect 23532 3720 23538 3732
rect 24029 3723 24087 3729
rect 24029 3720 24041 3723
rect 23532 3692 24041 3720
rect 23532 3680 23538 3692
rect 24029 3689 24041 3692
rect 24075 3689 24087 3723
rect 24029 3683 24087 3689
rect 24118 3680 24124 3732
rect 24176 3720 24182 3732
rect 24489 3723 24547 3729
rect 24489 3720 24501 3723
rect 24176 3692 24501 3720
rect 24176 3680 24182 3692
rect 24489 3689 24501 3692
rect 24535 3720 24547 3723
rect 24670 3720 24676 3732
rect 24535 3692 24676 3720
rect 24535 3689 24547 3692
rect 24489 3683 24547 3689
rect 24670 3680 24676 3692
rect 24728 3680 24734 3732
rect 24762 3680 24768 3732
rect 24820 3720 24826 3732
rect 25038 3720 25044 3732
rect 24820 3692 25044 3720
rect 24820 3680 24826 3692
rect 25038 3680 25044 3692
rect 25096 3680 25102 3732
rect 25590 3680 25596 3732
rect 25648 3720 25654 3732
rect 25777 3723 25835 3729
rect 25777 3720 25789 3723
rect 25648 3692 25789 3720
rect 25648 3680 25654 3692
rect 25777 3689 25789 3692
rect 25823 3689 25835 3723
rect 25777 3683 25835 3689
rect 11514 3612 11520 3664
rect 11572 3652 11578 3664
rect 11762 3655 11820 3661
rect 11762 3652 11774 3655
rect 11572 3624 11774 3652
rect 11572 3612 11578 3624
rect 11762 3621 11774 3624
rect 11808 3621 11820 3655
rect 11762 3615 11820 3621
rect 12986 3612 12992 3664
rect 13044 3652 13050 3664
rect 13449 3655 13507 3661
rect 13449 3652 13461 3655
rect 13044 3624 13461 3652
rect 13044 3612 13050 3624
rect 13449 3621 13461 3624
rect 13495 3621 13507 3655
rect 19518 3652 19524 3664
rect 19431 3624 19524 3652
rect 13449 3615 13507 3621
rect 19518 3612 19524 3624
rect 19576 3652 19582 3664
rect 20533 3655 20591 3661
rect 20533 3652 20545 3655
rect 19576 3624 20545 3652
rect 19576 3612 19582 3624
rect 20533 3621 20545 3624
rect 20579 3621 20591 3655
rect 20533 3615 20591 3621
rect 22186 3612 22192 3664
rect 22244 3652 22250 3664
rect 22244 3624 22416 3652
rect 22244 3612 22250 3624
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 14001 3587 14059 3593
rect 14001 3584 14013 3587
rect 13780 3556 14013 3584
rect 13780 3544 13786 3556
rect 14001 3553 14013 3556
rect 14047 3584 14059 3587
rect 14274 3584 14280 3596
rect 14047 3556 14280 3584
rect 14047 3553 14059 3556
rect 14001 3547 14059 3553
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 15470 3584 15476 3596
rect 15335 3556 15476 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 16574 3544 16580 3596
rect 16632 3584 16638 3596
rect 16741 3587 16799 3593
rect 16741 3584 16753 3587
rect 16632 3556 16753 3584
rect 16632 3544 16638 3556
rect 16741 3553 16753 3556
rect 16787 3553 16799 3587
rect 16741 3547 16799 3553
rect 19061 3587 19119 3593
rect 19061 3553 19073 3587
rect 19107 3584 19119 3587
rect 19613 3587 19671 3593
rect 19613 3584 19625 3587
rect 19107 3556 19625 3584
rect 19107 3553 19119 3556
rect 19061 3547 19119 3553
rect 19613 3553 19625 3556
rect 19659 3584 19671 3587
rect 20622 3584 20628 3596
rect 19659 3556 20628 3584
rect 19659 3553 19671 3556
rect 19613 3547 19671 3553
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 21542 3584 21548 3596
rect 21503 3556 21548 3584
rect 21542 3544 21548 3556
rect 21600 3544 21606 3596
rect 21812 3587 21870 3593
rect 21812 3553 21824 3587
rect 21858 3584 21870 3587
rect 22278 3584 22284 3596
rect 21858 3556 22284 3584
rect 21858 3553 21870 3556
rect 21812 3547 21870 3553
rect 22278 3544 22284 3556
rect 22336 3544 22342 3596
rect 22388 3584 22416 3624
rect 23198 3612 23204 3664
rect 23256 3652 23262 3664
rect 23661 3655 23719 3661
rect 23661 3652 23673 3655
rect 23256 3624 23673 3652
rect 23256 3612 23262 3624
rect 23661 3621 23673 3624
rect 23707 3652 23719 3655
rect 23842 3652 23848 3664
rect 23707 3624 23848 3652
rect 23707 3621 23719 3624
rect 23661 3615 23719 3621
rect 23842 3612 23848 3624
rect 23900 3612 23906 3664
rect 23934 3612 23940 3664
rect 23992 3652 23998 3664
rect 25409 3655 25467 3661
rect 25409 3652 25421 3655
rect 23992 3624 25421 3652
rect 23992 3612 23998 3624
rect 25409 3621 25421 3624
rect 25455 3652 25467 3655
rect 26142 3652 26148 3664
rect 25455 3624 26148 3652
rect 25455 3621 25467 3624
rect 25409 3615 25467 3621
rect 26142 3612 26148 3624
rect 26200 3612 26206 3664
rect 24397 3587 24455 3593
rect 24397 3584 24409 3587
rect 22388 3556 24409 3584
rect 24397 3553 24409 3556
rect 24443 3584 24455 3587
rect 25038 3584 25044 3596
rect 24443 3556 25044 3584
rect 24443 3553 24455 3556
rect 24397 3547 24455 3553
rect 25038 3544 25044 3556
rect 25096 3544 25102 3596
rect 11517 3519 11575 3525
rect 11517 3516 11529 3519
rect 11440 3488 11529 3516
rect 11517 3485 11529 3488
rect 11563 3485 11575 3519
rect 16485 3519 16543 3525
rect 16485 3516 16497 3519
rect 11517 3479 11575 3485
rect 16316 3488 16497 3516
rect 14645 3451 14703 3457
rect 8680 3420 9536 3448
rect 9508 3392 9536 3420
rect 14645 3417 14657 3451
rect 14691 3448 14703 3451
rect 14918 3448 14924 3460
rect 14691 3420 14924 3448
rect 14691 3417 14703 3420
rect 14645 3411 14703 3417
rect 14918 3408 14924 3420
rect 14976 3448 14982 3460
rect 15562 3448 15568 3460
rect 14976 3420 15568 3448
rect 14976 3408 14982 3420
rect 15562 3408 15568 3420
rect 15620 3408 15626 3460
rect 7929 3383 7987 3389
rect 7929 3349 7941 3383
rect 7975 3380 7987 3383
rect 8570 3380 8576 3392
rect 7975 3352 8576 3380
rect 7975 3349 7987 3352
rect 7929 3343 7987 3349
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 9490 3380 9496 3392
rect 9451 3352 9496 3380
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 11425 3383 11483 3389
rect 11425 3349 11437 3383
rect 11471 3380 11483 3383
rect 11514 3380 11520 3392
rect 11471 3352 11520 3380
rect 11471 3349 11483 3352
rect 11425 3343 11483 3349
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 12897 3383 12955 3389
rect 12897 3380 12909 3383
rect 11756 3352 12909 3380
rect 11756 3340 11762 3352
rect 12897 3349 12909 3352
rect 12943 3349 12955 3383
rect 12897 3343 12955 3349
rect 13906 3340 13912 3392
rect 13964 3380 13970 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 13964 3352 14197 3380
rect 13964 3340 13970 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 14185 3343 14243 3349
rect 15286 3340 15292 3392
rect 15344 3380 15350 3392
rect 15473 3383 15531 3389
rect 15473 3380 15485 3383
rect 15344 3352 15485 3380
rect 15344 3340 15350 3352
rect 15473 3349 15485 3352
rect 15519 3349 15531 3383
rect 15473 3343 15531 3349
rect 16206 3340 16212 3392
rect 16264 3380 16270 3392
rect 16316 3389 16344 3488
rect 16485 3485 16497 3488
rect 16531 3485 16543 3519
rect 19794 3516 19800 3528
rect 19755 3488 19800 3516
rect 16485 3479 16543 3485
rect 19794 3476 19800 3488
rect 19852 3476 19858 3528
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3516 24731 3519
rect 25130 3516 25136 3528
rect 24719 3488 25136 3516
rect 24719 3485 24731 3488
rect 24673 3479 24731 3485
rect 25130 3476 25136 3488
rect 25188 3516 25194 3528
rect 26234 3516 26240 3528
rect 25188 3488 26240 3516
rect 25188 3476 25194 3488
rect 26234 3476 26240 3488
rect 26292 3476 26298 3528
rect 19150 3448 19156 3460
rect 19111 3420 19156 3448
rect 19150 3408 19156 3420
rect 19208 3408 19214 3460
rect 23934 3408 23940 3460
rect 23992 3448 23998 3460
rect 24578 3448 24584 3460
rect 23992 3420 24584 3448
rect 23992 3408 23998 3420
rect 24578 3408 24584 3420
rect 24636 3408 24642 3460
rect 16301 3383 16359 3389
rect 16301 3380 16313 3383
rect 16264 3352 16313 3380
rect 16264 3340 16270 3352
rect 16301 3349 16313 3352
rect 16347 3349 16359 3383
rect 17862 3380 17868 3392
rect 17823 3352 17868 3380
rect 16301 3343 16359 3349
rect 17862 3340 17868 3352
rect 17920 3380 17926 3392
rect 18417 3383 18475 3389
rect 18417 3380 18429 3383
rect 17920 3352 18429 3380
rect 17920 3340 17926 3352
rect 18417 3349 18429 3352
rect 18463 3380 18475 3383
rect 18598 3380 18604 3392
rect 18463 3352 18604 3380
rect 18463 3349 18475 3352
rect 18417 3343 18475 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 21082 3340 21088 3392
rect 21140 3380 21146 3392
rect 21910 3380 21916 3392
rect 21140 3352 21916 3380
rect 21140 3340 21146 3352
rect 21910 3340 21916 3352
rect 21968 3340 21974 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 7466 3176 7472 3188
rect 7427 3148 7472 3176
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 8018 3176 8024 3188
rect 7883 3148 8024 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 8018 3136 8024 3148
rect 8076 3176 8082 3188
rect 8386 3176 8392 3188
rect 8076 3148 8392 3176
rect 8076 3136 8082 3148
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 9033 3179 9091 3185
rect 9033 3145 9045 3179
rect 9079 3176 9091 3179
rect 9490 3176 9496 3188
rect 9079 3148 9496 3176
rect 9079 3145 9091 3148
rect 9033 3139 9091 3145
rect 9490 3136 9496 3148
rect 9548 3176 9554 3188
rect 10873 3179 10931 3185
rect 10873 3176 10885 3179
rect 9548 3148 10885 3176
rect 9548 3136 9554 3148
rect 10873 3145 10885 3148
rect 10919 3145 10931 3179
rect 10873 3139 10931 3145
rect 11054 3136 11060 3188
rect 11112 3176 11118 3188
rect 11517 3179 11575 3185
rect 11517 3176 11529 3179
rect 11112 3148 11529 3176
rect 11112 3136 11118 3148
rect 11517 3145 11529 3148
rect 11563 3176 11575 3179
rect 11698 3176 11704 3188
rect 11563 3148 11704 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 12618 3176 12624 3188
rect 12579 3148 12624 3176
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 13722 3176 13728 3188
rect 13683 3148 13728 3176
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 15470 3136 15476 3188
rect 15528 3176 15534 3188
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 15528 3148 16129 3176
rect 15528 3136 15534 3148
rect 16117 3145 16129 3148
rect 16163 3145 16175 3179
rect 16117 3139 16175 3145
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 19794 3176 19800 3188
rect 19576 3148 19800 3176
rect 19576 3136 19582 3148
rect 19794 3136 19800 3148
rect 19852 3176 19858 3188
rect 20073 3179 20131 3185
rect 20073 3176 20085 3179
rect 19852 3148 20085 3176
rect 19852 3136 19858 3148
rect 20073 3145 20085 3148
rect 20119 3176 20131 3179
rect 21913 3179 21971 3185
rect 21913 3176 21925 3179
rect 20119 3148 21925 3176
rect 20119 3145 20131 3148
rect 20073 3139 20131 3145
rect 21913 3145 21925 3148
rect 21959 3145 21971 3179
rect 21913 3139 21971 3145
rect 22278 3136 22284 3188
rect 22336 3176 22342 3188
rect 22465 3179 22523 3185
rect 22465 3176 22477 3179
rect 22336 3148 22477 3176
rect 22336 3136 22342 3148
rect 22465 3145 22477 3148
rect 22511 3176 22523 3179
rect 23293 3179 23351 3185
rect 23293 3176 23305 3179
rect 22511 3148 23305 3176
rect 22511 3145 22523 3148
rect 22465 3139 22523 3145
rect 23293 3145 23305 3148
rect 23339 3145 23351 3179
rect 23658 3176 23664 3188
rect 23619 3148 23664 3176
rect 23293 3139 23351 3145
rect 23658 3136 23664 3148
rect 23716 3136 23722 3188
rect 24670 3176 24676 3188
rect 24631 3148 24676 3176
rect 24670 3136 24676 3148
rect 24728 3136 24734 3188
rect 25130 3176 25136 3188
rect 25091 3148 25136 3176
rect 25130 3136 25136 3148
rect 25188 3136 25194 3188
rect 26142 3176 26148 3188
rect 26103 3148 26148 3176
rect 26142 3136 26148 3148
rect 26200 3136 26206 3188
rect 7926 3108 7932 3120
rect 7887 3080 7932 3108
rect 7926 3068 7932 3080
rect 7984 3068 7990 3120
rect 19429 3111 19487 3117
rect 19429 3077 19441 3111
rect 19475 3077 19487 3111
rect 19429 3071 19487 3077
rect 25869 3111 25927 3117
rect 25869 3077 25881 3111
rect 25915 3108 25927 3111
rect 26234 3108 26240 3120
rect 25915 3080 26240 3108
rect 25915 3077 25927 3080
rect 25869 3071 25927 3077
rect 8570 3040 8576 3052
rect 8531 3012 8576 3040
rect 8570 3000 8576 3012
rect 8628 3000 8634 3052
rect 9490 3040 9496 3052
rect 9451 3012 9496 3040
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 13078 3040 13084 3052
rect 13039 3012 13084 3040
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3040 13323 3043
rect 13354 3040 13360 3052
rect 13311 3012 13360 3040
rect 13311 3009 13323 3012
rect 13265 3003 13323 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 17770 3040 17776 3052
rect 17731 3012 17776 3040
rect 17770 3000 17776 3012
rect 17828 3040 17834 3052
rect 19444 3040 19472 3071
rect 26234 3068 26240 3080
rect 26292 3068 26298 3120
rect 19797 3043 19855 3049
rect 19797 3040 19809 3043
rect 17828 3012 18184 3040
rect 19444 3012 19809 3040
rect 17828 3000 17834 3012
rect 6917 2975 6975 2981
rect 6917 2941 6929 2975
rect 6963 2972 6975 2975
rect 9306 2972 9312 2984
rect 6963 2944 9312 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 9582 2932 9588 2984
rect 9640 2972 9646 2984
rect 9760 2975 9818 2981
rect 9760 2972 9772 2975
rect 9640 2944 9772 2972
rect 9640 2932 9646 2944
rect 9760 2941 9772 2944
rect 9806 2972 9818 2975
rect 11054 2972 11060 2984
rect 9806 2944 11060 2972
rect 9806 2941 9818 2944
rect 9760 2935 9818 2941
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 11790 2932 11796 2984
rect 11848 2972 11854 2984
rect 12161 2975 12219 2981
rect 12161 2972 12173 2975
rect 11848 2944 12173 2972
rect 11848 2932 11854 2944
rect 12161 2941 12173 2944
rect 12207 2972 12219 2975
rect 14185 2975 14243 2981
rect 12207 2944 12388 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 8389 2907 8447 2913
rect 8389 2873 8401 2907
rect 8435 2904 8447 2907
rect 8478 2904 8484 2916
rect 8435 2876 8484 2904
rect 8435 2873 8447 2876
rect 8389 2867 8447 2873
rect 8478 2864 8484 2876
rect 8536 2864 8542 2916
rect 11885 2907 11943 2913
rect 11885 2873 11897 2907
rect 11931 2904 11943 2907
rect 12360 2904 12388 2944
rect 14185 2941 14197 2975
rect 14231 2972 14243 2975
rect 16206 2972 16212 2984
rect 14231 2944 16212 2972
rect 14231 2941 14243 2944
rect 14185 2935 14243 2941
rect 16206 2932 16212 2944
rect 16264 2932 16270 2984
rect 16574 2972 16580 2984
rect 16487 2944 16580 2972
rect 16574 2932 16580 2944
rect 16632 2932 16638 2984
rect 16669 2975 16727 2981
rect 16669 2941 16681 2975
rect 16715 2972 16727 2975
rect 16758 2972 16764 2984
rect 16715 2944 16764 2972
rect 16715 2941 16727 2944
rect 16669 2935 16727 2941
rect 16758 2932 16764 2944
rect 16816 2972 16822 2984
rect 17221 2975 17279 2981
rect 17221 2972 17233 2975
rect 16816 2944 17233 2972
rect 16816 2932 16822 2944
rect 17221 2941 17233 2944
rect 17267 2941 17279 2975
rect 18046 2972 18052 2984
rect 18007 2944 18052 2972
rect 17221 2935 17279 2941
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18156 2972 18184 3012
rect 19797 3009 19809 3012
rect 19843 3040 19855 3043
rect 23109 3043 23167 3049
rect 19843 3012 20668 3040
rect 19843 3009 19855 3012
rect 19797 3003 19855 3009
rect 18305 2975 18363 2981
rect 18305 2972 18317 2975
rect 18156 2944 18317 2972
rect 18305 2941 18317 2944
rect 18351 2972 18363 2975
rect 20070 2972 20076 2984
rect 18351 2944 20076 2972
rect 18351 2941 18363 2944
rect 18305 2935 18363 2941
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 20530 2972 20536 2984
rect 20491 2944 20536 2972
rect 20530 2932 20536 2944
rect 20588 2932 20594 2984
rect 20640 2972 20668 3012
rect 23109 3009 23121 3043
rect 23155 3040 23167 3043
rect 24213 3043 24271 3049
rect 24213 3040 24225 3043
rect 23155 3012 24225 3040
rect 23155 3009 23167 3012
rect 23109 3003 23167 3009
rect 24213 3009 24225 3012
rect 24259 3009 24271 3043
rect 24213 3003 24271 3009
rect 23124 2972 23152 3003
rect 20640 2944 23152 2972
rect 23293 2975 23351 2981
rect 23293 2941 23305 2975
rect 23339 2972 23351 2975
rect 23566 2972 23572 2984
rect 23339 2944 23572 2972
rect 23339 2941 23351 2944
rect 23293 2935 23351 2941
rect 23566 2932 23572 2944
rect 23624 2932 23630 2984
rect 23842 2932 23848 2984
rect 23900 2972 23906 2984
rect 24029 2975 24087 2981
rect 24029 2972 24041 2975
rect 23900 2944 24041 2972
rect 23900 2932 23906 2944
rect 24029 2941 24041 2944
rect 24075 2941 24087 2975
rect 24029 2935 24087 2941
rect 12989 2907 13047 2913
rect 12989 2904 13001 2907
rect 11931 2876 12296 2904
rect 12360 2876 13001 2904
rect 11931 2873 11943 2876
rect 11885 2867 11943 2873
rect 6641 2839 6699 2845
rect 6641 2805 6653 2839
rect 6687 2836 6699 2839
rect 6822 2836 6828 2848
rect 6687 2808 6828 2836
rect 6687 2805 6699 2808
rect 6641 2799 6699 2805
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 8202 2796 8208 2848
rect 8260 2836 8266 2848
rect 8297 2839 8355 2845
rect 8297 2836 8309 2839
rect 8260 2808 8309 2836
rect 8260 2796 8266 2808
rect 8297 2805 8309 2808
rect 8343 2805 8355 2839
rect 12268 2836 12296 2876
rect 12989 2873 13001 2876
rect 13035 2873 13047 2907
rect 12989 2867 13047 2873
rect 14093 2907 14151 2913
rect 14093 2873 14105 2907
rect 14139 2904 14151 2907
rect 14430 2907 14488 2913
rect 14430 2904 14442 2907
rect 14139 2876 14442 2904
rect 14139 2873 14151 2876
rect 14093 2867 14151 2873
rect 14430 2873 14442 2876
rect 14476 2904 14488 2907
rect 15102 2904 15108 2916
rect 14476 2876 15108 2904
rect 14476 2873 14488 2876
rect 14430 2867 14488 2873
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 16592 2904 16620 2932
rect 17678 2904 17684 2916
rect 16592 2876 17684 2904
rect 17678 2864 17684 2876
rect 17736 2904 17742 2916
rect 19797 2907 19855 2913
rect 19797 2904 19809 2907
rect 17736 2876 19809 2904
rect 17736 2864 17742 2876
rect 19797 2873 19809 2876
rect 19843 2873 19855 2907
rect 19797 2867 19855 2873
rect 20254 2864 20260 2916
rect 20312 2904 20318 2916
rect 20441 2907 20499 2913
rect 20441 2904 20453 2907
rect 20312 2876 20453 2904
rect 20312 2864 20318 2876
rect 20441 2873 20453 2876
rect 20487 2904 20499 2907
rect 20800 2907 20858 2913
rect 20800 2904 20812 2907
rect 20487 2876 20812 2904
rect 20487 2873 20499 2876
rect 20441 2867 20499 2873
rect 20800 2873 20812 2876
rect 20846 2904 20858 2907
rect 21818 2904 21824 2916
rect 20846 2876 21824 2904
rect 20846 2873 20858 2876
rect 20800 2867 20858 2873
rect 21818 2864 21824 2876
rect 21876 2864 21882 2916
rect 23474 2904 23480 2916
rect 23387 2876 23480 2904
rect 23474 2864 23480 2876
rect 23532 2904 23538 2916
rect 24121 2907 24179 2913
rect 24121 2904 24133 2907
rect 23532 2876 24133 2904
rect 23532 2864 23538 2876
rect 24121 2873 24133 2876
rect 24167 2873 24179 2907
rect 24121 2867 24179 2873
rect 12434 2836 12440 2848
rect 12268 2808 12440 2836
rect 8297 2799 8355 2805
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 15562 2836 15568 2848
rect 15523 2808 15568 2836
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 16574 2796 16580 2848
rect 16632 2836 16638 2848
rect 16853 2839 16911 2845
rect 16853 2836 16865 2839
rect 16632 2808 16865 2836
rect 16632 2796 16638 2808
rect 16853 2805 16865 2808
rect 16899 2805 16911 2839
rect 16853 2799 16911 2805
rect 17310 2796 17316 2848
rect 17368 2836 17374 2848
rect 17770 2836 17776 2848
rect 17368 2808 17776 2836
rect 17368 2796 17374 2808
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 25406 2836 25412 2848
rect 25367 2808 25412 2836
rect 25406 2796 25412 2808
rect 25464 2796 25470 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 7098 2632 7104 2644
rect 7059 2604 7104 2632
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 8113 2635 8171 2641
rect 8113 2601 8125 2635
rect 8159 2632 8171 2635
rect 8202 2632 8208 2644
rect 8159 2604 8208 2632
rect 8159 2601 8171 2604
rect 8113 2595 8171 2601
rect 6914 2524 6920 2576
rect 6972 2564 6978 2576
rect 8128 2564 8156 2595
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 10505 2635 10563 2641
rect 10505 2601 10517 2635
rect 10551 2632 10563 2635
rect 10778 2632 10784 2644
rect 10551 2604 10784 2632
rect 10551 2601 10563 2604
rect 10505 2595 10563 2601
rect 6972 2536 8156 2564
rect 6972 2524 6978 2536
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 8478 2496 8484 2508
rect 7699 2468 8484 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 10520 2496 10548 2595
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 10962 2632 10968 2644
rect 10923 2604 10968 2632
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 11425 2635 11483 2641
rect 11425 2601 11437 2635
rect 11471 2632 11483 2635
rect 12066 2632 12072 2644
rect 11471 2604 12072 2632
rect 11471 2601 11483 2604
rect 11425 2595 11483 2601
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 15289 2635 15347 2641
rect 15289 2601 15301 2635
rect 15335 2632 15347 2635
rect 15562 2632 15568 2644
rect 15335 2604 15568 2632
rect 15335 2601 15347 2604
rect 15289 2595 15347 2601
rect 15562 2592 15568 2604
rect 15620 2592 15626 2644
rect 16850 2632 16856 2644
rect 16811 2604 16856 2632
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 19705 2635 19763 2641
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 20070 2632 20076 2644
rect 19751 2604 20076 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 20622 2592 20628 2644
rect 20680 2632 20686 2644
rect 21177 2635 21235 2641
rect 21177 2632 21189 2635
rect 20680 2604 21189 2632
rect 20680 2592 20686 2604
rect 21177 2601 21189 2604
rect 21223 2601 21235 2635
rect 21634 2632 21640 2644
rect 21595 2604 21640 2632
rect 21177 2595 21235 2601
rect 21634 2592 21640 2604
rect 21692 2592 21698 2644
rect 22278 2632 22284 2644
rect 22239 2604 22284 2632
rect 22278 2592 22284 2604
rect 22336 2592 22342 2644
rect 22649 2635 22707 2641
rect 22649 2601 22661 2635
rect 22695 2632 22707 2635
rect 23290 2632 23296 2644
rect 22695 2604 23296 2632
rect 22695 2601 22707 2604
rect 22649 2595 22707 2601
rect 12434 2564 12440 2576
rect 12347 2536 12440 2564
rect 12434 2524 12440 2536
rect 12492 2564 12498 2576
rect 12888 2567 12946 2573
rect 12888 2564 12900 2567
rect 12492 2536 12900 2564
rect 12492 2524 12498 2536
rect 12888 2533 12900 2536
rect 12934 2564 12946 2567
rect 13354 2564 13360 2576
rect 12934 2536 13360 2564
rect 12934 2533 12946 2536
rect 12888 2527 12946 2533
rect 13354 2524 13360 2536
rect 13412 2524 13418 2576
rect 15580 2564 15608 2592
rect 15718 2567 15776 2573
rect 15718 2564 15730 2567
rect 15580 2536 15730 2564
rect 15718 2533 15730 2536
rect 15764 2533 15776 2567
rect 15718 2527 15776 2533
rect 16206 2524 16212 2576
rect 16264 2564 16270 2576
rect 17405 2567 17463 2573
rect 17405 2564 17417 2567
rect 16264 2536 17417 2564
rect 16264 2524 16270 2536
rect 17405 2533 17417 2536
rect 17451 2533 17463 2567
rect 17405 2527 17463 2533
rect 19426 2524 19432 2576
rect 19484 2564 19490 2576
rect 20993 2567 21051 2573
rect 19484 2536 20668 2564
rect 19484 2524 19490 2536
rect 9907 2468 10548 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 10778 2456 10784 2508
rect 10836 2496 10842 2508
rect 11333 2499 11391 2505
rect 11333 2496 11345 2499
rect 10836 2468 11345 2496
rect 10836 2456 10842 2468
rect 11333 2465 11345 2468
rect 11379 2465 11391 2499
rect 11333 2459 11391 2465
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12584 2468 12633 2496
rect 12584 2456 12590 2468
rect 12621 2465 12633 2468
rect 12667 2496 12679 2499
rect 14553 2499 14611 2505
rect 14553 2496 14565 2499
rect 12667 2468 14565 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 14553 2465 14565 2468
rect 14599 2465 14611 2499
rect 14553 2459 14611 2465
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 16224 2496 16252 2524
rect 18581 2499 18639 2505
rect 18581 2496 18593 2499
rect 15519 2468 16252 2496
rect 18064 2468 18593 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 18064 2440 18092 2468
rect 18581 2465 18593 2468
rect 18627 2496 18639 2499
rect 19518 2496 19524 2508
rect 18627 2468 19524 2496
rect 18627 2465 18639 2468
rect 18581 2459 18639 2465
rect 19518 2456 19524 2468
rect 19576 2456 19582 2508
rect 20640 2505 20668 2536
rect 20993 2533 21005 2567
rect 21039 2564 21051 2567
rect 21652 2564 21680 2592
rect 21039 2536 21680 2564
rect 21039 2533 21051 2536
rect 20993 2527 21051 2533
rect 22002 2524 22008 2576
rect 22060 2564 22066 2576
rect 22664 2564 22692 2595
rect 23290 2592 23296 2604
rect 23348 2592 23354 2644
rect 23382 2592 23388 2644
rect 23440 2632 23446 2644
rect 23845 2635 23903 2641
rect 23845 2632 23857 2635
rect 23440 2604 23857 2632
rect 23440 2592 23446 2604
rect 23845 2601 23857 2604
rect 23891 2632 23903 2635
rect 23891 2604 24072 2632
rect 23891 2601 23903 2604
rect 23845 2595 23903 2601
rect 22060 2536 22692 2564
rect 23477 2567 23535 2573
rect 22060 2524 22066 2536
rect 23477 2533 23489 2567
rect 23523 2564 23535 2567
rect 23934 2564 23940 2576
rect 23523 2536 23940 2564
rect 23523 2533 23535 2536
rect 23477 2527 23535 2533
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 21542 2496 21548 2508
rect 20671 2468 21548 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 21542 2456 21548 2468
rect 21600 2496 21606 2508
rect 22094 2496 22100 2508
rect 21600 2468 22100 2496
rect 21600 2456 21606 2468
rect 22094 2456 22100 2468
rect 22152 2456 22158 2508
rect 22833 2499 22891 2505
rect 22833 2465 22845 2499
rect 22879 2496 22891 2499
rect 23492 2496 23520 2527
rect 23934 2524 23940 2536
rect 23992 2524 23998 2576
rect 24044 2564 24072 2604
rect 24210 2592 24216 2644
rect 24268 2632 24274 2644
rect 24397 2635 24455 2641
rect 24397 2632 24409 2635
rect 24268 2604 24409 2632
rect 24268 2592 24274 2604
rect 24397 2601 24409 2604
rect 24443 2632 24455 2635
rect 25133 2635 25191 2641
rect 25133 2632 25145 2635
rect 24443 2604 25145 2632
rect 24443 2601 24455 2604
rect 24397 2595 24455 2601
rect 25133 2601 25145 2604
rect 25179 2632 25191 2635
rect 25866 2632 25872 2644
rect 25179 2604 25872 2632
rect 25179 2601 25191 2604
rect 25133 2595 25191 2601
rect 25866 2592 25872 2604
rect 25924 2592 25930 2644
rect 24489 2567 24547 2573
rect 24489 2564 24501 2567
rect 24044 2536 24501 2564
rect 24489 2533 24501 2536
rect 24535 2564 24547 2567
rect 25038 2564 25044 2576
rect 24535 2536 25044 2564
rect 24535 2533 24547 2536
rect 24489 2527 24547 2533
rect 25038 2524 25044 2536
rect 25096 2524 25102 2576
rect 22879 2468 23520 2496
rect 22879 2465 22891 2468
rect 22833 2459 22891 2465
rect 23566 2456 23572 2508
rect 23624 2496 23630 2508
rect 23624 2468 24624 2496
rect 23624 2456 23630 2468
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2428 8079 2431
rect 8570 2428 8576 2440
rect 8067 2400 8576 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 8754 2428 8760 2440
rect 8715 2400 8760 2428
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 11514 2388 11520 2440
rect 11572 2428 11578 2440
rect 11609 2431 11667 2437
rect 11609 2428 11621 2431
rect 11572 2400 11621 2428
rect 11572 2388 11578 2400
rect 11609 2397 11621 2400
rect 11655 2428 11667 2431
rect 18046 2428 18052 2440
rect 11655 2400 12112 2428
rect 18007 2400 18052 2428
rect 11655 2397 11667 2400
rect 11609 2391 11667 2397
rect 6733 2363 6791 2369
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 8772 2360 8800 2388
rect 6779 2332 8800 2360
rect 9217 2363 9275 2369
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 9217 2329 9229 2363
rect 9263 2360 9275 2363
rect 11532 2360 11560 2388
rect 9263 2332 11560 2360
rect 9263 2329 9275 2332
rect 9217 2323 9275 2329
rect 10042 2292 10048 2304
rect 10003 2264 10048 2292
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 10778 2292 10784 2304
rect 10739 2264 10784 2292
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 12084 2292 12112 2400
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 18138 2388 18144 2440
rect 18196 2428 18202 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 18196 2400 18337 2428
rect 18196 2388 18202 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 21818 2428 21824 2440
rect 21731 2400 21824 2428
rect 18325 2391 18383 2397
rect 21818 2388 21824 2400
rect 21876 2428 21882 2440
rect 22278 2428 22284 2440
rect 21876 2400 22284 2428
rect 21876 2388 21882 2400
rect 22278 2388 22284 2400
rect 22336 2388 22342 2440
rect 24596 2437 24624 2468
rect 24854 2456 24860 2508
rect 24912 2496 24918 2508
rect 25593 2499 25651 2505
rect 25593 2496 25605 2499
rect 24912 2468 25605 2496
rect 24912 2456 24918 2468
rect 25593 2465 25605 2468
rect 25639 2465 25651 2499
rect 25593 2459 25651 2465
rect 24581 2431 24639 2437
rect 24581 2397 24593 2431
rect 24627 2428 24639 2431
rect 25409 2431 25467 2437
rect 25409 2428 25421 2431
rect 24627 2400 25421 2428
rect 24627 2397 24639 2400
rect 24581 2391 24639 2397
rect 25409 2397 25421 2400
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 23750 2320 23756 2372
rect 23808 2360 23814 2372
rect 24029 2363 24087 2369
rect 24029 2360 24041 2363
rect 23808 2332 24041 2360
rect 23808 2320 23814 2332
rect 24029 2329 24041 2332
rect 24075 2329 24087 2363
rect 24029 2323 24087 2329
rect 14001 2295 14059 2301
rect 14001 2292 14013 2295
rect 12084 2264 14013 2292
rect 14001 2261 14013 2264
rect 14047 2261 14059 2295
rect 14001 2255 14059 2261
rect 22646 2252 22652 2304
rect 22704 2292 22710 2304
rect 23017 2295 23075 2301
rect 23017 2292 23029 2295
rect 22704 2264 23029 2292
rect 22704 2252 22710 2264
rect 23017 2261 23029 2264
rect 23063 2261 23075 2295
rect 23017 2255 23075 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 23658 1368 23664 1420
rect 23716 1408 23722 1420
rect 24026 1408 24032 1420
rect 23716 1380 24032 1408
rect 23716 1368 23722 1380
rect 24026 1368 24032 1380
rect 24084 1368 24090 1420
rect 22830 1232 22836 1284
rect 22888 1272 22894 1284
rect 24302 1272 24308 1284
rect 22888 1244 24308 1272
rect 22888 1232 22894 1244
rect 24302 1232 24308 1244
rect 24360 1232 24366 1284
rect 15838 552 15844 604
rect 15896 592 15902 604
rect 16114 592 16120 604
rect 15896 564 16120 592
rect 15896 552 15902 564
rect 16114 552 16120 564
rect 16172 552 16178 604
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 12992 24828 13044 24880
rect 24768 24828 24820 24880
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 24216 24352 24268 24404
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 10140 23808 10192 23860
rect 12992 23851 13044 23860
rect 12992 23817 13001 23851
rect 13001 23817 13035 23851
rect 13035 23817 13044 23851
rect 12992 23808 13044 23817
rect 17500 23808 17552 23860
rect 12348 23604 12400 23656
rect 24676 23808 24728 23860
rect 18144 23604 18196 23656
rect 23940 23604 23992 23656
rect 3516 23468 3568 23520
rect 4068 23468 4120 23520
rect 10692 23511 10744 23520
rect 10692 23477 10701 23511
rect 10701 23477 10735 23511
rect 10735 23477 10744 23511
rect 10692 23468 10744 23477
rect 19432 23511 19484 23520
rect 19432 23477 19441 23511
rect 19441 23477 19475 23511
rect 19475 23477 19484 23511
rect 19432 23468 19484 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 24860 23264 24912 23316
rect 12348 23196 12400 23248
rect 23940 23239 23992 23248
rect 23940 23205 23949 23239
rect 23949 23205 23983 23239
rect 23983 23205 23992 23239
rect 23940 23196 23992 23205
rect 11796 23171 11848 23180
rect 11796 23137 11805 23171
rect 11805 23137 11839 23171
rect 11839 23137 11848 23171
rect 11796 23128 11848 23137
rect 23848 23128 23900 23180
rect 24952 23171 25004 23180
rect 24952 23137 24961 23171
rect 24961 23137 24995 23171
rect 24995 23137 25004 23171
rect 24952 23128 25004 23137
rect 18236 22924 18288 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 24216 22720 24268 22772
rect 24032 22584 24084 22636
rect 24216 22584 24268 22636
rect 24584 22559 24636 22568
rect 24584 22525 24593 22559
rect 24593 22525 24627 22559
rect 24627 22525 24636 22559
rect 24584 22516 24636 22525
rect 24952 22448 25004 22500
rect 11796 22423 11848 22432
rect 11796 22389 11805 22423
rect 11805 22389 11839 22423
rect 11839 22389 11848 22423
rect 11796 22380 11848 22389
rect 23848 22423 23900 22432
rect 23848 22389 23857 22423
rect 23857 22389 23891 22423
rect 23891 22389 23900 22423
rect 23848 22380 23900 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 10048 22083 10100 22092
rect 10048 22049 10057 22083
rect 10057 22049 10091 22083
rect 10091 22049 10100 22083
rect 10048 22040 10100 22049
rect 17040 22083 17092 22092
rect 17040 22049 17049 22083
rect 17049 22049 17083 22083
rect 17083 22049 17092 22083
rect 17040 22040 17092 22049
rect 10324 22015 10376 22024
rect 10324 21981 10333 22015
rect 10333 21981 10367 22015
rect 10367 21981 10376 22015
rect 10324 21972 10376 21981
rect 17224 21947 17276 21956
rect 17224 21913 17233 21947
rect 17233 21913 17267 21947
rect 17267 21913 17276 21947
rect 17224 21904 17276 21913
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 17040 21675 17092 21684
rect 17040 21641 17049 21675
rect 17049 21641 17083 21675
rect 17083 21641 17092 21675
rect 17040 21632 17092 21641
rect 24676 21632 24728 21684
rect 13728 21539 13780 21548
rect 13728 21505 13737 21539
rect 13737 21505 13771 21539
rect 13771 21505 13780 21539
rect 13728 21496 13780 21505
rect 12992 21428 13044 21480
rect 23940 21428 23992 21480
rect 9680 21292 9732 21344
rect 10048 21335 10100 21344
rect 10048 21301 10057 21335
rect 10057 21301 10091 21335
rect 10091 21301 10100 21335
rect 10048 21292 10100 21301
rect 16212 21292 16264 21344
rect 17040 21292 17092 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 24768 21131 24820 21140
rect 24768 21097 24777 21131
rect 24777 21097 24811 21131
rect 24811 21097 24820 21131
rect 24768 21088 24820 21097
rect 16212 21063 16264 21072
rect 16212 21029 16221 21063
rect 16221 21029 16255 21063
rect 16255 21029 16264 21063
rect 16212 21020 16264 21029
rect 15844 20952 15896 21004
rect 24676 20952 24728 21004
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 25136 20587 25188 20596
rect 25136 20553 25145 20587
rect 25145 20553 25179 20587
rect 25179 20553 25188 20587
rect 25136 20544 25188 20553
rect 23940 20451 23992 20460
rect 23940 20417 23949 20451
rect 23949 20417 23983 20451
rect 23983 20417 23992 20451
rect 23940 20408 23992 20417
rect 24860 20340 24912 20392
rect 15844 20204 15896 20256
rect 23480 20247 23532 20256
rect 23480 20213 23489 20247
rect 23489 20213 23523 20247
rect 23523 20213 23532 20247
rect 23480 20204 23532 20213
rect 24584 20247 24636 20256
rect 24584 20213 24593 20247
rect 24593 20213 24627 20247
rect 24627 20213 24636 20247
rect 24584 20204 24636 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 24032 20000 24084 20052
rect 21456 19975 21508 19984
rect 21456 19941 21465 19975
rect 21465 19941 21499 19975
rect 21499 19941 21508 19975
rect 21456 19932 21508 19941
rect 20904 19864 20956 19916
rect 24032 19864 24084 19916
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 24860 19320 24912 19372
rect 24952 19295 25004 19304
rect 24952 19261 24961 19295
rect 24961 19261 24995 19295
rect 24995 19261 25004 19295
rect 24952 19252 25004 19261
rect 20904 19116 20956 19168
rect 23480 19159 23532 19168
rect 23480 19125 23489 19159
rect 23489 19125 23523 19159
rect 23523 19125 23532 19159
rect 23480 19116 23532 19125
rect 24584 19159 24636 19168
rect 24584 19125 24593 19159
rect 24593 19125 24627 19159
rect 24627 19125 24636 19159
rect 24584 19116 24636 19125
rect 24860 19116 24912 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 11060 18776 11112 18828
rect 16028 18819 16080 18828
rect 16028 18785 16037 18819
rect 16037 18785 16071 18819
rect 16071 18785 16080 18819
rect 16028 18776 16080 18785
rect 16304 18819 16356 18828
rect 16304 18785 16313 18819
rect 16313 18785 16347 18819
rect 16347 18785 16356 18819
rect 16304 18776 16356 18785
rect 11336 18683 11388 18692
rect 11336 18649 11345 18683
rect 11345 18649 11379 18683
rect 11379 18649 11388 18683
rect 11336 18640 11388 18649
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 13268 18164 13320 18216
rect 13452 18139 13504 18148
rect 13452 18105 13461 18139
rect 13461 18105 13495 18139
rect 13495 18105 13504 18139
rect 13452 18096 13504 18105
rect 11060 18028 11112 18080
rect 15292 18028 15344 18080
rect 16028 18071 16080 18080
rect 16028 18037 16037 18071
rect 16037 18037 16071 18071
rect 16071 18037 16080 18071
rect 16028 18028 16080 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 24676 17824 24728 17876
rect 10968 17756 11020 17808
rect 10140 17688 10192 17740
rect 25136 17688 25188 17740
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 24768 17323 24820 17332
rect 24768 17289 24777 17323
rect 24777 17289 24811 17323
rect 24811 17289 24820 17323
rect 24768 17280 24820 17289
rect 16028 17255 16080 17264
rect 16028 17221 16037 17255
rect 16037 17221 16071 17255
rect 16071 17221 16080 17255
rect 16028 17212 16080 17221
rect 12348 17076 12400 17128
rect 15568 17076 15620 17128
rect 12716 17051 12768 17060
rect 12716 17017 12725 17051
rect 12725 17017 12759 17051
rect 12759 17017 12768 17051
rect 12716 17008 12768 17017
rect 25136 17119 25188 17128
rect 25136 17085 25145 17119
rect 25145 17085 25179 17119
rect 25179 17085 25188 17119
rect 25136 17076 25188 17085
rect 10140 16940 10192 16992
rect 24400 16983 24452 16992
rect 24400 16949 24409 16983
rect 24409 16949 24443 16983
rect 24443 16949 24452 16983
rect 24400 16940 24452 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 24032 16736 24084 16788
rect 15568 16711 15620 16720
rect 15568 16677 15577 16711
rect 15577 16677 15611 16711
rect 15611 16677 15620 16711
rect 15568 16668 15620 16677
rect 15384 16600 15436 16652
rect 24676 16600 24728 16652
rect 24216 16396 24268 16448
rect 24952 16396 25004 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 24768 16235 24820 16244
rect 24768 16201 24777 16235
rect 24777 16201 24811 16235
rect 24811 16201 24820 16235
rect 24768 16192 24820 16201
rect 24676 16124 24728 16176
rect 18328 16099 18380 16108
rect 18328 16065 18337 16099
rect 18337 16065 18371 16099
rect 18371 16065 18380 16099
rect 18328 16056 18380 16065
rect 24216 15988 24268 16040
rect 15200 15852 15252 15904
rect 15384 15852 15436 15904
rect 18696 15852 18748 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 25044 15691 25096 15700
rect 25044 15657 25053 15691
rect 25053 15657 25087 15691
rect 25087 15657 25096 15691
rect 25044 15648 25096 15657
rect 24676 15580 24728 15632
rect 23480 15512 23532 15564
rect 24860 15555 24912 15564
rect 24860 15521 24869 15555
rect 24869 15521 24903 15555
rect 24903 15521 24912 15555
rect 24860 15512 24912 15521
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 25504 15147 25556 15156
rect 25504 15113 25513 15147
rect 25513 15113 25547 15147
rect 25547 15113 25556 15147
rect 25504 15104 25556 15113
rect 24216 15011 24268 15020
rect 24216 14977 24225 15011
rect 24225 14977 24259 15011
rect 24259 14977 24268 15011
rect 24216 14968 24268 14977
rect 23480 14943 23532 14952
rect 23480 14909 23489 14943
rect 23489 14909 23523 14943
rect 23523 14909 23532 14943
rect 23480 14900 23532 14909
rect 23664 14764 23716 14816
rect 25412 14900 25464 14952
rect 24860 14807 24912 14816
rect 24860 14773 24869 14807
rect 24869 14773 24903 14807
rect 24903 14773 24912 14807
rect 24860 14764 24912 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 23388 14535 23440 14544
rect 23388 14501 23397 14535
rect 23397 14501 23431 14535
rect 23431 14501 23440 14535
rect 23388 14492 23440 14501
rect 23112 14467 23164 14476
rect 23112 14433 23121 14467
rect 23121 14433 23155 14467
rect 23155 14433 23164 14467
rect 23112 14424 23164 14433
rect 24768 14424 24820 14476
rect 21272 14356 21324 14408
rect 24768 14263 24820 14272
rect 24768 14229 24777 14263
rect 24777 14229 24811 14263
rect 24811 14229 24820 14263
rect 24768 14220 24820 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 24124 14016 24176 14068
rect 24860 14016 24912 14068
rect 21824 13812 21876 13864
rect 23112 13855 23164 13864
rect 23112 13821 23121 13855
rect 23121 13821 23155 13855
rect 23155 13821 23164 13855
rect 23112 13812 23164 13821
rect 20444 13676 20496 13728
rect 21732 13676 21784 13728
rect 22284 13719 22336 13728
rect 22284 13685 22293 13719
rect 22293 13685 22327 13719
rect 22327 13685 22336 13719
rect 22284 13676 22336 13685
rect 24124 13676 24176 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 20904 13515 20956 13524
rect 20904 13481 20913 13515
rect 20913 13481 20947 13515
rect 20947 13481 20956 13515
rect 20904 13472 20956 13481
rect 21272 13515 21324 13524
rect 21272 13481 21281 13515
rect 21281 13481 21315 13515
rect 21315 13481 21324 13515
rect 21272 13472 21324 13481
rect 23388 13472 23440 13524
rect 23572 13472 23624 13524
rect 16304 13379 16356 13388
rect 16304 13345 16313 13379
rect 16313 13345 16347 13379
rect 16347 13345 16356 13379
rect 16304 13336 16356 13345
rect 21548 13336 21600 13388
rect 22928 13336 22980 13388
rect 24032 13336 24084 13388
rect 18144 13311 18196 13320
rect 18144 13277 18153 13311
rect 18153 13277 18187 13311
rect 18187 13277 18196 13311
rect 18144 13268 18196 13277
rect 18788 13268 18840 13320
rect 21640 13268 21692 13320
rect 23204 13311 23256 13320
rect 23204 13277 23213 13311
rect 23213 13277 23247 13311
rect 23247 13277 23256 13311
rect 23204 13268 23256 13277
rect 17776 13175 17828 13184
rect 17776 13141 17785 13175
rect 17785 13141 17819 13175
rect 17819 13141 17828 13175
rect 17776 13132 17828 13141
rect 20536 13132 20588 13184
rect 22652 13175 22704 13184
rect 22652 13141 22661 13175
rect 22661 13141 22695 13175
rect 22695 13141 22704 13175
rect 22652 13132 22704 13141
rect 23848 13175 23900 13184
rect 23848 13141 23857 13175
rect 23857 13141 23891 13175
rect 23891 13141 23900 13175
rect 23848 13132 23900 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 16304 12971 16356 12980
rect 16304 12937 16313 12971
rect 16313 12937 16347 12971
rect 16347 12937 16356 12971
rect 16304 12928 16356 12937
rect 21272 12928 21324 12980
rect 23204 12928 23256 12980
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 24032 12928 24084 12980
rect 25780 12971 25832 12980
rect 25780 12937 25789 12971
rect 25789 12937 25823 12971
rect 25823 12937 25832 12971
rect 25780 12928 25832 12937
rect 18420 12903 18472 12912
rect 18420 12869 18429 12903
rect 18429 12869 18463 12903
rect 18463 12869 18472 12903
rect 18420 12860 18472 12869
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 19524 12792 19576 12844
rect 20536 12835 20588 12844
rect 18788 12767 18840 12776
rect 18788 12733 18797 12767
rect 18797 12733 18831 12767
rect 18831 12733 18840 12767
rect 18788 12724 18840 12733
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 24124 12835 24176 12844
rect 24124 12801 24133 12835
rect 24133 12801 24167 12835
rect 24167 12801 24176 12835
rect 24124 12792 24176 12801
rect 23848 12767 23900 12776
rect 23848 12733 23857 12767
rect 23857 12733 23891 12767
rect 23891 12733 23900 12767
rect 23848 12724 23900 12733
rect 25780 12724 25832 12776
rect 19340 12656 19392 12708
rect 21640 12656 21692 12708
rect 18604 12588 18656 12640
rect 19984 12631 20036 12640
rect 19984 12597 19993 12631
rect 19993 12597 20027 12631
rect 20027 12597 20036 12631
rect 19984 12588 20036 12597
rect 21272 12588 21324 12640
rect 21548 12588 21600 12640
rect 22744 12588 22796 12640
rect 22928 12631 22980 12640
rect 22928 12597 22937 12631
rect 22937 12597 22971 12631
rect 22971 12597 22980 12631
rect 22928 12588 22980 12597
rect 25320 12631 25372 12640
rect 25320 12597 25329 12631
rect 25329 12597 25363 12631
rect 25363 12597 25372 12631
rect 25320 12588 25372 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 18972 12384 19024 12436
rect 19248 12427 19300 12436
rect 19248 12393 19257 12427
rect 19257 12393 19291 12427
rect 19291 12393 19300 12427
rect 19248 12384 19300 12393
rect 20720 12384 20772 12436
rect 21916 12384 21968 12436
rect 23756 12384 23808 12436
rect 24308 12384 24360 12436
rect 17408 12359 17460 12368
rect 17408 12325 17417 12359
rect 17417 12325 17451 12359
rect 17451 12325 17460 12359
rect 17408 12316 17460 12325
rect 17500 12248 17552 12300
rect 19340 12248 19392 12300
rect 17040 12180 17092 12232
rect 19708 12223 19760 12232
rect 19708 12189 19717 12223
rect 19717 12189 19751 12223
rect 19751 12189 19760 12223
rect 19708 12180 19760 12189
rect 24032 12291 24084 12300
rect 24032 12257 24041 12291
rect 24041 12257 24075 12291
rect 24075 12257 24084 12291
rect 24032 12248 24084 12257
rect 25688 12248 25740 12300
rect 20812 12112 20864 12164
rect 20260 12087 20312 12096
rect 20260 12053 20269 12087
rect 20269 12053 20303 12087
rect 20303 12053 20312 12087
rect 24216 12223 24268 12232
rect 24216 12189 24225 12223
rect 24225 12189 24259 12223
rect 24259 12189 24268 12223
rect 24216 12180 24268 12189
rect 20260 12044 20312 12053
rect 22468 12044 22520 12096
rect 22652 12044 22704 12096
rect 23204 12044 23256 12096
rect 23480 12087 23532 12096
rect 23480 12053 23489 12087
rect 23489 12053 23523 12087
rect 23523 12053 23532 12087
rect 23480 12044 23532 12053
rect 23572 12044 23624 12096
rect 24124 12044 24176 12096
rect 24860 12044 24912 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 19708 11840 19760 11892
rect 20812 11883 20864 11892
rect 20812 11849 20821 11883
rect 20821 11849 20855 11883
rect 20855 11849 20864 11883
rect 20812 11840 20864 11849
rect 22928 11840 22980 11892
rect 23940 11840 23992 11892
rect 25688 11883 25740 11892
rect 25688 11849 25697 11883
rect 25697 11849 25731 11883
rect 25731 11849 25740 11883
rect 25688 11840 25740 11849
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 22468 11747 22520 11756
rect 22468 11713 22477 11747
rect 22477 11713 22511 11747
rect 22511 11713 22520 11747
rect 22468 11704 22520 11713
rect 23112 11704 23164 11756
rect 16764 11568 16816 11620
rect 18236 11636 18288 11688
rect 20260 11636 20312 11688
rect 22284 11636 22336 11688
rect 17408 11568 17460 11620
rect 18972 11568 19024 11620
rect 19524 11568 19576 11620
rect 22744 11568 22796 11620
rect 23480 11568 23532 11620
rect 24032 11568 24084 11620
rect 17500 11543 17552 11552
rect 17500 11509 17509 11543
rect 17509 11509 17543 11543
rect 17543 11509 17552 11543
rect 17500 11500 17552 11509
rect 19340 11543 19392 11552
rect 19340 11509 19349 11543
rect 19349 11509 19383 11543
rect 19383 11509 19392 11543
rect 19340 11500 19392 11509
rect 20720 11500 20772 11552
rect 23112 11543 23164 11552
rect 23112 11509 23121 11543
rect 23121 11509 23155 11543
rect 23155 11509 23164 11543
rect 23112 11500 23164 11509
rect 25044 11543 25096 11552
rect 25044 11509 25053 11543
rect 25053 11509 25087 11543
rect 25087 11509 25096 11543
rect 25044 11500 25096 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 17500 11296 17552 11348
rect 19524 11296 19576 11348
rect 22744 11339 22796 11348
rect 22744 11305 22753 11339
rect 22753 11305 22787 11339
rect 22787 11305 22796 11339
rect 22744 11296 22796 11305
rect 23756 11339 23808 11348
rect 23756 11305 23765 11339
rect 23765 11305 23799 11339
rect 23799 11305 23808 11339
rect 23756 11296 23808 11305
rect 23848 11296 23900 11348
rect 24032 11296 24084 11348
rect 17040 11271 17092 11280
rect 17040 11237 17049 11271
rect 17049 11237 17083 11271
rect 17083 11237 17092 11271
rect 17040 11228 17092 11237
rect 22008 11228 22060 11280
rect 23112 11228 23164 11280
rect 23480 11228 23532 11280
rect 25044 11228 25096 11280
rect 13912 11203 13964 11212
rect 13912 11169 13921 11203
rect 13921 11169 13955 11203
rect 13955 11169 13964 11203
rect 13912 11160 13964 11169
rect 15384 11160 15436 11212
rect 18236 11160 18288 11212
rect 18420 11160 18472 11212
rect 20260 11160 20312 11212
rect 14280 11092 14332 11144
rect 15476 11135 15528 11144
rect 15476 11101 15485 11135
rect 15485 11101 15519 11135
rect 15519 11101 15528 11135
rect 15476 11092 15528 11101
rect 17316 11135 17368 11144
rect 16580 11067 16632 11076
rect 16580 11033 16589 11067
rect 16589 11033 16623 11067
rect 16623 11033 16632 11067
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 21456 11160 21508 11212
rect 21916 11160 21968 11212
rect 23756 11092 23808 11144
rect 16580 11024 16632 11033
rect 18144 10999 18196 11008
rect 18144 10965 18153 10999
rect 18153 10965 18187 10999
rect 18187 10965 18196 10999
rect 18144 10956 18196 10965
rect 23848 10956 23900 11008
rect 24216 10956 24268 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 13912 10752 13964 10804
rect 17040 10752 17092 10804
rect 17316 10752 17368 10804
rect 20260 10752 20312 10804
rect 14188 10548 14240 10600
rect 14740 10591 14792 10600
rect 14740 10557 14749 10591
rect 14749 10557 14783 10591
rect 14783 10557 14792 10591
rect 14740 10548 14792 10557
rect 21548 10752 21600 10804
rect 21824 10752 21876 10804
rect 23480 10795 23532 10804
rect 23480 10761 23489 10795
rect 23489 10761 23523 10795
rect 23523 10761 23532 10795
rect 23480 10752 23532 10761
rect 21916 10616 21968 10668
rect 22468 10659 22520 10668
rect 22468 10625 22477 10659
rect 22477 10625 22511 10659
rect 22511 10625 22520 10659
rect 22468 10616 22520 10625
rect 22100 10548 22152 10600
rect 23756 10548 23808 10600
rect 18144 10480 18196 10532
rect 23848 10480 23900 10532
rect 13728 10455 13780 10464
rect 13728 10421 13737 10455
rect 13737 10421 13771 10455
rect 13771 10421 13780 10455
rect 13728 10412 13780 10421
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 18420 10412 18472 10464
rect 20996 10455 21048 10464
rect 20996 10421 21005 10455
rect 21005 10421 21039 10455
rect 21039 10421 21048 10455
rect 20996 10412 21048 10421
rect 22100 10412 22152 10464
rect 24032 10412 24084 10464
rect 25320 10412 25372 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 13636 10251 13688 10260
rect 13636 10217 13645 10251
rect 13645 10217 13679 10251
rect 13679 10217 13688 10251
rect 13636 10208 13688 10217
rect 15384 10208 15436 10260
rect 17316 10208 17368 10260
rect 18420 10251 18472 10260
rect 18420 10217 18429 10251
rect 18429 10217 18463 10251
rect 18463 10217 18472 10251
rect 18420 10208 18472 10217
rect 18604 10251 18656 10260
rect 18604 10217 18613 10251
rect 18613 10217 18647 10251
rect 18647 10217 18656 10251
rect 18604 10208 18656 10217
rect 20260 10251 20312 10260
rect 20260 10217 20269 10251
rect 20269 10217 20303 10251
rect 20303 10217 20312 10251
rect 20260 10208 20312 10217
rect 16120 10140 16172 10192
rect 21180 10208 21232 10260
rect 22468 10208 22520 10260
rect 22928 10251 22980 10260
rect 22928 10217 22937 10251
rect 22937 10217 22971 10251
rect 22971 10217 22980 10251
rect 22928 10208 22980 10217
rect 23388 10251 23440 10260
rect 23388 10217 23397 10251
rect 23397 10217 23431 10251
rect 23431 10217 23440 10251
rect 23388 10208 23440 10217
rect 24032 10251 24084 10260
rect 24032 10217 24041 10251
rect 24041 10217 24075 10251
rect 24075 10217 24084 10251
rect 24032 10208 24084 10217
rect 24492 10251 24544 10260
rect 24492 10217 24501 10251
rect 24501 10217 24535 10251
rect 24535 10217 24544 10251
rect 24492 10208 24544 10217
rect 13360 10072 13412 10124
rect 13728 10072 13780 10124
rect 14096 10115 14148 10124
rect 14096 10081 14105 10115
rect 14105 10081 14139 10115
rect 14139 10081 14148 10115
rect 14096 10072 14148 10081
rect 18328 10072 18380 10124
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 12808 9868 12860 9920
rect 13544 9911 13596 9920
rect 13544 9877 13553 9911
rect 13553 9877 13587 9911
rect 13587 9877 13596 9911
rect 13544 9868 13596 9877
rect 14740 9868 14792 9920
rect 15384 9868 15436 9920
rect 17960 10004 18012 10056
rect 19064 10047 19116 10056
rect 19064 10013 19073 10047
rect 19073 10013 19107 10047
rect 19107 10013 19116 10047
rect 19064 10004 19116 10013
rect 21364 10140 21416 10192
rect 21732 10140 21784 10192
rect 23020 10140 23072 10192
rect 24860 10115 24912 10124
rect 24860 10081 24869 10115
rect 24869 10081 24903 10115
rect 24903 10081 24912 10115
rect 24860 10072 24912 10081
rect 25780 10072 25832 10124
rect 21548 10047 21600 10056
rect 21548 10013 21557 10047
rect 21557 10013 21591 10047
rect 21591 10013 21600 10047
rect 21548 10004 21600 10013
rect 23480 10004 23532 10056
rect 24032 10004 24084 10056
rect 22100 9936 22152 9988
rect 24308 9979 24360 9988
rect 24308 9945 24317 9979
rect 24317 9945 24351 9979
rect 24351 9945 24360 9979
rect 24308 9936 24360 9945
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 20720 9911 20772 9920
rect 20720 9877 20729 9911
rect 20729 9877 20763 9911
rect 20763 9877 20772 9911
rect 20720 9868 20772 9877
rect 21916 9911 21968 9920
rect 21916 9877 21925 9911
rect 21925 9877 21959 9911
rect 21959 9877 21968 9911
rect 21916 9868 21968 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 13360 9707 13412 9716
rect 13360 9673 13369 9707
rect 13369 9673 13403 9707
rect 13403 9673 13412 9707
rect 13360 9664 13412 9673
rect 20260 9664 20312 9716
rect 17960 9596 18012 9648
rect 19892 9639 19944 9648
rect 19892 9605 19901 9639
rect 19901 9605 19935 9639
rect 19935 9605 19944 9639
rect 19892 9596 19944 9605
rect 21180 9664 21232 9716
rect 23020 9707 23072 9716
rect 23020 9673 23029 9707
rect 23029 9673 23063 9707
rect 23063 9673 23072 9707
rect 23020 9664 23072 9673
rect 23480 9664 23532 9716
rect 24860 9664 24912 9716
rect 25780 9664 25832 9716
rect 20996 9596 21048 9648
rect 16120 9528 16172 9580
rect 16672 9571 16724 9580
rect 16672 9537 16681 9571
rect 16681 9537 16715 9571
rect 16715 9537 16724 9571
rect 16672 9528 16724 9537
rect 12808 9460 12860 9512
rect 13544 9460 13596 9512
rect 14740 9460 14792 9512
rect 18144 9460 18196 9512
rect 19524 9460 19576 9512
rect 21456 9460 21508 9512
rect 21732 9460 21784 9512
rect 23480 9460 23532 9512
rect 14188 9392 14240 9444
rect 13084 9324 13136 9376
rect 18788 9435 18840 9444
rect 18788 9401 18822 9435
rect 18822 9401 18840 9435
rect 18788 9392 18840 9401
rect 16028 9324 16080 9376
rect 16396 9324 16448 9376
rect 18328 9367 18380 9376
rect 18328 9333 18337 9367
rect 18337 9333 18371 9367
rect 18371 9333 18380 9367
rect 18328 9324 18380 9333
rect 20904 9324 20956 9376
rect 21272 9324 21324 9376
rect 21916 9324 21968 9376
rect 25044 9367 25096 9376
rect 25044 9333 25053 9367
rect 25053 9333 25087 9367
rect 25087 9333 25096 9367
rect 25044 9324 25096 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 10692 9120 10744 9172
rect 13544 9120 13596 9172
rect 14004 9163 14056 9172
rect 14004 9129 14013 9163
rect 14013 9129 14047 9163
rect 14047 9129 14056 9163
rect 14004 9120 14056 9129
rect 14096 9120 14148 9172
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 16672 9163 16724 9172
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 18788 9120 18840 9172
rect 21548 9120 21600 9172
rect 23388 9120 23440 9172
rect 24860 9163 24912 9172
rect 24860 9129 24869 9163
rect 24869 9129 24903 9163
rect 24903 9129 24912 9163
rect 24860 9120 24912 9129
rect 21272 9052 21324 9104
rect 21824 9052 21876 9104
rect 10692 8984 10744 9036
rect 12164 8984 12216 9036
rect 14832 8984 14884 9036
rect 16856 8984 16908 9036
rect 20996 8984 21048 9036
rect 25044 8984 25096 9036
rect 10784 8916 10836 8968
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 15752 8959 15804 8968
rect 11520 8823 11572 8832
rect 11520 8789 11529 8823
rect 11529 8789 11563 8823
rect 11563 8789 11572 8823
rect 11520 8780 11572 8789
rect 15752 8925 15761 8959
rect 15761 8925 15795 8959
rect 15795 8925 15804 8959
rect 15752 8916 15804 8925
rect 12808 8780 12860 8832
rect 20628 8916 20680 8968
rect 23480 8959 23532 8968
rect 23480 8925 23489 8959
rect 23489 8925 23523 8959
rect 23523 8925 23532 8959
rect 23480 8916 23532 8925
rect 19524 8848 19576 8900
rect 16488 8780 16540 8832
rect 17040 8823 17092 8832
rect 17040 8789 17049 8823
rect 17049 8789 17083 8823
rect 17083 8789 17092 8823
rect 17040 8780 17092 8789
rect 19800 8780 19852 8832
rect 22284 8823 22336 8832
rect 22284 8789 22293 8823
rect 22293 8789 22327 8823
rect 22327 8789 22336 8823
rect 22284 8780 22336 8789
rect 24860 8780 24912 8832
rect 25320 8780 25372 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 10784 8619 10836 8628
rect 10784 8585 10793 8619
rect 10793 8585 10827 8619
rect 10827 8585 10836 8619
rect 10784 8576 10836 8585
rect 13176 8576 13228 8628
rect 11060 8508 11112 8560
rect 12164 8508 12216 8560
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 11520 8440 11572 8492
rect 12532 8372 12584 8424
rect 14096 8576 14148 8628
rect 16856 8619 16908 8628
rect 16856 8585 16865 8619
rect 16865 8585 16899 8619
rect 16899 8585 16908 8619
rect 16856 8576 16908 8585
rect 19156 8619 19208 8628
rect 19156 8585 19165 8619
rect 19165 8585 19199 8619
rect 19199 8585 19208 8619
rect 19156 8576 19208 8585
rect 19800 8576 19852 8628
rect 21272 8619 21324 8628
rect 13360 8508 13412 8560
rect 14832 8551 14884 8560
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 14832 8517 14841 8551
rect 14841 8517 14875 8551
rect 14875 8517 14884 8551
rect 14832 8508 14884 8517
rect 17868 8508 17920 8560
rect 15108 8372 15160 8424
rect 12440 8347 12492 8356
rect 12440 8313 12449 8347
rect 12449 8313 12483 8347
rect 12483 8313 12492 8347
rect 12440 8304 12492 8313
rect 13360 8304 13412 8356
rect 13452 8304 13504 8356
rect 15292 8372 15344 8424
rect 18512 8440 18564 8492
rect 21272 8585 21281 8619
rect 21281 8585 21315 8619
rect 21315 8585 21324 8619
rect 21272 8576 21324 8585
rect 21456 8508 21508 8560
rect 22652 8551 22704 8560
rect 22652 8517 22661 8551
rect 22661 8517 22695 8551
rect 22695 8517 22704 8551
rect 22652 8508 22704 8517
rect 16488 8372 16540 8424
rect 19800 8415 19852 8424
rect 16396 8304 16448 8356
rect 15108 8236 15160 8288
rect 18420 8279 18472 8288
rect 18420 8245 18429 8279
rect 18429 8245 18463 8279
rect 18463 8245 18472 8279
rect 18420 8236 18472 8245
rect 19800 8381 19809 8415
rect 19809 8381 19843 8415
rect 19843 8381 19852 8415
rect 19800 8372 19852 8381
rect 23204 8576 23256 8628
rect 23480 8508 23532 8560
rect 24124 8440 24176 8492
rect 25044 8576 25096 8628
rect 25412 8483 25464 8492
rect 25412 8449 25421 8483
rect 25421 8449 25455 8483
rect 25455 8449 25464 8483
rect 25412 8440 25464 8449
rect 23940 8372 23992 8424
rect 25228 8415 25280 8424
rect 25228 8381 25237 8415
rect 25237 8381 25271 8415
rect 25271 8381 25280 8415
rect 25228 8372 25280 8381
rect 18604 8236 18656 8288
rect 19524 8236 19576 8288
rect 19984 8304 20036 8356
rect 24216 8236 24268 8288
rect 24860 8236 24912 8288
rect 25688 8236 25740 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 10784 8032 10836 8084
rect 12164 8075 12216 8084
rect 12164 8041 12173 8075
rect 12173 8041 12207 8075
rect 12207 8041 12216 8075
rect 12164 8032 12216 8041
rect 13268 8075 13320 8084
rect 13268 8041 13277 8075
rect 13277 8041 13311 8075
rect 13311 8041 13320 8075
rect 13268 8032 13320 8041
rect 16580 8032 16632 8084
rect 16856 8032 16908 8084
rect 19248 8032 19300 8084
rect 19432 8032 19484 8084
rect 22008 8032 22060 8084
rect 22560 8032 22612 8084
rect 23020 8075 23072 8084
rect 23020 8041 23029 8075
rect 23029 8041 23063 8075
rect 23063 8041 23072 8075
rect 23020 8032 23072 8041
rect 23388 8032 23440 8084
rect 24124 8075 24176 8084
rect 24124 8041 24133 8075
rect 24133 8041 24167 8075
rect 24167 8041 24176 8075
rect 24124 8032 24176 8041
rect 10692 7964 10744 8016
rect 11520 7964 11572 8016
rect 13084 7964 13136 8016
rect 18604 7964 18656 8016
rect 21640 7964 21692 8016
rect 24216 7964 24268 8016
rect 24768 7964 24820 8016
rect 15108 7939 15160 7948
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 12808 7803 12860 7812
rect 12808 7769 12817 7803
rect 12817 7769 12851 7803
rect 12851 7769 12860 7803
rect 12808 7760 12860 7769
rect 13452 7760 13504 7812
rect 13544 7760 13596 7812
rect 13176 7735 13228 7744
rect 13176 7701 13185 7735
rect 13185 7701 13219 7735
rect 13219 7701 13228 7735
rect 13176 7692 13228 7701
rect 14648 7692 14700 7744
rect 15108 7905 15117 7939
rect 15117 7905 15151 7939
rect 15151 7905 15160 7939
rect 15108 7896 15160 7905
rect 16396 7896 16448 7948
rect 18420 7939 18472 7948
rect 18420 7905 18429 7939
rect 18429 7905 18463 7939
rect 18463 7905 18472 7939
rect 18420 7896 18472 7905
rect 15292 7871 15344 7880
rect 14832 7692 14884 7744
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 17684 7828 17736 7880
rect 20352 7828 20404 7880
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 19616 7760 19668 7812
rect 20904 7760 20956 7812
rect 23480 7896 23532 7948
rect 22376 7828 22428 7880
rect 24216 7828 24268 7880
rect 23296 7760 23348 7812
rect 17040 7692 17092 7744
rect 17960 7692 18012 7744
rect 19432 7735 19484 7744
rect 19432 7701 19441 7735
rect 19441 7701 19475 7735
rect 19475 7701 19484 7735
rect 19432 7692 19484 7701
rect 20168 7692 20220 7744
rect 20720 7735 20772 7744
rect 20720 7701 20729 7735
rect 20729 7701 20763 7735
rect 20763 7701 20772 7735
rect 20720 7692 20772 7701
rect 22100 7735 22152 7744
rect 22100 7701 22109 7735
rect 22109 7701 22143 7735
rect 22143 7701 22152 7735
rect 22652 7735 22704 7744
rect 22100 7692 22152 7701
rect 22652 7701 22661 7735
rect 22661 7701 22695 7735
rect 22695 7701 22704 7735
rect 22652 7692 22704 7701
rect 24124 7692 24176 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 10968 7488 11020 7540
rect 11520 7488 11572 7540
rect 13084 7531 13136 7540
rect 13084 7497 13093 7531
rect 13093 7497 13127 7531
rect 13127 7497 13136 7531
rect 13084 7488 13136 7497
rect 13176 7488 13228 7540
rect 14832 7488 14884 7540
rect 15752 7531 15804 7540
rect 15752 7497 15761 7531
rect 15761 7497 15795 7531
rect 15795 7497 15804 7531
rect 15752 7488 15804 7497
rect 21364 7531 21416 7540
rect 21364 7497 21373 7531
rect 21373 7497 21407 7531
rect 21407 7497 21416 7531
rect 21364 7488 21416 7497
rect 22376 7488 22428 7540
rect 23020 7531 23072 7540
rect 23020 7497 23029 7531
rect 23029 7497 23063 7531
rect 23063 7497 23072 7531
rect 23020 7488 23072 7497
rect 23664 7531 23716 7540
rect 23664 7497 23673 7531
rect 23673 7497 23707 7531
rect 23707 7497 23716 7531
rect 23664 7488 23716 7497
rect 23848 7488 23900 7540
rect 24216 7488 24268 7540
rect 26240 7488 26292 7540
rect 26884 7488 26936 7540
rect 21456 7420 21508 7472
rect 21732 7420 21784 7472
rect 16396 7395 16448 7404
rect 16396 7361 16405 7395
rect 16405 7361 16439 7395
rect 16439 7361 16448 7395
rect 16396 7352 16448 7361
rect 21272 7395 21324 7404
rect 21272 7361 21281 7395
rect 21281 7361 21315 7395
rect 21315 7361 21324 7395
rect 21272 7352 21324 7361
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 9036 7148 9088 7200
rect 13544 7327 13596 7336
rect 10048 7216 10100 7268
rect 13544 7293 13578 7327
rect 13578 7293 13596 7327
rect 13544 7284 13596 7293
rect 15292 7327 15344 7336
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 14648 7191 14700 7200
rect 14648 7157 14657 7191
rect 14657 7157 14691 7191
rect 14691 7157 14700 7191
rect 14648 7148 14700 7157
rect 15568 7191 15620 7200
rect 15568 7157 15577 7191
rect 15577 7157 15611 7191
rect 15611 7157 15620 7191
rect 15568 7148 15620 7157
rect 18052 7284 18104 7336
rect 19432 7284 19484 7336
rect 20720 7284 20772 7336
rect 23664 7284 23716 7336
rect 25228 7327 25280 7336
rect 25228 7293 25237 7327
rect 25237 7293 25271 7327
rect 25271 7293 25280 7327
rect 25228 7284 25280 7293
rect 18420 7216 18472 7268
rect 16304 7148 16356 7200
rect 17592 7148 17644 7200
rect 17684 7148 17736 7200
rect 18604 7191 18656 7200
rect 18604 7157 18613 7191
rect 18613 7157 18647 7191
rect 18647 7157 18656 7191
rect 18604 7148 18656 7157
rect 19248 7216 19300 7268
rect 20536 7216 20588 7268
rect 22100 7216 22152 7268
rect 25504 7259 25556 7268
rect 25504 7225 25513 7259
rect 25513 7225 25547 7259
rect 25547 7225 25556 7259
rect 25504 7216 25556 7225
rect 19432 7148 19484 7200
rect 20260 7191 20312 7200
rect 20260 7157 20269 7191
rect 20269 7157 20303 7191
rect 20303 7157 20312 7191
rect 20260 7148 20312 7157
rect 24768 7148 24820 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 13544 6944 13596 6996
rect 14648 6944 14700 6996
rect 16396 6944 16448 6996
rect 19248 6944 19300 6996
rect 20168 6944 20220 6996
rect 22836 6944 22888 6996
rect 23388 6944 23440 6996
rect 23480 6987 23532 6996
rect 23480 6953 23489 6987
rect 23489 6953 23523 6987
rect 23523 6953 23532 6987
rect 23480 6944 23532 6953
rect 24216 6944 24268 6996
rect 14740 6876 14792 6928
rect 17592 6919 17644 6928
rect 17592 6885 17601 6919
rect 17601 6885 17635 6919
rect 17635 6885 17644 6919
rect 17592 6876 17644 6885
rect 9864 6808 9916 6860
rect 10968 6808 11020 6860
rect 11888 6808 11940 6860
rect 16212 6808 16264 6860
rect 17868 6808 17920 6860
rect 19616 6919 19668 6928
rect 19616 6885 19625 6919
rect 19625 6885 19659 6919
rect 19659 6885 19668 6919
rect 19616 6876 19668 6885
rect 20444 6876 20496 6928
rect 23848 6919 23900 6928
rect 23848 6885 23882 6919
rect 23882 6885 23900 6919
rect 23848 6876 23900 6885
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 9680 6715 9732 6724
rect 9680 6681 9689 6715
rect 9689 6681 9723 6715
rect 9723 6681 9732 6715
rect 9680 6672 9732 6681
rect 10048 6672 10100 6724
rect 10784 6740 10836 6792
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 16856 6740 16908 6792
rect 17776 6783 17828 6792
rect 17776 6749 17785 6783
rect 17785 6749 17819 6783
rect 17819 6749 17828 6783
rect 17776 6740 17828 6749
rect 19524 6740 19576 6792
rect 20812 6808 20864 6860
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 23572 6783 23624 6792
rect 15660 6715 15712 6724
rect 15660 6681 15669 6715
rect 15669 6681 15703 6715
rect 15703 6681 15712 6715
rect 15660 6672 15712 6681
rect 17224 6715 17276 6724
rect 17224 6681 17233 6715
rect 17233 6681 17267 6715
rect 17267 6681 17276 6715
rect 17224 6672 17276 6681
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 9036 6604 9088 6613
rect 11152 6647 11204 6656
rect 11152 6613 11161 6647
rect 11161 6613 11195 6647
rect 11195 6613 11204 6647
rect 11152 6604 11204 6613
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 14740 6604 14792 6656
rect 18052 6604 18104 6656
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 18788 6604 18840 6613
rect 20352 6647 20404 6656
rect 20352 6613 20361 6647
rect 20361 6613 20395 6647
rect 20395 6613 20404 6647
rect 20352 6604 20404 6613
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 20904 6604 20956 6656
rect 23572 6749 23581 6783
rect 23581 6749 23615 6783
rect 23615 6749 23624 6783
rect 23572 6740 23624 6749
rect 22284 6647 22336 6656
rect 22284 6613 22293 6647
rect 22293 6613 22327 6647
rect 22327 6613 22336 6647
rect 22284 6604 22336 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 10048 6400 10100 6452
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 13728 6400 13780 6452
rect 14096 6400 14148 6452
rect 15844 6400 15896 6452
rect 16856 6400 16908 6452
rect 18880 6443 18932 6452
rect 18880 6409 18889 6443
rect 18889 6409 18923 6443
rect 18923 6409 18932 6443
rect 18880 6400 18932 6409
rect 20536 6400 20588 6452
rect 23848 6400 23900 6452
rect 16120 6332 16172 6384
rect 19064 6332 19116 6384
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 18788 6264 18840 6316
rect 19340 6264 19392 6316
rect 20260 6264 20312 6316
rect 20536 6264 20588 6316
rect 20812 6264 20864 6316
rect 8668 6196 8720 6248
rect 9036 6239 9088 6248
rect 9036 6205 9045 6239
rect 9045 6205 9079 6239
rect 9079 6205 9088 6239
rect 9036 6196 9088 6205
rect 16212 6239 16264 6248
rect 16212 6205 16221 6239
rect 16221 6205 16255 6239
rect 16255 6205 16264 6239
rect 16212 6196 16264 6205
rect 9128 6128 9180 6180
rect 18880 6196 18932 6248
rect 20628 6196 20680 6248
rect 23572 6264 23624 6316
rect 21272 6239 21324 6248
rect 21272 6205 21306 6239
rect 21306 6205 21324 6239
rect 20904 6128 20956 6180
rect 21272 6196 21324 6205
rect 22284 6196 22336 6248
rect 21364 6128 21416 6180
rect 22652 6128 22704 6180
rect 24584 6128 24636 6180
rect 10692 6060 10744 6112
rect 11152 6060 11204 6112
rect 12256 6103 12308 6112
rect 12256 6069 12265 6103
rect 12265 6069 12299 6103
rect 12299 6069 12308 6103
rect 12256 6060 12308 6069
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 13452 6060 13504 6069
rect 14188 6103 14240 6112
rect 14188 6069 14197 6103
rect 14197 6069 14231 6103
rect 14231 6069 14240 6103
rect 14188 6060 14240 6069
rect 14648 6103 14700 6112
rect 14648 6069 14657 6103
rect 14657 6069 14691 6103
rect 14691 6069 14700 6103
rect 14648 6060 14700 6069
rect 15936 6060 15988 6112
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 17500 6103 17552 6112
rect 17500 6069 17509 6103
rect 17509 6069 17543 6103
rect 17543 6069 17552 6103
rect 17500 6060 17552 6069
rect 17776 6103 17828 6112
rect 17776 6069 17785 6103
rect 17785 6069 17819 6103
rect 17819 6069 17828 6103
rect 17776 6060 17828 6069
rect 18972 6060 19024 6112
rect 19524 6060 19576 6112
rect 20444 6103 20496 6112
rect 20444 6069 20453 6103
rect 20453 6069 20487 6103
rect 20487 6069 20496 6103
rect 20444 6060 20496 6069
rect 22192 6060 22244 6112
rect 22376 6103 22428 6112
rect 22376 6069 22385 6103
rect 22385 6069 22419 6103
rect 22419 6069 22428 6103
rect 22376 6060 22428 6069
rect 25044 6060 25096 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 9128 5899 9180 5908
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 9864 5899 9916 5908
rect 9864 5865 9873 5899
rect 9873 5865 9907 5899
rect 9907 5865 9916 5899
rect 9864 5856 9916 5865
rect 10140 5856 10192 5908
rect 11888 5899 11940 5908
rect 11888 5865 11897 5899
rect 11897 5865 11931 5899
rect 11931 5865 11940 5899
rect 11888 5856 11940 5865
rect 12992 5899 13044 5908
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 13268 5856 13320 5908
rect 18328 5856 18380 5908
rect 19064 5856 19116 5908
rect 19248 5856 19300 5908
rect 19432 5856 19484 5908
rect 20352 5899 20404 5908
rect 12532 5831 12584 5840
rect 12532 5797 12541 5831
rect 12541 5797 12575 5831
rect 12575 5797 12584 5831
rect 12532 5788 12584 5797
rect 12900 5788 12952 5840
rect 17224 5788 17276 5840
rect 10600 5720 10652 5772
rect 10784 5763 10836 5772
rect 10784 5729 10818 5763
rect 10818 5729 10836 5763
rect 10784 5720 10836 5729
rect 12348 5720 12400 5772
rect 15660 5763 15712 5772
rect 15660 5729 15669 5763
rect 15669 5729 15703 5763
rect 15703 5729 15712 5763
rect 15660 5720 15712 5729
rect 12440 5652 12492 5704
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 12900 5627 12952 5636
rect 12900 5593 12909 5627
rect 12909 5593 12943 5627
rect 12943 5593 12952 5627
rect 15752 5652 15804 5704
rect 16396 5652 16448 5704
rect 16672 5652 16724 5704
rect 19432 5720 19484 5772
rect 20352 5865 20361 5899
rect 20361 5865 20395 5899
rect 20395 5865 20404 5899
rect 20352 5856 20404 5865
rect 20536 5856 20588 5908
rect 20720 5856 20772 5908
rect 21180 5856 21232 5908
rect 23664 5899 23716 5908
rect 23664 5865 23673 5899
rect 23673 5865 23707 5899
rect 23707 5865 23716 5899
rect 23664 5856 23716 5865
rect 23756 5856 23808 5908
rect 23848 5788 23900 5840
rect 20168 5720 20220 5772
rect 20720 5720 20772 5772
rect 19892 5652 19944 5704
rect 23112 5720 23164 5772
rect 23296 5720 23348 5772
rect 23664 5720 23716 5772
rect 12900 5584 12952 5593
rect 15936 5584 15988 5636
rect 21088 5584 21140 5636
rect 22008 5652 22060 5704
rect 24676 5720 24728 5772
rect 25596 5720 25648 5772
rect 21916 5584 21968 5636
rect 23572 5584 23624 5636
rect 25044 5627 25096 5636
rect 25044 5593 25053 5627
rect 25053 5593 25087 5627
rect 25087 5593 25096 5627
rect 25044 5584 25096 5593
rect 15844 5559 15896 5568
rect 15844 5525 15853 5559
rect 15853 5525 15887 5559
rect 15887 5525 15896 5559
rect 15844 5516 15896 5525
rect 16580 5516 16632 5568
rect 17776 5516 17828 5568
rect 22100 5559 22152 5568
rect 22100 5525 22109 5559
rect 22109 5525 22143 5559
rect 22143 5525 22152 5559
rect 22100 5516 22152 5525
rect 22652 5516 22704 5568
rect 25412 5559 25464 5568
rect 25412 5525 25421 5559
rect 25421 5525 25455 5559
rect 25455 5525 25464 5559
rect 25412 5516 25464 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 10784 5312 10836 5364
rect 12348 5312 12400 5364
rect 17224 5312 17276 5364
rect 18512 5312 18564 5364
rect 16672 5244 16724 5296
rect 12348 5176 12400 5228
rect 8668 5151 8720 5160
rect 8668 5117 8677 5151
rect 8677 5117 8711 5151
rect 8711 5117 8720 5151
rect 8668 5108 8720 5117
rect 12900 5151 12952 5160
rect 12900 5117 12934 5151
rect 12934 5117 12952 5151
rect 9496 5040 9548 5092
rect 12348 5040 12400 5092
rect 12900 5108 12952 5117
rect 14740 5108 14792 5160
rect 15108 5151 15160 5160
rect 15108 5117 15117 5151
rect 15117 5117 15151 5151
rect 15151 5117 15160 5151
rect 15108 5108 15160 5117
rect 16488 5108 16540 5160
rect 19156 5312 19208 5364
rect 19340 5355 19392 5364
rect 19340 5321 19349 5355
rect 19349 5321 19383 5355
rect 19383 5321 19392 5355
rect 19340 5312 19392 5321
rect 21180 5312 21232 5364
rect 22008 5355 22060 5364
rect 21732 5244 21784 5296
rect 22008 5321 22017 5355
rect 22017 5321 22051 5355
rect 22051 5321 22060 5355
rect 22008 5312 22060 5321
rect 23112 5355 23164 5364
rect 23112 5321 23121 5355
rect 23121 5321 23155 5355
rect 23155 5321 23164 5355
rect 23112 5312 23164 5321
rect 23664 5312 23716 5364
rect 25596 5355 25648 5364
rect 25596 5321 25605 5355
rect 25605 5321 25639 5355
rect 25639 5321 25648 5355
rect 25596 5312 25648 5321
rect 22100 5244 22152 5296
rect 19892 5219 19944 5228
rect 19892 5185 19901 5219
rect 19901 5185 19935 5219
rect 19935 5185 19944 5219
rect 19892 5176 19944 5185
rect 20904 5151 20956 5160
rect 20904 5117 20913 5151
rect 20913 5117 20947 5151
rect 20947 5117 20956 5151
rect 20904 5108 20956 5117
rect 21824 5151 21876 5160
rect 21824 5117 21833 5151
rect 21833 5117 21867 5151
rect 21867 5117 21876 5151
rect 22652 5219 22704 5228
rect 22652 5185 22661 5219
rect 22661 5185 22695 5219
rect 22695 5185 22704 5219
rect 22652 5176 22704 5185
rect 21824 5108 21876 5117
rect 23388 5108 23440 5160
rect 23664 5151 23716 5160
rect 23664 5117 23673 5151
rect 23673 5117 23707 5151
rect 23707 5117 23716 5151
rect 23664 5108 23716 5117
rect 13452 5040 13504 5092
rect 18604 5040 18656 5092
rect 9128 4972 9180 5024
rect 10692 4972 10744 5024
rect 12992 4972 13044 5024
rect 15016 5015 15068 5024
rect 15016 4981 15025 5015
rect 15025 4981 15059 5015
rect 15059 4981 15068 5015
rect 15016 4972 15068 4981
rect 16488 5015 16540 5024
rect 16488 4981 16497 5015
rect 16497 4981 16531 5015
rect 16531 4981 16540 5015
rect 16488 4972 16540 4981
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 18052 4972 18104 5024
rect 18420 5015 18472 5024
rect 18420 4981 18429 5015
rect 18429 4981 18463 5015
rect 18463 4981 18472 5015
rect 18420 4972 18472 4981
rect 19156 5015 19208 5024
rect 19156 4981 19165 5015
rect 19165 4981 19199 5015
rect 19199 4981 19208 5015
rect 19156 4972 19208 4981
rect 20076 5040 20128 5092
rect 20168 5040 20220 5092
rect 23112 5040 23164 5092
rect 25044 5108 25096 5160
rect 23940 5083 23992 5092
rect 23940 5049 23974 5083
rect 23974 5049 23992 5083
rect 23940 5040 23992 5049
rect 24676 5040 24728 5092
rect 20812 5015 20864 5024
rect 20812 4981 20821 5015
rect 20821 4981 20855 5015
rect 20855 4981 20864 5015
rect 20812 4972 20864 4981
rect 25136 4972 25188 5024
rect 25596 4972 25648 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 9128 4768 9180 4820
rect 10140 4768 10192 4820
rect 11612 4811 11664 4820
rect 11612 4777 11621 4811
rect 11621 4777 11655 4811
rect 11655 4777 11664 4811
rect 11612 4768 11664 4777
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 13544 4768 13596 4820
rect 16396 4768 16448 4820
rect 17592 4768 17644 4820
rect 19248 4768 19300 4820
rect 20720 4811 20772 4820
rect 20720 4777 20729 4811
rect 20729 4777 20763 4811
rect 20763 4777 20772 4811
rect 20720 4768 20772 4777
rect 22468 4768 22520 4820
rect 23940 4811 23992 4820
rect 23940 4777 23949 4811
rect 23949 4777 23983 4811
rect 23983 4777 23992 4811
rect 23940 4768 23992 4777
rect 24216 4768 24268 4820
rect 24768 4768 24820 4820
rect 25228 4768 25280 4820
rect 9680 4632 9732 4684
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 12992 4700 13044 4752
rect 17868 4700 17920 4752
rect 21456 4700 21508 4752
rect 23020 4700 23072 4752
rect 25044 4700 25096 4752
rect 15568 4675 15620 4684
rect 15568 4641 15602 4675
rect 15602 4641 15620 4675
rect 15568 4632 15620 4641
rect 17408 4632 17460 4684
rect 19524 4632 19576 4684
rect 19984 4632 20036 4684
rect 20996 4632 21048 4684
rect 21548 4632 21600 4684
rect 23664 4632 23716 4684
rect 9772 4496 9824 4548
rect 10692 4564 10744 4616
rect 12348 4564 12400 4616
rect 12532 4564 12584 4616
rect 15108 4607 15160 4616
rect 15108 4573 15117 4607
rect 15117 4573 15151 4607
rect 15151 4573 15160 4607
rect 15108 4564 15160 4573
rect 10968 4496 11020 4548
rect 8208 4471 8260 4480
rect 8208 4437 8217 4471
rect 8217 4437 8251 4471
rect 8251 4437 8260 4471
rect 8208 4428 8260 4437
rect 8668 4428 8720 4480
rect 9036 4471 9088 4480
rect 9036 4437 9045 4471
rect 9045 4437 9079 4471
rect 9079 4437 9088 4471
rect 9036 4428 9088 4437
rect 10692 4471 10744 4480
rect 10692 4437 10701 4471
rect 10701 4437 10735 4471
rect 10735 4437 10744 4471
rect 10692 4428 10744 4437
rect 17960 4564 18012 4616
rect 18512 4564 18564 4616
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 20076 4564 20128 4616
rect 25136 4607 25188 4616
rect 25136 4573 25145 4607
rect 25145 4573 25179 4607
rect 25179 4573 25188 4607
rect 25136 4564 25188 4573
rect 19984 4496 20036 4548
rect 16212 4428 16264 4480
rect 16672 4428 16724 4480
rect 17868 4428 17920 4480
rect 19892 4471 19944 4480
rect 19892 4437 19901 4471
rect 19901 4437 19935 4471
rect 19935 4437 19944 4471
rect 19892 4428 19944 4437
rect 20260 4471 20312 4480
rect 20260 4437 20269 4471
rect 20269 4437 20303 4471
rect 20303 4437 20312 4471
rect 20260 4428 20312 4437
rect 22008 4428 22060 4480
rect 23664 4428 23716 4480
rect 25596 4471 25648 4480
rect 25596 4437 25605 4471
rect 25605 4437 25639 4471
rect 25639 4437 25648 4471
rect 25596 4428 25648 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 8208 4156 8260 4208
rect 10784 4224 10836 4276
rect 15936 4267 15988 4276
rect 15936 4233 15945 4267
rect 15945 4233 15979 4267
rect 15979 4233 15988 4267
rect 15936 4224 15988 4233
rect 17224 4224 17276 4276
rect 19524 4267 19576 4276
rect 19524 4233 19533 4267
rect 19533 4233 19567 4267
rect 19567 4233 19576 4267
rect 19524 4224 19576 4233
rect 20996 4267 21048 4276
rect 20996 4233 21005 4267
rect 21005 4233 21039 4267
rect 21039 4233 21048 4267
rect 20996 4224 21048 4233
rect 23020 4224 23072 4276
rect 25228 4224 25280 4276
rect 9496 4131 9548 4140
rect 9496 4097 9505 4131
rect 9505 4097 9539 4131
rect 9539 4097 9548 4131
rect 9496 4088 9548 4097
rect 12072 4088 12124 4140
rect 8576 4020 8628 4072
rect 9036 4020 9088 4072
rect 9588 4020 9640 4072
rect 10692 4020 10744 4072
rect 12992 4088 13044 4140
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 15568 4088 15620 4140
rect 16488 4131 16540 4140
rect 16488 4097 16497 4131
rect 16497 4097 16531 4131
rect 16531 4097 16540 4131
rect 16488 4088 16540 4097
rect 17408 4131 17460 4140
rect 17408 4097 17417 4131
rect 17417 4097 17451 4131
rect 17451 4097 17460 4131
rect 17408 4088 17460 4097
rect 18052 4088 18104 4140
rect 18604 4131 18656 4140
rect 18604 4097 18613 4131
rect 18613 4097 18647 4131
rect 18647 4097 18656 4131
rect 23388 4156 23440 4208
rect 18604 4088 18656 4097
rect 15936 4020 15988 4072
rect 18144 4020 18196 4072
rect 18696 4020 18748 4072
rect 7656 3927 7708 3936
rect 7656 3893 7665 3927
rect 7665 3893 7699 3927
rect 7699 3893 7708 3927
rect 7656 3884 7708 3893
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 9496 3952 9548 4004
rect 12072 3952 12124 4004
rect 13084 3952 13136 4004
rect 8760 3884 8812 3936
rect 9772 3884 9824 3936
rect 12440 3884 12492 3936
rect 14188 3927 14240 3936
rect 14188 3893 14197 3927
rect 14197 3893 14231 3927
rect 14231 3893 14240 3927
rect 14188 3884 14240 3893
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 15660 3884 15712 3936
rect 17868 3952 17920 4004
rect 19156 3995 19208 4004
rect 19156 3961 19165 3995
rect 19165 3961 19199 3995
rect 19199 3961 19208 3995
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 22376 4131 22428 4140
rect 22376 4097 22385 4131
rect 22385 4097 22419 4131
rect 22419 4097 22428 4131
rect 22376 4088 22428 4097
rect 20168 4020 20220 4072
rect 23296 4020 23348 4072
rect 23940 4063 23992 4072
rect 23940 4029 23949 4063
rect 23949 4029 23983 4063
rect 23983 4029 23992 4063
rect 23940 4020 23992 4029
rect 24216 4063 24268 4072
rect 24216 4029 24250 4063
rect 24250 4029 24268 4063
rect 24216 4020 24268 4029
rect 19156 3952 19208 3961
rect 17592 3884 17644 3936
rect 17960 3884 18012 3936
rect 18144 3884 18196 3936
rect 18420 3927 18472 3936
rect 18420 3893 18429 3927
rect 18429 3893 18463 3927
rect 18463 3893 18472 3927
rect 18420 3884 18472 3893
rect 19524 3884 19576 3936
rect 21456 3884 21508 3936
rect 21640 3884 21692 3936
rect 22008 3884 22060 3936
rect 22100 3927 22152 3936
rect 22100 3893 22109 3927
rect 22109 3893 22143 3927
rect 22143 3893 22152 3927
rect 25320 3927 25372 3936
rect 22100 3884 22152 3893
rect 25320 3893 25329 3927
rect 25329 3893 25363 3927
rect 25363 3893 25372 3927
rect 25320 3884 25372 3893
rect 26240 3927 26292 3936
rect 26240 3893 26249 3927
rect 26249 3893 26283 3927
rect 26283 3893 26292 3927
rect 26240 3884 26292 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 7012 3723 7064 3732
rect 7012 3689 7021 3723
rect 7021 3689 7055 3723
rect 7055 3689 7064 3723
rect 7012 3680 7064 3689
rect 7656 3680 7708 3732
rect 9956 3723 10008 3732
rect 9956 3689 9965 3723
rect 9965 3689 9999 3723
rect 9999 3689 10008 3723
rect 9956 3680 10008 3689
rect 10692 3680 10744 3732
rect 8484 3612 8536 3664
rect 8392 3587 8444 3596
rect 8392 3553 8401 3587
rect 8401 3553 8435 3587
rect 8435 3553 8444 3587
rect 8392 3544 8444 3553
rect 7472 3476 7524 3528
rect 8760 3544 8812 3596
rect 9312 3544 9364 3596
rect 10968 3544 11020 3596
rect 11060 3476 11112 3528
rect 13084 3680 13136 3732
rect 14372 3680 14424 3732
rect 15568 3680 15620 3732
rect 15936 3723 15988 3732
rect 15936 3689 15945 3723
rect 15945 3689 15979 3723
rect 15979 3689 15988 3723
rect 15936 3680 15988 3689
rect 20168 3723 20220 3732
rect 20168 3689 20177 3723
rect 20177 3689 20211 3723
rect 20211 3689 20220 3723
rect 20168 3680 20220 3689
rect 21088 3723 21140 3732
rect 21088 3689 21097 3723
rect 21097 3689 21131 3723
rect 21131 3689 21140 3723
rect 21088 3680 21140 3689
rect 23020 3680 23072 3732
rect 23480 3680 23532 3732
rect 24124 3680 24176 3732
rect 24676 3680 24728 3732
rect 24768 3680 24820 3732
rect 25044 3723 25096 3732
rect 25044 3689 25053 3723
rect 25053 3689 25087 3723
rect 25087 3689 25096 3723
rect 25044 3680 25096 3689
rect 25596 3680 25648 3732
rect 11520 3612 11572 3664
rect 12992 3612 13044 3664
rect 19524 3655 19576 3664
rect 19524 3621 19533 3655
rect 19533 3621 19567 3655
rect 19567 3621 19576 3655
rect 19524 3612 19576 3621
rect 22192 3612 22244 3664
rect 13728 3544 13780 3596
rect 14280 3544 14332 3596
rect 15476 3544 15528 3596
rect 16580 3544 16632 3596
rect 20628 3544 20680 3596
rect 21548 3587 21600 3596
rect 21548 3553 21557 3587
rect 21557 3553 21591 3587
rect 21591 3553 21600 3587
rect 21548 3544 21600 3553
rect 22284 3544 22336 3596
rect 23204 3612 23256 3664
rect 23848 3612 23900 3664
rect 23940 3612 23992 3664
rect 26148 3612 26200 3664
rect 25044 3544 25096 3596
rect 14924 3408 14976 3460
rect 15568 3408 15620 3460
rect 8576 3340 8628 3392
rect 9496 3383 9548 3392
rect 9496 3349 9505 3383
rect 9505 3349 9539 3383
rect 9539 3349 9548 3383
rect 9496 3340 9548 3349
rect 11520 3340 11572 3392
rect 11704 3340 11756 3392
rect 13912 3340 13964 3392
rect 15292 3340 15344 3392
rect 16212 3340 16264 3392
rect 19800 3519 19852 3528
rect 19800 3485 19809 3519
rect 19809 3485 19843 3519
rect 19843 3485 19852 3519
rect 19800 3476 19852 3485
rect 25136 3476 25188 3528
rect 26240 3476 26292 3528
rect 19156 3451 19208 3460
rect 19156 3417 19165 3451
rect 19165 3417 19199 3451
rect 19199 3417 19208 3451
rect 19156 3408 19208 3417
rect 23940 3408 23992 3460
rect 24584 3408 24636 3460
rect 17868 3383 17920 3392
rect 17868 3349 17877 3383
rect 17877 3349 17911 3383
rect 17911 3349 17920 3383
rect 17868 3340 17920 3349
rect 18604 3340 18656 3392
rect 21088 3340 21140 3392
rect 21916 3340 21968 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 7472 3179 7524 3188
rect 7472 3145 7481 3179
rect 7481 3145 7515 3179
rect 7515 3145 7524 3179
rect 7472 3136 7524 3145
rect 8024 3136 8076 3188
rect 8392 3136 8444 3188
rect 9496 3136 9548 3188
rect 11060 3136 11112 3188
rect 11704 3136 11756 3188
rect 12624 3179 12676 3188
rect 12624 3145 12633 3179
rect 12633 3145 12667 3179
rect 12667 3145 12676 3179
rect 12624 3136 12676 3145
rect 13728 3179 13780 3188
rect 13728 3145 13737 3179
rect 13737 3145 13771 3179
rect 13771 3145 13780 3179
rect 13728 3136 13780 3145
rect 15476 3136 15528 3188
rect 19524 3136 19576 3188
rect 19800 3136 19852 3188
rect 22284 3136 22336 3188
rect 23664 3179 23716 3188
rect 23664 3145 23673 3179
rect 23673 3145 23707 3179
rect 23707 3145 23716 3179
rect 23664 3136 23716 3145
rect 24676 3179 24728 3188
rect 24676 3145 24685 3179
rect 24685 3145 24719 3179
rect 24719 3145 24728 3179
rect 24676 3136 24728 3145
rect 25136 3179 25188 3188
rect 25136 3145 25145 3179
rect 25145 3145 25179 3179
rect 25179 3145 25188 3179
rect 25136 3136 25188 3145
rect 26148 3179 26200 3188
rect 26148 3145 26157 3179
rect 26157 3145 26191 3179
rect 26191 3145 26200 3179
rect 26148 3136 26200 3145
rect 7932 3111 7984 3120
rect 7932 3077 7941 3111
rect 7941 3077 7975 3111
rect 7975 3077 7984 3111
rect 7932 3068 7984 3077
rect 8576 3043 8628 3052
rect 8576 3009 8585 3043
rect 8585 3009 8619 3043
rect 8619 3009 8628 3043
rect 8576 3000 8628 3009
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 13360 3000 13412 3052
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 26240 3068 26292 3120
rect 17776 3000 17828 3009
rect 9312 2975 9364 2984
rect 9312 2941 9321 2975
rect 9321 2941 9355 2975
rect 9355 2941 9364 2975
rect 9312 2932 9364 2941
rect 9588 2932 9640 2984
rect 11060 2932 11112 2984
rect 11796 2932 11848 2984
rect 8484 2864 8536 2916
rect 16212 2932 16264 2984
rect 16580 2975 16632 2984
rect 16580 2941 16589 2975
rect 16589 2941 16623 2975
rect 16623 2941 16632 2975
rect 16580 2932 16632 2941
rect 16764 2932 16816 2984
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 20076 2932 20128 2984
rect 20536 2975 20588 2984
rect 20536 2941 20545 2975
rect 20545 2941 20579 2975
rect 20579 2941 20588 2975
rect 20536 2932 20588 2941
rect 23572 2932 23624 2984
rect 23848 2932 23900 2984
rect 6828 2796 6880 2848
rect 8208 2796 8260 2848
rect 15108 2864 15160 2916
rect 17684 2864 17736 2916
rect 20260 2864 20312 2916
rect 21824 2864 21876 2916
rect 23480 2907 23532 2916
rect 23480 2873 23489 2907
rect 23489 2873 23523 2907
rect 23523 2873 23532 2907
rect 23480 2864 23532 2873
rect 12440 2796 12492 2848
rect 15568 2839 15620 2848
rect 15568 2805 15577 2839
rect 15577 2805 15611 2839
rect 15611 2805 15620 2839
rect 15568 2796 15620 2805
rect 16580 2796 16632 2848
rect 17316 2796 17368 2848
rect 17776 2796 17828 2848
rect 25412 2839 25464 2848
rect 25412 2805 25421 2839
rect 25421 2805 25455 2839
rect 25455 2805 25464 2839
rect 25412 2796 25464 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 7104 2635 7156 2644
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 6920 2524 6972 2576
rect 8208 2592 8260 2644
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 10784 2592 10836 2644
rect 10968 2635 11020 2644
rect 10968 2601 10977 2635
rect 10977 2601 11011 2635
rect 11011 2601 11020 2635
rect 10968 2592 11020 2601
rect 12072 2635 12124 2644
rect 12072 2601 12081 2635
rect 12081 2601 12115 2635
rect 12115 2601 12124 2635
rect 12072 2592 12124 2601
rect 15568 2592 15620 2644
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 20076 2592 20128 2644
rect 20628 2592 20680 2644
rect 21640 2635 21692 2644
rect 21640 2601 21649 2635
rect 21649 2601 21683 2635
rect 21683 2601 21692 2635
rect 21640 2592 21692 2601
rect 22284 2635 22336 2644
rect 22284 2601 22293 2635
rect 22293 2601 22327 2635
rect 22327 2601 22336 2635
rect 22284 2592 22336 2601
rect 12440 2567 12492 2576
rect 12440 2533 12449 2567
rect 12449 2533 12483 2567
rect 12483 2533 12492 2567
rect 12440 2524 12492 2533
rect 13360 2524 13412 2576
rect 16212 2524 16264 2576
rect 19432 2524 19484 2576
rect 10784 2456 10836 2508
rect 12532 2456 12584 2508
rect 19524 2456 19576 2508
rect 22008 2524 22060 2576
rect 23296 2592 23348 2644
rect 23388 2592 23440 2644
rect 21548 2499 21600 2508
rect 21548 2465 21557 2499
rect 21557 2465 21591 2499
rect 21591 2465 21600 2499
rect 21548 2456 21600 2465
rect 22100 2456 22152 2508
rect 23940 2524 23992 2576
rect 24216 2592 24268 2644
rect 25872 2592 25924 2644
rect 25044 2524 25096 2576
rect 23572 2456 23624 2508
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 11520 2388 11572 2440
rect 18052 2431 18104 2440
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 10784 2295 10836 2304
rect 10784 2261 10793 2295
rect 10793 2261 10827 2295
rect 10827 2261 10836 2295
rect 10784 2252 10836 2261
rect 18052 2397 18061 2431
rect 18061 2397 18095 2431
rect 18095 2397 18104 2431
rect 18052 2388 18104 2397
rect 18144 2388 18196 2440
rect 21824 2431 21876 2440
rect 21824 2397 21833 2431
rect 21833 2397 21867 2431
rect 21867 2397 21876 2431
rect 21824 2388 21876 2397
rect 22284 2388 22336 2440
rect 24860 2456 24912 2508
rect 23756 2320 23808 2372
rect 22652 2252 22704 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 23664 1368 23716 1420
rect 24032 1368 24084 1420
rect 22836 1232 22888 1284
rect 24308 1232 24360 1284
rect 15844 552 15896 604
rect 16120 552 16172 604
<< metal2 >>
rect 3514 27520 3570 28000
rect 10506 27520 10562 28000
rect 17498 27520 17554 28000
rect 24030 27704 24086 27713
rect 24030 27639 24086 27648
rect 3528 23526 3556 27520
rect 10520 27418 10548 27520
rect 10152 27390 10548 27418
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 10152 23866 10180 27390
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 12992 24880 13044 24886
rect 12992 24822 13044 24828
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 13004 23866 13032 24822
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 17512 23866 17540 27520
rect 23570 26616 23626 26625
rect 23570 26551 23626 26560
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17222 23760 17278 23769
rect 17222 23695 17278 23704
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 3516 23520 3568 23526
rect 3516 23462 3568 23468
rect 4068 23520 4120 23526
rect 10692 23520 10744 23526
rect 4068 23462 4120 23468
rect 10690 23488 10692 23497
rect 10744 23488 10746 23497
rect 4080 13433 4108 23462
rect 10289 23420 10585 23440
rect 10690 23423 10746 23432
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 12360 23254 12388 23598
rect 12348 23248 12400 23254
rect 12348 23190 12400 23196
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 11808 22438 11836 23122
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 13726 22672 13782 22681
rect 13726 22607 13782 22616
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 10060 21350 10088 22034
rect 10324 22024 10376 22030
rect 10322 21992 10324 22001
rect 10376 21992 10378 22001
rect 10322 21927 10378 21936
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 8114 16960 8170 16969
rect 8114 16895 8170 16904
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 4066 13424 4122 13433
rect 4066 13359 4122 13368
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 7930 10976 7986 10985
rect 5622 10908 5918 10928
rect 7930 10911 7986 10920
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 1582 9480 1638 9489
rect 1582 9415 1638 9424
rect 294 8120 350 8129
rect 294 8055 350 8064
rect 308 480 336 8055
rect 938 7440 994 7449
rect 938 7375 994 7384
rect 952 480 980 7375
rect 1596 480 1624 9415
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 2226 8528 2282 8537
rect 2226 8463 2282 8472
rect 2240 480 2268 8463
rect 7010 7984 7066 7993
rect 7010 7919 7066 7928
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5446 7304 5502 7313
rect 5446 7239 5502 7248
rect 3514 4584 3570 4593
rect 3514 4519 3570 4528
rect 2870 4176 2926 4185
rect 2870 4111 2926 4120
rect 2884 480 2912 4111
rect 3528 480 3556 4519
rect 4802 1728 4858 1737
rect 4802 1663 4858 1672
rect 4158 1592 4214 1601
rect 4158 1527 4214 1536
rect 4172 480 4200 1527
rect 4816 480 4844 1663
rect 5460 480 5488 7239
rect 6734 6896 6790 6905
rect 6734 6831 6790 6840
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6090 6216 6146 6225
rect 6090 6151 6146 6160
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6104 480 6132 6151
rect 6748 480 6776 6831
rect 7024 3738 7052 7919
rect 7378 5808 7434 5817
rect 7378 5743 7434 5752
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7102 2952 7158 2961
rect 7102 2887 7158 2896
rect 6828 2848 6880 2854
rect 6880 2808 6960 2836
rect 6828 2790 6880 2796
rect 6932 2582 6960 2808
rect 7116 2650 7144 2887
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 7392 480 7420 5743
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7668 3738 7696 3878
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 3194 7512 3470
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7944 3126 7972 10911
rect 8128 3942 8156 16895
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8574 6760 8630 6769
rect 8574 6695 8630 6704
rect 8588 5914 8616 6695
rect 9048 6662 9076 7142
rect 9692 6730 9720 21286
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11072 18086 11100 18770
rect 11334 18728 11390 18737
rect 11334 18663 11336 18672
rect 11388 18663 11390 18672
rect 11336 18634 11388 18640
rect 11060 18080 11112 18086
rect 10980 18028 11060 18034
rect 10980 18022 11112 18028
rect 10980 18006 11100 18022
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10980 17814 11008 18006
rect 10968 17808 11020 17814
rect 10968 17750 11020 17756
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10152 16998 10180 17682
rect 10140 16992 10192 16998
rect 10138 16960 10140 16969
rect 10192 16960 10194 16969
rect 10138 16895 10194 16904
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 9954 15328 10010 15337
rect 9954 15263 10010 15272
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 6254 9076 6598
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8680 5166 8708 6190
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9140 5914 9168 6122
rect 9876 5914 9904 6802
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8220 4214 8248 4422
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8588 4078 8616 4558
rect 8680 4486 8708 5102
rect 9140 5030 9168 5850
rect 9494 5128 9550 5137
rect 9494 5063 9496 5072
rect 9548 5063 9550 5072
rect 9496 5034 9548 5040
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9140 4826 9168 4966
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 9048 4078 9076 4422
rect 9494 4176 9550 4185
rect 9692 4162 9720 4626
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9550 4134 9720 4162
rect 9494 4111 9496 4120
rect 9548 4111 9550 4120
rect 9496 4082 9548 4088
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8404 3194 8432 3538
rect 8496 3505 8524 3606
rect 8772 3602 8800 3878
rect 9402 3632 9458 3641
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 9312 3596 9364 3602
rect 9402 3567 9458 3576
rect 9312 3538 9364 3544
rect 8482 3496 8538 3505
rect 8482 3431 8538 3440
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 8036 480 8064 3130
rect 8496 2922 8524 3431
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8588 3097 8616 3334
rect 8574 3088 8630 3097
rect 8574 3023 8576 3032
rect 8628 3023 8630 3032
rect 8576 2994 8628 3000
rect 9324 2990 9352 3538
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 8208 2848 8260 2854
rect 9416 2836 9444 3567
rect 9508 3398 9536 3946
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9508 3194 9536 3334
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9600 3074 9628 4014
rect 9784 3942 9812 4490
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9968 3738 9996 15263
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 11150 9616 11206 9625
rect 11150 9551 11206 9560
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10690 9208 10746 9217
rect 10690 9143 10692 9152
rect 10744 9143 10746 9152
rect 10692 9114 10744 9120
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10598 8528 10654 8537
rect 10598 8463 10600 8472
rect 10652 8463 10654 8472
rect 10600 8434 10652 8440
rect 10704 8401 10732 8978
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10796 8634 10824 8910
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 11072 8566 11100 8910
rect 11060 8560 11112 8566
rect 10782 8528 10838 8537
rect 11060 8502 11112 8508
rect 10782 8463 10838 8472
rect 10690 8392 10746 8401
rect 10690 8327 10746 8336
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8022 10732 8327
rect 10796 8090 10824 8463
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10060 6730 10088 7210
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10796 6798 10824 7822
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10874 7304 10930 7313
rect 10874 7239 10930 7248
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 10060 6458 10088 6666
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10152 5914 10180 6734
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10152 4826 10180 5850
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10612 5658 10640 5714
rect 10704 5658 10732 6054
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10612 5630 10732 5658
rect 10704 5030 10732 5630
rect 10796 5370 10824 5714
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10704 4622 10732 4966
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10704 4486 10732 4558
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10704 4078 10732 4422
rect 10796 4282 10824 5306
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3738 10732 4014
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 9508 3058 9628 3074
rect 9496 3052 9628 3058
rect 9548 3046 9628 3052
rect 9496 2994 9548 3000
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 8208 2790 8260 2796
rect 9324 2808 9444 2836
rect 8220 2650 8248 2790
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8482 2544 8538 2553
rect 8482 2479 8484 2488
rect 8536 2479 8538 2488
rect 8484 2450 8536 2456
rect 8576 2440 8628 2446
rect 8760 2440 8812 2446
rect 8576 2382 8628 2388
rect 8758 2408 8760 2417
rect 8812 2408 8814 2417
rect 8588 2281 8616 2382
rect 8758 2343 8814 2352
rect 8574 2272 8630 2281
rect 8574 2207 8630 2216
rect 8666 2136 8722 2145
rect 8666 2071 8722 2080
rect 8680 480 8708 2071
rect 9324 480 9352 2808
rect 9600 2650 9628 2926
rect 10888 2802 10916 7239
rect 10980 6866 11008 7482
rect 11164 7449 11192 9551
rect 11808 9217 11836 22374
rect 13740 21554 13768 22607
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 17052 21690 17080 22034
rect 17236 21962 17264 23695
rect 18144 23656 18196 23662
rect 18196 23604 18276 23610
rect 18144 23598 18276 23604
rect 18156 23582 18276 23598
rect 18248 22982 18276 23582
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 17224 21956 17276 21962
rect 17224 21898 17276 21904
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 12992 21480 13044 21486
rect 12992 21422 13044 21428
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12714 17096 12770 17105
rect 12360 15337 12388 17070
rect 12714 17031 12716 17040
rect 12768 17031 12770 17040
rect 12716 17002 12768 17008
rect 12622 15872 12678 15881
rect 12622 15807 12678 15816
rect 12346 15328 12402 15337
rect 12346 15263 12402 15272
rect 11794 9208 11850 9217
rect 11794 9143 11850 9152
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11532 8498 11560 8774
rect 12176 8566 12204 8978
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11532 8022 11560 8434
rect 12176 8090 12204 8502
rect 12532 8424 12584 8430
rect 12438 8392 12494 8401
rect 12532 8366 12584 8372
rect 12438 8327 12440 8336
rect 12492 8327 12494 8336
rect 12440 8298 12492 8304
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11532 7546 11560 7958
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11150 7440 11206 7449
rect 11150 7375 11206 7384
rect 11978 7440 12034 7449
rect 11978 7375 12034 7384
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 6118 11192 6598
rect 11900 6458 11928 6802
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11610 6080 11666 6089
rect 11610 6015 11666 6024
rect 11334 5264 11390 5273
rect 11334 5199 11390 5208
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10980 3777 11008 4490
rect 10966 3768 11022 3777
rect 10966 3703 11022 3712
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10796 2774 10916 2802
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10796 2650 10824 2774
rect 10980 2650 11008 3538
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11072 3194 11100 3470
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11072 2990 11100 3130
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10796 2310 10824 2450
rect 10048 2304 10100 2310
rect 10784 2304 10836 2310
rect 10048 2246 10100 2252
rect 10690 2272 10746 2281
rect 10060 2009 10088 2246
rect 10784 2246 10836 2252
rect 10690 2207 10746 2216
rect 10046 2000 10102 2009
rect 10046 1935 10102 1944
rect 10046 1864 10102 1873
rect 10046 1799 10102 1808
rect 10060 480 10088 1799
rect 10704 480 10732 2207
rect 10796 2145 10824 2246
rect 10782 2136 10838 2145
rect 10782 2071 10838 2080
rect 11348 480 11376 5199
rect 11624 4826 11652 6015
rect 11900 5914 11928 6394
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11532 3398 11560 3606
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11532 2446 11560 3334
rect 11716 3194 11744 3334
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11796 2984 11848 2990
rect 11794 2952 11796 2961
rect 11848 2952 11850 2961
rect 11794 2887 11850 2896
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 11992 480 12020 7375
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12268 5817 12296 6054
rect 12544 5846 12572 8366
rect 12532 5840 12584 5846
rect 12254 5808 12310 5817
rect 12532 5782 12584 5788
rect 12254 5743 12310 5752
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12360 5370 12388 5714
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12452 5250 12480 5646
rect 12360 5234 12572 5250
rect 12348 5228 12572 5234
rect 12400 5222 12572 5228
rect 12348 5170 12400 5176
rect 12438 5128 12494 5137
rect 12348 5092 12400 5098
rect 12438 5063 12494 5072
rect 12348 5034 12400 5040
rect 12360 4622 12388 5034
rect 12452 4826 12480 5063
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12544 4706 12572 5222
rect 12452 4678 12572 4706
rect 12348 4616 12400 4622
rect 12070 4584 12126 4593
rect 12348 4558 12400 4564
rect 12070 4519 12126 4528
rect 12084 4146 12112 4519
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 12084 2650 12112 3946
rect 12452 3942 12480 4678
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12452 2582 12480 2790
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12544 2514 12572 4558
rect 12636 3194 12664 15807
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12820 9518 12848 9862
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12820 8838 12848 9454
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12820 7818 12848 8774
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12912 5846 12940 6054
rect 13004 5914 13032 21422
rect 17052 21350 17080 21626
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 16224 21078 16252 21286
rect 16212 21072 16264 21078
rect 16212 21014 16264 21020
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15856 20262 15884 20946
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13450 18184 13506 18193
rect 13174 9480 13230 9489
rect 13174 9415 13230 9424
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13096 8022 13124 9318
rect 13188 8634 13216 9415
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13280 8090 13308 18158
rect 13450 18119 13452 18128
rect 13504 18119 13506 18128
rect 13452 18090 13504 18096
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 13634 16144 13690 16153
rect 13634 16079 13690 16088
rect 13648 10266 13676 16079
rect 15200 15904 15252 15910
rect 15198 15872 15200 15881
rect 15252 15872 15254 15881
rect 15198 15807 15254 15816
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 13818 14920 13874 14929
rect 13818 14855 13874 14864
rect 13832 10985 13860 14855
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14554 12744 14610 12753
rect 14554 12679 14610 12688
rect 13910 11656 13966 11665
rect 13910 11591 13966 11600
rect 13924 11218 13952 11591
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13818 10976 13874 10985
rect 13818 10911 13874 10920
rect 13924 10810 13952 11154
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13740 10130 13768 10406
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 13372 9722 13400 10066
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13556 9518 13584 9862
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13556 9178 13584 9454
rect 14108 9178 14136 10066
rect 14200 10062 14228 10542
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14200 9450 14228 9998
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13372 8362 13400 8502
rect 14016 8498 14044 9114
rect 14108 8634 14136 9114
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 13096 7546 13124 7958
rect 13464 7818 13492 8298
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13188 7546 13216 7686
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13464 6118 13492 7754
rect 13556 7342 13584 7754
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13556 7002 13584 7278
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13740 6458 13768 7822
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6458 14136 6598
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 12900 5840 12952 5846
rect 12898 5808 12900 5817
rect 12952 5808 12954 5817
rect 12898 5743 12954 5752
rect 12912 5717 12940 5743
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12912 5166 12940 5578
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12992 5024 13044 5030
rect 12714 4992 12770 5001
rect 12992 4966 13044 4972
rect 12714 4927 12770 4936
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12728 2394 12756 4927
rect 13004 4758 13032 4966
rect 12992 4752 13044 4758
rect 12992 4694 13044 4700
rect 13004 4146 13032 4694
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13004 3670 13032 4082
rect 13082 4040 13138 4049
rect 13082 3975 13084 3984
rect 13136 3975 13138 3984
rect 13084 3946 13136 3952
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 13096 3058 13124 3674
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 12636 2366 12756 2394
rect 12636 480 12664 2366
rect 13280 480 13308 5850
rect 13464 5098 13492 6054
rect 13544 5704 13596 5710
rect 14200 5681 14228 6054
rect 13544 5646 13596 5652
rect 14186 5672 14242 5681
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 13556 4826 13584 5646
rect 14186 5607 14242 5616
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14200 3641 14228 3878
rect 14186 3632 14242 3641
rect 13728 3596 13780 3602
rect 14292 3602 14320 11086
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 3738 14412 3878
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14186 3567 14242 3576
rect 14280 3596 14332 3602
rect 13728 3538 13780 3544
rect 14280 3538 14332 3544
rect 13740 3194 13768 3538
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13372 2689 13400 2994
rect 13358 2680 13414 2689
rect 13358 2615 13414 2624
rect 13372 2582 13400 2615
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 13924 480 13952 3334
rect 14568 480 14596 12679
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14752 9926 14780 10542
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14648 7744 14700 7750
rect 14752 7721 14780 9454
rect 15304 9178 15332 18022
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15580 16726 15608 17070
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15396 15910 15424 16594
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15382 11248 15438 11257
rect 15382 11183 15384 11192
rect 15436 11183 15438 11192
rect 15384 11154 15436 11160
rect 15396 10266 15424 11154
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15396 9058 15424 9862
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 15304 9030 15424 9058
rect 14844 8566 14872 8978
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14832 8560 14884 8566
rect 14830 8528 14832 8537
rect 14884 8528 14886 8537
rect 14830 8463 14886 8472
rect 15304 8430 15332 9030
rect 15108 8424 15160 8430
rect 15292 8424 15344 8430
rect 15160 8372 15240 8378
rect 15108 8366 15240 8372
rect 15292 8366 15344 8372
rect 15120 8350 15240 8366
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15120 7954 15148 8230
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 14832 7744 14884 7750
rect 14648 7686 14700 7692
rect 14738 7712 14794 7721
rect 14660 7562 14688 7686
rect 15212 7732 15240 8350
rect 15304 7886 15332 8366
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15212 7704 15332 7732
rect 14832 7686 14884 7692
rect 14738 7647 14794 7656
rect 14660 7534 14780 7562
rect 14844 7546 14872 7686
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14660 7002 14688 7142
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14752 6934 14780 7534
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14740 6656 14792 6662
rect 14844 6644 14872 7482
rect 15304 7342 15332 7704
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 14792 6616 14872 6644
rect 14740 6598 14792 6604
rect 14648 6112 14700 6118
rect 14646 6080 14648 6089
rect 14700 6080 14702 6089
rect 14646 6015 14702 6024
rect 14752 5166 14780 6598
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 15108 5160 15160 5166
rect 15108 5102 15160 5108
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 15028 4593 15056 4966
rect 15120 4622 15148 5102
rect 15108 4616 15160 4622
rect 15014 4584 15070 4593
rect 15108 4558 15160 4564
rect 15014 4519 15070 4528
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14936 3466 14964 4082
rect 15488 3602 15516 11086
rect 15658 9480 15714 9489
rect 15658 9415 15714 9424
rect 15568 7200 15620 7206
rect 15566 7168 15568 7177
rect 15620 7168 15622 7177
rect 15566 7103 15622 7112
rect 15672 6730 15700 9415
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15764 7546 15792 8910
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15856 6458 15884 20198
rect 17222 19952 17278 19961
rect 17222 19887 17278 19896
rect 16302 18864 16358 18873
rect 16028 18828 16080 18834
rect 16302 18799 16304 18808
rect 16028 18770 16080 18776
rect 16356 18799 16358 18808
rect 16304 18770 16356 18776
rect 16040 18086 16068 18770
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16028 17264 16080 17270
rect 16026 17232 16028 17241
rect 16080 17232 16082 17241
rect 16026 17167 16082 17176
rect 16302 13424 16358 13433
rect 16302 13359 16304 13368
rect 16356 13359 16358 13368
rect 16304 13330 16356 13336
rect 16316 12986 16344 13330
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 16764 11620 16816 11626
rect 16764 11562 16816 11568
rect 16408 11082 16620 11098
rect 16408 11076 16632 11082
rect 16408 11070 16580 11076
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16132 10198 16160 10406
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 15934 9888 15990 9897
rect 15934 9823 15990 9832
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15580 4146 15608 4626
rect 15672 4593 15700 5714
rect 15764 5710 15792 6258
rect 15948 6236 15976 9823
rect 16132 9586 16160 10134
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16408 9382 16436 11070
rect 16580 11018 16632 11024
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16040 6882 16068 9318
rect 16684 9178 16712 9522
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16488 8832 16540 8838
rect 16540 8792 16620 8820
rect 16488 8774 16540 8780
rect 16394 8664 16450 8673
rect 16394 8599 16450 8608
rect 16408 8362 16436 8599
rect 16488 8424 16540 8430
rect 16592 8378 16620 8792
rect 16540 8372 16620 8378
rect 16488 8366 16620 8372
rect 16396 8356 16448 8362
rect 16500 8350 16620 8366
rect 16396 8298 16448 8304
rect 16592 8090 16620 8350
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16408 7410 16436 7890
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16118 6896 16174 6905
rect 16040 6854 16118 6882
rect 16118 6831 16174 6840
rect 16212 6860 16264 6866
rect 16132 6798 16160 6831
rect 16212 6802 16264 6808
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16132 6390 16160 6734
rect 16120 6384 16172 6390
rect 16120 6326 16172 6332
rect 16224 6254 16252 6802
rect 16212 6248 16264 6254
rect 15948 6208 16160 6236
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15948 5642 15976 6054
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 15844 5568 15896 5574
rect 15842 5536 15844 5545
rect 15896 5536 15898 5545
rect 15842 5471 15898 5480
rect 15658 4584 15714 4593
rect 15658 4519 15714 4528
rect 15948 4282 15976 5578
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15580 3738 15608 4082
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 14924 3460 14976 3466
rect 14924 3402 14976 3408
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15106 2952 15162 2961
rect 15106 2887 15108 2896
rect 15160 2887 15162 2896
rect 15108 2858 15160 2864
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15304 1714 15332 3334
rect 15488 3194 15516 3538
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15580 2854 15608 3402
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15580 2650 15608 2790
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 15212 1686 15332 1714
rect 15212 480 15240 1686
rect 15672 1601 15700 3878
rect 15948 3738 15976 4014
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15948 3369 15976 3674
rect 15934 3360 15990 3369
rect 15934 3295 15990 3304
rect 15658 1592 15714 1601
rect 15658 1527 15714 1536
rect 16132 610 16160 6208
rect 16210 6216 16212 6225
rect 16264 6216 16266 6225
rect 16210 6151 16266 6160
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16224 3398 16252 4422
rect 16316 3913 16344 7142
rect 16408 7002 16436 7346
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16408 4826 16436 5646
rect 16580 5568 16632 5574
rect 16500 5528 16580 5556
rect 16500 5166 16528 5528
rect 16580 5510 16632 5516
rect 16684 5302 16712 5646
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16500 4146 16528 4966
rect 16684 4486 16712 5238
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16302 3904 16358 3913
rect 16302 3839 16358 3848
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16224 2990 16252 3334
rect 16592 2990 16620 3538
rect 16776 2990 16804 11562
rect 17052 11286 17080 12174
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 17052 10810 17080 11222
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17130 9752 17186 9761
rect 17130 9687 17186 9696
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16868 8634 16896 8978
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16868 8090 16896 8570
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16868 6798 16896 8026
rect 17052 7750 17080 8774
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16868 6458 16896 6734
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 17052 5137 17080 6054
rect 17038 5128 17094 5137
rect 17038 5063 17094 5072
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16224 2582 16252 2926
rect 16580 2848 16632 2854
rect 16500 2796 16580 2802
rect 16500 2790 16632 2796
rect 16500 2774 16620 2790
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 15844 604 15896 610
rect 15844 546 15896 552
rect 16120 604 16172 610
rect 16120 546 16172 552
rect 15856 480 15884 546
rect 16500 480 16528 2774
rect 16854 2680 16910 2689
rect 16854 2615 16856 2624
rect 16908 2615 16910 2624
rect 16856 2586 16908 2592
rect 17144 480 17172 9687
rect 17236 6730 17264 19887
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 17776 13184 17828 13190
rect 18156 13161 18184 13262
rect 17776 13126 17828 13132
rect 18142 13152 18198 13161
rect 17406 13016 17462 13025
rect 17406 12951 17462 12960
rect 17420 12374 17448 12951
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17316 11144 17368 11150
rect 17420 11121 17448 11562
rect 17512 11558 17540 12242
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 11354 17540 11494
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17316 11086 17368 11092
rect 17406 11112 17462 11121
rect 17328 10810 17356 11086
rect 17406 11047 17462 11056
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17328 10266 17356 10746
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17788 8673 17816 13126
rect 18142 13087 18198 13096
rect 18248 11694 18276 22918
rect 18326 16688 18382 16697
rect 18326 16623 18382 16632
rect 18340 16114 18368 16623
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18420 12912 18472 12918
rect 18418 12880 18420 12889
rect 18472 12880 18474 12889
rect 18418 12815 18474 12824
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18418 11792 18474 11801
rect 18418 11727 18420 11736
rect 18472 11727 18474 11736
rect 18420 11698 18472 11704
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18248 11218 18276 11630
rect 18236 11212 18288 11218
rect 18236 11154 18288 11160
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18156 10538 18184 10950
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9654 18000 9998
rect 18156 9926 18184 10474
rect 18432 10470 18460 11154
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18432 10266 18460 10406
rect 18616 10266 18644 12582
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 18156 9518 18184 9862
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18340 9382 18368 10066
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 17774 8664 17830 8673
rect 17774 8599 17830 8608
rect 17868 8560 17920 8566
rect 17314 8528 17370 8537
rect 17868 8502 17920 8508
rect 17314 8463 17370 8472
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17236 5370 17264 5782
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17236 4282 17264 5306
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17328 2854 17356 8463
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17696 7206 17724 7822
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17604 6934 17632 7142
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17406 6760 17462 6769
rect 17406 6695 17462 6704
rect 17420 4690 17448 6695
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17512 5409 17540 6054
rect 17498 5400 17554 5409
rect 17498 5335 17554 5344
rect 17604 4826 17632 6870
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17420 4146 17448 4626
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17604 1737 17632 3878
rect 17696 2922 17724 7142
rect 17880 6866 17908 8502
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17788 6118 17816 6734
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17788 5574 17816 6054
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 3754 17816 4966
rect 17868 4752 17920 4758
rect 17972 4740 18000 7686
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 6662 18092 7278
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18064 5030 18092 6598
rect 18340 5914 18368 9318
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18432 7954 18460 8230
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18432 7274 18460 7890
rect 18420 7268 18472 7274
rect 18420 7210 18472 7216
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18524 5370 18552 8434
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18616 8022 18644 8230
rect 18604 8016 18656 8022
rect 18604 7958 18656 7964
rect 18616 7206 18644 7958
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18512 5364 18564 5370
rect 18512 5306 18564 5312
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 17920 4712 18092 4740
rect 17868 4694 17920 4700
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17880 4010 17908 4422
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17972 3942 18000 4558
rect 18064 4146 18092 4712
rect 18432 4321 18460 4966
rect 18524 4622 18552 5306
rect 18616 5098 18644 7142
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18418 4312 18474 4321
rect 18418 4247 18474 4256
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18156 3942 18184 4014
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 17788 3726 18092 3754
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17774 3088 17830 3097
rect 17774 3023 17776 3032
rect 17828 3023 17830 3032
rect 17776 2994 17828 3000
rect 17880 2961 17908 3334
rect 18064 2990 18092 3726
rect 18432 3641 18460 3878
rect 18418 3632 18474 3641
rect 18418 3567 18474 3576
rect 18616 3398 18644 4082
rect 18708 4078 18736 15846
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18800 12782 18828 13262
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18984 12442 19012 12786
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19352 12458 19380 12650
rect 19260 12442 19380 12458
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 19248 12436 19380 12442
rect 19300 12430 19380 12436
rect 19248 12378 19300 12384
rect 18984 11626 19012 12378
rect 19260 12347 19288 12378
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19352 12073 19380 12242
rect 19338 12064 19394 12073
rect 19338 11999 19394 12008
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 19352 11558 19380 11999
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18800 9178 18828 9386
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 19076 8401 19104 9998
rect 19154 8800 19210 8809
rect 19154 8735 19210 8744
rect 19168 8634 19196 8735
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19062 8392 19118 8401
rect 19062 8327 19118 8336
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19154 7304 19210 7313
rect 19260 7274 19288 8026
rect 19352 7857 19380 11494
rect 19444 8090 19472 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19982 22128 20038 22137
rect 19982 22063 20038 22072
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19996 16153 20024 22063
rect 23480 20256 23532 20262
rect 21454 20224 21510 20233
rect 23480 20198 23532 20204
rect 21454 20159 21510 20168
rect 21468 19990 21496 20159
rect 21456 19984 21508 19990
rect 23492 19961 23520 20198
rect 21456 19926 21508 19932
rect 23478 19952 23534 19961
rect 20904 19916 20956 19922
rect 23478 19887 23534 19896
rect 20904 19858 20956 19864
rect 20916 19174 20944 19858
rect 20904 19168 20956 19174
rect 23480 19168 23532 19174
rect 20904 19110 20956 19116
rect 21362 19136 21418 19145
rect 19982 16144 20038 16153
rect 19982 16079 20038 16088
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19536 11801 19564 12786
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19708 12232 19760 12238
rect 19706 12200 19708 12209
rect 19760 12200 19762 12209
rect 19706 12135 19762 12144
rect 19720 11898 19748 12135
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19522 11792 19578 11801
rect 19522 11727 19578 11736
rect 19996 11665 20024 12582
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20272 11694 20300 12038
rect 20260 11688 20312 11694
rect 19982 11656 20038 11665
rect 19524 11620 19576 11626
rect 20260 11630 20312 11636
rect 19982 11591 20038 11600
rect 19524 11562 19576 11568
rect 19536 11354 19564 11562
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 20074 11384 20130 11393
rect 19524 11348 19576 11354
rect 20074 11319 20130 11328
rect 19524 11290 19576 11296
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19890 10024 19946 10033
rect 19890 9959 19946 9968
rect 19904 9654 19932 9959
rect 20088 9897 20116 11319
rect 20272 11218 20300 11630
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20272 10810 20300 11154
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 20272 10266 20300 10746
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20074 9888 20130 9897
rect 20074 9823 20130 9832
rect 20272 9722 20300 10202
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 19892 9648 19944 9654
rect 19892 9590 19944 9596
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19904 9466 19932 9590
rect 19536 8906 19564 9454
rect 19904 9438 20024 9466
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19536 8294 19564 8842
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19812 8673 19840 8774
rect 19798 8664 19854 8673
rect 19798 8599 19800 8608
rect 19852 8599 19854 8608
rect 19800 8570 19852 8576
rect 19812 8430 19840 8570
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19996 8362 20024 9438
rect 20074 8392 20130 8401
rect 19984 8356 20036 8362
rect 20074 8327 20130 8336
rect 19984 8298 20036 8304
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19338 7848 19394 7857
rect 19338 7783 19394 7792
rect 19432 7744 19484 7750
rect 19536 7732 19564 8230
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19982 7984 20038 7993
rect 19982 7919 20038 7928
rect 19616 7812 19668 7818
rect 19616 7754 19668 7760
rect 19484 7704 19564 7732
rect 19432 7686 19484 7692
rect 19444 7342 19472 7686
rect 19628 7585 19656 7754
rect 19614 7576 19670 7585
rect 19614 7511 19670 7520
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19154 7239 19210 7248
rect 19248 7268 19300 7274
rect 18878 6760 18934 6769
rect 18878 6695 18934 6704
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18800 6322 18828 6598
rect 18892 6458 18920 6695
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18892 6254 18920 6394
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18984 4185 19012 6054
rect 19076 5914 19104 6326
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 19168 5370 19196 7239
rect 19248 7210 19300 7216
rect 19260 7002 19288 7210
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19260 5914 19288 6938
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19156 5024 19208 5030
rect 19154 4992 19156 5001
rect 19208 4992 19210 5001
rect 19154 4927 19210 4936
rect 19260 4826 19288 5850
rect 19352 5370 19380 6258
rect 19444 5914 19472 7142
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19616 6928 19668 6934
rect 19614 6896 19616 6905
rect 19668 6896 19670 6905
rect 19614 6831 19670 6840
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19536 6118 19564 6734
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19536 5817 19564 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19522 5808 19578 5817
rect 19432 5772 19484 5778
rect 19522 5743 19578 5752
rect 19432 5714 19484 5720
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19444 5001 19472 5714
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 19904 5234 19932 5646
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19430 4992 19486 5001
rect 19430 4927 19486 4936
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19996 4690 20024 7919
rect 20088 6066 20116 8327
rect 20352 7880 20404 7886
rect 20456 7857 20484 13670
rect 20916 13530 20944 19110
rect 21362 19071 21418 19080
rect 23478 19136 23480 19145
rect 23532 19136 23534 19145
rect 23478 19071 23534 19080
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21284 13530 21312 14350
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 21178 13152 21234 13161
rect 20548 12850 20576 13126
rect 21178 13087 21234 13096
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20548 12458 20576 12786
rect 20548 12442 20760 12458
rect 20548 12436 20772 12442
rect 20548 12430 20720 12436
rect 20720 12378 20772 12384
rect 20732 12347 20760 12378
rect 20812 12164 20864 12170
rect 20812 12106 20864 12112
rect 20824 11898 20852 12106
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20732 11257 20760 11494
rect 20718 11248 20774 11257
rect 20718 11183 20774 11192
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20732 9489 20760 9862
rect 21008 9761 21036 10406
rect 21192 10266 21220 13087
rect 21284 12986 21312 13466
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21284 10713 21312 12582
rect 21270 10704 21326 10713
rect 21270 10639 21326 10648
rect 21180 10260 21232 10266
rect 21180 10202 21232 10208
rect 20994 9752 21050 9761
rect 21192 9722 21220 10202
rect 21376 10198 21404 19071
rect 23480 15564 23532 15570
rect 23480 15506 23532 15512
rect 23492 14958 23520 15506
rect 23480 14952 23532 14958
rect 23478 14920 23480 14929
rect 23532 14920 23534 14929
rect 23478 14855 23534 14864
rect 23386 14784 23442 14793
rect 23386 14719 23442 14728
rect 23400 14550 23428 14719
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 23112 14476 23164 14482
rect 23112 14418 23164 14424
rect 23124 13870 23152 14418
rect 23478 13968 23534 13977
rect 23478 13903 23534 13912
rect 21824 13864 21876 13870
rect 23112 13864 23164 13870
rect 21824 13806 21876 13812
rect 22374 13832 22430 13841
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21560 12646 21588 13330
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21652 12714 21680 13262
rect 21640 12708 21692 12714
rect 21640 12650 21692 12656
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21652 12458 21680 12650
rect 21643 12430 21680 12458
rect 21546 12336 21602 12345
rect 21643 12322 21671 12430
rect 21643 12294 21680 12322
rect 21546 12271 21602 12280
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 21364 10192 21416 10198
rect 21364 10134 21416 10140
rect 20994 9687 21050 9696
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 20996 9648 21048 9654
rect 21468 9636 21496 11154
rect 21560 10810 21588 12271
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21548 10056 21600 10062
rect 21652 10044 21680 12294
rect 21744 10198 21772 13670
rect 21836 10810 21864 13806
rect 23112 13806 23164 13812
rect 22374 13767 22430 13776
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 21928 11218 21956 12378
rect 22296 11694 22324 13670
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 21824 10804 21876 10810
rect 21824 10746 21876 10752
rect 21928 10674 21956 11154
rect 22020 10690 22048 11222
rect 21916 10668 21968 10674
rect 22020 10662 22140 10690
rect 21916 10610 21968 10616
rect 22112 10606 22140 10662
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 21732 10192 21784 10198
rect 21732 10134 21784 10140
rect 21652 10016 21772 10044
rect 21548 9998 21600 10004
rect 20996 9590 21048 9596
rect 21284 9608 21496 9636
rect 20718 9480 20774 9489
rect 20718 9415 20774 9424
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20352 7822 20404 7828
rect 20442 7848 20498 7857
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 20180 7002 20208 7686
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 20272 6322 20300 7142
rect 20364 6662 20392 7822
rect 20442 7783 20498 7792
rect 20640 7721 20668 8910
rect 20916 7818 20944 9318
rect 21008 9042 21036 9590
rect 21284 9382 21312 9608
rect 21456 9512 21508 9518
rect 21456 9454 21508 9460
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 20996 9036 21048 9042
rect 20996 8978 21048 8984
rect 21284 8634 21312 9046
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21468 8566 21496 9454
rect 21560 9178 21588 9998
rect 21744 9874 21772 10016
rect 22112 9994 22140 10406
rect 22100 9988 22152 9994
rect 22100 9930 22152 9936
rect 21652 9846 21772 9874
rect 21916 9920 21968 9926
rect 22112 9874 22140 9930
rect 21916 9862 21968 9868
rect 21652 9602 21680 9846
rect 21652 9574 21864 9602
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21456 8560 21508 8566
rect 21456 8502 21508 8508
rect 21362 8120 21418 8129
rect 21362 8055 21418 8064
rect 21178 7848 21234 7857
rect 20904 7812 20956 7818
rect 21178 7783 21234 7792
rect 20904 7754 20956 7760
rect 20720 7744 20772 7750
rect 20626 7712 20682 7721
rect 20720 7686 20772 7692
rect 20626 7647 20682 7656
rect 20732 7342 20760 7686
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 20444 6928 20496 6934
rect 20444 6870 20496 6876
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20364 6089 20392 6598
rect 20456 6118 20484 6870
rect 20548 6458 20576 7210
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20444 6112 20496 6118
rect 20350 6080 20406 6089
rect 20088 6038 20300 6066
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 20180 5098 20208 5714
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 20168 5092 20220 5098
rect 20168 5034 20220 5040
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 18970 4176 19026 4185
rect 18970 4111 19026 4120
rect 18696 4072 18748 4078
rect 19444 4049 19472 4558
rect 19536 4282 19564 4626
rect 20088 4622 20116 5034
rect 20076 4616 20128 4622
rect 20272 4570 20300 6038
rect 20444 6054 20496 6060
rect 20350 6015 20406 6024
rect 20350 5944 20406 5953
rect 20548 5914 20576 6258
rect 20640 6254 20668 6598
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20732 5914 20760 7278
rect 20994 7032 21050 7041
rect 20994 6967 21050 6976
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20824 6322 20852 6802
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20916 6662 20944 6734
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20916 6186 20944 6598
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20902 5944 20958 5953
rect 20350 5879 20352 5888
rect 20404 5879 20406 5888
rect 20536 5908 20588 5914
rect 20352 5850 20404 5856
rect 20536 5850 20588 5856
rect 20720 5908 20772 5914
rect 20902 5879 20958 5888
rect 20720 5850 20772 5856
rect 20548 5794 20576 5850
rect 20548 5778 20760 5794
rect 20548 5772 20772 5778
rect 20548 5766 20720 5772
rect 20720 5714 20772 5720
rect 20732 4826 20760 5714
rect 20916 5166 20944 5879
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 20812 5024 20864 5030
rect 20810 4992 20812 5001
rect 20864 4992 20866 5001
rect 20810 4927 20866 4936
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 21008 4690 21036 6967
rect 21192 5914 21220 7783
rect 21376 7546 21404 8055
rect 21640 8016 21692 8022
rect 21640 7958 21692 7964
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21456 7472 21508 7478
rect 21456 7414 21508 7420
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21284 6254 21312 7346
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 21364 6180 21416 6186
rect 21364 6122 21416 6128
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 21088 5636 21140 5642
rect 21088 5578 21140 5584
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 20076 4558 20128 4564
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19904 4049 19932 4422
rect 18696 4014 18748 4020
rect 19430 4040 19486 4049
rect 19156 4004 19208 4010
rect 19430 3975 19486 3984
rect 19890 4040 19946 4049
rect 19890 3975 19946 3984
rect 19156 3946 19208 3952
rect 19168 3913 19196 3946
rect 19524 3936 19576 3942
rect 19154 3904 19210 3913
rect 19524 3878 19576 3884
rect 19154 3839 19210 3848
rect 19430 3768 19486 3777
rect 19430 3703 19486 3712
rect 19154 3496 19210 3505
rect 19154 3431 19156 3440
rect 19208 3431 19210 3440
rect 19156 3402 19208 3408
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18418 3088 18474 3097
rect 18418 3023 18474 3032
rect 18052 2984 18104 2990
rect 17866 2952 17922 2961
rect 17684 2916 17736 2922
rect 18142 2952 18198 2961
rect 18104 2932 18142 2938
rect 18052 2926 18142 2932
rect 18064 2910 18142 2926
rect 17866 2887 17922 2896
rect 18142 2887 18198 2896
rect 17684 2858 17736 2864
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17590 1728 17646 1737
rect 17590 1663 17646 1672
rect 17788 480 17816 2790
rect 18156 2446 18184 2887
rect 18052 2440 18104 2446
rect 18050 2408 18052 2417
rect 18144 2440 18196 2446
rect 18104 2408 18106 2417
rect 18144 2382 18196 2388
rect 18050 2343 18106 2352
rect 18432 480 18460 3023
rect 19444 2582 19472 3703
rect 19536 3670 19564 3878
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19524 3664 19576 3670
rect 19524 3606 19576 3612
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19812 3194 19840 3470
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19536 2514 19564 3130
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19524 2508 19576 2514
rect 19524 2450 19576 2456
rect 19996 2258 20024 4490
rect 20088 3913 20116 4558
rect 20180 4542 20300 4570
rect 20180 4078 20208 4542
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20272 4146 20300 4422
rect 21008 4282 21036 4626
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20074 3904 20130 3913
rect 20074 3839 20130 3848
rect 20180 3738 20208 4014
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20180 3505 20208 3674
rect 20166 3496 20222 3505
rect 20166 3431 20222 3440
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 20088 2650 20116 2926
rect 20272 2922 20300 4082
rect 21100 3738 21128 5578
rect 21192 5370 21220 5850
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20536 2984 20588 2990
rect 20534 2952 20536 2961
rect 20588 2952 20590 2961
rect 20260 2916 20312 2922
rect 20534 2887 20590 2896
rect 20260 2858 20312 2864
rect 20640 2650 20668 3538
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 19812 2230 20024 2258
rect 19154 1456 19210 1465
rect 19154 1391 19210 1400
rect 19168 480 19196 1391
rect 19812 480 19840 2230
rect 20442 2000 20498 2009
rect 20442 1935 20498 1944
rect 20456 480 20484 1935
rect 21100 480 21128 3334
rect 21376 2961 21404 6122
rect 21468 4758 21496 7414
rect 21456 4752 21508 4758
rect 21456 4694 21508 4700
rect 21548 4684 21600 4690
rect 21548 4626 21600 4632
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21468 3369 21496 3878
rect 21560 3602 21588 4626
rect 21652 3942 21680 7958
rect 21744 7886 21772 9454
rect 21836 9110 21864 9574
rect 21928 9382 21956 9862
rect 22020 9846 22140 9874
rect 21916 9376 21968 9382
rect 21916 9318 21968 9324
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21744 7478 21772 7822
rect 21928 7585 21956 9318
rect 22020 8090 22048 9846
rect 22190 9480 22246 9489
rect 22190 9415 22246 9424
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 21914 7576 21970 7585
rect 21914 7511 21970 7520
rect 21732 7472 21784 7478
rect 21732 7414 21784 7420
rect 22112 7274 22140 7686
rect 22204 7449 22232 9415
rect 22388 9217 22416 13767
rect 23492 13546 23520 13903
rect 23400 13530 23520 13546
rect 23584 13530 23612 26551
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 23952 23254 23980 23598
rect 23940 23248 23992 23254
rect 23940 23190 23992 23196
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23860 22438 23888 23122
rect 24044 22642 24072 27639
rect 24490 27520 24546 28000
rect 24122 27160 24178 27169
rect 24122 27095 24178 27104
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 23848 22432 23900 22438
rect 23848 22374 23900 22380
rect 23860 22137 23888 22374
rect 23846 22128 23902 22137
rect 23846 22063 23902 22072
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 24030 21448 24086 21457
rect 23952 20466 23980 21422
rect 24030 21383 24086 21392
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 23754 20360 23810 20369
rect 23754 20295 23810 20304
rect 23662 19136 23718 19145
rect 23662 19071 23718 19080
rect 23676 17241 23704 19071
rect 23768 18737 23796 20295
rect 24044 20058 24072 21383
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 24032 19916 24084 19922
rect 24032 19858 24084 19864
rect 24044 18873 24072 19858
rect 24030 18864 24086 18873
rect 24030 18799 24086 18808
rect 23754 18728 23810 18737
rect 23754 18663 23810 18672
rect 24030 18048 24086 18057
rect 24030 17983 24086 17992
rect 23662 17232 23718 17241
rect 23662 17167 23718 17176
rect 24044 16794 24072 17983
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 23938 15056 23994 15065
rect 23938 14991 23994 15000
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23388 13524 23520 13530
rect 23440 13518 23520 13524
rect 23572 13524 23624 13530
rect 23388 13466 23440 13472
rect 23572 13466 23624 13472
rect 22928 13388 22980 13394
rect 22928 13330 22980 13336
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22664 12102 22692 13126
rect 22940 12646 22968 13330
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23216 12986 23244 13262
rect 23400 12986 23428 13466
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22480 11762 22508 12038
rect 22756 11778 22784 12582
rect 22940 12073 22968 12582
rect 23216 12102 23244 12922
rect 23204 12096 23256 12102
rect 22926 12064 22982 12073
rect 23204 12038 23256 12044
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 22926 11999 22982 12008
rect 22940 11898 22968 11999
rect 22928 11892 22980 11898
rect 22928 11834 22980 11840
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22572 11750 22784 11778
rect 23202 11792 23258 11801
rect 23112 11756 23164 11762
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22480 10266 22508 10610
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22374 9208 22430 9217
rect 22374 9143 22430 9152
rect 22284 8832 22336 8838
rect 22282 8800 22284 8809
rect 22336 8800 22338 8809
rect 22282 8735 22338 8744
rect 22388 7886 22416 9143
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22388 7546 22416 7822
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22190 7440 22246 7449
rect 22190 7375 22246 7384
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22284 6656 22336 6662
rect 22284 6598 22336 6604
rect 22296 6254 22324 6598
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22008 5704 22060 5710
rect 22008 5646 22060 5652
rect 21916 5636 21968 5642
rect 21916 5578 21968 5584
rect 21732 5296 21784 5302
rect 21732 5238 21784 5244
rect 21822 5264 21878 5273
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 21548 3596 21600 3602
rect 21548 3538 21600 3544
rect 21454 3360 21510 3369
rect 21454 3295 21510 3304
rect 21362 2952 21418 2961
rect 21362 2887 21418 2896
rect 21468 2825 21496 3295
rect 21454 2816 21510 2825
rect 21454 2751 21510 2760
rect 21638 2816 21694 2825
rect 21638 2751 21694 2760
rect 21652 2650 21680 2751
rect 21640 2644 21692 2650
rect 21640 2586 21692 2592
rect 21548 2508 21600 2514
rect 21548 2450 21600 2456
rect 21560 1601 21588 2450
rect 21546 1592 21602 1601
rect 21546 1527 21602 1536
rect 21744 480 21772 5238
rect 21822 5199 21878 5208
rect 21836 5166 21864 5199
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 21928 3398 21956 5578
rect 22020 5370 22048 5646
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 22112 5302 22140 5510
rect 22100 5296 22152 5302
rect 22100 5238 22152 5244
rect 22008 4480 22060 4486
rect 22008 4422 22060 4428
rect 22020 3942 22048 4422
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 22006 2952 22062 2961
rect 21824 2916 21876 2922
rect 22006 2887 22062 2896
rect 21824 2858 21876 2864
rect 21836 2446 21864 2858
rect 22020 2582 22048 2887
rect 22008 2576 22060 2582
rect 22008 2518 22060 2524
rect 22112 2514 22140 3878
rect 22204 3670 22232 6054
rect 22388 4162 22416 6054
rect 22480 4826 22508 10202
rect 22572 8090 22600 11750
rect 23202 11727 23258 11736
rect 23112 11698 23164 11704
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22756 11354 22784 11562
rect 23124 11558 23152 11698
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 23124 11286 23152 11494
rect 23112 11280 23164 11286
rect 23112 11222 23164 11228
rect 22926 11112 22982 11121
rect 22926 11047 22982 11056
rect 22940 10266 22968 11047
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 23020 10192 23072 10198
rect 23020 10134 23072 10140
rect 23032 9722 23060 10134
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23216 8634 23244 11727
rect 23492 11626 23520 12038
rect 23480 11620 23532 11626
rect 23480 11562 23532 11568
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23492 10810 23520 11222
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23584 10282 23612 12038
rect 23400 10266 23612 10282
rect 23388 10260 23612 10266
rect 23440 10254 23612 10260
rect 23388 10202 23440 10208
rect 23400 9178 23428 10202
rect 23570 10160 23626 10169
rect 23570 10095 23626 10104
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23492 9722 23520 9998
rect 23480 9716 23532 9722
rect 23480 9658 23532 9664
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23492 8974 23520 9454
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 22652 8560 22704 8566
rect 22650 8528 22652 8537
rect 23480 8560 23532 8566
rect 22704 8528 22706 8537
rect 23480 8502 23532 8508
rect 22650 8463 22706 8472
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 23388 8084 23440 8090
rect 23492 8072 23520 8502
rect 23440 8044 23520 8072
rect 23388 8026 23440 8032
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22664 7449 22692 7686
rect 23032 7546 23060 8026
rect 23296 7812 23348 7818
rect 23296 7754 23348 7760
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 22650 7440 22706 7449
rect 22650 7375 22706 7384
rect 22836 6996 22888 7002
rect 22836 6938 22888 6944
rect 22652 6180 22704 6186
rect 22652 6122 22704 6128
rect 22664 5574 22692 6122
rect 22652 5568 22704 5574
rect 22652 5510 22704 5516
rect 22664 5234 22692 5510
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22468 4820 22520 4826
rect 22468 4762 22520 4768
rect 22296 4146 22416 4162
rect 22296 4140 22428 4146
rect 22296 4134 22376 4140
rect 22192 3664 22244 3670
rect 22192 3606 22244 3612
rect 22296 3602 22324 4134
rect 22376 4082 22428 4088
rect 22374 4040 22430 4049
rect 22374 3975 22430 3984
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 22296 3194 22324 3538
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 22282 3088 22338 3097
rect 22282 3023 22338 3032
rect 22296 2650 22324 3023
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 22296 2446 22324 2586
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22388 480 22416 3975
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 22664 1465 22692 2246
rect 22650 1456 22706 1465
rect 22650 1391 22706 1400
rect 22848 1290 22876 6938
rect 22926 6216 22982 6225
rect 22926 6151 22982 6160
rect 22940 5817 22968 6151
rect 22926 5808 22982 5817
rect 22926 5743 22982 5752
rect 23110 5808 23166 5817
rect 23308 5778 23336 7754
rect 23400 7002 23428 8026
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23492 7002 23520 7890
rect 23584 7041 23612 10095
rect 23676 7546 23704 14758
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23860 12889 23888 13126
rect 23846 12880 23902 12889
rect 23846 12815 23902 12824
rect 23860 12782 23888 12815
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23768 11354 23796 12378
rect 23952 12209 23980 14991
rect 24136 14074 24164 27095
rect 24504 25242 24532 27520
rect 24674 26072 24730 26081
rect 24674 26007 24730 26016
rect 24228 25214 24532 25242
rect 24228 24410 24256 25214
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24216 24404 24268 24410
rect 24216 24346 24268 24352
rect 24214 24304 24270 24313
rect 24214 24239 24270 24248
rect 24228 22778 24256 24239
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23866 24716 26007
rect 24766 25392 24822 25401
rect 24766 25327 24822 25336
rect 24780 24886 24808 25327
rect 24768 24880 24820 24886
rect 24768 24822 24820 24828
rect 24766 24712 24822 24721
rect 24766 24647 24822 24656
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 24780 23338 24808 24647
rect 24780 23322 24900 23338
rect 24780 23316 24912 23322
rect 24780 23310 24860 23316
rect 24860 23258 24912 23264
rect 24674 23216 24730 23225
rect 24674 23151 24730 23160
rect 24952 23180 25004 23186
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24216 22772 24268 22778
rect 24216 22714 24268 22720
rect 24582 22672 24638 22681
rect 24216 22636 24268 22642
rect 24582 22607 24638 22616
rect 24216 22578 24268 22584
rect 24228 16454 24256 22578
rect 24596 22574 24624 22607
rect 24584 22568 24636 22574
rect 24584 22510 24636 22516
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21690 24716 23151
rect 24952 23122 25004 23128
rect 24766 22536 24822 22545
rect 24964 22506 24992 23122
rect 24766 22471 24822 22480
rect 24952 22500 25004 22506
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24780 21146 24808 22471
rect 24952 22442 25004 22448
rect 24964 22001 24992 22442
rect 24950 21992 25006 22001
rect 24950 21927 25006 21936
rect 25134 21992 25190 22001
rect 25134 21927 25190 21936
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20482 24716 20946
rect 24766 20904 24822 20913
rect 24766 20839 24822 20848
rect 24596 20454 24716 20482
rect 24596 20262 24624 20454
rect 24584 20256 24636 20262
rect 24582 20224 24584 20233
rect 24636 20224 24638 20233
rect 24582 20159 24638 20168
rect 24674 19680 24730 19689
rect 24289 19612 24585 19632
rect 24674 19615 24730 19624
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24584 19168 24636 19174
rect 24584 19110 24636 19116
rect 24596 18873 24624 19110
rect 24582 18864 24638 18873
rect 24582 18799 24638 18808
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 17882 24716 19615
rect 24780 19258 24808 20839
rect 25148 20602 25176 21927
rect 26238 21040 26294 21049
rect 26238 20975 26294 20984
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 24872 19378 24900 20334
rect 24860 19372 24912 19378
rect 24860 19314 24912 19320
rect 24952 19304 25004 19310
rect 24780 19230 24900 19258
rect 24952 19246 25004 19252
rect 24872 19174 24900 19230
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24766 18592 24822 18601
rect 24766 18527 24822 18536
rect 24676 17876 24728 17882
rect 24676 17818 24728 17824
rect 24674 17504 24730 17513
rect 24289 17436 24585 17456
rect 24674 17439 24730 17448
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17082 24716 17439
rect 24780 17338 24808 18527
rect 24964 18193 24992 19246
rect 24950 18184 25006 18193
rect 24950 18119 25006 18128
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 25148 17134 25176 17682
rect 25136 17128 25188 17134
rect 25134 17096 25136 17105
rect 25188 17096 25190 17105
rect 24688 17054 24808 17082
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24412 16697 24440 16934
rect 24398 16688 24454 16697
rect 24398 16623 24454 16632
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24216 16448 24268 16454
rect 24216 16390 24268 16396
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16182 24716 16594
rect 24780 16250 24808 17054
rect 25134 17031 25190 17040
rect 25042 16824 25098 16833
rect 25042 16759 25098 16768
rect 24952 16448 25004 16454
rect 24952 16390 25004 16396
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24216 16040 24268 16046
rect 24216 15982 24268 15988
rect 24228 15026 24256 15982
rect 24688 15638 24716 16118
rect 24766 15736 24822 15745
rect 24766 15671 24822 15680
rect 24676 15632 24728 15638
rect 24676 15574 24728 15580
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24780 14482 24808 15671
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24872 14822 24900 15506
rect 24860 14816 24912 14822
rect 24858 14784 24860 14793
rect 24912 14784 24914 14793
rect 24858 14719 24914 14728
rect 24768 14476 24820 14482
rect 24768 14418 24820 14424
rect 24780 14362 24808 14418
rect 24780 14334 24900 14362
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 24780 13841 24808 14214
rect 24872 14074 24900 14334
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24766 13832 24822 13841
rect 24766 13767 24822 13776
rect 24124 13728 24176 13734
rect 24124 13670 24176 13676
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 24044 13025 24072 13330
rect 24030 13016 24086 13025
rect 24030 12951 24032 12960
rect 24084 12951 24086 12960
rect 24032 12922 24084 12928
rect 24136 12850 24164 13670
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24306 12880 24362 12889
rect 24124 12844 24176 12850
rect 24306 12815 24362 12824
rect 24124 12786 24176 12792
rect 24320 12442 24348 12815
rect 24308 12436 24360 12442
rect 24308 12378 24360 12384
rect 24032 12300 24084 12306
rect 24032 12242 24084 12248
rect 23938 12200 23994 12209
rect 23938 12135 23994 12144
rect 24044 11914 24072 12242
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 24124 12096 24176 12102
rect 24124 12038 24176 12044
rect 23952 11898 24072 11914
rect 23940 11892 24072 11898
rect 23992 11886 24072 11892
rect 23940 11834 23992 11840
rect 23756 11348 23808 11354
rect 23756 11290 23808 11296
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23860 11234 23888 11290
rect 23768 11206 23888 11234
rect 23768 11150 23796 11206
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23768 10606 23796 11086
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 23860 10538 23888 10950
rect 23848 10532 23900 10538
rect 23848 10474 23900 10480
rect 23952 8430 23980 11834
rect 24136 11778 24164 12038
rect 24044 11750 24164 11778
rect 24044 11626 24072 11750
rect 24032 11620 24084 11626
rect 24032 11562 24084 11568
rect 24044 11354 24072 11562
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 24228 11014 24256 12174
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24872 11393 24900 12038
rect 24858 11384 24914 11393
rect 24858 11319 24914 11328
rect 24674 11112 24730 11121
rect 24674 11047 24730 11056
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24490 10704 24546 10713
rect 24490 10639 24546 10648
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 24044 10266 24072 10406
rect 24504 10266 24532 10639
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 24044 10062 24072 10202
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 24306 10024 24362 10033
rect 24306 9959 24308 9968
rect 24360 9959 24362 9968
rect 24308 9930 24360 9936
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24030 8936 24086 8945
rect 24030 8871 24086 8880
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 23754 7712 23810 7721
rect 23754 7647 23810 7656
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23664 7336 23716 7342
rect 23664 7278 23716 7284
rect 23570 7032 23626 7041
rect 23388 6996 23440 7002
rect 23388 6938 23440 6944
rect 23480 6996 23532 7002
rect 23570 6967 23626 6976
rect 23480 6938 23532 6944
rect 23110 5743 23112 5752
rect 23164 5743 23166 5752
rect 23296 5772 23348 5778
rect 23112 5714 23164 5720
rect 23296 5714 23348 5720
rect 23124 5370 23152 5714
rect 23202 5672 23258 5681
rect 23202 5607 23258 5616
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23112 5092 23164 5098
rect 23112 5034 23164 5040
rect 23124 5001 23152 5034
rect 23110 4992 23166 5001
rect 23110 4927 23166 4936
rect 23020 4752 23072 4758
rect 23020 4694 23072 4700
rect 23032 4282 23060 4694
rect 23110 4312 23166 4321
rect 23020 4276 23072 4282
rect 23110 4247 23166 4256
rect 23020 4218 23072 4224
rect 23032 3738 23060 4218
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 22836 1284 22888 1290
rect 22836 1226 22888 1232
rect 23124 626 23152 4247
rect 23216 3670 23244 5607
rect 23492 5522 23520 6938
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23584 6322 23612 6734
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 23584 5642 23612 6258
rect 23676 5914 23704 7278
rect 23768 5914 23796 7647
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 23860 6934 23888 7482
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 23860 6458 23888 6870
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23664 5772 23716 5778
rect 23664 5714 23716 5720
rect 23572 5636 23624 5642
rect 23572 5578 23624 5584
rect 23676 5522 23704 5714
rect 23400 5494 23520 5522
rect 23584 5494 23704 5522
rect 23400 5284 23428 5494
rect 23400 5256 23520 5284
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 23400 5001 23428 5102
rect 23386 4992 23442 5001
rect 23386 4927 23442 4936
rect 23388 4208 23440 4214
rect 23388 4150 23440 4156
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 23204 3664 23256 3670
rect 23204 3606 23256 3612
rect 23308 2650 23336 4014
rect 23400 2650 23428 4150
rect 23492 3738 23520 5256
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23584 3074 23612 5494
rect 23664 5364 23716 5370
rect 23768 5352 23796 5850
rect 23860 5846 23888 6394
rect 23848 5840 23900 5846
rect 24044 5817 24072 8871
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24124 8492 24176 8498
rect 24124 8434 24176 8440
rect 24136 8090 24164 8434
rect 24216 8288 24268 8294
rect 24214 8256 24216 8265
rect 24268 8256 24270 8265
rect 24214 8191 24270 8200
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 24228 8022 24256 8191
rect 24216 8016 24268 8022
rect 24216 7958 24268 7964
rect 24216 7880 24268 7886
rect 24216 7822 24268 7828
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24136 7410 24164 7686
rect 24228 7546 24256 7822
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24228 7002 24256 7346
rect 24216 6996 24268 7002
rect 24216 6938 24268 6944
rect 24122 6216 24178 6225
rect 24122 6151 24178 6160
rect 23848 5782 23900 5788
rect 24030 5808 24086 5817
rect 24030 5743 24086 5752
rect 23716 5324 23796 5352
rect 23664 5306 23716 5312
rect 23664 5160 23716 5166
rect 23664 5102 23716 5108
rect 23676 4690 23704 5102
rect 23940 5092 23992 5098
rect 23940 5034 23992 5040
rect 23952 4826 23980 5034
rect 23940 4820 23992 4826
rect 23940 4762 23992 4768
rect 23664 4684 23716 4690
rect 23664 4626 23716 4632
rect 23676 4486 23704 4626
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 24030 4176 24086 4185
rect 24030 4111 24086 4120
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23952 3670 23980 4014
rect 23848 3664 23900 3670
rect 23662 3632 23718 3641
rect 23848 3606 23900 3612
rect 23940 3664 23992 3670
rect 23940 3606 23992 3612
rect 23662 3567 23718 3576
rect 23676 3194 23704 3567
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23584 3046 23704 3074
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23480 2916 23532 2922
rect 23480 2858 23532 2864
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 23492 1873 23520 2858
rect 23584 2514 23612 2926
rect 23676 2564 23704 3046
rect 23860 2990 23888 3606
rect 23940 3460 23992 3466
rect 23940 3402 23992 3408
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 23846 2816 23902 2825
rect 23846 2751 23902 2760
rect 23676 2536 23796 2564
rect 23572 2508 23624 2514
rect 23572 2450 23624 2456
rect 23768 2378 23796 2536
rect 23756 2372 23808 2378
rect 23756 2314 23808 2320
rect 23478 1864 23534 1873
rect 23478 1799 23534 1808
rect 23664 1420 23716 1426
rect 23664 1362 23716 1368
rect 23032 598 23152 626
rect 23032 480 23060 598
rect 23676 480 23704 1362
rect 294 0 350 480
rect 938 0 994 480
rect 1582 0 1638 480
rect 2226 0 2282 480
rect 2870 0 2926 480
rect 3514 0 3570 480
rect 4158 0 4214 480
rect 4802 0 4858 480
rect 5446 0 5502 480
rect 6090 0 6146 480
rect 6734 0 6790 480
rect 7378 0 7434 480
rect 8022 0 8078 480
rect 8666 0 8722 480
rect 9310 0 9366 480
rect 10046 0 10102 480
rect 10690 0 10746 480
rect 11334 0 11390 480
rect 11978 0 12034 480
rect 12622 0 12678 480
rect 13266 0 13322 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15198 0 15254 480
rect 15842 0 15898 480
rect 16486 0 16542 480
rect 17130 0 17186 480
rect 17774 0 17830 480
rect 18418 0 18474 480
rect 19154 0 19210 480
rect 19798 0 19854 480
rect 20442 0 20498 480
rect 21086 0 21142 480
rect 21730 0 21786 480
rect 22374 0 22430 480
rect 23018 0 23074 480
rect 23662 0 23718 480
rect 23860 377 23888 2751
rect 23952 2582 23980 3402
rect 23940 2576 23992 2582
rect 23940 2518 23992 2524
rect 24044 1426 24072 4111
rect 24136 3738 24164 6151
rect 24228 4826 24256 6938
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24584 6180 24636 6186
rect 24584 6122 24636 6128
rect 24596 5658 24624 6122
rect 24688 5778 24716 11047
rect 24766 10568 24822 10577
rect 24766 10503 24822 10512
rect 24780 8106 24808 10503
rect 24860 10124 24912 10130
rect 24860 10066 24912 10072
rect 24872 9722 24900 10066
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24872 9625 24900 9658
rect 24858 9616 24914 9625
rect 24858 9551 24914 9560
rect 24858 9208 24914 9217
rect 24858 9143 24860 9152
rect 24912 9143 24914 9152
rect 24860 9114 24912 9120
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 24872 8294 24900 8774
rect 24860 8288 24912 8294
rect 24860 8230 24912 8236
rect 24780 8078 24900 8106
rect 24768 8016 24820 8022
rect 24768 7958 24820 7964
rect 24780 7206 24808 7958
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24596 5630 24716 5658
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5098 24716 5630
rect 24676 5092 24728 5098
rect 24676 5034 24728 5040
rect 24674 4992 24730 5001
rect 24674 4927 24730 4936
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24228 4078 24256 4762
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4321 24716 4927
rect 24780 4826 24808 7142
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24872 4706 24900 8078
rect 24964 5250 24992 16390
rect 25056 15706 25084 16759
rect 25502 16280 25558 16289
rect 25502 16215 25558 16224
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 25516 15162 25544 16215
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25412 14952 25464 14958
rect 25412 14894 25464 14900
rect 25318 12744 25374 12753
rect 25318 12679 25374 12688
rect 25332 12646 25360 12679
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 25056 11286 25084 11494
rect 25044 11280 25096 11286
rect 25044 11222 25096 11228
rect 25320 10464 25372 10470
rect 25320 10406 25372 10412
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 25056 9042 25084 9318
rect 25044 9036 25096 9042
rect 25044 8978 25096 8984
rect 25056 8634 25084 8978
rect 25332 8838 25360 10406
rect 25320 8832 25372 8838
rect 25320 8774 25372 8780
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 25424 8498 25452 14894
rect 25778 14648 25834 14657
rect 25778 14583 25834 14592
rect 25686 13424 25742 13433
rect 25686 13359 25742 13368
rect 25700 12306 25728 13359
rect 25792 12986 25820 14583
rect 25780 12980 25832 12986
rect 25780 12922 25832 12928
rect 25792 12782 25820 12922
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 25688 12300 25740 12306
rect 25688 12242 25740 12248
rect 25700 11898 25728 12242
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 25780 10124 25832 10130
rect 25780 10066 25832 10072
rect 25792 9722 25820 10066
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25228 8424 25280 8430
rect 25228 8366 25280 8372
rect 25240 8129 25268 8366
rect 25688 8288 25740 8294
rect 25688 8230 25740 8236
rect 25226 8120 25282 8129
rect 25226 8055 25282 8064
rect 25226 7440 25282 7449
rect 25226 7375 25282 7384
rect 25240 7342 25268 7375
rect 25228 7336 25280 7342
rect 25228 7278 25280 7284
rect 25504 7268 25556 7274
rect 25504 7210 25556 7216
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 25056 5642 25084 6054
rect 25516 5953 25544 7210
rect 25502 5944 25558 5953
rect 25502 5879 25558 5888
rect 25596 5772 25648 5778
rect 25596 5714 25648 5720
rect 25044 5636 25096 5642
rect 25044 5578 25096 5584
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 25502 5536 25558 5545
rect 24964 5222 25268 5250
rect 25056 5166 25084 5222
rect 25044 5160 25096 5166
rect 24950 5128 25006 5137
rect 25044 5102 25096 5108
rect 24950 5063 25006 5072
rect 24780 4678 24900 4706
rect 24674 4312 24730 4321
rect 24674 4247 24730 4256
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 24780 3890 24808 4678
rect 24596 3862 24808 3890
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24214 3496 24270 3505
rect 24596 3466 24624 3862
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 24768 3732 24820 3738
rect 24768 3674 24820 3680
rect 24214 3431 24270 3440
rect 24584 3460 24636 3466
rect 24228 2650 24256 3431
rect 24584 3402 24636 3408
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3194 24716 3674
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 2009 24716 3130
rect 24674 2000 24730 2009
rect 24674 1935 24730 1944
rect 24032 1420 24084 1426
rect 24032 1362 24084 1368
rect 24308 1284 24360 1290
rect 24308 1226 24360 1232
rect 24320 480 24348 1226
rect 24780 921 24808 3674
rect 24858 2544 24914 2553
rect 24858 2479 24860 2488
rect 24912 2479 24914 2488
rect 24860 2450 24912 2456
rect 24766 912 24822 921
rect 24766 847 24822 856
rect 24964 480 24992 5063
rect 25136 5024 25188 5030
rect 25136 4966 25188 4972
rect 25044 4752 25096 4758
rect 25044 4694 25096 4700
rect 25056 3913 25084 4694
rect 25148 4622 25176 4966
rect 25240 4826 25268 5222
rect 25228 4820 25280 4826
rect 25228 4762 25280 4768
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 25042 3904 25098 3913
rect 25042 3839 25098 3848
rect 25056 3738 25084 3839
rect 25044 3732 25096 3738
rect 25044 3674 25096 3680
rect 25044 3596 25096 3602
rect 25044 3538 25096 3544
rect 25056 3210 25084 3538
rect 25148 3534 25176 4558
rect 25240 4282 25268 4762
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 25136 3528 25188 3534
rect 25136 3470 25188 3476
rect 25134 3224 25190 3233
rect 25056 3182 25134 3210
rect 25134 3159 25136 3168
rect 25188 3159 25190 3168
rect 25136 3130 25188 3136
rect 25332 3097 25360 3878
rect 25318 3088 25374 3097
rect 25318 3023 25374 3032
rect 25424 2961 25452 5510
rect 25502 5471 25558 5480
rect 25410 2952 25466 2961
rect 25410 2887 25466 2896
rect 25412 2848 25464 2854
rect 25410 2816 25412 2825
rect 25464 2816 25466 2825
rect 25410 2751 25466 2760
rect 25044 2576 25096 2582
rect 25042 2544 25044 2553
rect 25096 2544 25098 2553
rect 25042 2479 25098 2488
rect 25516 626 25544 5471
rect 25608 5370 25636 5714
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 25596 5024 25648 5030
rect 25700 5012 25728 8230
rect 25648 4984 25728 5012
rect 25596 4966 25648 4972
rect 25608 4486 25636 4966
rect 25596 4480 25648 4486
rect 25596 4422 25648 4428
rect 25608 3738 25636 4422
rect 25792 3777 25820 9658
rect 26252 7546 26280 20975
rect 26330 13832 26386 13841
rect 26330 13767 26386 13776
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26240 3936 26292 3942
rect 26240 3878 26292 3884
rect 25778 3768 25834 3777
rect 25596 3732 25648 3738
rect 25778 3703 25834 3712
rect 25596 3674 25648 3680
rect 25792 2802 25820 3703
rect 26148 3664 26200 3670
rect 26148 3606 26200 3612
rect 26160 3194 26188 3606
rect 26252 3534 26280 3878
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 26148 3188 26200 3194
rect 26148 3130 26200 3136
rect 26252 3126 26280 3470
rect 26240 3120 26292 3126
rect 26240 3062 26292 3068
rect 26344 2972 26372 13767
rect 26884 7540 26936 7546
rect 26884 7482 26936 7488
rect 26252 2944 26372 2972
rect 25792 2774 25912 2802
rect 25884 2650 25912 2774
rect 25872 2644 25924 2650
rect 25872 2586 25924 2592
rect 25516 598 25636 626
rect 25608 480 25636 598
rect 26252 480 26280 2944
rect 26896 480 26924 7482
rect 27526 2816 27582 2825
rect 27526 2751 27582 2760
rect 27540 480 27568 2751
rect 23846 368 23902 377
rect 23846 303 23902 312
rect 24306 0 24362 480
rect 24950 0 25006 480
rect 25594 0 25650 480
rect 26238 0 26294 480
rect 26882 0 26938 480
rect 27526 0 27582 480
<< via2 >>
rect 24030 27648 24086 27704
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 23570 26560 23626 26616
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 17222 23704 17278 23760
rect 10690 23468 10692 23488
rect 10692 23468 10744 23488
rect 10744 23468 10746 23488
rect 10690 23432 10746 23468
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 13726 22616 13782 22672
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 10322 21972 10324 21992
rect 10324 21972 10376 21992
rect 10376 21972 10378 21992
rect 10322 21936 10378 21972
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 8114 16904 8170 16960
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 4066 13368 4122 13424
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 7930 10920 7986 10976
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 1582 9424 1638 9480
rect 294 8064 350 8120
rect 938 7384 994 7440
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 2226 8472 2282 8528
rect 7010 7928 7066 7984
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5446 7248 5502 7304
rect 3514 4528 3570 4584
rect 2870 4120 2926 4176
rect 4802 1672 4858 1728
rect 4158 1536 4214 1592
rect 6734 6840 6790 6896
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 6090 6160 6146 6216
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7378 5752 7434 5808
rect 7102 2896 7158 2952
rect 8574 6704 8630 6760
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 11334 18692 11390 18728
rect 11334 18672 11336 18692
rect 11336 18672 11388 18692
rect 11388 18672 11390 18692
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10138 16940 10140 16960
rect 10140 16940 10192 16960
rect 10192 16940 10194 16960
rect 10138 16904 10194 16940
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 9954 15272 10010 15328
rect 9494 5092 9550 5128
rect 9494 5072 9496 5092
rect 9496 5072 9548 5092
rect 9548 5072 9550 5092
rect 9494 4140 9550 4176
rect 9494 4120 9496 4140
rect 9496 4120 9548 4140
rect 9548 4120 9550 4140
rect 9402 3576 9458 3632
rect 8482 3440 8538 3496
rect 8574 3052 8630 3088
rect 8574 3032 8576 3052
rect 8576 3032 8628 3052
rect 8628 3032 8630 3052
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 11150 9560 11206 9616
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10690 9172 10746 9208
rect 10690 9152 10692 9172
rect 10692 9152 10744 9172
rect 10744 9152 10746 9172
rect 10598 8492 10654 8528
rect 10598 8472 10600 8492
rect 10600 8472 10652 8492
rect 10652 8472 10654 8492
rect 10782 8472 10838 8528
rect 10690 8336 10746 8392
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10874 7248 10930 7304
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 8482 2508 8538 2544
rect 8482 2488 8484 2508
rect 8484 2488 8536 2508
rect 8536 2488 8538 2508
rect 8758 2388 8760 2408
rect 8760 2388 8812 2408
rect 8812 2388 8814 2408
rect 8758 2352 8814 2388
rect 8574 2216 8630 2272
rect 8666 2080 8722 2136
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 12714 17060 12770 17096
rect 12714 17040 12716 17060
rect 12716 17040 12768 17060
rect 12768 17040 12770 17060
rect 12622 15816 12678 15872
rect 12346 15272 12402 15328
rect 11794 9152 11850 9208
rect 12438 8356 12494 8392
rect 12438 8336 12440 8356
rect 12440 8336 12492 8356
rect 12492 8336 12494 8356
rect 11150 7384 11206 7440
rect 11978 7384 12034 7440
rect 11610 6024 11666 6080
rect 11334 5208 11390 5264
rect 10966 3712 11022 3768
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10690 2216 10746 2272
rect 10046 1944 10102 2000
rect 10046 1808 10102 1864
rect 10782 2080 10838 2136
rect 11794 2932 11796 2952
rect 11796 2932 11848 2952
rect 11848 2932 11850 2952
rect 11794 2896 11850 2932
rect 12254 5752 12310 5808
rect 12438 5072 12494 5128
rect 12070 4528 12126 4584
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 13174 9424 13230 9480
rect 13450 18148 13506 18184
rect 13450 18128 13452 18148
rect 13452 18128 13504 18148
rect 13504 18128 13506 18148
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 13634 16088 13690 16144
rect 15198 15852 15200 15872
rect 15200 15852 15252 15872
rect 15252 15852 15254 15872
rect 15198 15816 15254 15852
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 13818 14864 13874 14920
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14554 12688 14610 12744
rect 13910 11600 13966 11656
rect 13818 10920 13874 10976
rect 12898 5788 12900 5808
rect 12900 5788 12952 5808
rect 12952 5788 12954 5808
rect 12898 5752 12954 5788
rect 12714 4936 12770 4992
rect 13082 4004 13138 4040
rect 13082 3984 13084 4004
rect 13084 3984 13136 4004
rect 13136 3984 13138 4004
rect 14186 5616 14242 5672
rect 14186 3576 14242 3632
rect 13358 2624 13414 2680
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15382 11212 15438 11248
rect 15382 11192 15384 11212
rect 15384 11192 15436 11212
rect 15436 11192 15438 11212
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14830 8508 14832 8528
rect 14832 8508 14884 8528
rect 14884 8508 14886 8528
rect 14830 8472 14886 8508
rect 14738 7656 14794 7712
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14646 6060 14648 6080
rect 14648 6060 14700 6080
rect 14700 6060 14702 6080
rect 14646 6024 14702 6060
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15014 4528 15070 4584
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15658 9424 15714 9480
rect 15566 7148 15568 7168
rect 15568 7148 15620 7168
rect 15620 7148 15622 7168
rect 15566 7112 15622 7148
rect 17222 19896 17278 19952
rect 16302 18828 16358 18864
rect 16302 18808 16304 18828
rect 16304 18808 16356 18828
rect 16356 18808 16358 18828
rect 16026 17212 16028 17232
rect 16028 17212 16080 17232
rect 16080 17212 16082 17232
rect 16026 17176 16082 17212
rect 16302 13388 16358 13424
rect 16302 13368 16304 13388
rect 16304 13368 16356 13388
rect 16356 13368 16358 13388
rect 15934 9832 15990 9888
rect 16394 8608 16450 8664
rect 16118 6840 16174 6896
rect 15842 5516 15844 5536
rect 15844 5516 15896 5536
rect 15896 5516 15898 5536
rect 15842 5480 15898 5516
rect 15658 4528 15714 4584
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15106 2916 15162 2952
rect 15106 2896 15108 2916
rect 15108 2896 15160 2916
rect 15160 2896 15162 2916
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15934 3304 15990 3360
rect 15658 1536 15714 1592
rect 16210 6196 16212 6216
rect 16212 6196 16264 6216
rect 16264 6196 16266 6216
rect 16210 6160 16266 6196
rect 16302 3848 16358 3904
rect 17130 9696 17186 9752
rect 17038 5072 17094 5128
rect 16854 2644 16910 2680
rect 16854 2624 16856 2644
rect 16856 2624 16908 2644
rect 16908 2624 16910 2644
rect 17406 12960 17462 13016
rect 17406 11056 17462 11112
rect 18142 13096 18198 13152
rect 18326 16632 18382 16688
rect 18418 12860 18420 12880
rect 18420 12860 18472 12880
rect 18472 12860 18474 12880
rect 18418 12824 18474 12860
rect 18418 11756 18474 11792
rect 18418 11736 18420 11756
rect 18420 11736 18472 11756
rect 18472 11736 18474 11756
rect 17774 8608 17830 8664
rect 17314 8472 17370 8528
rect 17406 6704 17462 6760
rect 17498 5344 17554 5400
rect 18418 4256 18474 4312
rect 17774 3052 17830 3088
rect 17774 3032 17776 3052
rect 17776 3032 17828 3052
rect 17828 3032 17830 3052
rect 18418 3576 18474 3632
rect 19338 12008 19394 12064
rect 19154 8744 19210 8800
rect 19062 8336 19118 8392
rect 19154 7248 19210 7304
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19982 22072 20038 22128
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 21454 20168 21510 20224
rect 23478 19896 23534 19952
rect 19982 16088 20038 16144
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19706 12180 19708 12200
rect 19708 12180 19760 12200
rect 19760 12180 19762 12200
rect 19706 12144 19762 12180
rect 19522 11736 19578 11792
rect 19982 11600 20038 11656
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 20074 11328 20130 11384
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19890 9968 19946 10024
rect 20074 9832 20130 9888
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19798 8628 19854 8664
rect 19798 8608 19800 8628
rect 19800 8608 19852 8628
rect 19852 8608 19854 8628
rect 20074 8336 20130 8392
rect 19338 7792 19394 7848
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19982 7928 20038 7984
rect 19614 7520 19670 7576
rect 18878 6704 18934 6760
rect 19154 4972 19156 4992
rect 19156 4972 19208 4992
rect 19208 4972 19210 4992
rect 19154 4936 19210 4972
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19614 6876 19616 6896
rect 19616 6876 19668 6896
rect 19668 6876 19670 6896
rect 19614 6840 19670 6876
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19522 5752 19578 5808
rect 19430 4936 19486 4992
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 21362 19080 21418 19136
rect 23478 19116 23480 19136
rect 23480 19116 23532 19136
rect 23532 19116 23534 19136
rect 23478 19080 23534 19116
rect 21178 13096 21234 13152
rect 20718 11192 20774 11248
rect 21270 10648 21326 10704
rect 20994 9696 21050 9752
rect 23478 14900 23480 14920
rect 23480 14900 23532 14920
rect 23532 14900 23534 14920
rect 23478 14864 23534 14900
rect 23386 14728 23442 14784
rect 23478 13912 23534 13968
rect 21546 12280 21602 12336
rect 22374 13776 22430 13832
rect 20718 9424 20774 9480
rect 20442 7792 20498 7848
rect 21362 8064 21418 8120
rect 21178 7792 21234 7848
rect 20626 7656 20682 7712
rect 18970 4120 19026 4176
rect 20350 6024 20406 6080
rect 20350 5908 20406 5944
rect 20994 6976 21050 7032
rect 20350 5888 20352 5908
rect 20352 5888 20404 5908
rect 20404 5888 20406 5908
rect 20902 5888 20958 5944
rect 20810 4972 20812 4992
rect 20812 4972 20864 4992
rect 20864 4972 20866 4992
rect 20810 4936 20866 4972
rect 19430 3984 19486 4040
rect 19890 3984 19946 4040
rect 19154 3848 19210 3904
rect 19430 3712 19486 3768
rect 19154 3460 19210 3496
rect 19154 3440 19156 3460
rect 19156 3440 19208 3460
rect 19208 3440 19210 3460
rect 18418 3032 18474 3088
rect 17866 2896 17922 2952
rect 18142 2896 18198 2952
rect 17590 1672 17646 1728
rect 18050 2388 18052 2408
rect 18052 2388 18104 2408
rect 18104 2388 18106 2408
rect 18050 2352 18106 2388
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20074 3848 20130 3904
rect 20166 3440 20222 3496
rect 20534 2932 20536 2952
rect 20536 2932 20588 2952
rect 20588 2932 20590 2952
rect 20534 2896 20590 2932
rect 19154 1400 19210 1456
rect 20442 1944 20498 2000
rect 22190 9424 22246 9480
rect 21914 7520 21970 7576
rect 24122 27104 24178 27160
rect 23846 22072 23902 22128
rect 24030 21392 24086 21448
rect 23754 20304 23810 20360
rect 23662 19080 23718 19136
rect 24030 18808 24086 18864
rect 23754 18672 23810 18728
rect 24030 17992 24086 18048
rect 23662 17176 23718 17232
rect 23938 15000 23994 15056
rect 22926 12008 22982 12064
rect 22374 9152 22430 9208
rect 22282 8780 22284 8800
rect 22284 8780 22336 8800
rect 22336 8780 22338 8800
rect 22282 8744 22338 8780
rect 22190 7384 22246 7440
rect 21454 3304 21510 3360
rect 21362 2896 21418 2952
rect 21454 2760 21510 2816
rect 21638 2760 21694 2816
rect 21546 1536 21602 1592
rect 21822 5208 21878 5264
rect 22006 2896 22062 2952
rect 23202 11736 23258 11792
rect 22926 11056 22982 11112
rect 23570 10104 23626 10160
rect 22650 8508 22652 8528
rect 22652 8508 22704 8528
rect 22704 8508 22706 8528
rect 22650 8472 22706 8508
rect 22650 7384 22706 7440
rect 22374 3984 22430 4040
rect 22282 3032 22338 3088
rect 22650 1400 22706 1456
rect 22926 6160 22982 6216
rect 22926 5752 22982 5808
rect 23110 5772 23166 5808
rect 23846 12824 23902 12880
rect 24674 26016 24730 26072
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24214 24248 24270 24304
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 25336 24822 25392
rect 24766 24656 24822 24712
rect 24674 23160 24730 23216
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24582 22616 24638 22672
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24766 22480 24822 22536
rect 24950 21936 25006 21992
rect 25134 21936 25190 21992
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24766 20848 24822 20904
rect 24582 20204 24584 20224
rect 24584 20204 24636 20224
rect 24636 20204 24638 20224
rect 24582 20168 24638 20204
rect 24674 19624 24730 19680
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24582 18808 24638 18864
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 26238 20984 26294 21040
rect 24766 18536 24822 18592
rect 24674 17448 24730 17504
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24950 18128 25006 18184
rect 24398 16632 24454 16688
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 25134 17076 25136 17096
rect 25136 17076 25188 17096
rect 25188 17076 25190 17096
rect 25134 17040 25190 17076
rect 25042 16768 25098 16824
rect 24766 15680 24822 15736
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24858 14764 24860 14784
rect 24860 14764 24912 14784
rect 24912 14764 24914 14784
rect 24858 14728 24914 14764
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24766 13776 24822 13832
rect 24030 12980 24086 13016
rect 24030 12960 24032 12980
rect 24032 12960 24084 12980
rect 24084 12960 24086 12980
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24306 12824 24362 12880
rect 23938 12144 23994 12200
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24858 11328 24914 11384
rect 24674 11056 24730 11112
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24490 10648 24546 10704
rect 24306 9988 24362 10024
rect 24306 9968 24308 9988
rect 24308 9968 24360 9988
rect 24360 9968 24362 9988
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24030 8880 24086 8936
rect 23754 7656 23810 7712
rect 23570 6976 23626 7032
rect 23110 5752 23112 5772
rect 23112 5752 23164 5772
rect 23164 5752 23166 5772
rect 23202 5616 23258 5672
rect 23110 4936 23166 4992
rect 23110 4256 23166 4312
rect 23386 4936 23442 4992
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24214 8236 24216 8256
rect 24216 8236 24268 8256
rect 24268 8236 24270 8256
rect 24214 8200 24270 8236
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24122 6160 24178 6216
rect 24030 5752 24086 5808
rect 24030 4120 24086 4176
rect 23662 3576 23718 3632
rect 23846 2760 23902 2816
rect 23478 1808 23534 1864
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24766 10512 24822 10568
rect 24858 9560 24914 9616
rect 24858 9172 24914 9208
rect 24858 9152 24860 9172
rect 24860 9152 24912 9172
rect 24912 9152 24914 9172
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24674 4936 24730 4992
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 25502 16224 25558 16280
rect 25318 12688 25374 12744
rect 25778 14592 25834 14648
rect 25686 13368 25742 13424
rect 25226 8064 25282 8120
rect 25226 7384 25282 7440
rect 25502 5888 25558 5944
rect 24950 5072 25006 5128
rect 24674 4256 24730 4312
rect 24214 3440 24270 3496
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24674 1944 24730 2000
rect 24858 2508 24914 2544
rect 24858 2488 24860 2508
rect 24860 2488 24912 2508
rect 24912 2488 24914 2508
rect 24766 856 24822 912
rect 25042 3848 25098 3904
rect 25134 3188 25190 3224
rect 25134 3168 25136 3188
rect 25136 3168 25188 3188
rect 25188 3168 25190 3188
rect 25318 3032 25374 3088
rect 25502 5480 25558 5536
rect 25410 2896 25466 2952
rect 25410 2796 25412 2816
rect 25412 2796 25464 2816
rect 25464 2796 25466 2816
rect 25410 2760 25466 2796
rect 25042 2524 25044 2544
rect 25044 2524 25096 2544
rect 25096 2524 25098 2544
rect 25042 2488 25098 2524
rect 26330 13776 26386 13832
rect 25778 3712 25834 3768
rect 27526 2760 27582 2816
rect 23846 312 23902 368
<< metal3 >>
rect 24025 27706 24091 27709
rect 27520 27706 28000 27736
rect 24025 27704 28000 27706
rect 24025 27648 24030 27704
rect 24086 27648 28000 27704
rect 24025 27646 28000 27648
rect 24025 27643 24091 27646
rect 27520 27616 28000 27646
rect 24117 27162 24183 27165
rect 27520 27162 28000 27192
rect 24117 27160 28000 27162
rect 24117 27104 24122 27160
rect 24178 27104 28000 27160
rect 24117 27102 28000 27104
rect 24117 27099 24183 27102
rect 27520 27072 28000 27102
rect 23565 26618 23631 26621
rect 27520 26618 28000 26648
rect 23565 26616 28000 26618
rect 23565 26560 23570 26616
rect 23626 26560 28000 26616
rect 23565 26558 28000 26560
rect 23565 26555 23631 26558
rect 27520 26528 28000 26558
rect 24669 26074 24735 26077
rect 27520 26074 28000 26104
rect 24669 26072 28000 26074
rect 24669 26016 24674 26072
rect 24730 26016 28000 26072
rect 24669 26014 28000 26016
rect 24669 26011 24735 26014
rect 27520 25984 28000 26014
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 24761 25394 24827 25397
rect 27520 25394 28000 25424
rect 24761 25392 28000 25394
rect 24761 25336 24766 25392
rect 24822 25336 28000 25392
rect 24761 25334 28000 25336
rect 24761 25331 24827 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 27520 24850 28000 24880
rect 24902 24790 28000 24850
rect 24761 24714 24827 24717
rect 24902 24714 24962 24790
rect 27520 24760 28000 24790
rect 24761 24712 24962 24714
rect 24761 24656 24766 24712
rect 24822 24656 24962 24712
rect 24761 24654 24962 24656
rect 24761 24651 24827 24654
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 24209 24306 24275 24309
rect 27520 24306 28000 24336
rect 24209 24304 28000 24306
rect 24209 24248 24214 24304
rect 24270 24248 28000 24304
rect 24209 24246 28000 24248
rect 24209 24243 24275 24246
rect 27520 24216 28000 24246
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 17217 23762 17283 23765
rect 27520 23762 28000 23792
rect 17217 23760 28000 23762
rect 17217 23704 17222 23760
rect 17278 23704 28000 23760
rect 17217 23702 28000 23704
rect 17217 23699 17283 23702
rect 27520 23672 28000 23702
rect 10685 23490 10751 23493
rect 10685 23488 12634 23490
rect 10685 23432 10690 23488
rect 10746 23432 12634 23488
rect 10685 23430 12634 23432
rect 10685 23427 10751 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 12574 23218 12634 23430
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 19374 23218 19380 23220
rect 12574 23158 19380 23218
rect 19374 23156 19380 23158
rect 19444 23156 19450 23220
rect 24669 23218 24735 23221
rect 27520 23218 28000 23248
rect 24669 23216 28000 23218
rect 24669 23160 24674 23216
rect 24730 23160 28000 23216
rect 24669 23158 28000 23160
rect 24669 23155 24735 23158
rect 27520 23128 28000 23158
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 13721 22674 13787 22677
rect 24577 22674 24643 22677
rect 13721 22672 24643 22674
rect 13721 22616 13726 22672
rect 13782 22616 24582 22672
rect 24638 22616 24643 22672
rect 13721 22614 24643 22616
rect 13721 22611 13787 22614
rect 24577 22611 24643 22614
rect 24761 22538 24827 22541
rect 27520 22538 28000 22568
rect 24761 22536 28000 22538
rect 24761 22480 24766 22536
rect 24822 22480 28000 22536
rect 24761 22478 28000 22480
rect 24761 22475 24827 22478
rect 27520 22448 28000 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 19977 22130 20043 22133
rect 23841 22130 23907 22133
rect 19977 22128 23907 22130
rect 19977 22072 19982 22128
rect 20038 22072 23846 22128
rect 23902 22072 23907 22128
rect 19977 22070 23907 22072
rect 19977 22067 20043 22070
rect 23841 22067 23907 22070
rect 10317 21994 10383 21997
rect 24945 21994 25011 21997
rect 10317 21992 25011 21994
rect 10317 21936 10322 21992
rect 10378 21936 24950 21992
rect 25006 21936 25011 21992
rect 10317 21934 25011 21936
rect 10317 21931 10383 21934
rect 24945 21931 25011 21934
rect 25129 21994 25195 21997
rect 27520 21994 28000 22024
rect 25129 21992 28000 21994
rect 25129 21936 25134 21992
rect 25190 21936 28000 21992
rect 25129 21934 28000 21936
rect 25129 21931 25195 21934
rect 27520 21904 28000 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 24025 21450 24091 21453
rect 27520 21450 28000 21480
rect 24025 21448 28000 21450
rect 24025 21392 24030 21448
rect 24086 21392 28000 21448
rect 24025 21390 28000 21392
rect 24025 21387 24091 21390
rect 27520 21360 28000 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 19374 20980 19380 21044
rect 19444 21042 19450 21044
rect 26233 21042 26299 21045
rect 19444 21040 26299 21042
rect 19444 20984 26238 21040
rect 26294 20984 26299 21040
rect 19444 20982 26299 20984
rect 19444 20980 19450 20982
rect 26233 20979 26299 20982
rect 24761 20906 24827 20909
rect 27520 20906 28000 20936
rect 24761 20904 28000 20906
rect 24761 20848 24766 20904
rect 24822 20848 28000 20904
rect 24761 20846 28000 20848
rect 24761 20843 24827 20846
rect 27520 20816 28000 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 23749 20362 23815 20365
rect 27520 20362 28000 20392
rect 23749 20360 28000 20362
rect 23749 20304 23754 20360
rect 23810 20304 28000 20360
rect 23749 20302 28000 20304
rect 23749 20299 23815 20302
rect 27520 20272 28000 20302
rect 21449 20226 21515 20229
rect 24577 20226 24643 20229
rect 21449 20224 24643 20226
rect 21449 20168 21454 20224
rect 21510 20168 24582 20224
rect 24638 20168 24643 20224
rect 21449 20166 24643 20168
rect 21449 20163 21515 20166
rect 24577 20163 24643 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 17217 19954 17283 19957
rect 23473 19954 23539 19957
rect 17217 19952 23539 19954
rect 17217 19896 17222 19952
rect 17278 19896 23478 19952
rect 23534 19896 23539 19952
rect 17217 19894 23539 19896
rect 17217 19891 17283 19894
rect 23473 19891 23539 19894
rect 24669 19682 24735 19685
rect 27520 19682 28000 19712
rect 24669 19680 28000 19682
rect 24669 19624 24674 19680
rect 24730 19624 28000 19680
rect 24669 19622 28000 19624
rect 24669 19619 24735 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 27520 19592 28000 19622
rect 24277 19551 24597 19552
rect 21357 19138 21423 19141
rect 23473 19138 23539 19141
rect 21357 19136 23539 19138
rect 21357 19080 21362 19136
rect 21418 19080 23478 19136
rect 23534 19080 23539 19136
rect 21357 19078 23539 19080
rect 21357 19075 21423 19078
rect 23473 19075 23539 19078
rect 23657 19138 23723 19141
rect 27520 19138 28000 19168
rect 23657 19136 28000 19138
rect 23657 19080 23662 19136
rect 23718 19080 28000 19136
rect 23657 19078 28000 19080
rect 23657 19075 23723 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 16297 18866 16363 18869
rect 24025 18866 24091 18869
rect 24577 18866 24643 18869
rect 16297 18864 24643 18866
rect 16297 18808 16302 18864
rect 16358 18808 24030 18864
rect 24086 18808 24582 18864
rect 24638 18808 24643 18864
rect 16297 18806 24643 18808
rect 16297 18803 16363 18806
rect 24025 18803 24091 18806
rect 24577 18803 24643 18806
rect 11329 18730 11395 18733
rect 23749 18730 23815 18733
rect 11329 18728 23815 18730
rect 11329 18672 11334 18728
rect 11390 18672 23754 18728
rect 23810 18672 23815 18728
rect 11329 18670 23815 18672
rect 11329 18667 11395 18670
rect 23749 18667 23815 18670
rect 24761 18594 24827 18597
rect 27520 18594 28000 18624
rect 24761 18592 28000 18594
rect 24761 18536 24766 18592
rect 24822 18536 28000 18592
rect 24761 18534 28000 18536
rect 24761 18531 24827 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 27520 18504 28000 18534
rect 24277 18463 24597 18464
rect 13445 18186 13511 18189
rect 24945 18186 25011 18189
rect 13445 18184 25011 18186
rect 13445 18128 13450 18184
rect 13506 18128 24950 18184
rect 25006 18128 25011 18184
rect 13445 18126 25011 18128
rect 13445 18123 13511 18126
rect 24945 18123 25011 18126
rect 24025 18050 24091 18053
rect 27520 18050 28000 18080
rect 24025 18048 28000 18050
rect 24025 17992 24030 18048
rect 24086 17992 28000 18048
rect 24025 17990 28000 17992
rect 24025 17987 24091 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 17990
rect 19610 17919 19930 17920
rect 24669 17506 24735 17509
rect 27520 17506 28000 17536
rect 24669 17504 28000 17506
rect 24669 17448 24674 17504
rect 24730 17448 28000 17504
rect 24669 17446 28000 17448
rect 24669 17443 24735 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17446
rect 24277 17375 24597 17376
rect 16021 17234 16087 17237
rect 23657 17234 23723 17237
rect 16021 17232 23723 17234
rect 16021 17176 16026 17232
rect 16082 17176 23662 17232
rect 23718 17176 23723 17232
rect 16021 17174 23723 17176
rect 16021 17171 16087 17174
rect 23657 17171 23723 17174
rect 12709 17098 12775 17101
rect 25129 17098 25195 17101
rect 12709 17096 25195 17098
rect 12709 17040 12714 17096
rect 12770 17040 25134 17096
rect 25190 17040 25195 17096
rect 12709 17038 25195 17040
rect 12709 17035 12775 17038
rect 25129 17035 25195 17038
rect 8109 16962 8175 16965
rect 10133 16962 10199 16965
rect 8109 16960 10199 16962
rect 8109 16904 8114 16960
rect 8170 16904 10138 16960
rect 10194 16904 10199 16960
rect 8109 16902 10199 16904
rect 8109 16899 8175 16902
rect 10133 16899 10199 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 25037 16826 25103 16829
rect 27520 16826 28000 16856
rect 25037 16824 28000 16826
rect 25037 16768 25042 16824
rect 25098 16768 28000 16824
rect 25037 16766 28000 16768
rect 25037 16763 25103 16766
rect 27520 16736 28000 16766
rect 18321 16690 18387 16693
rect 24393 16690 24459 16693
rect 18321 16688 24459 16690
rect 18321 16632 18326 16688
rect 18382 16632 24398 16688
rect 24454 16632 24459 16688
rect 18321 16630 24459 16632
rect 18321 16627 18387 16630
rect 24393 16627 24459 16630
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 25497 16282 25563 16285
rect 27520 16282 28000 16312
rect 25497 16280 28000 16282
rect 25497 16224 25502 16280
rect 25558 16224 28000 16280
rect 25497 16222 28000 16224
rect 25497 16219 25563 16222
rect 27520 16192 28000 16222
rect 13629 16146 13695 16149
rect 19977 16146 20043 16149
rect 13629 16144 20043 16146
rect 13629 16088 13634 16144
rect 13690 16088 19982 16144
rect 20038 16088 20043 16144
rect 13629 16086 20043 16088
rect 13629 16083 13695 16086
rect 19977 16083 20043 16086
rect 12617 15874 12683 15877
rect 15193 15874 15259 15877
rect 12617 15872 15259 15874
rect 12617 15816 12622 15872
rect 12678 15816 15198 15872
rect 15254 15816 15259 15872
rect 12617 15814 15259 15816
rect 12617 15811 12683 15814
rect 15193 15811 15259 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 24761 15738 24827 15741
rect 27520 15738 28000 15768
rect 24761 15736 28000 15738
rect 24761 15680 24766 15736
rect 24822 15680 28000 15736
rect 24761 15678 28000 15680
rect 24761 15675 24827 15678
rect 27520 15648 28000 15678
rect 9949 15330 10015 15333
rect 12341 15330 12407 15333
rect 9949 15328 12407 15330
rect 9949 15272 9954 15328
rect 10010 15272 12346 15328
rect 12402 15272 12407 15328
rect 9949 15270 12407 15272
rect 9949 15267 10015 15270
rect 12341 15267 12407 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 27520 15194 28000 15224
rect 27478 15104 28000 15194
rect 23933 15058 23999 15061
rect 27478 15058 27538 15104
rect 23933 15056 27538 15058
rect 23933 15000 23938 15056
rect 23994 15000 27538 15056
rect 23933 14998 27538 15000
rect 23933 14995 23999 14998
rect 13813 14922 13879 14925
rect 23473 14922 23539 14925
rect 13813 14920 23539 14922
rect 13813 14864 13818 14920
rect 13874 14864 23478 14920
rect 23534 14864 23539 14920
rect 13813 14862 23539 14864
rect 13813 14859 13879 14862
rect 23473 14859 23539 14862
rect 23381 14786 23447 14789
rect 24853 14786 24919 14789
rect 23381 14784 24919 14786
rect 23381 14728 23386 14784
rect 23442 14728 24858 14784
rect 24914 14728 24919 14784
rect 23381 14726 24919 14728
rect 23381 14723 23447 14726
rect 24853 14723 24919 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 25773 14650 25839 14653
rect 27520 14650 28000 14680
rect 25773 14648 28000 14650
rect 25773 14592 25778 14648
rect 25834 14592 28000 14648
rect 25773 14590 28000 14592
rect 25773 14587 25839 14590
rect 27520 14560 28000 14590
rect 5610 14176 5930 14177
rect 0 14106 480 14136
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 14046 2698 14106
rect 0 14016 480 14046
rect 2638 13834 2698 14046
rect 23473 13970 23539 13973
rect 27520 13970 28000 14000
rect 23473 13968 28000 13970
rect 23473 13912 23478 13968
rect 23534 13912 28000 13968
rect 23473 13910 28000 13912
rect 23473 13907 23539 13910
rect 27520 13880 28000 13910
rect 22369 13834 22435 13837
rect 2638 13832 22435 13834
rect 2638 13776 22374 13832
rect 22430 13776 22435 13832
rect 2638 13774 22435 13776
rect 22369 13771 22435 13774
rect 24761 13834 24827 13837
rect 26325 13834 26391 13837
rect 24761 13832 26391 13834
rect 24761 13776 24766 13832
rect 24822 13776 26330 13832
rect 26386 13776 26391 13832
rect 24761 13774 26391 13776
rect 24761 13771 24827 13774
rect 26325 13771 26391 13774
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 4061 13426 4127 13429
rect 16297 13426 16363 13429
rect 4061 13424 16363 13426
rect 4061 13368 4066 13424
rect 4122 13368 16302 13424
rect 16358 13368 16363 13424
rect 4061 13366 16363 13368
rect 4061 13363 4127 13366
rect 16297 13363 16363 13366
rect 25681 13426 25747 13429
rect 27520 13426 28000 13456
rect 25681 13424 28000 13426
rect 25681 13368 25686 13424
rect 25742 13368 28000 13424
rect 25681 13366 28000 13368
rect 25681 13363 25747 13366
rect 27520 13336 28000 13366
rect 18137 13154 18203 13157
rect 21173 13154 21239 13157
rect 18137 13152 21239 13154
rect 18137 13096 18142 13152
rect 18198 13096 21178 13152
rect 21234 13096 21239 13152
rect 18137 13094 21239 13096
rect 18137 13091 18203 13094
rect 21173 13091 21239 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 17401 13018 17467 13021
rect 24025 13018 24091 13021
rect 17401 13016 24091 13018
rect 17401 12960 17406 13016
rect 17462 12960 24030 13016
rect 24086 12960 24091 13016
rect 17401 12958 24091 12960
rect 17401 12955 17467 12958
rect 24025 12955 24091 12958
rect 18413 12882 18479 12885
rect 23841 12882 23907 12885
rect 18413 12880 23907 12882
rect 18413 12824 18418 12880
rect 18474 12824 23846 12880
rect 23902 12824 23907 12880
rect 18413 12822 23907 12824
rect 18413 12819 18479 12822
rect 23841 12819 23907 12822
rect 24301 12882 24367 12885
rect 27520 12882 28000 12912
rect 24301 12880 28000 12882
rect 24301 12824 24306 12880
rect 24362 12824 28000 12880
rect 24301 12822 28000 12824
rect 24301 12819 24367 12822
rect 27520 12792 28000 12822
rect 14549 12746 14615 12749
rect 25313 12746 25379 12749
rect 14549 12744 25379 12746
rect 14549 12688 14554 12744
rect 14610 12688 25318 12744
rect 25374 12688 25379 12744
rect 14549 12686 25379 12688
rect 14549 12683 14615 12686
rect 25313 12683 25379 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 21541 12338 21607 12341
rect 27520 12338 28000 12368
rect 21541 12336 28000 12338
rect 21541 12280 21546 12336
rect 21602 12280 28000 12336
rect 21541 12278 28000 12280
rect 21541 12275 21607 12278
rect 27520 12248 28000 12278
rect 19701 12202 19767 12205
rect 23933 12202 23999 12205
rect 19701 12200 23999 12202
rect 19701 12144 19706 12200
rect 19762 12144 23938 12200
rect 23994 12144 23999 12200
rect 19701 12142 23999 12144
rect 19701 12139 19767 12142
rect 23933 12139 23999 12142
rect 19333 12066 19399 12069
rect 22921 12066 22987 12069
rect 19333 12064 22987 12066
rect 19333 12008 19338 12064
rect 19394 12008 22926 12064
rect 22982 12008 22987 12064
rect 19333 12006 22987 12008
rect 19333 12003 19399 12006
rect 22921 12003 22987 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 18413 11794 18479 11797
rect 19517 11794 19583 11797
rect 18413 11792 19583 11794
rect 18413 11736 18418 11792
rect 18474 11736 19522 11792
rect 19578 11736 19583 11792
rect 18413 11734 19583 11736
rect 18413 11731 18479 11734
rect 19517 11731 19583 11734
rect 23197 11794 23263 11797
rect 27520 11794 28000 11824
rect 23197 11792 28000 11794
rect 23197 11736 23202 11792
rect 23258 11736 28000 11792
rect 23197 11734 28000 11736
rect 23197 11731 23263 11734
rect 27520 11704 28000 11734
rect 13905 11658 13971 11661
rect 19977 11658 20043 11661
rect 13905 11656 20043 11658
rect 13905 11600 13910 11656
rect 13966 11600 19982 11656
rect 20038 11600 20043 11656
rect 13905 11598 20043 11600
rect 13905 11595 13971 11598
rect 19977 11595 20043 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 20069 11386 20135 11389
rect 24853 11386 24919 11389
rect 20069 11384 24919 11386
rect 20069 11328 20074 11384
rect 20130 11328 24858 11384
rect 24914 11328 24919 11384
rect 20069 11326 24919 11328
rect 20069 11323 20135 11326
rect 24853 11323 24919 11326
rect 15377 11250 15443 11253
rect 20713 11250 20779 11253
rect 15377 11248 20779 11250
rect 15377 11192 15382 11248
rect 15438 11192 20718 11248
rect 20774 11192 20779 11248
rect 15377 11190 20779 11192
rect 15377 11187 15443 11190
rect 20713 11187 20779 11190
rect 17401 11114 17467 11117
rect 22921 11114 22987 11117
rect 17401 11112 22987 11114
rect 17401 11056 17406 11112
rect 17462 11056 22926 11112
rect 22982 11056 22987 11112
rect 17401 11054 22987 11056
rect 17401 11051 17467 11054
rect 22921 11051 22987 11054
rect 24669 11114 24735 11117
rect 27520 11114 28000 11144
rect 24669 11112 28000 11114
rect 24669 11056 24674 11112
rect 24730 11056 28000 11112
rect 24669 11054 28000 11056
rect 24669 11051 24735 11054
rect 27520 11024 28000 11054
rect 7925 10978 7991 10981
rect 13813 10978 13879 10981
rect 7925 10976 13879 10978
rect 7925 10920 7930 10976
rect 7986 10920 13818 10976
rect 13874 10920 13879 10976
rect 7925 10918 13879 10920
rect 7925 10915 7991 10918
rect 13813 10915 13879 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 21265 10706 21331 10709
rect 24485 10706 24551 10709
rect 21265 10704 24551 10706
rect 21265 10648 21270 10704
rect 21326 10648 24490 10704
rect 24546 10648 24551 10704
rect 21265 10646 24551 10648
rect 21265 10643 21331 10646
rect 24485 10643 24551 10646
rect 24761 10570 24827 10573
rect 27520 10570 28000 10600
rect 24761 10568 28000 10570
rect 24761 10512 24766 10568
rect 24822 10512 28000 10568
rect 24761 10510 28000 10512
rect 24761 10507 24827 10510
rect 27520 10480 28000 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 23565 10162 23631 10165
rect 23565 10160 24916 10162
rect 23565 10104 23570 10160
rect 23626 10104 24916 10160
rect 23565 10102 24916 10104
rect 23565 10099 23631 10102
rect 19885 10026 19951 10029
rect 24301 10026 24367 10029
rect 19885 10024 24367 10026
rect 19885 9968 19890 10024
rect 19946 9968 24306 10024
rect 24362 9968 24367 10024
rect 19885 9966 24367 9968
rect 24856 10026 24916 10102
rect 27520 10026 28000 10056
rect 24856 9966 28000 10026
rect 19885 9963 19951 9966
rect 24301 9963 24367 9966
rect 27520 9936 28000 9966
rect 15929 9890 15995 9893
rect 20069 9890 20135 9893
rect 15929 9888 20135 9890
rect 15929 9832 15934 9888
rect 15990 9832 20074 9888
rect 20130 9832 20135 9888
rect 15929 9830 20135 9832
rect 15929 9827 15995 9830
rect 20069 9827 20135 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 17125 9754 17191 9757
rect 20989 9754 21055 9757
rect 17125 9752 21055 9754
rect 17125 9696 17130 9752
rect 17186 9696 20994 9752
rect 21050 9696 21055 9752
rect 17125 9694 21055 9696
rect 17125 9691 17191 9694
rect 20989 9691 21055 9694
rect 11145 9618 11211 9621
rect 24853 9618 24919 9621
rect 11145 9616 24919 9618
rect 11145 9560 11150 9616
rect 11206 9560 24858 9616
rect 24914 9560 24919 9616
rect 11145 9558 24919 9560
rect 11145 9555 11211 9558
rect 24853 9555 24919 9558
rect 1577 9482 1643 9485
rect 13169 9482 13235 9485
rect 1577 9480 13235 9482
rect 1577 9424 1582 9480
rect 1638 9424 13174 9480
rect 13230 9424 13235 9480
rect 1577 9422 13235 9424
rect 1577 9419 1643 9422
rect 13169 9419 13235 9422
rect 15653 9482 15719 9485
rect 20713 9482 20779 9485
rect 15653 9480 20779 9482
rect 15653 9424 15658 9480
rect 15714 9424 20718 9480
rect 20774 9424 20779 9480
rect 15653 9422 20779 9424
rect 15653 9419 15719 9422
rect 20713 9419 20779 9422
rect 22185 9482 22251 9485
rect 27520 9482 28000 9512
rect 22185 9480 28000 9482
rect 22185 9424 22190 9480
rect 22246 9424 28000 9480
rect 22185 9422 28000 9424
rect 22185 9419 22251 9422
rect 27520 9392 28000 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 10685 9210 10751 9213
rect 11789 9210 11855 9213
rect 10685 9208 11855 9210
rect 10685 9152 10690 9208
rect 10746 9152 11794 9208
rect 11850 9152 11855 9208
rect 10685 9150 11855 9152
rect 10685 9147 10751 9150
rect 11789 9147 11855 9150
rect 22369 9210 22435 9213
rect 24853 9210 24919 9213
rect 22369 9208 24919 9210
rect 22369 9152 22374 9208
rect 22430 9152 24858 9208
rect 24914 9152 24919 9208
rect 22369 9150 24919 9152
rect 22369 9147 22435 9150
rect 24853 9147 24919 9150
rect 24025 8938 24091 8941
rect 27520 8938 28000 8968
rect 24025 8936 28000 8938
rect 24025 8880 24030 8936
rect 24086 8880 28000 8936
rect 24025 8878 28000 8880
rect 24025 8875 24091 8878
rect 27520 8848 28000 8878
rect 19149 8802 19215 8805
rect 22277 8802 22343 8805
rect 19149 8800 22343 8802
rect 19149 8744 19154 8800
rect 19210 8744 22282 8800
rect 22338 8744 22343 8800
rect 19149 8742 22343 8744
rect 19149 8739 19215 8742
rect 22277 8739 22343 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 16389 8666 16455 8669
rect 17769 8666 17835 8669
rect 19793 8666 19859 8669
rect 16389 8664 19859 8666
rect 16389 8608 16394 8664
rect 16450 8608 17774 8664
rect 17830 8608 19798 8664
rect 19854 8608 19859 8664
rect 16389 8606 19859 8608
rect 16389 8603 16455 8606
rect 17769 8603 17835 8606
rect 19793 8603 19859 8606
rect 2221 8530 2287 8533
rect 10593 8530 10659 8533
rect 2221 8528 10659 8530
rect 2221 8472 2226 8528
rect 2282 8472 10598 8528
rect 10654 8472 10659 8528
rect 2221 8470 10659 8472
rect 2221 8467 2287 8470
rect 10593 8467 10659 8470
rect 10777 8530 10843 8533
rect 14825 8530 14891 8533
rect 10777 8528 14891 8530
rect 10777 8472 10782 8528
rect 10838 8472 14830 8528
rect 14886 8472 14891 8528
rect 10777 8470 14891 8472
rect 10777 8467 10843 8470
rect 14825 8467 14891 8470
rect 17309 8530 17375 8533
rect 22645 8530 22711 8533
rect 17309 8528 22711 8530
rect 17309 8472 17314 8528
rect 17370 8472 22650 8528
rect 22706 8472 22711 8528
rect 17309 8470 22711 8472
rect 17309 8467 17375 8470
rect 22645 8467 22711 8470
rect 10685 8394 10751 8397
rect 12433 8394 12499 8397
rect 10685 8392 12499 8394
rect 10685 8336 10690 8392
rect 10746 8336 12438 8392
rect 12494 8336 12499 8392
rect 10685 8334 12499 8336
rect 10685 8331 10751 8334
rect 12433 8331 12499 8334
rect 19057 8394 19123 8397
rect 20069 8394 20135 8397
rect 19057 8392 20135 8394
rect 19057 8336 19062 8392
rect 19118 8336 20074 8392
rect 20130 8336 20135 8392
rect 19057 8334 20135 8336
rect 19057 8331 19123 8334
rect 20069 8331 20135 8334
rect 24209 8258 24275 8261
rect 27520 8258 28000 8288
rect 24209 8256 28000 8258
rect 24209 8200 24214 8256
rect 24270 8200 28000 8256
rect 24209 8198 28000 8200
rect 24209 8195 24275 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8198
rect 19610 8127 19930 8128
rect 289 8122 355 8125
rect 21357 8122 21423 8125
rect 25221 8122 25287 8125
rect 289 8120 6930 8122
rect 289 8064 294 8120
rect 350 8064 6930 8120
rect 289 8062 6930 8064
rect 289 8059 355 8062
rect 6870 7850 6930 8062
rect 21357 8120 25287 8122
rect 21357 8064 21362 8120
rect 21418 8064 25226 8120
rect 25282 8064 25287 8120
rect 21357 8062 25287 8064
rect 21357 8059 21423 8062
rect 25221 8059 25287 8062
rect 7005 7986 7071 7989
rect 19977 7986 20043 7989
rect 7005 7984 19810 7986
rect 7005 7928 7010 7984
rect 7066 7928 19810 7984
rect 7005 7926 19810 7928
rect 7005 7923 7071 7926
rect 19333 7850 19399 7853
rect 6870 7848 19399 7850
rect 6870 7792 19338 7848
rect 19394 7792 19399 7848
rect 6870 7790 19399 7792
rect 19333 7787 19399 7790
rect 14733 7714 14799 7717
rect 7606 7712 14799 7714
rect 7606 7656 14738 7712
rect 14794 7656 14799 7712
rect 7606 7654 14799 7656
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 933 7442 999 7445
rect 7606 7442 7666 7654
rect 14733 7651 14799 7654
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 19609 7578 19675 7581
rect 16990 7576 19675 7578
rect 16990 7520 19614 7576
rect 19670 7520 19675 7576
rect 16990 7518 19675 7520
rect 19750 7578 19810 7926
rect 19977 7984 24916 7986
rect 19977 7928 19982 7984
rect 20038 7928 24916 7984
rect 19977 7926 24916 7928
rect 19977 7923 20043 7926
rect 20437 7850 20503 7853
rect 21173 7850 21239 7853
rect 20437 7848 21239 7850
rect 20437 7792 20442 7848
rect 20498 7792 21178 7848
rect 21234 7792 21239 7848
rect 20437 7790 21239 7792
rect 20437 7787 20503 7790
rect 21173 7787 21239 7790
rect 20621 7714 20687 7717
rect 23749 7714 23815 7717
rect 20621 7712 23815 7714
rect 20621 7656 20626 7712
rect 20682 7656 23754 7712
rect 23810 7656 23815 7712
rect 20621 7654 23815 7656
rect 24856 7714 24916 7926
rect 27520 7714 28000 7744
rect 24856 7654 28000 7714
rect 20621 7651 20687 7654
rect 23749 7651 23815 7654
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7654
rect 24277 7583 24597 7584
rect 21909 7578 21975 7581
rect 19750 7576 21975 7578
rect 19750 7520 21914 7576
rect 21970 7520 21975 7576
rect 19750 7518 21975 7520
rect 11145 7442 11211 7445
rect 933 7440 7666 7442
rect 933 7384 938 7440
rect 994 7384 7666 7440
rect 933 7382 7666 7384
rect 7790 7440 11211 7442
rect 7790 7384 11150 7440
rect 11206 7384 11211 7440
rect 7790 7382 11211 7384
rect 933 7379 999 7382
rect 5441 7306 5507 7309
rect 7790 7306 7850 7382
rect 11145 7379 11211 7382
rect 11973 7442 12039 7445
rect 16990 7442 17050 7518
rect 19609 7515 19675 7518
rect 21909 7515 21975 7518
rect 22185 7442 22251 7445
rect 11973 7440 17050 7442
rect 11973 7384 11978 7440
rect 12034 7384 17050 7440
rect 11973 7382 17050 7384
rect 17174 7440 22251 7442
rect 17174 7384 22190 7440
rect 22246 7384 22251 7440
rect 17174 7382 22251 7384
rect 11973 7379 12039 7382
rect 10869 7306 10935 7309
rect 17174 7306 17234 7382
rect 22185 7379 22251 7382
rect 22645 7442 22711 7445
rect 25221 7442 25287 7445
rect 22645 7440 25287 7442
rect 22645 7384 22650 7440
rect 22706 7384 25226 7440
rect 25282 7384 25287 7440
rect 22645 7382 25287 7384
rect 22645 7379 22711 7382
rect 25221 7379 25287 7382
rect 5441 7304 7850 7306
rect 5441 7248 5446 7304
rect 5502 7248 7850 7304
rect 5441 7246 7850 7248
rect 8342 7246 10794 7306
rect 5441 7243 5507 7246
rect 6729 6898 6795 6901
rect 8342 6898 8402 7246
rect 10734 7170 10794 7246
rect 10869 7304 17234 7306
rect 10869 7248 10874 7304
rect 10930 7248 17234 7304
rect 10869 7246 17234 7248
rect 19149 7306 19215 7309
rect 19149 7304 24916 7306
rect 19149 7248 19154 7304
rect 19210 7248 24916 7304
rect 19149 7246 24916 7248
rect 10869 7243 10935 7246
rect 19149 7243 19215 7246
rect 15561 7170 15627 7173
rect 10734 7168 15627 7170
rect 10734 7112 15566 7168
rect 15622 7112 15627 7168
rect 10734 7110 15627 7112
rect 24856 7170 24916 7246
rect 27520 7170 28000 7200
rect 24856 7110 28000 7170
rect 15561 7107 15627 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 27520 7080 28000 7110
rect 19610 7039 19930 7040
rect 20989 7034 21055 7037
rect 23565 7034 23631 7037
rect 20989 7032 23631 7034
rect 20989 6976 20994 7032
rect 21050 6976 23570 7032
rect 23626 6976 23631 7032
rect 20989 6974 23631 6976
rect 20989 6971 21055 6974
rect 23565 6971 23631 6974
rect 6729 6896 8402 6898
rect 6729 6840 6734 6896
rect 6790 6840 8402 6896
rect 6729 6838 8402 6840
rect 16113 6898 16179 6901
rect 19609 6898 19675 6901
rect 16113 6896 19675 6898
rect 16113 6840 16118 6896
rect 16174 6840 19614 6896
rect 19670 6840 19675 6896
rect 16113 6838 19675 6840
rect 6729 6835 6795 6838
rect 16113 6835 16179 6838
rect 19609 6835 19675 6838
rect 8569 6762 8635 6765
rect 17401 6762 17467 6765
rect 8569 6760 17467 6762
rect 8569 6704 8574 6760
rect 8630 6704 17406 6760
rect 17462 6704 17467 6760
rect 8569 6702 17467 6704
rect 8569 6699 8635 6702
rect 17401 6699 17467 6702
rect 18873 6762 18939 6765
rect 18873 6760 24916 6762
rect 18873 6704 18878 6760
rect 18934 6704 24916 6760
rect 18873 6702 24916 6704
rect 18873 6699 18939 6702
rect 24856 6626 24916 6702
rect 27520 6626 28000 6656
rect 24856 6566 28000 6626
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6566
rect 24277 6495 24597 6496
rect 6085 6218 6151 6221
rect 16205 6218 16271 6221
rect 6085 6216 16271 6218
rect 6085 6160 6090 6216
rect 6146 6160 16210 6216
rect 16266 6160 16271 6216
rect 6085 6158 16271 6160
rect 6085 6155 6151 6158
rect 16205 6155 16271 6158
rect 22921 6218 22987 6221
rect 24117 6218 24183 6221
rect 22921 6216 24183 6218
rect 22921 6160 22926 6216
rect 22982 6160 24122 6216
rect 24178 6160 24183 6216
rect 22921 6158 24183 6160
rect 22921 6155 22987 6158
rect 24117 6155 24183 6158
rect 11605 6082 11671 6085
rect 14641 6082 14707 6085
rect 11605 6080 14707 6082
rect 11605 6024 11610 6080
rect 11666 6024 14646 6080
rect 14702 6024 14707 6080
rect 11605 6022 14707 6024
rect 11605 6019 11671 6022
rect 14641 6019 14707 6022
rect 20345 6082 20411 6085
rect 27520 6082 28000 6112
rect 20345 6080 28000 6082
rect 20345 6024 20350 6080
rect 20406 6024 28000 6080
rect 20345 6022 28000 6024
rect 20345 6019 20411 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 20345 5946 20411 5949
rect 20897 5946 20963 5949
rect 25497 5946 25563 5949
rect 20345 5944 25563 5946
rect 20345 5888 20350 5944
rect 20406 5888 20902 5944
rect 20958 5888 25502 5944
rect 25558 5888 25563 5944
rect 20345 5886 25563 5888
rect 20345 5883 20411 5886
rect 20897 5883 20963 5886
rect 25497 5883 25563 5886
rect 7373 5810 7439 5813
rect 12249 5810 12315 5813
rect 7373 5808 12315 5810
rect 7373 5752 7378 5808
rect 7434 5752 12254 5808
rect 12310 5752 12315 5808
rect 7373 5750 12315 5752
rect 7373 5747 7439 5750
rect 12249 5747 12315 5750
rect 12893 5810 12959 5813
rect 19517 5810 19583 5813
rect 22921 5810 22987 5813
rect 12893 5808 22987 5810
rect 12893 5752 12898 5808
rect 12954 5752 19522 5808
rect 19578 5752 22926 5808
rect 22982 5752 22987 5808
rect 12893 5750 22987 5752
rect 12893 5747 12959 5750
rect 19517 5747 19583 5750
rect 22921 5747 22987 5750
rect 23105 5810 23171 5813
rect 24025 5810 24091 5813
rect 23105 5808 24091 5810
rect 23105 5752 23110 5808
rect 23166 5752 24030 5808
rect 24086 5752 24091 5808
rect 23105 5750 24091 5752
rect 23105 5747 23171 5750
rect 24025 5747 24091 5750
rect 14181 5674 14247 5677
rect 23197 5674 23263 5677
rect 14181 5672 23263 5674
rect 14181 5616 14186 5672
rect 14242 5616 23202 5672
rect 23258 5616 23263 5672
rect 14181 5614 23263 5616
rect 14181 5611 14247 5614
rect 23197 5611 23263 5614
rect 23982 5614 24778 5674
rect 15837 5538 15903 5541
rect 23982 5538 24042 5614
rect 15837 5536 24042 5538
rect 15837 5480 15842 5536
rect 15898 5480 24042 5536
rect 15837 5478 24042 5480
rect 24718 5538 24778 5614
rect 25497 5538 25563 5541
rect 24718 5536 25563 5538
rect 24718 5480 25502 5536
rect 25558 5480 25563 5536
rect 24718 5478 25563 5480
rect 15837 5475 15903 5478
rect 25497 5475 25563 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 17493 5402 17559 5405
rect 27520 5402 28000 5432
rect 17493 5400 22018 5402
rect 17493 5344 17498 5400
rect 17554 5344 22018 5400
rect 17493 5342 22018 5344
rect 17493 5339 17559 5342
rect 11329 5266 11395 5269
rect 21817 5266 21883 5269
rect 11329 5264 21883 5266
rect 11329 5208 11334 5264
rect 11390 5208 21822 5264
rect 21878 5208 21883 5264
rect 11329 5206 21883 5208
rect 21958 5266 22018 5342
rect 24672 5342 28000 5402
rect 24672 5266 24732 5342
rect 27520 5312 28000 5342
rect 21958 5232 22064 5266
rect 22142 5232 24732 5266
rect 21958 5206 24732 5232
rect 11329 5203 11395 5206
rect 21817 5203 21883 5206
rect 22004 5172 22202 5206
rect 9489 5130 9555 5133
rect 12433 5130 12499 5133
rect 9489 5128 12499 5130
rect 9489 5072 9494 5128
rect 9550 5072 12438 5128
rect 12494 5072 12499 5128
rect 9489 5070 12499 5072
rect 9489 5067 9555 5070
rect 12433 5067 12499 5070
rect 17033 5130 17099 5133
rect 24945 5130 25011 5133
rect 17033 5128 20132 5130
rect 17033 5072 17038 5128
rect 17094 5072 20132 5128
rect 17033 5070 20132 5072
rect 17033 5067 17099 5070
rect 12709 4994 12775 4997
rect 19149 4994 19215 4997
rect 19425 4994 19491 4997
rect 12709 4992 19491 4994
rect 12709 4936 12714 4992
rect 12770 4936 19154 4992
rect 19210 4936 19430 4992
rect 19486 4936 19491 4992
rect 12709 4934 19491 4936
rect 12709 4931 12775 4934
rect 19149 4931 19215 4934
rect 19425 4931 19491 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 20072 4858 20132 5070
rect 23246 5128 25011 5130
rect 23246 5072 24950 5128
rect 25006 5072 25011 5128
rect 23246 5070 25011 5072
rect 20805 4994 20871 4997
rect 23105 4994 23171 4997
rect 20805 4992 23171 4994
rect 20805 4936 20810 4992
rect 20866 4936 23110 4992
rect 23166 4936 23171 4992
rect 20805 4934 23171 4936
rect 20805 4931 20871 4934
rect 23105 4931 23171 4934
rect 23246 4858 23306 5070
rect 24945 5067 25011 5070
rect 23381 4994 23447 4997
rect 24669 4994 24735 4997
rect 23381 4992 24735 4994
rect 23381 4936 23386 4992
rect 23442 4936 24674 4992
rect 24730 4936 24735 4992
rect 23381 4934 24735 4936
rect 23381 4931 23447 4934
rect 24669 4931 24735 4934
rect 27520 4858 28000 4888
rect 20072 4798 23306 4858
rect 24856 4798 28000 4858
rect 3509 4586 3575 4589
rect 12065 4586 12131 4589
rect 3509 4584 12131 4586
rect 3509 4528 3514 4584
rect 3570 4528 12070 4584
rect 12126 4528 12131 4584
rect 3509 4526 12131 4528
rect 3509 4523 3575 4526
rect 12065 4523 12131 4526
rect 15009 4586 15075 4589
rect 15653 4586 15719 4589
rect 24856 4586 24916 4798
rect 27520 4768 28000 4798
rect 15009 4584 24916 4586
rect 15009 4528 15014 4584
rect 15070 4528 15658 4584
rect 15714 4528 24916 4584
rect 15009 4526 24916 4528
rect 15009 4523 15075 4526
rect 15653 4523 15719 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 18413 4314 18479 4317
rect 23105 4314 23171 4317
rect 18413 4312 23171 4314
rect 18413 4256 18418 4312
rect 18474 4256 23110 4312
rect 23166 4256 23171 4312
rect 18413 4254 23171 4256
rect 18413 4251 18479 4254
rect 23105 4251 23171 4254
rect 24669 4314 24735 4317
rect 27520 4314 28000 4344
rect 24669 4312 28000 4314
rect 24669 4256 24674 4312
rect 24730 4256 28000 4312
rect 24669 4254 28000 4256
rect 24669 4251 24735 4254
rect 27520 4224 28000 4254
rect 2865 4178 2931 4181
rect 9489 4178 9555 4181
rect 2865 4176 9555 4178
rect 2865 4120 2870 4176
rect 2926 4120 9494 4176
rect 9550 4120 9555 4176
rect 2865 4118 9555 4120
rect 2865 4115 2931 4118
rect 9489 4115 9555 4118
rect 18965 4178 19031 4181
rect 24025 4178 24091 4181
rect 18965 4176 24091 4178
rect 18965 4120 18970 4176
rect 19026 4120 24030 4176
rect 24086 4120 24091 4176
rect 18965 4118 24091 4120
rect 18965 4115 19031 4118
rect 24025 4115 24091 4118
rect 13077 4042 13143 4045
rect 19425 4042 19491 4045
rect 13077 4040 19491 4042
rect 13077 3984 13082 4040
rect 13138 3984 19430 4040
rect 19486 3984 19491 4040
rect 13077 3982 19491 3984
rect 13077 3979 13143 3982
rect 19425 3979 19491 3982
rect 19885 4042 19951 4045
rect 22369 4042 22435 4045
rect 19885 4040 22435 4042
rect 19885 3984 19890 4040
rect 19946 3984 22374 4040
rect 22430 3984 22435 4040
rect 19885 3982 22435 3984
rect 19885 3979 19951 3982
rect 22369 3979 22435 3982
rect 16297 3906 16363 3909
rect 19149 3906 19215 3909
rect 16297 3904 19215 3906
rect 16297 3848 16302 3904
rect 16358 3848 19154 3904
rect 19210 3848 19215 3904
rect 16297 3846 19215 3848
rect 16297 3843 16363 3846
rect 19149 3843 19215 3846
rect 20069 3906 20135 3909
rect 25037 3906 25103 3909
rect 20069 3904 25103 3906
rect 20069 3848 20074 3904
rect 20130 3848 25042 3904
rect 25098 3848 25103 3904
rect 20069 3846 25103 3848
rect 20069 3843 20135 3846
rect 25037 3843 25103 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 10961 3770 11027 3773
rect 19425 3770 19491 3773
rect 10961 3768 19491 3770
rect 10961 3712 10966 3768
rect 11022 3712 19430 3768
rect 19486 3712 19491 3768
rect 10961 3710 19491 3712
rect 10961 3707 11027 3710
rect 19425 3707 19491 3710
rect 25773 3770 25839 3773
rect 27520 3770 28000 3800
rect 25773 3768 28000 3770
rect 25773 3712 25778 3768
rect 25834 3712 28000 3768
rect 25773 3710 28000 3712
rect 25773 3707 25839 3710
rect 27520 3680 28000 3710
rect 9397 3634 9463 3637
rect 14181 3634 14247 3637
rect 9397 3632 14247 3634
rect 9397 3576 9402 3632
rect 9458 3576 14186 3632
rect 14242 3576 14247 3632
rect 9397 3574 14247 3576
rect 9397 3571 9463 3574
rect 14181 3571 14247 3574
rect 18413 3634 18479 3637
rect 23657 3634 23723 3637
rect 18413 3632 23723 3634
rect 18413 3576 18418 3632
rect 18474 3576 23662 3632
rect 23718 3576 23723 3632
rect 18413 3574 23723 3576
rect 18413 3571 18479 3574
rect 23657 3571 23723 3574
rect 8477 3498 8543 3501
rect 19149 3498 19215 3501
rect 8477 3496 19215 3498
rect 8477 3440 8482 3496
rect 8538 3440 19154 3496
rect 19210 3440 19215 3496
rect 8477 3438 19215 3440
rect 8477 3435 8543 3438
rect 19149 3435 19215 3438
rect 20161 3498 20227 3501
rect 24209 3498 24275 3501
rect 20161 3496 24275 3498
rect 20161 3440 20166 3496
rect 20222 3440 24214 3496
rect 24270 3440 24275 3496
rect 20161 3438 24275 3440
rect 20161 3435 20227 3438
rect 24209 3435 24275 3438
rect 15929 3362 15995 3365
rect 21449 3362 21515 3365
rect 15929 3360 21515 3362
rect 15929 3304 15934 3360
rect 15990 3304 21454 3360
rect 21510 3304 21515 3360
rect 15929 3302 21515 3304
rect 15929 3299 15995 3302
rect 21449 3299 21515 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 25129 3226 25195 3229
rect 27520 3226 28000 3256
rect 25129 3224 28000 3226
rect 25129 3168 25134 3224
rect 25190 3168 28000 3224
rect 25129 3166 28000 3168
rect 25129 3163 25195 3166
rect 27520 3136 28000 3166
rect 8569 3090 8635 3093
rect 17769 3090 17835 3093
rect 8569 3088 17835 3090
rect 8569 3032 8574 3088
rect 8630 3032 17774 3088
rect 17830 3032 17835 3088
rect 8569 3030 17835 3032
rect 8569 3027 8635 3030
rect 17769 3027 17835 3030
rect 18413 3090 18479 3093
rect 22277 3090 22343 3093
rect 25313 3090 25379 3093
rect 18413 3088 22202 3090
rect 18413 3032 18418 3088
rect 18474 3032 22202 3088
rect 18413 3030 22202 3032
rect 18413 3027 18479 3030
rect 7097 2954 7163 2957
rect 11789 2954 11855 2957
rect 7097 2952 11855 2954
rect 7097 2896 7102 2952
rect 7158 2896 11794 2952
rect 11850 2896 11855 2952
rect 7097 2894 11855 2896
rect 7097 2891 7163 2894
rect 11789 2891 11855 2894
rect 15101 2954 15167 2957
rect 17861 2954 17927 2957
rect 15101 2952 17927 2954
rect 15101 2896 15106 2952
rect 15162 2896 17866 2952
rect 17922 2896 17927 2952
rect 15101 2894 17927 2896
rect 15101 2891 15167 2894
rect 17861 2891 17927 2894
rect 18137 2954 18203 2957
rect 20529 2954 20595 2957
rect 21357 2954 21423 2957
rect 22001 2954 22067 2957
rect 18137 2952 22067 2954
rect 18137 2896 18142 2952
rect 18198 2896 20534 2952
rect 20590 2896 21362 2952
rect 21418 2896 22006 2952
rect 22062 2896 22067 2952
rect 18137 2894 22067 2896
rect 22142 2954 22202 3030
rect 22277 3088 25379 3090
rect 22277 3032 22282 3088
rect 22338 3032 25318 3088
rect 25374 3032 25379 3088
rect 22277 3030 25379 3032
rect 22277 3027 22343 3030
rect 25313 3027 25379 3030
rect 25405 2954 25471 2957
rect 22142 2952 25471 2954
rect 22142 2896 25410 2952
rect 25466 2896 25471 2952
rect 22142 2894 25471 2896
rect 18137 2891 18203 2894
rect 20529 2891 20595 2894
rect 21357 2891 21423 2894
rect 22001 2891 22067 2894
rect 25405 2891 25471 2894
rect 21449 2818 21515 2821
rect 21633 2818 21699 2821
rect 23841 2818 23907 2821
rect 21449 2816 23907 2818
rect 21449 2760 21454 2816
rect 21510 2760 21638 2816
rect 21694 2760 23846 2816
rect 23902 2760 23907 2816
rect 21449 2758 23907 2760
rect 21449 2755 21515 2758
rect 21633 2755 21699 2758
rect 23841 2755 23907 2758
rect 25405 2818 25471 2821
rect 27521 2818 27587 2821
rect 25405 2816 27587 2818
rect 25405 2760 25410 2816
rect 25466 2760 27526 2816
rect 27582 2760 27587 2816
rect 25405 2758 27587 2760
rect 25405 2755 25471 2758
rect 27521 2755 27587 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 13353 2682 13419 2685
rect 16849 2682 16915 2685
rect 13353 2680 16915 2682
rect 13353 2624 13358 2680
rect 13414 2624 16854 2680
rect 16910 2624 16915 2680
rect 13353 2622 16915 2624
rect 13353 2619 13419 2622
rect 16849 2619 16915 2622
rect 8477 2546 8543 2549
rect 24853 2546 24919 2549
rect 8477 2544 24919 2546
rect 8477 2488 8482 2544
rect 8538 2488 24858 2544
rect 24914 2488 24919 2544
rect 8477 2486 24919 2488
rect 8477 2483 8543 2486
rect 24853 2483 24919 2486
rect 25037 2546 25103 2549
rect 27520 2546 28000 2576
rect 25037 2544 28000 2546
rect 25037 2488 25042 2544
rect 25098 2488 28000 2544
rect 25037 2486 28000 2488
rect 25037 2483 25103 2486
rect 27520 2456 28000 2486
rect 8753 2410 8819 2413
rect 18045 2410 18111 2413
rect 8753 2408 18111 2410
rect 8753 2352 8758 2408
rect 8814 2352 18050 2408
rect 18106 2352 18111 2408
rect 8753 2350 18111 2352
rect 8753 2347 8819 2350
rect 18045 2347 18111 2350
rect 8569 2274 8635 2277
rect 10685 2274 10751 2277
rect 8569 2272 10751 2274
rect 8569 2216 8574 2272
rect 8630 2216 10690 2272
rect 10746 2216 10751 2272
rect 8569 2214 10751 2216
rect 8569 2211 8635 2214
rect 10685 2211 10751 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 8661 2138 8727 2141
rect 10777 2138 10843 2141
rect 8661 2136 10843 2138
rect 8661 2080 8666 2136
rect 8722 2080 10782 2136
rect 10838 2080 10843 2136
rect 8661 2078 10843 2080
rect 8661 2075 8727 2078
rect 10777 2075 10843 2078
rect 10041 2002 10107 2005
rect 20437 2002 20503 2005
rect 10041 2000 20503 2002
rect 10041 1944 10046 2000
rect 10102 1944 20442 2000
rect 20498 1944 20503 2000
rect 10041 1942 20503 1944
rect 10041 1939 10107 1942
rect 20437 1939 20503 1942
rect 24669 2002 24735 2005
rect 27520 2002 28000 2032
rect 24669 2000 28000 2002
rect 24669 1944 24674 2000
rect 24730 1944 28000 2000
rect 24669 1942 28000 1944
rect 24669 1939 24735 1942
rect 27520 1912 28000 1942
rect 10041 1866 10107 1869
rect 23473 1866 23539 1869
rect 10041 1864 23539 1866
rect 10041 1808 10046 1864
rect 10102 1808 23478 1864
rect 23534 1808 23539 1864
rect 10041 1806 23539 1808
rect 10041 1803 10107 1806
rect 23473 1803 23539 1806
rect 4797 1730 4863 1733
rect 17585 1730 17651 1733
rect 4797 1728 17651 1730
rect 4797 1672 4802 1728
rect 4858 1672 17590 1728
rect 17646 1672 17651 1728
rect 4797 1670 17651 1672
rect 4797 1667 4863 1670
rect 17585 1667 17651 1670
rect 4153 1594 4219 1597
rect 15653 1594 15719 1597
rect 4153 1592 15719 1594
rect 4153 1536 4158 1592
rect 4214 1536 15658 1592
rect 15714 1536 15719 1592
rect 4153 1534 15719 1536
rect 4153 1531 4219 1534
rect 15653 1531 15719 1534
rect 21541 1594 21607 1597
rect 21541 1592 24962 1594
rect 21541 1536 21546 1592
rect 21602 1536 24962 1592
rect 21541 1534 24962 1536
rect 21541 1531 21607 1534
rect 19149 1458 19215 1461
rect 22645 1458 22711 1461
rect 19149 1456 22711 1458
rect 19149 1400 19154 1456
rect 19210 1400 22650 1456
rect 22706 1400 22711 1456
rect 19149 1398 22711 1400
rect 24902 1458 24962 1534
rect 27520 1458 28000 1488
rect 24902 1398 28000 1458
rect 19149 1395 19215 1398
rect 22645 1395 22711 1398
rect 27520 1368 28000 1398
rect 24761 914 24827 917
rect 27520 914 28000 944
rect 24761 912 28000 914
rect 24761 856 24766 912
rect 24822 856 28000 912
rect 24761 854 28000 856
rect 24761 851 24827 854
rect 27520 824 28000 854
rect 23841 370 23907 373
rect 27520 370 28000 400
rect 23841 368 28000 370
rect 23841 312 23846 368
rect 23902 312 28000 368
rect 23841 310 28000 312
rect 23841 307 23907 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 19380 23156 19444 23220
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 19380 20980 19444 21044
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19379 23220 19445 23221
rect 19379 23156 19380 23220
rect 19444 23156 19445 23220
rect 19379 23155 19445 23156
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 19382 21045 19442 23155
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19379 21044 19445 21045
rect 19379 20980 19380 21044
rect 19444 20980 19445 21044
rect 19379 20979 19445 20980
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _40_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7084 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1604681595
transform 1 0 6900 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_66
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68
timestamp 1604681595
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_70
timestamp 1604681595
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1604681595
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_87
timestamp 1604681595
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1604681595
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1604681595
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1604681595
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _80_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9476 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12604 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14168 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__90__A
timestamp 1604681595
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_144
timestamp 1604681595
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_134
timestamp 1604681595
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1604681595
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__88__A
timestamp 1604681595
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1604681595
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152
timestamp 1604681595
transform 1 0 15088 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1604681595
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_165
timestamp 1604681595
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_177
timestamp 1604681595
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_173
timestamp 1604681595
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1604681595
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1604681595
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1604681595
transform 1 0 16652 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1604681595
transform 1 0 17940 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1604681595
transform 1 0 17572 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1604681595
transform 1 0 20056 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1604681595
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_207
timestamp 1604681595
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604681595
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_210
timestamp 1604681595
transform 1 0 20424 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_227
timestamp 1604681595
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20516 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1604681595
transform 1 0 22632 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_230
timestamp 1604681595
transform 1 0 22264 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_235
timestamp 1604681595
transform 1 0 22724 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_231
timestamp 1604681595
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1604681595
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_258
timestamp 1604681595
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_254
timestamp 1604681595
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1604681595
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_266
timestamp 1604681595
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_262
timestamp 1604681595
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_270
timestamp 1604681595
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_274
timestamp 1604681595
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604681595
transform 1 0 6992 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67
timestamp 1604681595
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_71
timestamp 1604681595
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9936 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604681595
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11500 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_109
timestamp 1604681595
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _90_
timestamp 1604681595
transform 1 0 13984 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_132
timestamp 1604681595
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_136
timestamp 1604681595
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_144
timestamp 1604681595
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15916 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_148
timestamp 1604681595
transform 1 0 14720 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_158
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1604681595
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16468 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_2_186
timestamp 1604681595
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19136 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_205
timestamp 1604681595
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 21528 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21068 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20516 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_209
timestamp 1604681595
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1604681595
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_219
timestamp 1604681595
transform 1 0 21252 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1604681595
transform 1 0 23276 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_247
timestamp 1604681595
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_258
timestamp 1604681595
transform 1 0 24840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_262
timestamp 1604681595
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_266
timestamp 1604681595
transform 1 0 25576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_270
timestamp 1604681595
transform 1 0 25944 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_274
timestamp 1604681595
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8096 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_72
timestamp 1604681595
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9660 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_85
timestamp 1604681595
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1604681595
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12512 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_112
timestamp 1604681595
transform 1 0 11408 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14352 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_133
timestamp 1604681595
transform 1 0 13340 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_137
timestamp 1604681595
transform 1 0 13708 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_140
timestamp 1604681595
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15916 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_153
timestamp 1604681595
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1604681595
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_170
timestamp 1604681595
transform 1 0 16744 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21712 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_210
timestamp 1604681595
transform 1 0 20424 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_214
timestamp 1604681595
transform 1 0 20792 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_217
timestamp 1604681595
transform 1 0 21068 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_221
timestamp 1604681595
transform 1 0 21436 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23920 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23092 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_233
timestamp 1604681595
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_237
timestamp 1604681595
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_241
timestamp 1604681595
transform 1 0 23276 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_267
timestamp 1604681595
transform 1 0 25668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 26220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_271
timestamp 1604681595
transform 1 0 26036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_275
timestamp 1604681595
transform 1 0 26404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604681595
transform 1 0 8556 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_78
timestamp 1604681595
transform 1 0 8280 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604681595
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 11592 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_106 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_121
timestamp 1604681595
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_144
timestamp 1604681595
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_148
timestamp 1604681595
transform 1 0 14720 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17756 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_173
timestamp 1604681595
transform 1 0 17020 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_177
timestamp 1604681595
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19320 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_196
timestamp 1604681595
transform 1 0 19136 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_200
timestamp 1604681595
transform 1 0 19504 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_210
timestamp 1604681595
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1604681595
transform 1 0 21252 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_223
timestamp 1604681595
transform 1 0 21620 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_226
timestamp 1604681595
transform 1 0 21896 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23920 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_246
timestamp 1604681595
transform 1 0 23736 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1604681595
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24472 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 24288 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_263
timestamp 1604681595
transform 1 0 25300 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_267
timestamp 1604681595
transform 1 0 25668 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8648 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1604681595
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1604681595
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_109
timestamp 1604681595
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_105
timestamp 1604681595
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12604 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_5_144
timestamp 1604681595
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1604681595
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19320 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 18768 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_190
timestamp 1604681595
transform 1 0 18584 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_194
timestamp 1604681595
transform 1 0 18952 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_207
timestamp 1604681595
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 20884 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 21988 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_211
timestamp 1604681595
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_219
timestamp 1604681595
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_223
timestamp 1604681595
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1604681595
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604681595
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1604681595
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1604681595
transform 1 0 25392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_268
timestamp 1604681595
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_272
timestamp 1604681595
transform 1 0 26128 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_276
timestamp 1604681595
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_82
timestamp 1604681595
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1604681595
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_101
timestamp 1604681595
transform 1 0 10396 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_97
timestamp 1604681595
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_105
timestamp 1604681595
transform 1 0 10764 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_121
timestamp 1604681595
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_125
timestamp 1604681595
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 14168 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_138
timestamp 1604681595
transform 1 0 13800 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1604681595
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_136
timestamp 1604681595
transform 1 0 13616 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_145
timestamp 1604681595
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp 1604681595
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_150
timestamp 1604681595
transform 1 0 14904 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15180 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1604681595
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_162
timestamp 1604681595
transform 1 0 16008 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1604681595
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_166
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_170
timestamp 1604681595
transform 1 0 16744 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_169
timestamp 1604681595
transform 1 0 16652 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16744 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_194
timestamp 1604681595
transform 1 0 18952 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_190
timestamp 1604681595
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_193
timestamp 1604681595
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1604681595
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_207
timestamp 1604681595
transform 1 0 20148 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19320 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_211
timestamp 1604681595
transform 1 0 20516 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_210
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20792 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_229
timestamp 1604681595
transform 1 0 22172 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_224
timestamp 1604681595
transform 1 0 21712 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20976 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_7_235
timestamp 1604681595
transform 1 0 22724 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_237
timestamp 1604681595
transform 1 0 22908 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22356 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 22540 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604681595
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_241
timestamp 1604681595
transform 1 0 23276 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23460 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23644 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1604681595
transform 1 0 25208 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24656 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_254
timestamp 1604681595
transform 1 0 24472 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_258
timestamp 1604681595
transform 1 0 24840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_266
timestamp 1604681595
transform 1 0 25576 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1604681595
transform 1 0 25392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_268
timestamp 1604681595
transform 1 0 25760 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1604681595
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_276
timestamp 1604681595
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11776 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_107
timestamp 1604681595
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_111
timestamp 1604681595
transform 1 0 11316 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_115
timestamp 1604681595
transform 1 0 11684 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_139
timestamp 1604681595
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_143
timestamp 1604681595
transform 1 0 14260 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15640 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 14904 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_148
timestamp 1604681595
transform 1 0 14720 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1604681595
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17204 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17020 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_167
timestamp 1604681595
transform 1 0 16468 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_184
timestamp 1604681595
transform 1 0 18032 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_189
timestamp 1604681595
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_193
timestamp 1604681595
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1604681595
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_210
timestamp 1604681595
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23552 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_234
timestamp 1604681595
transform 1 0 22632 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_238
timestamp 1604681595
transform 1 0 23000 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1604681595
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_128
timestamp 1604681595
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_151
timestamp 1604681595
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_155
timestamp 1604681595
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_168
timestamp 1604681595
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_172
timestamp 1604681595
transform 1 0 16928 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_177
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18860 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1604681595
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_192
timestamp 1604681595
transform 1 0 18768 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_212
timestamp 1604681595
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_216
timestamp 1604681595
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_229
timestamp 1604681595
transform 1 0 22172 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_233
timestamp 1604681595
transform 1 0 22540 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1604681595
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604681595
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25208 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_254
timestamp 1604681595
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_258
timestamp 1604681595
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_268
timestamp 1604681595
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 26312 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_272
timestamp 1604681595
transform 1 0 26128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_276
timestamp 1604681595
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604681595
transform 1 0 9752 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_101
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_104
timestamp 1604681595
transform 1 0 10672 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_10_124
timestamp 1604681595
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13248 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_128
timestamp 1604681595
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1604681595
transform 1 0 14076 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 14720 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_147
timestamp 1604681595
transform 1 0 14628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17572 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1604681595
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1604681595
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_181
timestamp 1604681595
transform 1 0 17756 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_193
timestamp 1604681595
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1604681595
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_201
timestamp 1604681595
transform 1 0 19596 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_206
timestamp 1604681595
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21068 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_210
timestamp 1604681595
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_226
timestamp 1604681595
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 22632 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22448 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_230
timestamp 1604681595
transform 1 0 22264 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_243
timestamp 1604681595
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_247
timestamp 1604681595
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 25208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_260
timestamp 1604681595
transform 1 0 25024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_264
timestamp 1604681595
transform 1 0 25392 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_272
timestamp 1604681595
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_94
timestamp 1604681595
transform 1 0 9752 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1604681595
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12052 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1604681595
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13432 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_126
timestamp 1604681595
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_130
timestamp 1604681595
transform 1 0 13064 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_143
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15456 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 14996 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1604681595
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604681595
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19872 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 19596 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1604681595
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_197
timestamp 1604681595
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21804 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_223
timestamp 1604681595
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_227
timestamp 1604681595
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_231
timestamp 1604681595
transform 1 0 22356 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1604681595
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_254
timestamp 1604681595
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_258
timestamp 1604681595
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_268
timestamp 1604681595
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_272
timestamp 1604681595
transform 1 0 26128 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_276
timestamp 1604681595
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_99
timestamp 1604681595
transform 1 0 10212 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12052 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_111
timestamp 1604681595
transform 1 0 11316 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1604681595
transform 1 0 11684 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_142
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_146
timestamp 1604681595
transform 1 0 14536 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_150
timestamp 1604681595
transform 1 0 14904 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1604681595
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17204 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_167
timestamp 1604681595
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_171
timestamp 1604681595
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 19780 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19136 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1604681595
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_198
timestamp 1604681595
transform 1 0 19320 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_210
timestamp 1604681595
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23460 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22908 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_234
timestamp 1604681595
transform 1 0 22632 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_262
timestamp 1604681595
transform 1 0 25208 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1604681595
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_132
timestamp 1604681595
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_130
timestamp 1604681595
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_126
timestamp 1604681595
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13432 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1604681595
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1604681595
transform 1 0 15180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_158
timestamp 1604681595
transform 1 0 15640 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_159
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 15916 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16100 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_13_176
timestamp 1604681595
transform 1 0 17296 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_172
timestamp 1604681595
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_180
timestamp 1604681595
transform 1 0 17664 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_186
timestamp 1604681595
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_182
timestamp 1604681595
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18492 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_199
timestamp 1604681595
transform 1 0 19412 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_207
timestamp 1604681595
transform 1 0 20148 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_210
timestamp 1604681595
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1604681595
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1604681595
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_228
timestamp 1604681595
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_224
timestamp 1604681595
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21620 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_236
timestamp 1604681595
transform 1 0 22816 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_232
timestamp 1604681595
transform 1 0 22448 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_239
timestamp 1604681595
transform 1 0 23092 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_236
timestamp 1604681595
transform 1 0 22816 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22632 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 22908 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1604681595
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_246
timestamp 1604681595
transform 1 0 23736 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1604681595
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23920 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23276 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24472 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24288 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1604681595
transform 1 0 25392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_268
timestamp 1604681595
transform 1 0 25760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_272
timestamp 1604681595
transform 1 0 26128 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_276
timestamp 1604681595
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604681595
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 13708 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_135
timestamp 1604681595
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_144
timestamp 1604681595
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14720 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_171
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_167
timestamp 1604681595
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_203
timestamp 1604681595
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_207
timestamp 1604681595
transform 1 0 20148 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1604681595
transform 1 0 20792 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 21896 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21712 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_211
timestamp 1604681595
transform 1 0 20516 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1604681595
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1604681595
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_235
timestamp 1604681595
transform 1 0 22724 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1604681595
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_268
timestamp 1604681595
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_272
timestamp 1604681595
transform 1 0 26128 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604681595
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_129
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_137
timestamp 1604681595
transform 1 0 13708 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_160
timestamp 1604681595
transform 1 0 15824 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18308 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16652 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_178
timestamp 1604681595
transform 1 0 17480 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_186
timestamp 1604681595
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21344 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_210
timestamp 1604681595
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23828 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23644 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23276 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_243
timestamp 1604681595
transform 1 0 23460 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_266
timestamp 1604681595
transform 1 0 25576 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604681595
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_165
timestamp 1604681595
transform 1 0 16284 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1604681595
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_176
timestamp 1604681595
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1604681595
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 18400 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19412 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_191
timestamp 1604681595
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_195
timestamp 1604681595
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1604681595
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_222
timestamp 1604681595
transform 1 0 21528 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__87__A
timestamp 1604681595
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1604681595
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_268
timestamp 1604681595
transform 1 0 25760 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_276
timestamp 1604681595
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1604681595
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1604681595
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_162
timestamp 1604681595
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_166
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17112 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_180
timestamp 1604681595
transform 1 0 17664 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_194
timestamp 1604681595
transform 1 0 18952 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1604681595
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23460 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22816 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_234
timestamp 1604681595
transform 1 0 22632 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_238
timestamp 1604681595
transform 1 0 23000 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_242
timestamp 1604681595
transform 1 0 23368 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1604681595
transform 1 0 25208 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 24656 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_254
timestamp 1604681595
transform 1 0 24472 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1604681595
transform 1 0 24840 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_266
timestamp 1604681595
transform 1 0 25576 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1604681595
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1604681595
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1604681595
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 16284 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_159
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_162
timestamp 1604681595
transform 1 0 16008 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604681595
transform 1 0 18124 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_167
timestamp 1604681595
transform 1 0 16468 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_196
timestamp 1604681595
transform 1 0 19136 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_192
timestamp 1604681595
transform 1 0 18768 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_188
timestamp 1604681595
transform 1 0 18400 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1604681595
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18400 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_207
timestamp 1604681595
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_204
timestamp 1604681595
transform 1 0 19872 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_201
timestamp 1604681595
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19964 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19964 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_218
timestamp 1604681595
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_214
timestamp 1604681595
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_224
timestamp 1604681595
transform 1 0 21712 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_226
timestamp 1604681595
transform 1 0 21896 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1604681595
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_232
timestamp 1604681595
transform 1 0 22448 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_239
timestamp 1604681595
transform 1 0 23092 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_235
timestamp 1604681595
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22632 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_243
timestamp 1604681595
transform 1 0 23460 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_243
timestamp 1604681595
transform 1 0 23460 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23276 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23828 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_249
timestamp 1604681595
transform 1 0 24012 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 24564 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _89_
timestamp 1604681595
transform 1 0 25116 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__89__A
timestamp 1604681595
transform 1 0 25668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_253
timestamp 1604681595
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_265
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_259
timestamp 1604681595
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1604681595
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1604681595
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1604681595
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 19320 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_201
timestamp 1604681595
transform 1 0 19596 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 21252 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_213
timestamp 1604681595
transform 1 0 20700 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_222
timestamp 1604681595
transform 1 0 21528 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 22264 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23092 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_233
timestamp 1604681595
transform 1 0 22540 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_241
timestamp 1604681595
transform 1 0 23276 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 24564 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 25116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_259
timestamp 1604681595
transform 1 0 24932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_263
timestamp 1604681595
transform 1 0 25300 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_275
timestamp 1604681595
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_218
timestamp 1604681595
transform 1 0 21160 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_230
timestamp 1604681595
transform 1 0 22264 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_238
timestamp 1604681595
transform 1 0 23000 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_245
timestamp 1604681595
transform 1 0 23644 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1604681595
transform 1 0 24380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_259
timestamp 1604681595
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1604681595
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23828 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 25300 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_255
timestamp 1604681595
transform 1 0 24564 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_260
timestamp 1604681595
transform 1 0 25024 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_267
timestamp 1604681595
transform 1 0 25668 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_271
timestamp 1604681595
transform 1 0 26036 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23552 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_243
timestamp 1604681595
transform 1 0 23460 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_250
timestamp 1604681595
transform 1 0 24104 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 24840 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_262
timestamp 1604681595
transform 1 0 25208 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1604681595
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_147
timestamp 1604681595
transform 1 0 14628 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp 1604681595
transform 1 0 15180 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_156
timestamp 1604681595
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_168
timestamp 1604681595
transform 1 0 16560 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1604681595
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18768 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_190
timestamp 1604681595
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_194
timestamp 1604681595
transform 1 0 18952 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_206
timestamp 1604681595
transform 1 0 20056 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_218
timestamp 1604681595
transform 1 0 21160 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_230
timestamp 1604681595
transform 1 0 22264 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_242
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 24564 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_259
timestamp 1604681595
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_263
timestamp 1604681595
transform 1 0 25300 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1604681595
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_101
timestamp 1604681595
transform 1 0 10396 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1604681595
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13156 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_129
timestamp 1604681595
transform 1 0 12972 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_133
timestamp 1604681595
transform 1 0 13340 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_145
timestamp 1604681595
transform 1 0 14444 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 15824 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_160
timestamp 1604681595
transform 1 0 15824 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_157
timestamp 1604681595
transform 1 0 15548 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_164
timestamp 1604681595
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_172
timestamp 1604681595
transform 1 0 16928 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_184
timestamp 1604681595
transform 1 0 18032 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_168
timestamp 1604681595
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1604681595
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_196
timestamp 1604681595
transform 1 0 19136 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_208
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 24564 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_259
timestamp 1604681595
transform 1 0 24932 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_259
timestamp 1604681595
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_263
timestamp 1604681595
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1604681595
transform 1 0 26036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_275
timestamp 1604681595
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_259
timestamp 1604681595
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1604681595
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_106
timestamp 1604681595
transform 1 0 10856 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_111
timestamp 1604681595
transform 1 0 11316 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1604681595
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13156 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_137
timestamp 1604681595
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_141
timestamp 1604681595
transform 1 0 14076 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_153
timestamp 1604681595
transform 1 0 15180 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_161
timestamp 1604681595
transform 1 0 15916 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_164
timestamp 1604681595
transform 1 0 16192 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_176
timestamp 1604681595
transform 1 0 17296 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1604681595
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 11132 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_105
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_113
timestamp 1604681595
transform 1 0 11500 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_125
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_137
timestamp 1604681595
transform 1 0 13708 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16008 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1604681595
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_180
timestamp 1604681595
transform 1 0 17664 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_192
timestamp 1604681595
transform 1 0 18768 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_204
timestamp 1604681595
transform 1 0 19872 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_216
timestamp 1604681595
transform 1 0 20976 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604681595
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 24932 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 25484 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 24564 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_251
timestamp 1604681595
transform 1 0 24196 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_263
timestamp 1604681595
transform 1 0 25300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_267
timestamp 1604681595
transform 1 0 25668 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_275
timestamp 1604681595
transform 1 0 26404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21160 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_224
timestamp 1604681595
transform 1 0 21712 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_236
timestamp 1604681595
transform 1 0 22816 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_248
timestamp 1604681595
transform 1 0 23920 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 24564 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_254
timestamp 1604681595
transform 1 0 24472 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_259
timestamp 1604681595
transform 1 0 24932 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_271
timestamp 1604681595
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15916 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_159
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_163
timestamp 1604681595
transform 1 0 16100 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_160
timestamp 1604681595
transform 1 0 15824 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_175
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_167
timestamp 1604681595
transform 1 0 16468 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_179
timestamp 1604681595
transform 1 0 17572 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_191
timestamp 1604681595
transform 1 0 18676 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_203
timestamp 1604681595
transform 1 0 19780 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_211
timestamp 1604681595
transform 1 0 20516 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604681595
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_251
timestamp 1604681595
transform 1 0 24196 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 24564 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 24932 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 24564 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_267
timestamp 1604681595
transform 1 0 25668 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_263
timestamp 1604681595
transform 1 0 25300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 25484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_259
timestamp 1604681595
transform 1 0 24932 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_275
timestamp 1604681595
transform 1 0 26404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_271
timestamp 1604681595
transform 1 0 26036 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604681595
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_86
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_94
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_99
timestamp 1604681595
transform 1 0 10212 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_111
timestamp 1604681595
transform 1 0 11316 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_119
timestamp 1604681595
transform 1 0 12052 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13432 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14168 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_131
timestamp 1604681595
transform 1 0 13156 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_140
timestamp 1604681595
transform 1 0 13984 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_144
timestamp 1604681595
transform 1 0 14352 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 17020 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_168
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_172
timestamp 1604681595
transform 1 0 16928 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_175
timestamp 1604681595
transform 1 0 17204 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_253
timestamp 1604681595
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_259
timestamp 1604681595
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_263
timestamp 1604681595
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_275
timestamp 1604681595
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10028 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_103
timestamp 1604681595
transform 1 0 10580 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_115
timestamp 1604681595
transform 1 0 11684 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_127
timestamp 1604681595
transform 1 0 12788 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_139
timestamp 1604681595
transform 1 0 13892 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_151
timestamp 1604681595
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_166
timestamp 1604681595
transform 1 0 16376 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 17020 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_172
timestamp 1604681595
transform 1 0 16928 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1604681595
transform 1 0 17388 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_189
timestamp 1604681595
transform 1 0 18492 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1604681595
transform 1 0 19596 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1604681595
transform 1 0 20700 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604681595
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604681595
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_110
timestamp 1604681595
transform 1 0 11224 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1604681595
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1604681595
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1604681595
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1604681595
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1604681595
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1604681595
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23828 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1604681595
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_249
timestamp 1604681595
transform 1 0 24012 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 24564 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 25116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 25484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_259
timestamp 1604681595
transform 1 0 24932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_263
timestamp 1604681595
transform 1 0 25300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_267
timestamp 1604681595
transform 1 0 25668 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_275
timestamp 1604681595
transform 1 0 26404 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11776 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_105
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_113
timestamp 1604681595
transform 1 0 11500 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_122
timestamp 1604681595
transform 1 0 12328 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_134
timestamp 1604681595
transform 1 0 13432 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_146
timestamp 1604681595
transform 1 0 14536 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_152
timestamp 1604681595
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1604681595
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_178
timestamp 1604681595
transform 1 0 17480 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_186
timestamp 1604681595
transform 1 0 18216 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_198
timestamp 1604681595
transform 1 0 19320 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_210
timestamp 1604681595
transform 1 0 20424 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1604681595
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_239
timestamp 1604681595
transform 1 0 23092 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 24932 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_251
timestamp 1604681595
transform 1 0 24196 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1604681595
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604681595
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 10028 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_86
timestamp 1604681595
transform 1 0 9016 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_94
timestamp 1604681595
transform 1 0 9752 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_101
timestamp 1604681595
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_105
timestamp 1604681595
transform 1 0 10764 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_117
timestamp 1604681595
transform 1 0 11868 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_121
timestamp 1604681595
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 12788 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 13340 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_131
timestamp 1604681595
transform 1 0 13156 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1604681595
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1604681595
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_171
timestamp 1604681595
transform 1 0 16836 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1604681595
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_203
timestamp 1604681595
transform 1 0 19780 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604681595
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_215
timestamp 1604681595
transform 1 0 20884 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_227
timestamp 1604681595
transform 1 0 21988 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1604681595
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 23276 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_239
timestamp 1604681595
transform 1 0 23092 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1604681595
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_239
timestamp 1604681595
transform 1 0 23092 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_245
timestamp 1604681595
transform 1 0 23644 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_253
timestamp 1604681595
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_259
timestamp 1604681595
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_263
timestamp 1604681595
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_257
timestamp 1604681595
transform 1 0 24748 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_269
timestamp 1604681595
transform 1 0 25852 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_275
timestamp 1604681595
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1604681595
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 26882 0 26938 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 27526 0 27582 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 24490 27520 24546 28000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 4 nsew default input
rlabel metal2 s 17498 27520 17554 28000 6 ccff_head
port 5 nsew default input
rlabel metal3 s 0 14016 480 14136 6 ccff_tail
port 6 nsew default tristate
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_in[0]
port 7 nsew default input
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[10]
port 8 nsew default input
rlabel metal3 s 27520 11024 28000 11144 6 chanx_right_in[11]
port 9 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_in[12]
port 10 nsew default input
rlabel metal3 s 27520 12248 28000 12368 6 chanx_right_in[13]
port 11 nsew default input
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_in[14]
port 12 nsew default input
rlabel metal3 s 27520 13336 28000 13456 6 chanx_right_in[15]
port 13 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_in[16]
port 14 nsew default input
rlabel metal3 s 27520 14560 28000 14680 6 chanx_right_in[17]
port 15 nsew default input
rlabel metal3 s 27520 15104 28000 15224 6 chanx_right_in[18]
port 16 nsew default input
rlabel metal3 s 27520 15648 28000 15768 6 chanx_right_in[19]
port 17 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_in[1]
port 18 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[2]
port 19 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_in[3]
port 20 nsew default input
rlabel metal3 s 27520 7080 28000 7200 6 chanx_right_in[4]
port 21 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[5]
port 22 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[6]
port 23 nsew default input
rlabel metal3 s 27520 8848 28000 8968 6 chanx_right_in[7]
port 24 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_in[8]
port 25 nsew default input
rlabel metal3 s 27520 9936 28000 10056 6 chanx_right_in[9]
port 26 nsew default input
rlabel metal3 s 27520 16192 28000 16312 6 chanx_right_out[0]
port 27 nsew default tristate
rlabel metal3 s 27520 21904 28000 22024 6 chanx_right_out[10]
port 28 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[11]
port 29 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[12]
port 30 nsew default tristate
rlabel metal3 s 27520 23672 28000 23792 6 chanx_right_out[13]
port 31 nsew default tristate
rlabel metal3 s 27520 24216 28000 24336 6 chanx_right_out[14]
port 32 nsew default tristate
rlabel metal3 s 27520 24760 28000 24880 6 chanx_right_out[15]
port 33 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[16]
port 34 nsew default tristate
rlabel metal3 s 27520 25984 28000 26104 6 chanx_right_out[17]
port 35 nsew default tristate
rlabel metal3 s 27520 26528 28000 26648 6 chanx_right_out[18]
port 36 nsew default tristate
rlabel metal3 s 27520 27072 28000 27192 6 chanx_right_out[19]
port 37 nsew default tristate
rlabel metal3 s 27520 16736 28000 16856 6 chanx_right_out[1]
port 38 nsew default tristate
rlabel metal3 s 27520 17416 28000 17536 6 chanx_right_out[2]
port 39 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_out[3]
port 40 nsew default tristate
rlabel metal3 s 27520 18504 28000 18624 6 chanx_right_out[4]
port 41 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[5]
port 42 nsew default tristate
rlabel metal3 s 27520 19592 28000 19712 6 chanx_right_out[6]
port 43 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[7]
port 44 nsew default tristate
rlabel metal3 s 27520 20816 28000 20936 6 chanx_right_out[8]
port 45 nsew default tristate
rlabel metal3 s 27520 21360 28000 21480 6 chanx_right_out[9]
port 46 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_in[0]
port 47 nsew default input
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_in[10]
port 48 nsew default input
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_in[11]
port 49 nsew default input
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[12]
port 50 nsew default input
rlabel metal2 s 9310 0 9366 480 6 chany_bottom_in[13]
port 51 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_in[14]
port 52 nsew default input
rlabel metal2 s 10690 0 10746 480 6 chany_bottom_in[15]
port 53 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[16]
port 54 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[17]
port 55 nsew default input
rlabel metal2 s 12622 0 12678 480 6 chany_bottom_in[18]
port 56 nsew default input
rlabel metal2 s 13266 0 13322 480 6 chany_bottom_in[19]
port 57 nsew default input
rlabel metal2 s 1582 0 1638 480 6 chany_bottom_in[1]
port 58 nsew default input
rlabel metal2 s 2226 0 2282 480 6 chany_bottom_in[2]
port 59 nsew default input
rlabel metal2 s 2870 0 2926 480 6 chany_bottom_in[3]
port 60 nsew default input
rlabel metal2 s 3514 0 3570 480 6 chany_bottom_in[4]
port 61 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_in[5]
port 62 nsew default input
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[6]
port 63 nsew default input
rlabel metal2 s 5446 0 5502 480 6 chany_bottom_in[7]
port 64 nsew default input
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_in[8]
port 65 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[9]
port 66 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_out[0]
port 67 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[10]
port 68 nsew default tristate
rlabel metal2 s 21086 0 21142 480 6 chany_bottom_out[11]
port 69 nsew default tristate
rlabel metal2 s 21730 0 21786 480 6 chany_bottom_out[12]
port 70 nsew default tristate
rlabel metal2 s 22374 0 22430 480 6 chany_bottom_out[13]
port 71 nsew default tristate
rlabel metal2 s 23018 0 23074 480 6 chany_bottom_out[14]
port 72 nsew default tristate
rlabel metal2 s 23662 0 23718 480 6 chany_bottom_out[15]
port 73 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[16]
port 74 nsew default tristate
rlabel metal2 s 24950 0 25006 480 6 chany_bottom_out[17]
port 75 nsew default tristate
rlabel metal2 s 25594 0 25650 480 6 chany_bottom_out[18]
port 76 nsew default tristate
rlabel metal2 s 26238 0 26294 480 6 chany_bottom_out[19]
port 77 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[1]
port 78 nsew default tristate
rlabel metal2 s 15198 0 15254 480 6 chany_bottom_out[2]
port 79 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[3]
port 80 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[4]
port 81 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[5]
port 82 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_out[6]
port 83 nsew default tristate
rlabel metal2 s 18418 0 18474 480 6 chany_bottom_out[7]
port 84 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_bottom_out[8]
port 85 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[9]
port 86 nsew default tristate
rlabel metal2 s 3514 27520 3570 28000 6 prog_clk
port 87 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_34_
port 88 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_35_
port 89 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_36_
port 90 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 right_bottom_grid_pin_37_
port 91 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 right_bottom_grid_pin_38_
port 92 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 right_bottom_grid_pin_39_
port 93 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 right_bottom_grid_pin_40_
port 94 nsew default input
rlabel metal3 s 27520 4224 28000 4344 6 right_bottom_grid_pin_41_
port 95 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 right_top_grid_pin_1_
port 96 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 97 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 98 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
