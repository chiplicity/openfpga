magic
tech EFS8A
magscale 1 2
timestamp 1604441278
<< locali >>
rect 53717 142495 53751 142665
rect 51325 142087 51359 142257
rect 52153 142155 52187 142393
rect 91253 138619 91287 141305
rect 91345 138551 91379 141305
rect 92725 138551 92759 141305
rect 93771 138517 94013 138551
rect 97049 138415 97083 138585
rect 132653 134471 132687 143413
rect 163105 138619 163139 141305
rect 222721 124815 222755 127501
rect 132653 113663 132687 117777
rect 222813 107951 222847 110229
rect 54821 86123 54855 90237
rect 132377 88775 132411 95745
rect 54821 76467 54855 79221
rect 36053 68715 36087 68817
rect 49393 68783 49427 69701
rect 96773 68715 96807 69769
rect 99567 68613 99659 68647
rect 99625 68511 99659 68613
rect 110055 68477 110239 68511
rect 110205 68375 110239 68477
rect 116185 68103 116219 68341
rect 124741 68103 124775 68273
rect 222537 28187 222571 37741
<< viali >>
rect 132653 143413 132687 143447
rect 53717 142665 53751 142699
rect 53717 142461 53751 142495
rect 52153 142393 52187 142427
rect 51325 142257 51359 142291
rect 52153 142121 52187 142155
rect 51325 142053 51359 142087
rect 91253 141305 91287 141339
rect 91253 138585 91287 138619
rect 91345 141305 91379 141339
rect 91345 138517 91379 138551
rect 92725 141305 92759 141339
rect 97049 138585 97083 138619
rect 92725 138517 92759 138551
rect 93737 138517 93771 138551
rect 94013 138517 94047 138551
rect 97049 138381 97083 138415
rect 163105 141305 163139 141339
rect 163105 138585 163139 138619
rect 132653 134437 132687 134471
rect 222721 127501 222755 127535
rect 222721 124781 222755 124815
rect 132653 117777 132687 117811
rect 132653 113629 132687 113663
rect 222813 110229 222847 110263
rect 222813 107917 222847 107951
rect 132377 95745 132411 95779
rect 54821 90237 54855 90271
rect 132377 88741 132411 88775
rect 54821 86089 54855 86123
rect 54821 79221 54855 79255
rect 54821 76433 54855 76467
rect 96773 69769 96807 69803
rect 49393 69701 49427 69735
rect 36053 68817 36087 68851
rect 49393 68749 49427 68783
rect 36053 68681 36087 68715
rect 96773 68681 96807 68715
rect 99533 68613 99567 68647
rect 99625 68477 99659 68511
rect 110021 68477 110055 68511
rect 110205 68341 110239 68375
rect 116185 68341 116219 68375
rect 116185 68069 116219 68103
rect 124741 68273 124775 68307
rect 124741 68069 124775 68103
rect 222537 37741 222571 37775
rect 222537 28153 222571 28187
<< metal1 >>
rect 23526 244860 23532 244912
rect 23584 244900 23590 244912
rect 70538 244900 70544 244912
rect 23584 244872 70544 244900
rect 23584 244860 23590 244872
rect 70538 244860 70544 244872
rect 70596 244860 70602 244912
rect 105222 244860 105228 244912
rect 105280 244900 105286 244912
rect 149658 244900 149664 244912
rect 105280 244872 149664 244900
rect 105280 244860 105286 244872
rect 149658 244860 149664 244872
rect 149716 244860 149722 244912
rect 50758 244792 50764 244844
rect 50816 244832 50822 244844
rect 142390 244832 142396 244844
rect 50816 244804 142396 244832
rect 50816 244792 50822 244804
rect 142390 244792 142396 244804
rect 142448 244792 142454 244844
rect 157478 244792 157484 244844
rect 157536 244832 157542 244844
rect 159778 244832 159784 244844
rect 157536 244804 159784 244832
rect 157536 244792 157542 244804
rect 159778 244792 159784 244804
rect 159836 244792 159842 244844
rect 85626 242412 85632 242464
rect 85684 242412 85690 242464
rect 85644 242180 85672 242412
rect 132546 242180 132552 242192
rect 85644 242152 132552 242180
rect 132546 242140 132552 242152
rect 132604 242140 132610 242192
rect 165298 242140 165304 242192
rect 165356 242180 165362 242192
rect 214242 242180 214248 242192
rect 165356 242152 214248 242180
rect 165356 242140 165362 242152
rect 214242 242140 214248 242152
rect 214300 242140 214306 242192
rect 93354 242072 93360 242124
rect 93412 242112 93418 242124
rect 187010 242112 187016 242124
rect 93412 242084 187016 242112
rect 93412 242072 93418 242084
rect 187010 242072 187016 242084
rect 187068 242072 187074 242124
rect 167782 229764 167788 229816
rect 167840 229804 167846 229816
rect 168518 229804 168524 229816
rect 167840 229776 168524 229804
rect 167840 229764 167846 229776
rect 168518 229764 168524 229776
rect 168576 229764 168582 229816
rect 207250 223372 207256 223424
rect 207308 223412 207314 223424
rect 223074 223412 223080 223424
rect 207308 223384 223080 223412
rect 207308 223372 207314 223384
rect 223074 223372 223080 223384
rect 223132 223372 223138 223424
rect 170082 222760 170088 222812
rect 170140 222800 170146 222812
rect 207250 222800 207256 222812
rect 170140 222772 207256 222800
rect 170140 222760 170146 222772
rect 207250 222760 207256 222772
rect 207308 222760 207314 222812
rect 71274 217932 71280 217984
rect 71332 217972 71338 217984
rect 71332 217944 98460 217972
rect 71332 217932 71338 217944
rect 98432 217916 98460 217944
rect 143678 217932 143684 217984
rect 143736 217972 143742 217984
rect 170082 217972 170088 217984
rect 143736 217944 170088 217972
rect 143736 217932 143742 217944
rect 170082 217932 170088 217944
rect 170140 217932 170146 217984
rect 46526 217864 46532 217916
rect 46584 217904 46590 217916
rect 98230 217904 98236 217916
rect 46584 217876 98236 217904
rect 46584 217864 46590 217876
rect 98230 217864 98236 217876
rect 98288 217864 98294 217916
rect 98414 217864 98420 217916
rect 98472 217904 98478 217916
rect 109270 217904 109276 217916
rect 98472 217876 109276 217904
rect 98472 217864 98478 217876
rect 109270 217864 109276 217876
rect 109328 217864 109334 217916
rect 118838 217864 118844 217916
rect 118896 217904 118902 217916
rect 169990 217904 169996 217916
rect 118896 217876 169996 217904
rect 118896 217864 118902 217876
rect 169990 217864 169996 217876
rect 170048 217864 170054 217916
rect 109270 217252 109276 217304
rect 109328 217292 109334 217304
rect 143678 217292 143684 217304
rect 109328 217264 143684 217292
rect 109328 217252 109334 217264
rect 143678 217252 143684 217264
rect 143736 217252 143742 217304
rect 37234 217184 37240 217236
rect 37292 217224 37298 217236
rect 71274 217224 71280 217236
rect 37292 217196 71280 217224
rect 37292 217184 37298 217196
rect 71274 217184 71280 217196
rect 71332 217184 71338 217236
rect 79370 217184 79376 217236
rect 79428 217224 79434 217236
rect 127762 217224 127768 217236
rect 79428 217196 127768 217224
rect 79428 217184 79434 217196
rect 127762 217184 127768 217196
rect 127820 217184 127826 217236
rect 81762 216572 81768 216624
rect 81820 216612 81826 216624
rect 93998 216612 94004 216624
rect 81820 216584 94004 216612
rect 81820 216572 81826 216584
rect 93998 216572 94004 216584
rect 94056 216572 94062 216624
rect 158582 216572 158588 216624
rect 158640 216612 158646 216624
rect 167230 216612 167236 216624
rect 158640 216584 167236 216612
rect 158640 216572 158646 216584
rect 167230 216572 167236 216584
rect 167288 216572 167294 216624
rect 91790 216504 91796 216556
rect 91848 216544 91854 216556
rect 102370 216544 102376 216556
rect 91848 216516 102376 216544
rect 91848 216504 91854 216516
rect 102370 216504 102376 216516
rect 102428 216504 102434 216556
rect 164102 216504 164108 216556
rect 164160 216544 164166 216556
rect 174222 216544 174228 216556
rect 164160 216516 174228 216544
rect 164160 216504 164166 216516
rect 174222 216504 174228 216516
rect 174280 216504 174286 216556
rect 86914 216436 86920 216488
rect 86972 216476 86978 216488
rect 98322 216476 98328 216488
rect 86972 216448 98328 216476
rect 86972 216436 86978 216448
rect 98322 216436 98328 216448
rect 98380 216436 98386 216488
rect 154074 216436 154080 216488
rect 154132 216476 154138 216488
rect 166034 216476 166040 216488
rect 154132 216448 166040 216476
rect 154132 216436 154138 216448
rect 166034 216436 166040 216448
rect 166092 216436 166098 216488
rect 62534 215756 62540 215808
rect 62592 215796 62598 215808
rect 71826 215796 71832 215808
rect 62592 215768 71832 215796
rect 62592 215756 62598 215768
rect 71826 215756 71832 215768
rect 71884 215756 71890 215808
rect 135398 215756 135404 215808
rect 135456 215796 135462 215808
rect 143770 215796 143776 215808
rect 135456 215768 143776 215796
rect 135456 215756 135462 215768
rect 143770 215756 143776 215768
rect 143828 215756 143834 215808
rect 100990 214600 100996 214652
rect 101048 214640 101054 214652
rect 102370 214640 102376 214652
rect 101048 214612 102376 214640
rect 101048 214600 101054 214612
rect 102370 214600 102376 214612
rect 102428 214600 102434 214652
rect 62626 214464 62632 214516
rect 62684 214504 62690 214516
rect 65018 214504 65024 214516
rect 62684 214476 65024 214504
rect 62684 214464 62690 214476
rect 65018 214464 65024 214476
rect 65076 214464 65082 214516
rect 135398 214464 135404 214516
rect 135456 214504 135462 214516
rect 136778 214504 136784 214516
rect 135456 214476 136784 214504
rect 135456 214464 135462 214476
rect 136778 214464 136784 214476
rect 136836 214464 136842 214516
rect 171830 213988 171836 214040
rect 171888 214028 171894 214040
rect 174038 214028 174044 214040
rect 171888 214000 174044 214028
rect 171888 213988 171894 214000
rect 174038 213988 174044 214000
rect 174096 213988 174102 214040
rect 100990 213308 100996 213360
rect 101048 213348 101054 213360
rect 102370 213348 102376 213360
rect 101048 213320 102376 213348
rect 101048 213308 101054 213320
rect 102370 213308 102376 213320
rect 102428 213308 102434 213360
rect 135030 213308 135036 213360
rect 135088 213348 135094 213360
rect 136778 213348 136784 213360
rect 135088 213320 136784 213348
rect 135088 213308 135094 213320
rect 136778 213308 136784 213320
rect 136836 213308 136842 213360
rect 62534 213240 62540 213292
rect 62592 213280 62598 213292
rect 65018 213280 65024 213292
rect 62592 213252 65024 213280
rect 62592 213240 62598 213252
rect 65018 213240 65024 213252
rect 65076 213240 65082 213292
rect 102462 213144 102468 213156
rect 102296 213116 102468 213144
rect 63730 213036 63736 213088
rect 63788 213076 63794 213088
rect 66214 213076 66220 213088
rect 63788 213048 66220 213076
rect 63788 213036 63794 213048
rect 66214 213036 66220 213048
rect 66272 213036 66278 213088
rect 100530 213036 100536 213088
rect 100588 213076 100594 213088
rect 102296 213076 102324 213116
rect 102462 213104 102468 213116
rect 102520 213104 102526 213156
rect 135398 213104 135404 213156
rect 135456 213144 135462 213156
rect 174222 213144 174228 213156
rect 135456 213116 135536 213144
rect 135456 213104 135462 213116
rect 100588 213048 102324 213076
rect 135508 213076 135536 213116
rect 172768 213116 174228 213144
rect 136870 213076 136876 213088
rect 135508 213048 136876 213076
rect 100588 213036 100594 213048
rect 136870 213036 136876 213048
rect 136928 213036 136934 213088
rect 172658 213036 172664 213088
rect 172716 213076 172722 213088
rect 172768 213076 172796 213116
rect 174222 213104 174228 213116
rect 174280 213104 174286 213156
rect 172716 213048 172796 213076
rect 172716 213036 172722 213048
rect 171738 212968 171744 213020
rect 171796 213008 171802 213020
rect 174038 213008 174044 213020
rect 171796 212980 174044 213008
rect 171796 212968 171802 212980
rect 174038 212968 174044 212980
rect 174096 212968 174102 213020
rect 101082 212220 101088 212272
rect 101140 212260 101146 212272
rect 102370 212260 102376 212272
rect 101140 212232 102376 212260
rect 101140 212220 101146 212232
rect 102370 212220 102376 212232
rect 102428 212220 102434 212272
rect 134662 212084 134668 212136
rect 134720 212124 134726 212136
rect 136962 212124 136968 212136
rect 134720 212096 136968 212124
rect 134720 212084 134726 212096
rect 136962 212084 136968 212096
rect 137020 212084 137026 212136
rect 100990 211880 100996 211932
rect 101048 211920 101054 211932
rect 102370 211920 102376 211932
rect 101048 211892 102376 211920
rect 101048 211880 101054 211892
rect 102370 211880 102376 211892
rect 102428 211880 102434 211932
rect 62626 211744 62632 211796
rect 62684 211784 62690 211796
rect 65018 211784 65024 211796
rect 62684 211756 65024 211784
rect 62684 211744 62690 211756
rect 65018 211744 65024 211756
rect 65076 211744 65082 211796
rect 134294 211744 134300 211796
rect 134352 211784 134358 211796
rect 136870 211784 136876 211796
rect 134352 211756 136876 211784
rect 134352 211744 134358 211756
rect 136870 211744 136876 211756
rect 136928 211744 136934 211796
rect 62350 211676 62356 211728
rect 62408 211716 62414 211728
rect 64926 211716 64932 211728
rect 62408 211688 64932 211716
rect 62408 211676 62414 211688
rect 64926 211676 64932 211688
rect 64984 211676 64990 211728
rect 174222 211716 174228 211728
rect 172768 211688 174228 211716
rect 172658 211608 172664 211660
rect 172716 211648 172722 211660
rect 172768 211648 172796 211688
rect 174222 211676 174228 211688
rect 174280 211676 174286 211728
rect 172716 211620 172796 211648
rect 172716 211608 172722 211620
rect 172566 211404 172572 211456
rect 172624 211444 172630 211456
rect 174038 211444 174044 211456
rect 172624 211416 174044 211444
rect 172624 211404 172630 211416
rect 174038 211404 174044 211416
rect 174096 211404 174102 211456
rect 62626 211064 62632 211116
rect 62684 211104 62690 211116
rect 65478 211104 65484 211116
rect 62684 211076 65484 211104
rect 62684 211064 62690 211076
rect 65478 211064 65484 211076
rect 65536 211064 65542 211116
rect 171830 210724 171836 210776
rect 171888 210764 171894 210776
rect 174130 210764 174136 210776
rect 171888 210736 174136 210764
rect 171888 210724 171894 210736
rect 174130 210724 174136 210736
rect 174188 210724 174194 210776
rect 62626 210384 62632 210436
rect 62684 210424 62690 210436
rect 65018 210424 65024 210436
rect 62684 210396 65024 210424
rect 62684 210384 62690 210396
rect 65018 210384 65024 210396
rect 65076 210384 65082 210436
rect 207894 210316 207900 210368
rect 207952 210356 207958 210368
rect 223534 210356 223540 210368
rect 207952 210328 223540 210356
rect 207952 210316 207958 210328
rect 223534 210316 223540 210328
rect 223592 210316 223598 210368
rect 171922 209636 171928 209688
rect 171980 209676 171986 209688
rect 174130 209676 174136 209688
rect 171980 209648 174136 209676
rect 171980 209636 171986 209648
rect 174130 209636 174136 209648
rect 174188 209636 174194 209688
rect 62626 209500 62632 209552
rect 62684 209540 62690 209552
rect 65478 209540 65484 209552
rect 62684 209512 65484 209540
rect 62684 209500 62690 209512
rect 65478 209500 65484 209512
rect 65536 209500 65542 209552
rect 62718 209024 62724 209076
rect 62776 209064 62782 209076
rect 65018 209064 65024 209076
rect 62776 209036 65024 209064
rect 62776 209024 62782 209036
rect 65018 209024 65024 209036
rect 65076 209024 65082 209076
rect 135306 209024 135312 209076
rect 135364 209064 135370 209076
rect 137698 209064 137704 209076
rect 135364 209036 137704 209064
rect 135364 209024 135370 209036
rect 137698 209024 137704 209036
rect 137756 209024 137762 209076
rect 174590 208996 174596 209008
rect 172768 208968 174596 208996
rect 171462 208888 171468 208940
rect 171520 208928 171526 208940
rect 172768 208928 172796 208968
rect 174590 208956 174596 208968
rect 174648 208956 174654 209008
rect 171520 208900 172796 208928
rect 171520 208888 171526 208900
rect 62534 208072 62540 208124
rect 62592 208112 62598 208124
rect 65662 208112 65668 208124
rect 62592 208084 65668 208112
rect 62592 208072 62598 208084
rect 65662 208072 65668 208084
rect 65720 208072 65726 208124
rect 135398 207664 135404 207716
rect 135456 207704 135462 207716
rect 136870 207704 136876 207716
rect 135456 207676 136876 207704
rect 135456 207664 135462 207676
rect 136870 207664 136876 207676
rect 136928 207664 136934 207716
rect 172566 207324 172572 207376
rect 172624 207364 172630 207376
rect 174038 207364 174044 207376
rect 172624 207336 174044 207364
rect 172624 207324 172630 207336
rect 174038 207324 174044 207336
rect 174096 207324 174102 207376
rect 62626 206848 62632 206900
rect 62684 206888 62690 206900
rect 65662 206888 65668 206900
rect 62684 206860 65668 206888
rect 62684 206848 62690 206860
rect 65662 206848 65668 206860
rect 65720 206848 65726 206900
rect 172658 202224 172664 202276
rect 172716 202264 172722 202276
rect 174222 202264 174228 202276
rect 172716 202236 174228 202264
rect 172716 202224 172722 202236
rect 174222 202224 174228 202236
rect 174280 202224 174286 202276
rect 62626 201884 62632 201936
rect 62684 201924 62690 201936
rect 65018 201924 65024 201936
rect 62684 201896 65024 201924
rect 62684 201884 62690 201896
rect 65018 201884 65024 201896
rect 65076 201884 65082 201936
rect 172658 200728 172664 200780
rect 172716 200768 172722 200780
rect 174130 200768 174136 200780
rect 172716 200740 174136 200768
rect 172716 200728 172722 200740
rect 174130 200728 174136 200740
rect 174188 200728 174194 200780
rect 100898 200660 100904 200712
rect 100956 200700 100962 200712
rect 102370 200700 102376 200712
rect 100956 200672 102376 200700
rect 100956 200660 100962 200672
rect 102370 200660 102376 200672
rect 102428 200660 102434 200712
rect 135398 200456 135404 200508
rect 135456 200496 135462 200508
rect 136778 200496 136784 200508
rect 135456 200468 136784 200496
rect 135456 200456 135462 200468
rect 136778 200456 136784 200468
rect 136836 200456 136842 200508
rect 62626 200388 62632 200440
rect 62684 200428 62690 200440
rect 65018 200428 65024 200440
rect 62684 200400 65024 200428
rect 62684 200388 62690 200400
rect 65018 200388 65024 200400
rect 65076 200388 65082 200440
rect 171646 199368 171652 199420
rect 171704 199408 171710 199420
rect 175234 199408 175240 199420
rect 171704 199380 175240 199408
rect 171704 199368 171710 199380
rect 175234 199368 175240 199380
rect 175292 199368 175298 199420
rect 100898 199300 100904 199352
rect 100956 199340 100962 199352
rect 102370 199340 102376 199352
rect 100956 199312 102376 199340
rect 100956 199300 100962 199312
rect 102370 199300 102376 199312
rect 102428 199300 102434 199352
rect 134754 199096 134760 199148
rect 134812 199136 134818 199148
rect 136778 199136 136784 199148
rect 134812 199108 136784 199136
rect 134812 199096 134818 199108
rect 136778 199096 136784 199108
rect 136836 199096 136842 199148
rect 62350 199028 62356 199080
rect 62408 199068 62414 199080
rect 65018 199068 65024 199080
rect 62408 199040 65024 199068
rect 62408 199028 62414 199040
rect 65018 199028 65024 199040
rect 65076 199028 65082 199080
rect 172658 198144 172664 198196
rect 172716 198184 172722 198196
rect 174130 198184 174136 198196
rect 172716 198156 174136 198184
rect 172716 198144 172722 198156
rect 174130 198144 174136 198156
rect 174188 198144 174194 198196
rect 100806 198008 100812 198060
rect 100864 198048 100870 198060
rect 102370 198048 102376 198060
rect 100864 198020 102376 198048
rect 100864 198008 100870 198020
rect 102370 198008 102376 198020
rect 102428 198008 102434 198060
rect 172658 198008 172664 198060
rect 172716 198048 172722 198060
rect 174222 198048 174228 198060
rect 172716 198020 174228 198048
rect 172716 198008 172722 198020
rect 174222 198008 174228 198020
rect 174280 198008 174286 198060
rect 65662 197912 65668 197924
rect 63748 197884 65668 197912
rect 62534 197804 62540 197856
rect 62592 197844 62598 197856
rect 63748 197844 63776 197884
rect 65662 197872 65668 197884
rect 65720 197872 65726 197924
rect 100898 197872 100904 197924
rect 100956 197912 100962 197924
rect 102462 197912 102468 197924
rect 100956 197884 102468 197912
rect 100956 197872 100962 197884
rect 102462 197872 102468 197884
rect 102520 197872 102526 197924
rect 62592 197816 63776 197844
rect 62592 197804 62598 197816
rect 62626 197736 62632 197788
rect 62684 197776 62690 197788
rect 65018 197776 65024 197788
rect 62684 197748 65024 197776
rect 62684 197736 62690 197748
rect 65018 197736 65024 197748
rect 65076 197736 65082 197788
rect 135398 197736 135404 197788
rect 135456 197776 135462 197788
rect 136778 197776 136784 197788
rect 135456 197748 136784 197776
rect 135456 197736 135462 197748
rect 136778 197736 136784 197748
rect 136836 197736 136842 197788
rect 135398 197396 135404 197448
rect 135456 197436 135462 197448
rect 136686 197436 136692 197448
rect 135456 197408 136692 197436
rect 135456 197396 135462 197408
rect 136686 197396 136692 197408
rect 136744 197396 136750 197448
rect 172566 196784 172572 196836
rect 172624 196824 172630 196836
rect 174130 196824 174136 196836
rect 172624 196796 174136 196824
rect 172624 196784 172630 196796
rect 174130 196784 174136 196796
rect 174188 196784 174194 196836
rect 100714 196648 100720 196700
rect 100772 196688 100778 196700
rect 102370 196688 102376 196700
rect 100772 196660 102376 196688
rect 100772 196648 100778 196660
rect 102370 196648 102376 196660
rect 102428 196648 102434 196700
rect 66214 196552 66220 196564
rect 63748 196524 66220 196552
rect 62626 196444 62632 196496
rect 62684 196484 62690 196496
rect 63748 196484 63776 196524
rect 66214 196512 66220 196524
rect 66272 196512 66278 196564
rect 100898 196512 100904 196564
rect 100956 196552 100962 196564
rect 102462 196552 102468 196564
rect 100956 196524 102468 196552
rect 100956 196512 100962 196524
rect 102462 196512 102468 196524
rect 102520 196512 102526 196564
rect 172658 196512 172664 196564
rect 172716 196552 172722 196564
rect 174222 196552 174228 196564
rect 172716 196524 174228 196552
rect 172716 196512 172722 196524
rect 174222 196512 174228 196524
rect 174280 196512 174286 196564
rect 62684 196456 63776 196484
rect 62684 196444 62690 196456
rect 135398 196376 135404 196428
rect 135456 196416 135462 196428
rect 136778 196416 136784 196428
rect 135456 196388 136784 196416
rect 135456 196376 135462 196388
rect 136778 196376 136784 196388
rect 136836 196376 136842 196428
rect 62534 196308 62540 196360
rect 62592 196348 62598 196360
rect 65018 196348 65024 196360
rect 62592 196320 65024 196348
rect 62592 196308 62598 196320
rect 65018 196308 65024 196320
rect 65076 196308 65082 196360
rect 135398 196172 135404 196224
rect 135456 196212 135462 196224
rect 136686 196212 136692 196224
rect 135456 196184 136692 196212
rect 135456 196172 135462 196184
rect 136686 196172 136692 196184
rect 136744 196172 136750 196224
rect 100898 195424 100904 195476
rect 100956 195464 100962 195476
rect 102554 195464 102560 195476
rect 100956 195436 102560 195464
rect 100956 195424 100962 195436
rect 102554 195424 102560 195436
rect 102612 195424 102618 195476
rect 172658 195288 172664 195340
rect 172716 195328 172722 195340
rect 174130 195328 174136 195340
rect 172716 195300 174136 195328
rect 172716 195288 172722 195300
rect 174130 195288 174136 195300
rect 174188 195288 174194 195340
rect 172382 195220 172388 195272
rect 172440 195260 172446 195272
rect 174222 195260 174228 195272
rect 172440 195232 174228 195260
rect 172440 195220 172446 195232
rect 174222 195220 174228 195232
rect 174280 195220 174286 195272
rect 66398 195192 66404 195204
rect 63748 195164 66404 195192
rect 62534 195084 62540 195136
rect 62592 195124 62598 195136
rect 63748 195124 63776 195164
rect 66398 195152 66404 195164
rect 66456 195152 66462 195204
rect 100898 195152 100904 195204
rect 100956 195192 100962 195204
rect 102370 195192 102376 195204
rect 100956 195164 102376 195192
rect 100956 195152 100962 195164
rect 102370 195152 102376 195164
rect 102428 195152 102434 195204
rect 136870 195192 136876 195204
rect 135508 195164 136876 195192
rect 62592 195096 63776 195124
rect 62592 195084 62598 195096
rect 135398 195084 135404 195136
rect 135456 195124 135462 195136
rect 135508 195124 135536 195164
rect 136870 195152 136876 195164
rect 136928 195152 136934 195204
rect 135456 195096 135536 195124
rect 135456 195084 135462 195096
rect 62626 195016 62632 195068
rect 62684 195056 62690 195068
rect 65018 195056 65024 195068
rect 62684 195028 65024 195056
rect 62684 195016 62690 195028
rect 65018 195016 65024 195028
rect 65076 195016 65082 195068
rect 135398 194812 135404 194864
rect 135456 194852 135462 194864
rect 136778 194852 136784 194864
rect 135456 194824 136784 194852
rect 135456 194812 135462 194824
rect 136778 194812 136784 194824
rect 136836 194812 136842 194864
rect 100622 194336 100628 194388
rect 100680 194376 100686 194388
rect 102462 194376 102468 194388
rect 100680 194348 102468 194376
rect 100680 194336 100686 194348
rect 102462 194336 102468 194348
rect 102520 194336 102526 194388
rect 171738 193928 171744 193980
rect 171796 193968 171802 193980
rect 174130 193968 174136 193980
rect 171796 193940 174136 193968
rect 171796 193928 171802 193940
rect 174130 193928 174136 193940
rect 174188 193928 174194 193980
rect 172658 193860 172664 193912
rect 172716 193900 172722 193912
rect 174222 193900 174228 193912
rect 172716 193872 174228 193900
rect 172716 193860 172722 193872
rect 174222 193860 174228 193872
rect 174280 193860 174286 193912
rect 100622 193792 100628 193844
rect 100680 193832 100686 193844
rect 102370 193832 102376 193844
rect 100680 193804 102376 193832
rect 100680 193792 100686 193804
rect 102370 193792 102376 193804
rect 102428 193792 102434 193844
rect 66398 193764 66404 193776
rect 63748 193736 66404 193764
rect 62626 193656 62632 193708
rect 62684 193696 62690 193708
rect 63748 193696 63776 193736
rect 66398 193724 66404 193736
rect 66456 193724 66462 193776
rect 62684 193668 63776 193696
rect 62684 193656 62690 193668
rect 135398 193656 135404 193708
rect 135456 193696 135462 193708
rect 136778 193696 136784 193708
rect 135456 193668 136784 193696
rect 135456 193656 135462 193668
rect 136778 193656 136784 193668
rect 136836 193656 136842 193708
rect 62534 193588 62540 193640
rect 62592 193628 62598 193640
rect 65018 193628 65024 193640
rect 62592 193600 65024 193628
rect 62592 193588 62598 193600
rect 65018 193588 65024 193600
rect 65076 193588 65082 193640
rect 135398 193452 135404 193504
rect 135456 193492 135462 193504
rect 136686 193492 136692 193504
rect 135456 193464 136692 193492
rect 135456 193452 135462 193464
rect 136686 193452 136692 193464
rect 136744 193452 136750 193504
rect 99886 192908 99892 192960
rect 99944 192948 99950 192960
rect 102462 192948 102468 192960
rect 99944 192920 102468 192948
rect 99944 192908 99950 192920
rect 102462 192908 102468 192920
rect 102520 192908 102526 192960
rect 172658 192704 172664 192756
rect 172716 192744 172722 192756
rect 174222 192744 174228 192756
rect 172716 192716 174228 192744
rect 172716 192704 172722 192716
rect 174222 192704 174228 192716
rect 174280 192704 174286 192756
rect 172014 192636 172020 192688
rect 172072 192676 172078 192688
rect 174130 192676 174136 192688
rect 172072 192648 174136 192676
rect 172072 192636 172078 192648
rect 174130 192636 174136 192648
rect 174188 192636 174194 192688
rect 171646 192568 171652 192620
rect 171704 192608 171710 192620
rect 174314 192608 174320 192620
rect 171704 192580 174320 192608
rect 171704 192568 171710 192580
rect 174314 192568 174320 192580
rect 174372 192568 174378 192620
rect 62626 192432 62632 192484
rect 62684 192472 62690 192484
rect 65662 192472 65668 192484
rect 62684 192444 65668 192472
rect 62684 192432 62690 192444
rect 65662 192432 65668 192444
rect 65720 192432 65726 192484
rect 100622 192432 100628 192484
rect 100680 192472 100686 192484
rect 102370 192472 102376 192484
rect 100680 192444 102376 192472
rect 100680 192432 100686 192444
rect 102370 192432 102376 192444
rect 102428 192432 102434 192484
rect 100530 192364 100536 192416
rect 100588 192404 100594 192416
rect 102646 192404 102652 192416
rect 100588 192376 102652 192404
rect 100588 192364 100594 192376
rect 102646 192364 102652 192376
rect 102704 192364 102710 192416
rect 135306 192364 135312 192416
rect 135364 192404 135370 192416
rect 136870 192404 136876 192416
rect 135364 192376 136876 192404
rect 135364 192364 135370 192376
rect 136870 192364 136876 192376
rect 136928 192364 136934 192416
rect 135398 192296 135404 192348
rect 135456 192336 135462 192348
rect 136778 192336 136784 192348
rect 135456 192308 136784 192336
rect 135456 192296 135462 192308
rect 136778 192296 136784 192308
rect 136836 192296 136842 192348
rect 62534 192228 62540 192280
rect 62592 192268 62598 192280
rect 64926 192268 64932 192280
rect 62592 192240 64932 192268
rect 62592 192228 62598 192240
rect 64926 192228 64932 192240
rect 64984 192228 64990 192280
rect 135214 192092 135220 192144
rect 135272 192132 135278 192144
rect 136686 192132 136692 192144
rect 135272 192104 136692 192132
rect 135272 192092 135278 192104
rect 136686 192092 136692 192104
rect 136744 192092 136750 192144
rect 62350 191616 62356 191668
rect 62408 191656 62414 191668
rect 65018 191656 65024 191668
rect 62408 191628 65024 191656
rect 62408 191616 62414 191628
rect 65018 191616 65024 191628
rect 65076 191616 65082 191668
rect 100622 191208 100628 191260
rect 100680 191248 100686 191260
rect 102278 191248 102284 191260
rect 100680 191220 102284 191248
rect 100680 191208 100686 191220
rect 102278 191208 102284 191220
rect 102336 191208 102342 191260
rect 172658 191208 172664 191260
rect 172716 191248 172722 191260
rect 174038 191248 174044 191260
rect 172716 191220 174044 191248
rect 172716 191208 172722 191220
rect 174038 191208 174044 191220
rect 174096 191208 174102 191260
rect 171830 191072 171836 191124
rect 171888 191112 171894 191124
rect 175326 191112 175332 191124
rect 171888 191084 175332 191112
rect 171888 191072 171894 191084
rect 175326 191072 175332 191084
rect 175384 191072 175390 191124
rect 100898 191004 100904 191056
rect 100956 191044 100962 191056
rect 102554 191044 102560 191056
rect 100956 191016 102560 191044
rect 100956 191004 100962 191016
rect 102554 191004 102560 191016
rect 102612 191004 102618 191056
rect 134202 191004 134208 191056
rect 134260 191044 134266 191056
rect 137146 191044 137152 191056
rect 134260 191016 137152 191044
rect 134260 191004 134266 191016
rect 137146 191004 137152 191016
rect 137204 191004 137210 191056
rect 62350 190800 62356 190852
rect 62408 190840 62414 190852
rect 65018 190840 65024 190852
rect 62408 190812 65024 190840
rect 62408 190800 62414 190812
rect 65018 190800 65024 190812
rect 65076 190800 65082 190852
rect 135398 190732 135404 190784
rect 135456 190772 135462 190784
rect 136778 190772 136784 190784
rect 135456 190744 136784 190772
rect 135456 190732 135462 190744
rect 136778 190732 136784 190744
rect 136836 190732 136842 190784
rect 100438 190120 100444 190172
rect 100496 190160 100502 190172
rect 102370 190160 102376 190172
rect 100496 190132 102376 190160
rect 100496 190120 100502 190132
rect 102370 190120 102376 190132
rect 102428 190120 102434 190172
rect 171646 189916 171652 189968
rect 171704 189956 171710 189968
rect 174406 189956 174412 189968
rect 171704 189928 174412 189956
rect 171704 189916 171710 189928
rect 174406 189916 174412 189928
rect 174464 189916 174470 189968
rect 99978 189848 99984 189900
rect 100036 189888 100042 189900
rect 102462 189888 102468 189900
rect 100036 189860 102468 189888
rect 100036 189848 100042 189860
rect 102462 189848 102468 189860
rect 102520 189848 102526 189900
rect 171830 189712 171836 189764
rect 171888 189752 171894 189764
rect 175418 189752 175424 189764
rect 171888 189724 175424 189752
rect 171888 189712 171894 189724
rect 175418 189712 175424 189724
rect 175476 189712 175482 189764
rect 63638 189644 63644 189696
rect 63696 189684 63702 189696
rect 66398 189684 66404 189696
rect 63696 189656 66404 189684
rect 63696 189644 63702 189656
rect 66398 189644 66404 189656
rect 66456 189644 66462 189696
rect 62626 189508 62632 189560
rect 62684 189548 62690 189560
rect 65202 189548 65208 189560
rect 62684 189520 65208 189548
rect 62684 189508 62690 189520
rect 65202 189508 65208 189520
rect 65260 189508 65266 189560
rect 134754 189236 134760 189288
rect 134812 189276 134818 189288
rect 136778 189276 136784 189288
rect 134812 189248 136784 189276
rect 134812 189236 134818 189248
rect 136778 189236 136784 189248
rect 136836 189236 136842 189288
rect 62626 189032 62632 189084
rect 62684 189072 62690 189084
rect 65018 189072 65024 189084
rect 62684 189044 65024 189072
rect 62684 189032 62690 189044
rect 65018 189032 65024 189044
rect 65076 189032 65082 189084
rect 134938 188148 134944 188200
rect 134996 188188 135002 188200
rect 137238 188188 137244 188200
rect 134996 188160 137244 188188
rect 134996 188148 135002 188160
rect 137238 188148 137244 188160
rect 137296 188148 137302 188200
rect 116446 187604 116452 187656
rect 116504 187644 116510 187656
rect 117412 187644 117418 187656
rect 116504 187616 117418 187644
rect 116504 187604 116510 187616
rect 117412 187604 117418 187616
rect 117470 187604 117476 187656
rect 183974 186856 183980 186908
rect 184032 186896 184038 186908
rect 184434 186896 184440 186908
rect 184032 186868 184440 186896
rect 184032 186856 184038 186868
rect 184434 186856 184440 186868
rect 184492 186856 184498 186908
rect 188482 186856 188488 186908
rect 188540 186896 188546 186908
rect 189126 186896 189132 186908
rect 188540 186868 189132 186896
rect 188540 186856 188546 186868
rect 189126 186856 189132 186868
rect 189184 186856 189190 186908
rect 36314 185428 36320 185480
rect 36372 185468 36378 185480
rect 40638 185468 40644 185480
rect 36372 185440 40644 185468
rect 36372 185428 36378 185440
rect 40638 185428 40644 185440
rect 40696 185428 40702 185480
rect 41006 185428 41012 185480
rect 41064 185468 41070 185480
rect 43398 185468 43404 185480
rect 41064 185440 43404 185468
rect 41064 185428 41070 185440
rect 43398 185428 43404 185440
rect 43456 185428 43462 185480
rect 43766 185428 43772 185480
rect 43824 185468 43830 185480
rect 44686 185468 44692 185480
rect 43824 185440 44692 185468
rect 43824 185428 43830 185440
rect 44686 185428 44692 185440
rect 44744 185428 44750 185480
rect 49010 185428 49016 185480
rect 49068 185468 49074 185480
rect 50574 185468 50580 185480
rect 49068 185440 50580 185468
rect 49068 185428 49074 185440
rect 50574 185428 50580 185440
rect 50632 185428 50638 185480
rect 50666 185428 50672 185480
rect 50724 185468 50730 185480
rect 53334 185468 53340 185480
rect 50724 185440 53340 185468
rect 50724 185428 50730 185440
rect 53334 185428 53340 185440
rect 53392 185428 53398 185480
rect 53426 185428 53432 185480
rect 53484 185468 53490 185480
rect 58118 185468 58124 185480
rect 53484 185440 58124 185468
rect 53484 185428 53490 185440
rect 58118 185428 58124 185440
rect 58176 185428 58182 185480
rect 110098 185428 110104 185480
rect 110156 185468 110162 185480
rect 111110 185468 111116 185480
rect 110156 185440 111116 185468
rect 110156 185428 110162 185440
rect 111110 185428 111116 185440
rect 111168 185428 111174 185480
rect 117550 185428 117556 185480
rect 117608 185468 117614 185480
rect 118930 185468 118936 185480
rect 117608 185440 118936 185468
rect 117608 185428 117614 185440
rect 118930 185428 118936 185440
rect 118988 185428 118994 185480
rect 120218 185428 120224 185480
rect 120276 185468 120282 185480
rect 122334 185468 122340 185480
rect 120276 185440 122340 185468
rect 120276 185428 120282 185440
rect 122334 185428 122340 185440
rect 122392 185428 122398 185480
rect 122426 185428 122432 185480
rect 122484 185468 122490 185480
rect 123438 185468 123444 185480
rect 122484 185440 123444 185468
rect 122484 185428 122490 185440
rect 123438 185428 123444 185440
rect 123496 185428 123502 185480
rect 124174 185428 124180 185480
rect 124232 185468 124238 185480
rect 128130 185468 128136 185480
rect 124232 185440 128136 185468
rect 124232 185428 124238 185440
rect 128130 185428 128136 185440
rect 128188 185428 128194 185480
rect 182226 185428 182232 185480
rect 182284 185468 182290 185480
rect 183238 185468 183244 185480
rect 182284 185440 183244 185468
rect 182284 185428 182290 185440
rect 183238 185428 183244 185440
rect 183296 185428 183302 185480
rect 188114 185428 188120 185480
rect 188172 185468 188178 185480
rect 188574 185468 188580 185480
rect 188172 185440 188580 185468
rect 188172 185428 188178 185440
rect 188574 185428 188580 185440
rect 188632 185428 188638 185480
rect 190598 185428 190604 185480
rect 190656 185468 190662 185480
rect 192530 185468 192536 185480
rect 190656 185440 192536 185468
rect 190656 185428 190662 185440
rect 192530 185428 192536 185440
rect 192588 185428 192594 185480
rect 192898 185428 192904 185480
rect 192956 185468 192962 185480
rect 195382 185468 195388 185480
rect 192956 185440 195388 185468
rect 192956 185428 192962 185440
rect 195382 185428 195388 185440
rect 195440 185428 195446 185480
rect 197314 185428 197320 185480
rect 197372 185468 197378 185480
rect 201638 185468 201644 185480
rect 197372 185440 201644 185468
rect 197372 185428 197378 185440
rect 201638 185428 201644 185440
rect 201696 185428 201702 185480
rect 40362 185360 40368 185412
rect 40420 185400 40426 185412
rect 43030 185400 43036 185412
rect 40420 185372 43036 185400
rect 40420 185360 40426 185372
rect 43030 185360 43036 185372
rect 43088 185360 43094 185412
rect 43122 185360 43128 185412
rect 43180 185400 43186 185412
rect 44594 185400 44600 185412
rect 43180 185372 44600 185400
rect 43180 185360 43186 185372
rect 44594 185360 44600 185372
rect 44652 185360 44658 185412
rect 49838 185360 49844 185412
rect 49896 185400 49902 185412
rect 51954 185400 51960 185412
rect 49896 185372 51960 185400
rect 49896 185360 49902 185372
rect 51954 185360 51960 185372
rect 52012 185360 52018 185412
rect 110742 185360 110748 185412
rect 110800 185400 110806 185412
rect 111478 185400 111484 185412
rect 110800 185372 111484 185400
rect 110800 185360 110806 185372
rect 111478 185360 111484 185372
rect 111536 185360 111542 185412
rect 118562 185360 118568 185412
rect 118620 185400 118626 185412
rect 120310 185400 120316 185412
rect 118620 185372 120316 185400
rect 118620 185360 118626 185372
rect 120310 185360 120316 185372
rect 120368 185360 120374 185412
rect 124542 185360 124548 185412
rect 124600 185400 124606 185412
rect 128682 185400 128688 185412
rect 124600 185372 128688 185400
rect 124600 185360 124606 185372
rect 128682 185360 128688 185372
rect 128740 185360 128746 185412
rect 191702 185360 191708 185412
rect 191760 185400 191766 185412
rect 193634 185400 193640 185412
rect 191760 185372 193640 185400
rect 191760 185360 191766 185372
rect 193634 185360 193640 185372
rect 193692 185360 193698 185412
rect 194094 185360 194100 185412
rect 194152 185400 194158 185412
rect 197130 185400 197136 185412
rect 194152 185372 197136 185400
rect 194152 185360 194158 185372
rect 197130 185360 197136 185372
rect 197188 185360 197194 185412
rect 37602 185292 37608 185344
rect 37660 185332 37666 185344
rect 41466 185332 41472 185344
rect 37660 185304 41472 185332
rect 37660 185292 37666 185304
rect 41466 185292 41472 185304
rect 41524 185292 41530 185344
rect 41742 185292 41748 185344
rect 41800 185332 41806 185344
rect 43858 185332 43864 185344
rect 41800 185304 43864 185332
rect 41800 185292 41806 185304
rect 43858 185292 43864 185304
rect 43916 185292 43922 185344
rect 52230 185292 52236 185344
rect 52288 185332 52294 185344
rect 56094 185332 56100 185344
rect 52288 185304 56100 185332
rect 52288 185292 52294 185304
rect 56094 185292 56100 185304
rect 56152 185292 56158 185344
rect 123806 185292 123812 185344
rect 123864 185332 123870 185344
rect 127578 185332 127584 185344
rect 123864 185304 127584 185332
rect 123864 185292 123870 185304
rect 127578 185292 127584 185304
rect 127636 185292 127642 185344
rect 176890 185292 176896 185344
rect 176948 185332 176954 185344
rect 177718 185332 177724 185344
rect 176948 185304 177724 185332
rect 176948 185292 176954 185304
rect 177718 185292 177724 185304
rect 177776 185292 177782 185344
rect 192530 185292 192536 185344
rect 192588 185332 192594 185344
rect 194830 185332 194836 185344
rect 192588 185304 194836 185332
rect 192588 185292 192594 185304
rect 194830 185292 194836 185304
rect 194888 185292 194894 185344
rect 195750 185292 195756 185344
rect 195808 185332 195814 185344
rect 199338 185332 199344 185344
rect 195808 185304 199344 185332
rect 195808 185292 195814 185304
rect 199338 185292 199344 185304
rect 199396 185292 199402 185344
rect 39718 185224 39724 185276
rect 39776 185264 39782 185276
rect 42662 185264 42668 185276
rect 39776 185236 42668 185264
rect 39776 185224 39782 185236
rect 42662 185224 42668 185236
rect 42720 185224 42726 185276
rect 49470 185224 49476 185276
rect 49528 185264 49534 185276
rect 51310 185264 51316 185276
rect 49528 185236 51316 185264
rect 49528 185224 49534 185236
rect 51310 185224 51316 185236
rect 51368 185224 51374 185276
rect 53058 185224 53064 185276
rect 53116 185264 53122 185276
rect 57382 185264 57388 185276
rect 53116 185236 57388 185264
rect 53116 185224 53122 185236
rect 57382 185224 57388 185236
rect 57440 185224 57446 185276
rect 105590 185224 105596 185276
rect 105648 185264 105654 185276
rect 109270 185264 109276 185276
rect 105648 185236 109276 185264
rect 105648 185224 105654 185236
rect 109270 185224 109276 185236
rect 109328 185224 109334 185276
rect 118930 185224 118936 185276
rect 118988 185264 118994 185276
rect 120586 185264 120592 185276
rect 118988 185236 120592 185264
rect 118988 185224 118994 185236
rect 120586 185224 120592 185236
rect 120644 185224 120650 185276
rect 123346 185224 123352 185276
rect 123404 185264 123410 185276
rect 127302 185264 127308 185276
rect 123404 185236 127308 185264
rect 123404 185224 123410 185236
rect 127302 185224 127308 185236
rect 127360 185224 127366 185276
rect 193358 185224 193364 185276
rect 193416 185264 193422 185276
rect 195934 185264 195940 185276
rect 193416 185236 195940 185264
rect 193416 185224 193422 185236
rect 195934 185224 195940 185236
rect 195992 185224 195998 185276
rect 196118 185224 196124 185276
rect 196176 185264 196182 185276
rect 199982 185264 199988 185276
rect 196176 185236 199988 185264
rect 196176 185224 196182 185236
rect 199982 185224 199988 185236
rect 200040 185224 200046 185276
rect 36958 185156 36964 185208
rect 37016 185196 37022 185208
rect 41006 185196 41012 185208
rect 37016 185168 41012 185196
rect 37016 185156 37022 185168
rect 41006 185156 41012 185168
rect 41064 185156 41070 185208
rect 50206 185156 50212 185208
rect 50264 185196 50270 185208
rect 52690 185196 52696 185208
rect 50264 185168 52696 185196
rect 50264 185156 50270 185168
rect 52690 185156 52696 185168
rect 52748 185156 52754 185208
rect 122610 185156 122616 185208
rect 122668 185196 122674 185208
rect 125830 185196 125836 185208
rect 122668 185168 125836 185196
rect 122668 185156 122674 185168
rect 125830 185156 125836 185168
rect 125888 185156 125894 185208
rect 177718 185156 177724 185208
rect 177776 185196 177782 185208
rect 181122 185196 181128 185208
rect 177776 185168 181128 185196
rect 177776 185156 177782 185168
rect 181122 185156 181128 185168
rect 181180 185156 181186 185208
rect 194554 185156 194560 185208
rect 194612 185196 194618 185208
rect 197682 185196 197688 185208
rect 194612 185168 197688 185196
rect 194612 185156 194618 185168
rect 197682 185156 197688 185168
rect 197740 185156 197746 185208
rect 34934 185088 34940 185140
rect 34992 185128 34998 185140
rect 39534 185128 39540 185140
rect 34992 185100 39540 185128
rect 34992 185088 34998 185100
rect 39534 185088 39540 185100
rect 39592 185088 39598 185140
rect 42386 185088 42392 185140
rect 42444 185128 42450 185140
rect 44226 185128 44232 185140
rect 42444 185100 44232 185128
rect 42444 185088 42450 185100
rect 44226 185088 44232 185100
rect 44284 185088 44290 185140
rect 52598 185088 52604 185140
rect 52656 185128 52662 185140
rect 56738 185128 56744 185140
rect 52656 185100 56744 185128
rect 52656 185088 52662 185100
rect 56738 185088 56744 185100
rect 56796 185088 56802 185140
rect 122978 185088 122984 185140
rect 123036 185128 123042 185140
rect 126382 185128 126388 185140
rect 123036 185100 126388 185128
rect 123036 185088 123042 185100
rect 126382 185088 126388 185100
rect 126440 185088 126446 185140
rect 190414 185088 190420 185140
rect 190472 185128 190478 185140
rect 191978 185128 191984 185140
rect 190472 185100 191984 185128
rect 190472 185088 190478 185100
rect 191978 185088 191984 185100
rect 192036 185088 192042 185140
rect 193726 185088 193732 185140
rect 193784 185128 193790 185140
rect 196486 185128 196492 185140
rect 193784 185100 196492 185128
rect 193784 185088 193790 185100
rect 196486 185088 196492 185100
rect 196544 185088 196550 185140
rect 38982 185020 38988 185072
rect 39040 185060 39046 185072
rect 42202 185060 42208 185072
rect 39040 185032 42208 185060
rect 39040 185020 39046 185032
rect 42202 185020 42208 185032
rect 42260 185020 42266 185072
rect 48642 185020 48648 185072
rect 48700 185060 48706 185072
rect 49930 185060 49936 185072
rect 48700 185032 49936 185060
rect 48700 185020 48706 185032
rect 49930 185020 49936 185032
rect 49988 185020 49994 185072
rect 51034 185020 51040 185072
rect 51092 185060 51098 185072
rect 53978 185060 53984 185072
rect 51092 185032 53984 185060
rect 51092 185020 51098 185032
rect 53978 185020 53984 185032
rect 54036 185020 54042 185072
rect 121322 185020 121328 185072
rect 121380 185060 121386 185072
rect 124450 185060 124456 185072
rect 121380 185032 124456 185060
rect 121380 185020 121386 185032
rect 124450 185020 124456 185032
rect 124508 185020 124514 185072
rect 194646 185020 194652 185072
rect 194704 185060 194710 185072
rect 198234 185060 198240 185072
rect 194704 185032 198240 185060
rect 194704 185020 194710 185032
rect 198234 185020 198240 185032
rect 198292 185020 198298 185072
rect 38338 184952 38344 185004
rect 38396 184992 38402 185004
rect 41834 184992 41840 185004
rect 38396 184964 41840 184992
rect 38396 184952 38402 184964
rect 41834 184952 41840 184964
rect 41892 184952 41898 185004
rect 51402 184952 51408 185004
rect 51460 184992 51466 185004
rect 54714 184992 54720 185004
rect 51460 184964 54720 184992
rect 51460 184952 51466 184964
rect 54714 184952 54720 184964
rect 54772 184952 54778 185004
rect 121782 184952 121788 185004
rect 121840 184992 121846 185004
rect 124634 184992 124640 185004
rect 121840 184964 124640 184992
rect 121840 184952 121846 184964
rect 124634 184952 124640 184964
rect 124692 184952 124698 185004
rect 181674 184952 181680 185004
rect 181732 184992 181738 185004
rect 183100 184992 183106 185004
rect 181732 184964 183106 184992
rect 181732 184952 181738 184964
rect 183100 184952 183106 184964
rect 183158 184952 183164 185004
rect 183422 184952 183428 185004
rect 183480 184992 183486 185004
rect 184296 184992 184302 185004
rect 183480 184964 184302 184992
rect 183480 184952 183486 184964
rect 184296 184952 184302 184964
rect 184354 184952 184360 185004
rect 188620 184952 188626 185004
rect 188678 184992 188684 185004
rect 189678 184992 189684 185004
rect 188678 184964 189684 184992
rect 188678 184952 188684 184964
rect 189678 184952 189684 184964
rect 189736 184952 189742 185004
rect 189816 184952 189822 185004
rect 189874 184992 189880 185004
rect 191426 184992 191432 185004
rect 189874 184964 191432 184992
rect 189874 184952 189880 184964
rect 191426 184952 191432 184964
rect 191484 184952 191490 185004
rect 191840 184952 191846 185004
rect 191898 184992 191904 185004
rect 194278 184992 194284 185004
rect 191898 184964 194284 184992
rect 191898 184952 191904 184964
rect 194278 184952 194284 184964
rect 194336 184952 194342 185004
rect 197820 184952 197826 185004
rect 197878 184992 197884 185004
rect 202834 184992 202840 185004
rect 197878 184964 202840 184992
rect 197878 184952 197884 184964
rect 202834 184952 202840 184964
rect 202892 184952 202898 185004
rect 51862 184884 51868 184936
rect 51920 184924 51926 184936
rect 55358 184924 55364 184936
rect 51920 184896 55364 184924
rect 51920 184884 51926 184896
rect 55358 184884 55364 184896
rect 55416 184884 55422 184936
rect 122150 184884 122156 184936
rect 122208 184924 122214 184936
rect 125186 184924 125192 184936
rect 122208 184896 125192 184924
rect 122208 184884 122214 184896
rect 125186 184884 125192 184896
rect 125244 184884 125250 184936
rect 182870 184884 182876 184936
rect 182928 184924 182934 184936
rect 183836 184924 183842 184936
rect 182928 184896 183842 184924
rect 182928 184884 182934 184896
rect 183836 184884 183842 184896
rect 183894 184884 183900 184936
rect 189080 184884 189086 184936
rect 189138 184924 189144 184936
rect 190230 184924 190236 184936
rect 189138 184896 190236 184924
rect 189138 184884 189144 184896
rect 190230 184884 190236 184896
rect 190288 184884 190294 184936
rect 191104 184884 191110 184936
rect 191162 184924 191168 184936
rect 193082 184924 193088 184936
rect 191162 184896 193088 184924
rect 191162 184884 191168 184896
rect 193082 184884 193088 184896
rect 193140 184884 193146 184936
rect 196624 184884 196630 184936
rect 196682 184924 196688 184936
rect 201086 184924 201092 184936
rect 196682 184896 201092 184924
rect 196682 184884 196688 184896
rect 201086 184884 201092 184896
rect 201144 184884 201150 184936
rect 189678 184816 189684 184868
rect 189736 184856 189742 184868
rect 190782 184856 190788 184868
rect 189736 184828 190788 184856
rect 189736 184816 189742 184828
rect 190782 184816 190788 184828
rect 190840 184816 190846 184868
rect 196486 184816 196492 184868
rect 196544 184856 196550 184868
rect 200534 184856 200540 184868
rect 196544 184828 200540 184856
rect 196544 184816 196550 184828
rect 200534 184816 200540 184828
rect 200592 184816 200598 184868
rect 195290 184748 195296 184800
rect 195348 184788 195354 184800
rect 198786 184788 198792 184800
rect 195348 184760 198792 184788
rect 195348 184748 195354 184760
rect 198786 184748 198792 184760
rect 198844 184748 198850 184800
rect 35578 184408 35584 184460
rect 35636 184448 35642 184460
rect 38154 184448 38160 184460
rect 35636 184420 38160 184448
rect 35636 184408 35642 184420
rect 38154 184408 38160 184420
rect 38212 184408 38218 184460
rect 39258 184408 39264 184460
rect 39316 184408 39322 184460
rect 53978 184408 53984 184460
rect 54036 184408 54042 184460
rect 54530 184408 54536 184460
rect 54588 184408 54594 184460
rect 34198 184272 34204 184324
rect 34256 184312 34262 184324
rect 39276 184312 39304 184408
rect 34256 184284 39304 184312
rect 34256 184272 34262 184284
rect 33554 184068 33560 184120
rect 33612 184108 33618 184120
rect 38890 184108 38896 184120
rect 33612 184080 38896 184108
rect 33612 184068 33618 184080
rect 38890 184068 38896 184080
rect 38948 184068 38954 184120
rect 53996 184108 54024 184408
rect 54548 184244 54576 184408
rect 106050 184340 106056 184392
rect 106108 184380 106114 184392
rect 107154 184380 107160 184392
rect 106108 184352 107160 184380
rect 106108 184340 106114 184352
rect 107154 184340 107160 184352
rect 107212 184340 107218 184392
rect 176982 184340 176988 184392
rect 177040 184380 177046 184392
rect 179374 184380 179380 184392
rect 177040 184352 179380 184380
rect 177040 184340 177046 184352
rect 179374 184340 179380 184352
rect 179432 184340 179438 184392
rect 59498 184244 59504 184256
rect 54548 184216 59504 184244
rect 59498 184204 59504 184216
rect 59556 184204 59562 184256
rect 177626 184136 177632 184188
rect 177684 184176 177690 184188
rect 178270 184176 178276 184188
rect 177684 184148 178276 184176
rect 177684 184136 177690 184148
rect 178270 184136 178276 184148
rect 178328 184136 178334 184188
rect 58762 184108 58768 184120
rect 53996 184080 58768 184108
rect 58762 184068 58768 184080
rect 58820 184068 58826 184120
rect 105958 184068 105964 184120
rect 106016 184108 106022 184120
rect 106602 184108 106608 184120
rect 106016 184080 106608 184108
rect 106016 184068 106022 184080
rect 106602 184068 106608 184080
rect 106660 184068 106666 184120
rect 108350 184108 108356 184120
rect 106712 184080 108356 184108
rect 106142 184000 106148 184052
rect 106200 184040 106206 184052
rect 106712 184040 106740 184080
rect 108350 184068 108356 184080
rect 108408 184068 108414 184120
rect 177810 184068 177816 184120
rect 177868 184108 177874 184120
rect 178822 184108 178828 184120
rect 177868 184080 178828 184108
rect 177868 184068 177874 184080
rect 178822 184068 178828 184080
rect 178880 184068 178886 184120
rect 180570 184108 180576 184120
rect 178932 184080 180576 184108
rect 106200 184012 106740 184040
rect 106200 184000 106206 184012
rect 177350 184000 177356 184052
rect 177408 184040 177414 184052
rect 178932 184040 178960 184080
rect 180570 184068 180576 184080
rect 180628 184068 180634 184120
rect 177408 184012 178960 184040
rect 177408 184000 177414 184012
rect 105590 182368 105596 182420
rect 105648 182408 105654 182420
rect 107890 182408 107896 182420
rect 105648 182380 107896 182408
rect 105648 182368 105654 182380
rect 107890 182368 107896 182380
rect 107948 182368 107954 182420
rect 177166 182164 177172 182216
rect 177224 182204 177230 182216
rect 180018 182204 180024 182216
rect 177224 182176 180024 182204
rect 177224 182164 177230 182176
rect 180018 182164 180024 182176
rect 180076 182164 180082 182216
rect 105406 180328 105412 180380
rect 105464 180368 105470 180380
rect 108074 180368 108080 180380
rect 105464 180340 108080 180368
rect 105464 180328 105470 180340
rect 108074 180328 108080 180340
rect 108132 180328 108138 180380
rect 178086 180328 178092 180380
rect 178144 180368 178150 180380
rect 179650 180368 179656 180380
rect 178144 180340 179656 180368
rect 178144 180328 178150 180340
rect 179650 180328 179656 180340
rect 179708 180328 179714 180380
rect 106326 178560 106332 178612
rect 106384 178600 106390 178612
rect 107890 178600 107896 178612
rect 106384 178572 107896 178600
rect 106384 178560 106390 178572
rect 107890 178560 107896 178572
rect 107948 178560 107954 178612
rect 177810 178560 177816 178612
rect 177868 178600 177874 178612
rect 179650 178600 179656 178612
rect 177868 178572 179656 178600
rect 177868 178560 177874 178572
rect 179650 178560 179656 178572
rect 179708 178560 179714 178612
rect 32634 177200 32640 177252
rect 32692 177240 32698 177252
rect 37418 177240 37424 177252
rect 32692 177212 37424 177240
rect 32692 177200 32698 177212
rect 37418 177200 37424 177212
rect 37476 177200 37482 177252
rect 106418 175840 106424 175892
rect 106476 175880 106482 175892
rect 107890 175880 107896 175892
rect 106476 175852 107896 175880
rect 106476 175840 106482 175852
rect 107890 175840 107896 175852
rect 107948 175840 107954 175892
rect 177718 175840 177724 175892
rect 177776 175880 177782 175892
rect 179650 175880 179656 175892
rect 177776 175852 179656 175880
rect 177776 175840 177782 175852
rect 179650 175840 179656 175852
rect 179708 175840 179714 175892
rect 57382 175772 57388 175824
rect 57440 175812 57446 175824
rect 59590 175812 59596 175824
rect 57440 175784 59596 175812
rect 57440 175772 57446 175784
rect 59590 175772 59596 175784
rect 59648 175772 59654 175824
rect 177166 175568 177172 175620
rect 177224 175608 177230 175620
rect 180294 175608 180300 175620
rect 177224 175580 180300 175608
rect 177224 175568 177230 175580
rect 180294 175568 180300 175580
rect 180352 175568 180358 175620
rect 106142 175364 106148 175416
rect 106200 175404 106206 175416
rect 108534 175404 108540 175416
rect 106200 175376 108540 175404
rect 106200 175364 106206 175376
rect 108534 175364 108540 175376
rect 108592 175364 108598 175416
rect 105958 173052 105964 173104
rect 106016 173092 106022 173104
rect 107890 173092 107896 173104
rect 106016 173064 107896 173092
rect 106016 173052 106022 173064
rect 107890 173052 107896 173064
rect 107948 173052 107954 173104
rect 177534 173052 177540 173104
rect 177592 173092 177598 173104
rect 179650 173092 179656 173104
rect 177592 173064 179656 173092
rect 177592 173052 177598 173064
rect 179650 173052 179656 173064
rect 179708 173052 179714 173104
rect 105682 171692 105688 171744
rect 105740 171732 105746 171744
rect 108074 171732 108080 171744
rect 105740 171704 108080 171732
rect 105740 171692 105746 171704
rect 108074 171692 108080 171704
rect 108132 171692 108138 171744
rect 178178 171692 178184 171744
rect 178236 171732 178242 171744
rect 179650 171732 179656 171744
rect 178236 171704 179656 171732
rect 178236 171692 178242 171704
rect 179650 171692 179656 171704
rect 179708 171692 179714 171744
rect 222798 169108 222804 169160
rect 222856 169148 222862 169160
rect 223534 169148 223540 169160
rect 222856 169120 223540 169148
rect 222856 169108 222862 169120
rect 223534 169108 223540 169120
rect 223592 169108 223598 169160
rect 201086 166116 201092 166168
rect 201144 166156 201150 166168
rect 204490 166156 204496 166168
rect 201144 166128 204496 166156
rect 201144 166116 201150 166128
rect 204490 166116 204496 166128
rect 204548 166116 204554 166168
rect 177166 165300 177172 165352
rect 177224 165340 177230 165352
rect 179558 165340 179564 165352
rect 177224 165312 179564 165340
rect 177224 165300 177230 165312
rect 179558 165300 179564 165312
rect 179616 165300 179622 165352
rect 105222 165232 105228 165284
rect 105280 165272 105286 165284
rect 107798 165272 107804 165284
rect 105280 165244 107804 165272
rect 105280 165232 105286 165244
rect 107798 165232 107804 165244
rect 107856 165232 107862 165284
rect 28862 164756 28868 164808
rect 28920 164796 28926 164808
rect 37418 164796 37424 164808
rect 28920 164768 37424 164796
rect 28920 164756 28926 164768
rect 37418 164756 37424 164768
rect 37476 164756 37482 164808
rect 54806 164756 54812 164808
rect 54864 164796 54870 164808
rect 59590 164796 59596 164808
rect 54864 164768 59596 164796
rect 54864 164756 54870 164768
rect 59590 164756 59596 164768
rect 59648 164756 59654 164808
rect 177534 163600 177540 163652
rect 177592 163640 177598 163652
rect 179558 163640 179564 163652
rect 177592 163612 179564 163640
rect 177592 163600 177598 163612
rect 179558 163600 179564 163612
rect 179616 163600 179622 163652
rect 105590 163464 105596 163516
rect 105648 163504 105654 163516
rect 107430 163504 107436 163516
rect 105648 163476 107436 163504
rect 105648 163464 105654 163476
rect 107430 163464 107436 163476
rect 107488 163464 107494 163516
rect 105774 163396 105780 163448
rect 105832 163436 105838 163448
rect 107798 163436 107804 163448
rect 105832 163408 107804 163436
rect 105832 163396 105838 163408
rect 107798 163396 107804 163408
rect 107856 163396 107862 163448
rect 176982 163396 176988 163448
rect 177040 163436 177046 163448
rect 179190 163436 179196 163448
rect 177040 163408 179196 163436
rect 177040 163396 177046 163408
rect 179190 163396 179196 163408
rect 179248 163396 179254 163448
rect 105682 162036 105688 162088
rect 105740 162076 105746 162088
rect 107798 162076 107804 162088
rect 105740 162048 107804 162076
rect 105740 162036 105746 162048
rect 107798 162036 107804 162048
rect 107856 162036 107862 162088
rect 176982 162036 176988 162088
rect 177040 162076 177046 162088
rect 179558 162076 179564 162088
rect 177040 162048 179564 162076
rect 177040 162036 177046 162048
rect 179558 162036 179564 162048
rect 179616 162036 179622 162088
rect 105222 161016 105228 161068
rect 105280 161056 105286 161068
rect 107706 161056 107712 161068
rect 105280 161028 107712 161056
rect 105280 161016 105286 161028
rect 107706 161016 107712 161028
rect 107764 161016 107770 161068
rect 177534 160880 177540 160932
rect 177592 160920 177598 160932
rect 179466 160920 179472 160932
rect 177592 160892 179472 160920
rect 177592 160880 177598 160892
rect 179466 160880 179472 160892
rect 179524 160880 179530 160932
rect 105590 159520 105596 159572
rect 105648 159560 105654 159572
rect 107614 159560 107620 159572
rect 105648 159532 107620 159560
rect 105648 159520 105654 159532
rect 107614 159520 107620 159532
rect 107672 159520 107678 159572
rect 177350 159248 177356 159300
rect 177408 159288 177414 159300
rect 179374 159288 179380 159300
rect 177408 159260 179380 159288
rect 177408 159248 177414 159260
rect 179374 159248 179380 159260
rect 179432 159248 179438 159300
rect 105774 158296 105780 158348
rect 105832 158336 105838 158348
rect 108718 158336 108724 158348
rect 105832 158308 108724 158336
rect 105832 158296 105838 158308
rect 108718 158296 108724 158308
rect 108776 158296 108782 158348
rect 177626 157956 177632 158008
rect 177684 157996 177690 158008
rect 180478 157996 180484 158008
rect 177684 157968 180484 157996
rect 177684 157956 177690 157968
rect 180478 157956 180484 157968
rect 180536 157956 180542 158008
rect 106142 157888 106148 157940
rect 106200 157928 106206 157940
rect 108626 157928 108632 157940
rect 106200 157900 108632 157928
rect 106200 157888 106206 157900
rect 108626 157888 108632 157900
rect 108684 157888 108690 157940
rect 178178 157888 178184 157940
rect 178236 157928 178242 157940
rect 180386 157928 180392 157940
rect 178236 157900 180392 157928
rect 178236 157888 178242 157900
rect 180386 157888 180392 157900
rect 180444 157888 180450 157940
rect 222798 156868 222804 156920
rect 222856 156908 222862 156920
rect 223534 156908 223540 156920
rect 222856 156880 223540 156908
rect 222856 156868 222862 156880
rect 223534 156868 223540 156880
rect 223592 156868 223598 156920
rect 106142 156664 106148 156716
rect 106200 156704 106206 156716
rect 108534 156704 108540 156716
rect 106200 156676 108540 156704
rect 106200 156664 106206 156676
rect 108534 156664 108540 156676
rect 108592 156664 108598 156716
rect 177350 156460 177356 156512
rect 177408 156500 177414 156512
rect 180294 156500 180300 156512
rect 177408 156472 180300 156500
rect 177408 156460 177414 156472
rect 180294 156460 180300 156472
rect 180352 156460 180358 156512
rect 105774 155304 105780 155356
rect 105832 155344 105838 155356
rect 107890 155344 107896 155356
rect 105832 155316 107896 155344
rect 105832 155304 105838 155316
rect 107890 155304 107896 155316
rect 107948 155304 107954 155356
rect 178086 155100 178092 155152
rect 178144 155140 178150 155152
rect 179650 155140 179656 155152
rect 178144 155112 179656 155140
rect 178144 155100 178150 155112
rect 179650 155100 179656 155112
rect 179708 155100 179714 155152
rect 57474 151496 57480 151548
rect 57532 151536 57538 151548
rect 59590 151536 59596 151548
rect 57532 151508 59596 151536
rect 57532 151496 57538 151508
rect 59590 151496 59596 151508
rect 59648 151496 59654 151548
rect 200534 151496 200540 151548
rect 200592 151536 200598 151548
rect 207342 151536 207348 151548
rect 200592 151508 207348 151536
rect 200592 151496 200598 151508
rect 207342 151496 207348 151508
rect 207400 151496 207406 151548
rect 105958 147008 105964 147060
rect 106016 147048 106022 147060
rect 108350 147048 108356 147060
rect 106016 147020 108356 147048
rect 106016 147008 106022 147020
rect 108350 147008 108356 147020
rect 108408 147008 108414 147060
rect 177350 146872 177356 146924
rect 177408 146912 177414 146924
rect 180570 146912 180576 146924
rect 177408 146884 180576 146912
rect 177408 146872 177414 146884
rect 180570 146872 180576 146884
rect 180628 146872 180634 146924
rect 178270 146124 178276 146176
rect 178328 146164 178334 146176
rect 179006 146164 179012 146176
rect 178328 146136 179012 146164
rect 178328 146124 178334 146136
rect 179006 146124 179012 146136
rect 179064 146124 179070 146176
rect 22238 145172 22244 145224
rect 22296 145212 22302 145224
rect 28678 145212 28684 145224
rect 22296 145184 28684 145212
rect 22296 145172 22302 145184
rect 28678 145172 28684 145184
rect 28736 145172 28742 145224
rect 207342 145172 207348 145224
rect 207400 145212 207406 145224
rect 210010 145212 210016 145224
rect 207400 145184 210016 145212
rect 207400 145172 207406 145184
rect 210010 145172 210016 145184
rect 210068 145212 210074 145224
rect 210286 145212 210292 145224
rect 210068 145184 210292 145212
rect 210068 145172 210074 145184
rect 210286 145172 210292 145184
rect 210344 145172 210350 145224
rect 178362 145104 178368 145156
rect 178420 145144 178426 145156
rect 181122 145144 181128 145156
rect 178420 145116 181128 145144
rect 178420 145104 178426 145116
rect 181122 145104 181128 145116
rect 181180 145104 181186 145156
rect 106694 144832 106700 144884
rect 106752 144872 106758 144884
rect 109270 144872 109276 144884
rect 106752 144844 109276 144872
rect 106752 144832 106758 144844
rect 109270 144832 109276 144844
rect 109328 144832 109334 144884
rect 191840 144696 191846 144748
rect 191898 144736 191904 144748
rect 194278 144736 194284 144748
rect 191898 144708 194284 144736
rect 191898 144696 191904 144708
rect 194278 144696 194284 144708
rect 194336 144696 194342 144748
rect 191472 144628 191478 144680
rect 191530 144668 191536 144680
rect 193634 144668 193640 144680
rect 191530 144640 193640 144668
rect 191530 144628 191536 144640
rect 193634 144628 193640 144640
rect 193692 144628 193698 144680
rect 197820 144628 197826 144680
rect 197878 144668 197884 144680
rect 202834 144668 202840 144680
rect 197878 144640 202840 144668
rect 197878 144628 197884 144640
rect 202834 144628 202840 144640
rect 202892 144628 202898 144680
rect 135490 144424 135496 144476
rect 135548 144464 135554 144476
rect 136318 144464 136324 144476
rect 135548 144436 136324 144464
rect 135548 144424 135554 144436
rect 136318 144424 136324 144436
rect 136376 144424 136382 144476
rect 125830 144220 125836 144272
rect 125888 144260 125894 144272
rect 131442 144260 131448 144272
rect 125888 144232 131448 144260
rect 125888 144220 125894 144232
rect 131442 144220 131448 144232
rect 131500 144220 131506 144272
rect 190598 144220 190604 144272
rect 190656 144260 190662 144272
rect 192530 144260 192536 144272
rect 190656 144232 192536 144260
rect 190656 144220 190662 144232
rect 192530 144220 192536 144232
rect 192588 144220 192594 144272
rect 198878 144220 198884 144272
rect 198936 144260 198942 144272
rect 203938 144260 203944 144272
rect 198936 144232 203944 144260
rect 198936 144220 198942 144232
rect 203938 144220 203944 144232
rect 203996 144220 204002 144272
rect 40638 144152 40644 144204
rect 40696 144192 40702 144204
rect 43030 144192 43036 144204
rect 40696 144164 43036 144192
rect 40696 144152 40702 144164
rect 43030 144152 43036 144164
rect 43088 144152 43094 144204
rect 54254 144152 54260 144204
rect 54312 144192 54318 144204
rect 59774 144192 59780 144204
rect 54312 144164 59780 144192
rect 54312 144152 54318 144164
rect 59774 144152 59780 144164
rect 59832 144152 59838 144204
rect 120218 144152 120224 144204
rect 120276 144192 120282 144204
rect 122334 144192 122340 144204
rect 120276 144164 122340 144192
rect 120276 144152 120282 144164
rect 122334 144152 122340 144164
rect 122392 144152 122398 144204
rect 126658 144152 126664 144204
rect 126716 144192 126722 144204
rect 132178 144192 132184 144204
rect 126716 144164 132184 144192
rect 126716 144152 126722 144164
rect 132178 144152 132184 144164
rect 132236 144152 132242 144204
rect 198510 144152 198516 144204
rect 198568 144192 198574 144204
rect 203386 144192 203392 144204
rect 198568 144164 203392 144192
rect 198568 144152 198574 144164
rect 203386 144152 203392 144164
rect 203444 144152 203450 144204
rect 41282 144084 41288 144136
rect 41340 144124 41346 144136
rect 43398 144124 43404 144136
rect 41340 144096 43404 144124
rect 41340 144084 41346 144096
rect 43398 144084 43404 144096
rect 43456 144084 43462 144136
rect 54622 144084 54628 144136
rect 54680 144124 54686 144136
rect 60418 144124 60424 144136
rect 54680 144096 60424 144124
rect 54680 144084 54686 144096
rect 60418 144084 60424 144096
rect 60476 144084 60482 144136
rect 105222 144084 105228 144136
rect 105280 144124 105286 144136
rect 105958 144124 105964 144136
rect 105280 144096 105964 144124
rect 105280 144084 105286 144096
rect 105958 144084 105964 144096
rect 106016 144084 106022 144136
rect 106510 144084 106516 144136
rect 106568 144124 106574 144136
rect 107154 144124 107160 144136
rect 106568 144096 107160 144124
rect 106568 144084 106574 144096
rect 107154 144084 107160 144096
rect 107212 144084 107218 144136
rect 118930 144084 118936 144136
rect 118988 144124 118994 144136
rect 120586 144124 120592 144136
rect 118988 144096 120592 144124
rect 118988 144084 118994 144096
rect 120586 144084 120592 144096
rect 120644 144084 120650 144136
rect 126290 144084 126296 144136
rect 126348 144124 126354 144136
rect 131626 144124 131632 144136
rect 126348 144096 131632 144124
rect 126348 144084 126354 144096
rect 131626 144084 131632 144096
rect 131684 144084 131690 144136
rect 132638 144084 132644 144136
rect 132696 144124 132702 144136
rect 174130 144124 174136 144136
rect 132696 144096 174136 144124
rect 132696 144084 132702 144096
rect 174130 144084 174136 144096
rect 174188 144084 174194 144136
rect 197498 144084 197504 144136
rect 197556 144124 197562 144136
rect 202190 144124 202196 144136
rect 197556 144096 202196 144124
rect 197556 144084 197562 144096
rect 202190 144084 202196 144096
rect 202248 144084 202254 144136
rect 132638 143444 132644 143456
rect 132599 143416 132644 143444
rect 132638 143404 132644 143416
rect 132696 143404 132702 143456
rect 34106 142656 34112 142708
rect 34164 142696 34170 142708
rect 39074 142696 39080 142708
rect 34164 142668 39080 142696
rect 34164 142656 34170 142668
rect 39074 142656 39080 142668
rect 39132 142656 39138 142708
rect 39258 142656 39264 142708
rect 39316 142696 39322 142708
rect 42202 142696 42208 142708
rect 39316 142668 42208 142696
rect 39316 142656 39322 142668
rect 42202 142656 42208 142668
rect 42260 142656 42266 142708
rect 43398 142656 43404 142708
rect 43456 142696 43462 142708
rect 44594 142696 44600 142708
rect 43456 142668 44600 142696
rect 43456 142656 43462 142668
rect 44594 142656 44600 142668
rect 44652 142656 44658 142708
rect 48274 142656 48280 142708
rect 48332 142696 48338 142708
rect 49470 142696 49476 142708
rect 48332 142668 49476 142696
rect 48332 142656 48338 142668
rect 49470 142656 49476 142668
rect 49528 142656 49534 142708
rect 51034 142656 51040 142708
rect 51092 142696 51098 142708
rect 53705 142699 53763 142705
rect 53705 142696 53717 142699
rect 51092 142668 53717 142696
rect 51092 142656 51098 142668
rect 53705 142665 53717 142668
rect 53751 142665 53763 142699
rect 53705 142659 53763 142665
rect 53794 142656 53800 142708
rect 53852 142696 53858 142708
rect 58670 142696 58676 142708
rect 53852 142668 58676 142696
rect 53852 142656 53858 142668
rect 58670 142656 58676 142668
rect 58728 142656 58734 142708
rect 62810 142656 62816 142708
rect 62868 142696 62874 142708
rect 62868 142668 65156 142696
rect 62868 142656 62874 142668
rect 16718 142588 16724 142640
rect 16776 142628 16782 142640
rect 31898 142628 31904 142640
rect 16776 142600 31904 142628
rect 16776 142588 16782 142600
rect 31898 142588 31904 142600
rect 31956 142588 31962 142640
rect 34658 142588 34664 142640
rect 34716 142628 34722 142640
rect 39442 142628 39448 142640
rect 34716 142600 39448 142628
rect 34716 142588 34722 142600
rect 39442 142588 39448 142600
rect 39500 142588 39506 142640
rect 42662 142588 42668 142640
rect 42720 142628 42726 142640
rect 44226 142628 44232 142640
rect 42720 142600 44232 142628
rect 42720 142588 42726 142600
rect 44226 142588 44232 142600
rect 44284 142588 44290 142640
rect 47814 142588 47820 142640
rect 47872 142628 47878 142640
rect 48826 142628 48832 142640
rect 47872 142600 48832 142628
rect 47872 142588 47878 142600
rect 48826 142588 48832 142600
rect 48884 142588 48890 142640
rect 49746 142588 49752 142640
rect 49804 142628 49810 142640
rect 51586 142628 51592 142640
rect 49804 142600 51592 142628
rect 49804 142588 49810 142600
rect 51586 142588 51592 142600
rect 51644 142588 51650 142640
rect 53058 142588 53064 142640
rect 53116 142628 53122 142640
rect 57658 142628 57664 142640
rect 53116 142600 57664 142628
rect 53116 142588 53122 142600
rect 57658 142588 57664 142600
rect 57716 142588 57722 142640
rect 37234 142520 37240 142572
rect 37292 142560 37298 142572
rect 41006 142560 41012 142572
rect 37292 142532 41012 142560
rect 37292 142520 37298 142532
rect 41006 142520 41012 142532
rect 41064 142520 41070 142572
rect 50206 142520 50212 142572
rect 50264 142560 50270 142572
rect 52966 142560 52972 142572
rect 50264 142532 52972 142560
rect 50264 142520 50270 142532
rect 52966 142520 52972 142532
rect 53024 142520 53030 142572
rect 53426 142520 53432 142572
rect 53484 142560 53490 142572
rect 58118 142560 58124 142572
rect 53484 142532 58124 142560
rect 53484 142520 53490 142532
rect 58118 142520 58124 142532
rect 58176 142520 58182 142572
rect 65128 142560 65156 142668
rect 66490 142656 66496 142708
rect 66548 142696 66554 142708
rect 67870 142696 67876 142708
rect 66548 142668 67876 142696
rect 66548 142656 66554 142668
rect 67870 142656 67876 142668
rect 67928 142656 67934 142708
rect 72838 142656 72844 142708
rect 72896 142696 72902 142708
rect 74494 142696 74500 142708
rect 72896 142668 74500 142696
rect 72896 142656 72902 142668
rect 74494 142656 74500 142668
rect 74552 142656 74558 142708
rect 74770 142656 74776 142708
rect 74828 142696 74834 142708
rect 75598 142696 75604 142708
rect 74828 142668 75604 142696
rect 74828 142656 74834 142668
rect 75598 142656 75604 142668
rect 75656 142656 75662 142708
rect 80106 142656 80112 142708
rect 80164 142696 80170 142708
rect 81670 142696 81676 142708
rect 80164 142668 81676 142696
rect 80164 142656 80170 142668
rect 81670 142656 81676 142668
rect 81728 142656 81734 142708
rect 84522 142656 84528 142708
rect 84580 142696 84586 142708
rect 89122 142696 89128 142708
rect 84580 142668 89128 142696
rect 84580 142656 84586 142668
rect 89122 142656 89128 142668
rect 89180 142656 89186 142708
rect 95470 142656 95476 142708
rect 95528 142696 95534 142708
rect 96758 142696 96764 142708
rect 95528 142668 96764 142696
rect 95528 142656 95534 142668
rect 96758 142656 96764 142668
rect 96816 142656 96822 142708
rect 110098 142656 110104 142708
rect 110156 142696 110162 142708
rect 111110 142696 111116 142708
rect 110156 142668 111116 142696
rect 110156 142656 110162 142668
rect 111110 142656 111116 142668
rect 111168 142656 111174 142708
rect 120678 142656 120684 142708
rect 120736 142696 120742 142708
rect 123438 142696 123444 142708
rect 120736 142668 123444 142696
rect 120736 142656 120742 142668
rect 123438 142656 123444 142668
rect 123496 142656 123502 142708
rect 125462 142656 125468 142708
rect 125520 142696 125526 142708
rect 130430 142696 130436 142708
rect 125520 142668 130436 142696
rect 125520 142656 125526 142668
rect 130430 142656 130436 142668
rect 130488 142656 130494 142708
rect 153246 142656 153252 142708
rect 153304 142696 153310 142708
rect 155822 142696 155828 142708
rect 153304 142668 155828 142696
rect 153304 142656 153310 142668
rect 155822 142656 155828 142668
rect 155880 142656 155886 142708
rect 156558 142656 156564 142708
rect 156616 142696 156622 142708
rect 161434 142696 161440 142708
rect 156616 142668 161440 142696
rect 156616 142656 156622 142668
rect 161434 142656 161440 142668
rect 161492 142656 161498 142708
rect 182226 142656 182232 142708
rect 182284 142696 182290 142708
rect 183238 142696 183244 142708
rect 182284 142668 183244 142696
rect 182284 142656 182290 142668
rect 183238 142656 183244 142668
rect 183296 142656 183302 142708
rect 189678 142656 189684 142708
rect 189736 142696 189742 142708
rect 190782 142696 190788 142708
rect 189736 142668 190788 142696
rect 189736 142656 189742 142668
rect 190782 142656 190788 142668
rect 190840 142656 190846 142708
rect 191334 142656 191340 142708
rect 191392 142696 191398 142708
rect 193082 142696 193088 142708
rect 191392 142668 193088 142696
rect 191392 142656 191398 142668
rect 193082 142656 193088 142668
rect 193140 142656 193146 142708
rect 196486 142656 196492 142708
rect 196544 142696 196550 142708
rect 200534 142696 200540 142708
rect 196544 142668 200540 142696
rect 196544 142656 196550 142668
rect 200534 142656 200540 142668
rect 200592 142656 200598 142708
rect 200994 142656 201000 142708
rect 201052 142696 201058 142708
rect 215898 142696 215904 142708
rect 201052 142668 215904 142696
rect 201052 142656 201058 142668
rect 215898 142656 215904 142668
rect 215956 142656 215962 142708
rect 81210 142588 81216 142640
rect 81268 142628 81274 142640
rect 83510 142628 83516 142640
rect 81268 142600 83516 142628
rect 81268 142588 81274 142600
rect 83510 142588 83516 142600
rect 83568 142588 83574 142640
rect 86730 142588 86736 142640
rect 86788 142628 86794 142640
rect 92802 142628 92808 142640
rect 86788 142600 92808 142628
rect 86788 142588 86794 142600
rect 92802 142588 92808 142600
rect 92860 142588 92866 142640
rect 119114 142588 119120 142640
rect 119172 142628 119178 142640
rect 121138 142628 121144 142640
rect 119172 142600 121144 142628
rect 119172 142588 119178 142600
rect 121138 142588 121144 142600
rect 121196 142588 121202 142640
rect 123898 142588 123904 142640
rect 123956 142628 123962 142640
rect 128130 142628 128136 142640
rect 123956 142600 128136 142628
rect 123956 142588 123962 142600
rect 128130 142588 128136 142600
rect 128188 142588 128194 142640
rect 154350 142588 154356 142640
rect 154408 142628 154414 142640
rect 157662 142628 157668 142640
rect 154408 142600 157668 142628
rect 154408 142588 154414 142600
rect 157662 142588 157668 142600
rect 157720 142588 157726 142640
rect 163274 142588 163280 142640
rect 163332 142628 163338 142640
rect 174406 142628 174412 142640
rect 163332 142600 174412 142628
rect 163332 142588 163338 142600
rect 174406 142588 174412 142600
rect 174464 142588 174470 142640
rect 189310 142588 189316 142640
rect 189368 142628 189374 142640
rect 190230 142628 190236 142640
rect 189368 142600 190236 142628
rect 189368 142588 189374 142600
rect 190230 142588 190236 142600
rect 190288 142588 190294 142640
rect 190506 142588 190512 142640
rect 190564 142628 190570 142640
rect 191978 142628 191984 142640
rect 190564 142600 191984 142628
rect 190564 142588 190570 142600
rect 191978 142588 191984 142600
rect 192036 142588 192042 142640
rect 194094 142588 194100 142640
rect 194152 142628 194158 142640
rect 197130 142628 197136 142640
rect 194152 142600 197136 142628
rect 194152 142588 194158 142600
rect 197130 142588 197136 142600
rect 197188 142588 197194 142640
rect 71182 142560 71188 142572
rect 65128 142532 71188 142560
rect 71182 142520 71188 142532
rect 71240 142520 71246 142572
rect 121046 142520 121052 142572
rect 121104 142560 121110 142572
rect 124450 142560 124456 142572
rect 121104 142532 124456 142560
rect 121104 142520 121110 142532
rect 124450 142520 124456 142532
rect 124508 142520 124514 142572
rect 124634 142520 124640 142572
rect 124692 142560 124698 142572
rect 129326 142560 129332 142572
rect 124692 142532 129332 142560
rect 124692 142520 124698 142532
rect 129326 142520 129332 142532
rect 129384 142520 129390 142572
rect 134110 142520 134116 142572
rect 134168 142560 134174 142572
rect 143218 142560 143224 142572
rect 134168 142532 143224 142560
rect 134168 142520 134174 142532
rect 143218 142520 143224 142532
rect 143276 142520 143282 142572
rect 155454 142520 155460 142572
rect 155512 142560 155518 142572
rect 159502 142560 159508 142572
rect 155512 142532 159508 142560
rect 155512 142520 155518 142532
rect 159502 142520 159508 142532
rect 159560 142520 159566 142572
rect 181674 142520 181680 142572
rect 181732 142560 181738 142572
rect 182778 142560 182784 142572
rect 181732 142532 182784 142560
rect 181732 142520 181738 142532
rect 182778 142520 182784 142532
rect 182836 142520 182842 142572
rect 193726 142520 193732 142572
rect 193784 142560 193790 142572
rect 196486 142560 196492 142572
rect 193784 142532 196492 142560
rect 193784 142520 193790 142532
rect 196486 142520 196492 142532
rect 196544 142520 196550 142572
rect 27574 142452 27580 142504
rect 27632 142492 27638 142504
rect 27632 142464 50344 142492
rect 27632 142452 27638 142464
rect 36590 142384 36596 142436
rect 36648 142424 36654 142436
rect 40362 142424 40368 142436
rect 36648 142396 40368 142424
rect 36648 142384 36654 142396
rect 40362 142384 40368 142396
rect 40420 142384 40426 142436
rect 48642 142384 48648 142436
rect 48700 142424 48706 142436
rect 50206 142424 50212 142436
rect 48700 142396 50212 142424
rect 48700 142384 48706 142396
rect 50206 142384 50212 142396
rect 50264 142384 50270 142436
rect 50316 142424 50344 142464
rect 50666 142452 50672 142504
rect 50724 142492 50730 142504
rect 53610 142492 53616 142504
rect 50724 142464 53616 142492
rect 50724 142452 50730 142464
rect 53610 142452 53616 142464
rect 53668 142452 53674 142504
rect 53705 142495 53763 142501
rect 53705 142461 53717 142495
rect 53751 142492 53763 142495
rect 54254 142492 54260 142504
rect 53751 142464 54260 142492
rect 53751 142461 53763 142464
rect 53705 142455 53763 142461
rect 54254 142452 54260 142464
rect 54312 142452 54318 142504
rect 102278 142452 102284 142504
rect 102336 142492 102342 142504
rect 174314 142492 174320 142504
rect 102336 142464 174320 142492
rect 102336 142452 102342 142464
rect 174314 142452 174320 142464
rect 174372 142452 174378 142504
rect 194554 142452 194560 142504
rect 194612 142492 194618 142504
rect 197682 142492 197688 142504
rect 194612 142464 197688 142492
rect 194612 142452 194618 142464
rect 197682 142452 197688 142464
rect 197740 142452 197746 142504
rect 52141 142427 52199 142433
rect 52141 142424 52153 142427
rect 50316 142396 52153 142424
rect 52141 142393 52153 142396
rect 52187 142393 52199 142427
rect 52141 142387 52199 142393
rect 52230 142384 52236 142436
rect 52288 142424 52294 142436
rect 56094 142424 56100 142436
rect 52288 142396 56100 142424
rect 52288 142384 52294 142396
rect 56094 142384 56100 142396
rect 56152 142384 56158 142436
rect 69158 142384 69164 142436
rect 69216 142424 69222 142436
rect 72286 142424 72292 142436
rect 69216 142396 72292 142424
rect 69216 142384 69222 142396
rect 72286 142384 72292 142396
rect 72344 142384 72350 142436
rect 85626 142384 85632 142436
rect 85684 142424 85690 142436
rect 90962 142424 90968 142436
rect 85684 142396 90968 142424
rect 85684 142384 85690 142396
rect 90962 142384 90968 142396
rect 91020 142384 91026 142436
rect 117458 142384 117464 142436
rect 117516 142424 117522 142436
rect 118838 142424 118844 142436
rect 117516 142396 118844 142424
rect 117516 142384 117522 142396
rect 118838 142384 118844 142396
rect 118896 142384 118902 142436
rect 119482 142384 119488 142436
rect 119540 142424 119546 142436
rect 121690 142424 121696 142436
rect 119540 142396 121696 142424
rect 119540 142384 119546 142396
rect 121690 142384 121696 142396
rect 121748 142384 121754 142436
rect 124266 142384 124272 142436
rect 124324 142424 124330 142436
rect 128682 142424 128688 142436
rect 124324 142396 128688 142424
rect 124324 142384 124330 142396
rect 128682 142384 128688 142396
rect 128740 142384 128746 142436
rect 159870 142384 159876 142436
rect 159928 142424 159934 142436
rect 167046 142424 167052 142436
rect 159928 142396 167052 142424
rect 159928 142384 159934 142396
rect 167046 142384 167052 142396
rect 167104 142384 167110 142436
rect 192898 142384 192904 142436
rect 192956 142424 192962 142436
rect 195382 142424 195388 142436
rect 192956 142396 195388 142424
rect 192956 142384 192962 142396
rect 195382 142384 195388 142396
rect 195440 142384 195446 142436
rect 195750 142384 195756 142436
rect 195808 142424 195814 142436
rect 199062 142424 199068 142436
rect 195808 142396 199068 142424
rect 195808 142384 195814 142396
rect 199062 142384 199068 142396
rect 199120 142384 199126 142436
rect 51862 142316 51868 142368
rect 51920 142356 51926 142368
rect 55358 142356 55364 142368
rect 51920 142328 55364 142356
rect 51920 142316 51926 142328
rect 55358 142316 55364 142328
rect 55416 142316 55422 142368
rect 98966 142316 98972 142368
rect 99024 142356 99030 142368
rect 102278 142356 102284 142368
rect 99024 142328 102284 142356
rect 99024 142316 99030 142328
rect 102278 142316 102284 142328
rect 102336 142316 102342 142368
rect 123714 142316 123720 142368
rect 123772 142356 123778 142368
rect 127578 142356 127584 142368
rect 123772 142328 127584 142356
rect 123772 142316 123778 142328
rect 127578 142316 127584 142328
rect 127636 142316 127642 142368
rect 160974 142316 160980 142368
rect 161032 142356 161038 142368
rect 168886 142356 168892 142368
rect 161032 142328 168892 142356
rect 161032 142316 161038 142328
rect 168886 142316 168892 142328
rect 168944 142316 168950 142368
rect 192438 142316 192444 142368
rect 192496 142356 192502 142368
rect 194830 142356 194836 142368
rect 192496 142328 194836 142356
rect 192496 142316 192502 142328
rect 194830 142316 194836 142328
rect 194888 142316 194894 142368
rect 196946 142316 196952 142368
rect 197004 142356 197010 142368
rect 201086 142356 201092 142368
rect 197004 142328 201092 142356
rect 197004 142316 197010 142328
rect 201086 142316 201092 142328
rect 201144 142316 201150 142368
rect 31898 142248 31904 142300
rect 31956 142288 31962 142300
rect 31956 142260 37832 142288
rect 31956 142248 31962 142260
rect 37804 142084 37832 142260
rect 39994 142248 40000 142300
rect 40052 142288 40058 142300
rect 42294 142288 42300 142300
rect 40052 142260 42300 142288
rect 40052 142248 40058 142260
rect 42294 142248 42300 142260
rect 42352 142248 42358 142300
rect 51313 142291 51371 142297
rect 51313 142288 51325 142291
rect 46452 142260 51325 142288
rect 38614 142180 38620 142232
rect 38672 142220 38678 142232
rect 41834 142220 41840 142232
rect 38672 142192 41840 142220
rect 38672 142180 38678 142192
rect 41834 142180 41840 142192
rect 41892 142180 41898 142232
rect 37878 142112 37884 142164
rect 37936 142152 37942 142164
rect 41466 142152 41472 142164
rect 37936 142124 41472 142152
rect 37936 142112 37942 142124
rect 41466 142112 41472 142124
rect 41524 142112 41530 142164
rect 42018 142112 42024 142164
rect 42076 142152 42082 142164
rect 43858 142152 43864 142164
rect 42076 142124 43864 142152
rect 42076 142112 42082 142124
rect 43858 142112 43864 142124
rect 43916 142112 43922 142164
rect 46452 142084 46480 142260
rect 51313 142257 51325 142260
rect 51359 142257 51371 142291
rect 51313 142251 51371 142257
rect 51402 142248 51408 142300
rect 51460 142288 51466 142300
rect 54990 142288 54996 142300
rect 51460 142260 54996 142288
rect 51460 142248 51466 142260
rect 54990 142248 54996 142260
rect 55048 142248 55054 142300
rect 62350 142248 62356 142300
rect 62408 142288 62414 142300
rect 63454 142288 63460 142300
rect 62408 142260 63460 142288
rect 62408 142248 62414 142260
rect 63454 142248 63460 142260
rect 63512 142248 63518 142300
rect 116630 142248 116636 142300
rect 116688 142288 116694 142300
rect 117642 142288 117648 142300
rect 116688 142260 117648 142288
rect 116688 142248 116694 142260
rect 117642 142248 117648 142260
rect 117700 142248 117706 142300
rect 120310 142248 120316 142300
rect 120368 142288 120374 142300
rect 123070 142288 123076 142300
rect 120368 142260 123076 142288
rect 120368 142248 120374 142260
rect 123070 142248 123076 142260
rect 123128 142248 123134 142300
rect 125094 142248 125100 142300
rect 125152 142288 125158 142300
rect 129878 142288 129884 142300
rect 125152 142260 129884 142288
rect 125152 142248 125158 142260
rect 129878 142248 129884 142260
rect 129936 142248 129942 142300
rect 167690 142248 167696 142300
rect 167748 142288 167754 142300
rect 174314 142288 174320 142300
rect 167748 142260 174320 142288
rect 167748 142248 167754 142260
rect 174314 142248 174320 142260
rect 174372 142248 174378 142300
rect 182870 142248 182876 142300
rect 182928 142288 182934 142300
rect 183606 142288 183612 142300
rect 182928 142260 183612 142288
rect 182928 142248 182934 142260
rect 183606 142248 183612 142260
rect 183664 142248 183670 142300
rect 193358 142248 193364 142300
rect 193416 142288 193422 142300
rect 195934 142288 195940 142300
rect 193416 142260 195940 142288
rect 193416 142248 193422 142260
rect 195934 142248 195940 142260
rect 195992 142248 195998 142300
rect 197314 142248 197320 142300
rect 197372 142288 197378 142300
rect 201638 142288 201644 142300
rect 197372 142260 201644 142288
rect 197372 142248 197378 142260
rect 201638 142248 201644 142260
rect 201696 142248 201702 142300
rect 49010 142180 49016 142232
rect 49068 142220 49074 142232
rect 50850 142220 50856 142232
rect 49068 142192 50856 142220
rect 49068 142180 49074 142192
rect 50850 142180 50856 142192
rect 50908 142180 50914 142232
rect 52230 142220 52236 142232
rect 51236 142192 52236 142220
rect 37804 142056 46480 142084
rect 49838 142044 49844 142096
rect 49896 142084 49902 142096
rect 51236 142084 51264 142192
rect 52230 142180 52236 142192
rect 52288 142180 52294 142232
rect 121506 142180 121512 142232
rect 121564 142220 121570 142232
rect 124634 142220 124640 142232
rect 121564 142192 124640 142220
rect 121564 142180 121570 142192
rect 124634 142180 124640 142192
rect 124692 142180 124698 142232
rect 134478 142180 134484 142232
rect 134536 142220 134542 142232
rect 135490 142220 135496 142232
rect 134536 142192 135496 142220
rect 134536 142180 134542 142192
rect 135490 142180 135496 142192
rect 135548 142180 135554 142232
rect 142666 142180 142672 142232
rect 142724 142220 142730 142232
rect 145426 142220 145432 142232
rect 142724 142192 145432 142220
rect 142724 142180 142730 142192
rect 145426 142180 145432 142192
rect 145484 142180 145490 142232
rect 172106 142180 172112 142232
rect 172164 142220 172170 142232
rect 175234 142220 175240 142232
rect 172164 142192 175240 142220
rect 172164 142180 172170 142192
rect 175234 142180 175240 142192
rect 175292 142180 175298 142232
rect 196118 142180 196124 142232
rect 196176 142220 196182 142232
rect 199614 142220 199620 142232
rect 196176 142192 199620 142220
rect 196176 142180 196182 142192
rect 199614 142180 199620 142192
rect 199672 142180 199678 142232
rect 52141 142155 52199 142161
rect 52141 142121 52153 142155
rect 52187 142152 52199 142155
rect 54898 142152 54904 142164
rect 52187 142124 54904 142152
rect 52187 142121 52199 142124
rect 52141 142115 52199 142121
rect 54898 142112 54904 142124
rect 54956 142112 54962 142164
rect 63454 142112 63460 142164
rect 63512 142152 63518 142164
rect 64558 142152 64564 142164
rect 63512 142124 64564 142152
rect 63512 142112 63518 142124
rect 64558 142112 64564 142124
rect 64616 142112 64622 142164
rect 87834 142112 87840 142164
rect 87892 142152 87898 142164
rect 94734 142152 94740 142164
rect 87892 142124 94740 142152
rect 87892 142112 87898 142124
rect 94734 142112 94740 142124
rect 94792 142112 94798 142164
rect 117090 142112 117096 142164
rect 117148 142152 117154 142164
rect 118194 142152 118200 142164
rect 117148 142124 118200 142152
rect 117148 142112 117154 142124
rect 118194 142112 118200 142124
rect 118252 142112 118258 142164
rect 118286 142112 118292 142164
rect 118344 142152 118350 142164
rect 119942 142152 119948 142164
rect 118344 142124 119948 142152
rect 118344 142112 118350 142124
rect 119942 142112 119948 142124
rect 120000 142112 120006 142164
rect 123346 142112 123352 142164
rect 123404 142152 123410 142164
rect 126934 142152 126940 142164
rect 123404 142124 126940 142152
rect 123404 142112 123410 142124
rect 126934 142112 126940 142124
rect 126992 142112 126998 142164
rect 158766 142112 158772 142164
rect 158824 142152 158830 142164
rect 165114 142152 165120 142164
rect 158824 142124 165120 142152
rect 158824 142112 158830 142124
rect 165114 142112 165120 142124
rect 165172 142112 165178 142164
rect 166586 142112 166592 142164
rect 166644 142152 166650 142164
rect 175418 142152 175424 142164
rect 166644 142124 175424 142152
rect 166644 142112 166650 142124
rect 175418 142112 175424 142124
rect 175476 142112 175482 142164
rect 194646 142112 194652 142164
rect 194704 142152 194710 142164
rect 198234 142152 198240 142164
rect 194704 142124 198240 142152
rect 194704 142112 194710 142124
rect 198234 142112 198240 142124
rect 198292 142112 198298 142164
rect 49896 142056 51264 142084
rect 51313 142087 51371 142093
rect 49896 142044 49902 142056
rect 51313 142053 51325 142087
rect 51359 142084 51371 142087
rect 57474 142084 57480 142096
rect 51359 142056 57480 142084
rect 51359 142053 51371 142056
rect 51313 142047 51371 142053
rect 57474 142044 57480 142056
rect 57532 142044 57538 142096
rect 134570 142044 134576 142096
rect 134628 142084 134634 142096
rect 135582 142084 135588 142096
rect 134628 142056 135588 142084
rect 134628 142044 134634 142056
rect 135582 142044 135588 142056
rect 135640 142044 135646 142096
rect 165482 142044 165488 142096
rect 165540 142084 165546 142096
rect 175142 142084 175148 142096
rect 165540 142056 175148 142084
rect 165540 142044 165546 142056
rect 175142 142044 175148 142056
rect 175200 142044 175206 142096
rect 195290 142044 195296 142096
rect 195348 142084 195354 142096
rect 198786 142084 198792 142096
rect 195348 142056 198792 142084
rect 195348 142044 195354 142056
rect 198786 142044 198792 142056
rect 198844 142044 198850 142096
rect 222522 142044 222528 142096
rect 222580 142084 222586 142096
rect 222798 142084 222804 142096
rect 222580 142056 222804 142084
rect 222580 142044 222586 142056
rect 222798 142044 222804 142056
rect 222856 142044 222862 142096
rect 52598 141976 52604 142028
rect 52656 142016 52662 142028
rect 57014 142016 57020 142028
rect 52656 141988 57020 142016
rect 52656 141976 52662 141988
rect 57014 141976 57020 141988
rect 57072 141976 57078 142028
rect 83418 141976 83424 142028
rect 83476 142016 83482 142028
rect 87282 142016 87288 142028
rect 83476 141988 87288 142016
rect 83476 141976 83482 141988
rect 87282 141976 87288 141988
rect 87340 141976 87346 142028
rect 88938 141976 88944 142028
rect 88996 142016 89002 142028
rect 96850 142016 96856 142028
rect 88996 141988 96856 142016
rect 88996 141976 89002 141988
rect 96850 141976 96856 141988
rect 96908 141976 96914 142028
rect 100070 141976 100076 142028
rect 100128 142016 100134 142028
rect 103106 142016 103112 142028
rect 100128 141988 103112 142016
rect 100128 141976 100134 141988
rect 103106 141976 103112 141988
rect 103164 141976 103170 142028
rect 110420 141976 110426 142028
rect 110478 142016 110484 142028
rect 111478 142016 111484 142028
rect 110478 141988 111484 142016
rect 110478 141976 110484 141988
rect 111478 141976 111484 141988
rect 111536 141976 111542 142028
rect 113272 141976 113278 142028
rect 113330 142016 113336 142028
rect 113502 142016 113508 142028
rect 113330 141988 113508 142016
rect 113330 141976 113336 141988
rect 113502 141976 113508 141988
rect 113560 141976 113566 142028
rect 116262 141976 116268 142028
rect 116320 142016 116326 142028
rect 117412 142016 117418 142028
rect 116320 141988 117418 142016
rect 116320 141976 116326 141988
rect 117412 141976 117418 141988
rect 117470 141976 117476 142028
rect 117826 141976 117832 142028
rect 117884 142016 117890 142028
rect 119712 142016 119718 142028
rect 117884 141988 119718 142016
rect 117884 141976 117890 141988
rect 119712 141976 119718 141988
rect 119770 141976 119776 142028
rect 121874 141976 121880 142028
rect 121932 142016 121938 142028
rect 125508 142016 125514 142028
rect 121932 141988 125514 142016
rect 121932 141976 121938 141988
rect 125508 141976 125514 141988
rect 125566 141976 125572 142028
rect 134294 141976 134300 142028
rect 134352 142016 134358 142028
rect 136870 142016 136876 142028
rect 134352 141988 136876 142016
rect 134352 141976 134358 141988
rect 136870 141976 136876 141988
rect 136928 141976 136934 142028
rect 168794 141976 168800 142028
rect 168852 142016 168858 142028
rect 172842 142016 172848 142028
rect 168852 141988 172848 142016
rect 168852 141976 168858 141988
rect 172842 141976 172848 141988
rect 172900 141976 172906 142028
rect 190138 141976 190144 142028
rect 190196 142016 190202 142028
rect 191426 142016 191432 142028
rect 190196 141988 191432 142016
rect 190196 141976 190202 141988
rect 191426 141976 191432 141988
rect 191484 141976 191490 142028
rect 207986 141976 207992 142028
rect 208044 142016 208050 142028
rect 221234 142016 221240 142028
rect 208044 141988 221240 142016
rect 208044 141976 208050 141988
rect 221234 141976 221240 141988
rect 221292 141976 221298 142028
rect 101174 141908 101180 141960
rect 101232 141948 101238 141960
rect 173210 141948 173216 141960
rect 101232 141920 173216 141948
rect 101232 141908 101238 141920
rect 173210 141908 173216 141920
rect 173268 141908 173274 141960
rect 207894 141908 207900 141960
rect 207952 141948 207958 141960
rect 210010 141948 210016 141960
rect 207952 141920 210016 141948
rect 207952 141908 207958 141920
rect 210010 141908 210016 141920
rect 210068 141908 210074 141960
rect 222522 141908 222528 141960
rect 222580 141948 222586 141960
rect 223534 141948 223540 141960
rect 222580 141920 223540 141948
rect 222580 141908 222586 141920
rect 223534 141908 223540 141920
rect 223592 141908 223598 141960
rect 70998 141840 71004 141892
rect 71056 141880 71062 141892
rect 73390 141880 73396 141892
rect 71056 141852 73396 141880
rect 71056 141840 71062 141852
rect 73390 141840 73396 141852
rect 73448 141840 73454 141892
rect 132362 141840 132368 141892
rect 132420 141880 132426 141892
rect 132420 141852 132684 141880
rect 132420 141840 132426 141852
rect 122886 141772 122892 141824
rect 122944 141812 122950 141824
rect 126382 141812 126388 141824
rect 122944 141784 126388 141812
rect 122944 141772 122950 141784
rect 126382 141772 126388 141784
rect 126440 141772 126446 141824
rect 35578 141704 35584 141756
rect 35636 141744 35642 141756
rect 39810 141744 39816 141756
rect 35636 141716 39816 141744
rect 35636 141704 35642 141716
rect 39810 141704 39816 141716
rect 39868 141704 39874 141756
rect 122242 141704 122248 141756
rect 122300 141744 122306 141756
rect 125830 141744 125836 141756
rect 122300 141716 125836 141744
rect 122300 141704 122306 141716
rect 125830 141704 125836 141716
rect 125888 141704 125894 141756
rect 35946 141636 35952 141688
rect 36004 141636 36010 141688
rect 40178 141636 40184 141688
rect 40236 141636 40242 141688
rect 35964 141336 35992 141636
rect 40196 141336 40224 141636
rect 82314 141500 82320 141552
rect 82372 141540 82378 141552
rect 85350 141540 85356 141552
rect 82372 141512 85356 141540
rect 82372 141500 82378 141512
rect 85350 141500 85356 141512
rect 85408 141500 85414 141552
rect 132656 141348 132684 141852
rect 152142 141772 152148 141824
rect 152200 141812 152206 141824
rect 153890 141812 153896 141824
rect 152200 141784 153896 141812
rect 152200 141772 152206 141784
rect 153890 141772 153896 141784
rect 153948 141772 153954 141824
rect 144506 141636 144512 141688
rect 144564 141676 144570 141688
rect 146530 141676 146536 141688
rect 144564 141648 146536 141676
rect 144564 141636 144570 141648
rect 146530 141636 146536 141648
rect 146588 141636 146594 141688
rect 157938 141568 157944 141620
rect 157996 141608 158002 141620
rect 163274 141608 163280 141620
rect 157996 141580 163280 141608
rect 157996 141568 158002 141580
rect 163274 141568 163280 141580
rect 163332 141568 163338 141620
rect 146438 141500 146444 141552
rect 146496 141540 146502 141552
rect 147634 141540 147640 141552
rect 146496 141512 147640 141540
rect 146496 141500 146502 141512
rect 147634 141500 147640 141512
rect 147692 141500 147698 141552
rect 151038 141500 151044 141552
rect 151096 141540 151102 141552
rect 152050 141540 152056 141552
rect 151096 141512 152056 141540
rect 151096 141500 151102 141512
rect 152050 141500 152056 141512
rect 152108 141500 152114 141552
rect 169898 141364 169904 141416
rect 169956 141404 169962 141416
rect 169956 141376 172888 141404
rect 169956 141364 169962 141376
rect 35964 141308 40224 141336
rect 90134 141296 90140 141348
rect 90192 141336 90198 141348
rect 91241 141339 91299 141345
rect 91241 141336 91253 141339
rect 90192 141308 91253 141336
rect 90192 141296 90198 141308
rect 91241 141305 91253 141308
rect 91287 141305 91299 141339
rect 91241 141299 91299 141305
rect 91333 141339 91391 141345
rect 91333 141305 91345 141339
rect 91379 141336 91391 141339
rect 92342 141336 92348 141348
rect 91379 141308 92348 141336
rect 91379 141305 91391 141308
rect 91333 141299 91391 141305
rect 92342 141296 92348 141308
rect 92400 141296 92406 141348
rect 92713 141339 92771 141345
rect 92713 141305 92725 141339
rect 92759 141336 92771 141339
rect 93446 141336 93452 141348
rect 92759 141308 93452 141336
rect 92759 141305 92771 141308
rect 92713 141299 92771 141305
rect 93446 141296 93452 141308
rect 93504 141296 93510 141348
rect 97862 141296 97868 141348
rect 97920 141336 97926 141348
rect 97920 141308 100944 141336
rect 97920 141296 97926 141308
rect 62810 141228 62816 141280
rect 62868 141268 62874 141280
rect 69250 141268 69256 141280
rect 62868 141240 69256 141268
rect 62868 141228 62874 141240
rect 69250 141228 69256 141240
rect 69308 141228 69314 141280
rect 62718 141160 62724 141212
rect 62776 141200 62782 141212
rect 68054 141200 68060 141212
rect 62776 141172 68060 141200
rect 62776 141160 62782 141172
rect 68054 141160 68060 141172
rect 68112 141160 68118 141212
rect 100916 141200 100944 141308
rect 132638 141296 132644 141348
rect 132696 141296 132702 141348
rect 140826 141296 140832 141348
rect 140884 141336 140890 141348
rect 144322 141336 144328 141348
rect 140884 141308 144328 141336
rect 140884 141296 140890 141308
rect 144322 141296 144328 141308
rect 144380 141296 144386 141348
rect 163093 141339 163151 141345
rect 163093 141305 163105 141339
rect 163139 141336 163151 141339
rect 164378 141336 164384 141348
rect 163139 141308 164384 141336
rect 163139 141305 163151 141308
rect 163093 141299 163151 141305
rect 164378 141296 164384 141308
rect 164436 141296 164442 141348
rect 171002 141296 171008 141348
rect 171060 141336 171066 141348
rect 171060 141308 172796 141336
rect 171060 141296 171066 141308
rect 102370 141200 102376 141212
rect 100916 141172 102376 141200
rect 102370 141160 102376 141172
rect 102428 141160 102434 141212
rect 172768 141200 172796 141308
rect 172860 141268 172888 141376
rect 174222 141268 174228 141280
rect 172860 141240 174228 141268
rect 174222 141228 174228 141240
rect 174280 141228 174286 141280
rect 174774 141200 174780 141212
rect 172768 141172 174780 141200
rect 174774 141160 174780 141172
rect 174832 141160 174838 141212
rect 135398 141092 135404 141144
rect 135456 141132 135462 141144
rect 141102 141132 141108 141144
rect 135456 141104 141108 141132
rect 135456 141092 135462 141104
rect 141102 141092 141108 141104
rect 141160 141092 141166 141144
rect 135398 140684 135404 140736
rect 135456 140724 135462 140736
rect 141010 140724 141016 140736
rect 135456 140696 141016 140724
rect 135456 140684 135462 140696
rect 141010 140684 141016 140696
rect 141068 140684 141074 140736
rect 62810 139868 62816 139920
rect 62868 139908 62874 139920
rect 66490 139908 66496 139920
rect 62868 139880 66496 139908
rect 62868 139868 62874 139880
rect 66490 139868 66496 139880
rect 66548 139868 66554 139920
rect 95470 139868 95476 139920
rect 95528 139908 95534 139920
rect 102370 139908 102376 139920
rect 95528 139880 102376 139908
rect 95528 139868 95534 139880
rect 102370 139868 102376 139880
rect 102428 139868 102434 139920
rect 172842 139868 172848 139920
rect 172900 139908 172906 139920
rect 174958 139908 174964 139920
rect 172900 139880 174964 139908
rect 172900 139868 172906 139880
rect 174958 139868 174964 139880
rect 175016 139868 175022 139920
rect 95562 139800 95568 139852
rect 95620 139840 95626 139852
rect 102462 139840 102468 139852
rect 95620 139812 102468 139840
rect 95620 139800 95626 139812
rect 102462 139800 102468 139812
rect 102520 139800 102526 139852
rect 135398 139800 135404 139852
rect 135456 139840 135462 139852
rect 139538 139840 139544 139852
rect 135456 139812 139544 139840
rect 135456 139800 135462 139812
rect 139538 139800 139544 139812
rect 139596 139800 139602 139852
rect 62718 139732 62724 139784
rect 62776 139772 62782 139784
rect 65110 139772 65116 139784
rect 62776 139744 65116 139772
rect 62776 139732 62782 139744
rect 65110 139732 65116 139744
rect 65168 139732 65174 139784
rect 94090 139732 94096 139784
rect 94148 139772 94154 139784
rect 102554 139772 102560 139784
rect 94148 139744 102560 139772
rect 94148 139732 94154 139744
rect 102554 139732 102560 139744
rect 102612 139732 102618 139784
rect 62810 139596 62816 139648
rect 62868 139636 62874 139648
rect 66582 139636 66588 139648
rect 62868 139608 66588 139636
rect 62868 139596 62874 139608
rect 66582 139596 66588 139608
rect 66640 139596 66646 139648
rect 135398 139460 135404 139512
rect 135456 139500 135462 139512
rect 138250 139500 138256 139512
rect 135456 139472 138256 139500
rect 135456 139460 135462 139472
rect 138250 139460 138256 139472
rect 138308 139460 138314 139512
rect 172474 138712 172480 138764
rect 172532 138752 172538 138764
rect 174222 138752 174228 138764
rect 172532 138724 174228 138752
rect 172532 138712 172538 138724
rect 174222 138712 174228 138724
rect 174280 138712 174286 138764
rect 62902 138644 62908 138696
rect 62960 138684 62966 138696
rect 66398 138684 66404 138696
rect 62960 138656 66404 138684
rect 62960 138644 62966 138656
rect 66398 138644 66404 138656
rect 66456 138644 66462 138696
rect 135122 138644 135128 138696
rect 135180 138684 135186 138696
rect 136962 138684 136968 138696
rect 135180 138656 136968 138684
rect 135180 138644 135186 138656
rect 136962 138644 136968 138656
rect 137020 138644 137026 138696
rect 172658 138644 172664 138696
rect 172716 138684 172722 138696
rect 174314 138684 174320 138696
rect 172716 138656 174320 138684
rect 172716 138644 172722 138656
rect 174314 138644 174320 138656
rect 174372 138644 174378 138696
rect 62810 138576 62816 138628
rect 62868 138616 62874 138628
rect 66214 138616 66220 138628
rect 62868 138588 66220 138616
rect 62868 138576 62874 138588
rect 66214 138576 66220 138588
rect 66272 138576 66278 138628
rect 91241 138619 91299 138625
rect 91241 138585 91253 138619
rect 91287 138616 91299 138619
rect 97037 138619 97095 138625
rect 97037 138616 97049 138619
rect 91287 138588 91468 138616
rect 91287 138585 91299 138588
rect 91241 138579 91299 138585
rect 91333 138551 91391 138557
rect 91333 138517 91345 138551
rect 91379 138517 91391 138551
rect 91440 138548 91468 138588
rect 92636 138588 97049 138616
rect 92636 138548 92664 138588
rect 97037 138585 97049 138588
rect 97083 138585 97095 138619
rect 97037 138579 97095 138585
rect 135398 138576 135404 138628
rect 135456 138616 135462 138628
rect 136870 138616 136876 138628
rect 135456 138588 136876 138616
rect 135456 138576 135462 138588
rect 136870 138576 136876 138588
rect 136928 138576 136934 138628
rect 163093 138619 163151 138625
rect 163093 138585 163105 138619
rect 163139 138585 163151 138619
rect 163093 138579 163151 138585
rect 91440 138520 92664 138548
rect 92713 138551 92771 138557
rect 91333 138511 91391 138517
rect 92713 138517 92725 138551
rect 92759 138548 92771 138551
rect 93725 138551 93783 138557
rect 93725 138548 93737 138551
rect 92759 138520 93737 138548
rect 92759 138517 92771 138520
rect 92713 138511 92771 138517
rect 93725 138517 93737 138520
rect 93771 138517 93783 138551
rect 93725 138511 93783 138517
rect 94001 138551 94059 138557
rect 94001 138517 94013 138551
rect 94047 138548 94059 138551
rect 102370 138548 102376 138560
rect 94047 138520 102376 138548
rect 94047 138517 94059 138520
rect 94001 138511 94059 138517
rect 91348 138480 91376 138511
rect 102370 138508 102376 138520
rect 102428 138508 102434 138560
rect 102462 138480 102468 138492
rect 91348 138452 102468 138480
rect 102462 138440 102468 138452
rect 102520 138440 102526 138492
rect 163108 138480 163136 138579
rect 174130 138480 174136 138492
rect 163108 138452 174136 138480
rect 174130 138440 174136 138452
rect 174188 138440 174194 138492
rect 97037 138415 97095 138421
rect 97037 138381 97049 138415
rect 97083 138412 97095 138415
rect 100990 138412 100996 138424
rect 97083 138384 100996 138412
rect 97083 138381 97095 138384
rect 97037 138375 97095 138381
rect 100990 138372 100996 138384
rect 101048 138372 101054 138424
rect 62718 137216 62724 137268
rect 62776 137256 62782 137268
rect 66214 137256 66220 137268
rect 62776 137228 66220 137256
rect 62776 137216 62782 137228
rect 66214 137216 66220 137228
rect 66272 137216 66278 137268
rect 135214 137216 135220 137268
rect 135272 137256 135278 137268
rect 136962 137256 136968 137268
rect 135272 137228 136968 137256
rect 135272 137216 135278 137228
rect 136962 137216 136968 137228
rect 137020 137216 137026 137268
rect 172658 137216 172664 137268
rect 172716 137256 172722 137268
rect 174038 137256 174044 137268
rect 172716 137228 174044 137256
rect 172716 137216 172722 137228
rect 174038 137216 174044 137228
rect 174096 137216 174102 137268
rect 62626 137148 62632 137200
rect 62684 137188 62690 137200
rect 66398 137188 66404 137200
rect 62684 137160 66404 137188
rect 62684 137148 62690 137160
rect 66398 137148 66404 137160
rect 66456 137148 66462 137200
rect 135306 137148 135312 137200
rect 135364 137188 135370 137200
rect 136870 137188 136876 137200
rect 135364 137160 136876 137188
rect 135364 137148 135370 137160
rect 136870 137148 136876 137160
rect 136928 137148 136934 137200
rect 172198 137148 172204 137200
rect 172256 137188 172262 137200
rect 173946 137188 173952 137200
rect 172256 137160 173952 137188
rect 172256 137148 172262 137160
rect 173946 137148 173952 137160
rect 174004 137148 174010 137200
rect 100622 137012 100628 137064
rect 100680 137052 100686 137064
rect 102830 137052 102836 137064
rect 100680 137024 102836 137052
rect 100680 137012 100686 137024
rect 102830 137012 102836 137024
rect 102888 137012 102894 137064
rect 100530 136672 100536 136724
rect 100588 136712 100594 136724
rect 102462 136712 102468 136724
rect 100588 136684 102468 136712
rect 100588 136672 100594 136684
rect 102462 136672 102468 136684
rect 102520 136672 102526 136724
rect 172566 136128 172572 136180
rect 172624 136168 172630 136180
rect 174130 136168 174136 136180
rect 172624 136140 174136 136168
rect 172624 136128 172630 136140
rect 174130 136128 174136 136140
rect 174188 136128 174194 136180
rect 100622 135992 100628 136044
rect 100680 136032 100686 136044
rect 102186 136032 102192 136044
rect 100680 136004 102192 136032
rect 100680 135992 100686 136004
rect 102186 135992 102192 136004
rect 102244 135992 102250 136044
rect 172658 135992 172664 136044
rect 172716 136032 172722 136044
rect 174498 136032 174504 136044
rect 172716 136004 174504 136032
rect 172716 135992 172722 136004
rect 174498 135992 174504 136004
rect 174556 135992 174562 136044
rect 62902 135856 62908 135908
rect 62960 135896 62966 135908
rect 66030 135896 66036 135908
rect 62960 135868 66036 135896
rect 62960 135856 62966 135868
rect 66030 135856 66036 135868
rect 66088 135856 66094 135908
rect 100898 135856 100904 135908
rect 100956 135896 100962 135908
rect 102094 135896 102100 135908
rect 100956 135868 102100 135896
rect 100956 135856 100962 135868
rect 102094 135856 102100 135868
rect 102152 135856 102158 135908
rect 134938 135856 134944 135908
rect 134996 135896 135002 135908
rect 136962 135896 136968 135908
rect 134996 135868 136968 135896
rect 134996 135856 135002 135868
rect 136962 135856 136968 135868
rect 137020 135856 137026 135908
rect 62994 135788 63000 135840
rect 63052 135828 63058 135840
rect 66398 135828 66404 135840
rect 63052 135800 66404 135828
rect 63052 135788 63058 135800
rect 66398 135788 66404 135800
rect 66456 135788 66462 135840
rect 135122 135788 135128 135840
rect 135180 135828 135186 135840
rect 136870 135828 136876 135840
rect 135180 135800 136876 135828
rect 135180 135788 135186 135800
rect 136870 135788 136876 135800
rect 136928 135788 136934 135840
rect 172014 135788 172020 135840
rect 172072 135828 172078 135840
rect 174314 135828 174320 135840
rect 172072 135800 174320 135828
rect 172072 135788 172078 135800
rect 174314 135788 174320 135800
rect 174372 135788 174378 135840
rect 100714 135720 100720 135772
rect 100772 135760 100778 135772
rect 102370 135760 102376 135772
rect 100772 135732 102376 135760
rect 100772 135720 100778 135732
rect 102370 135720 102376 135732
rect 102428 135720 102434 135772
rect 100990 135652 100996 135704
rect 101048 135692 101054 135704
rect 102462 135692 102468 135704
rect 101048 135664 102468 135692
rect 101048 135652 101054 135664
rect 102462 135652 102468 135664
rect 102520 135652 102526 135704
rect 100346 135584 100352 135636
rect 100404 135624 100410 135636
rect 102646 135624 102652 135636
rect 100404 135596 102652 135624
rect 100404 135584 100410 135596
rect 102646 135584 102652 135596
rect 102704 135584 102710 135636
rect 62718 134972 62724 135024
rect 62776 135012 62782 135024
rect 65018 135012 65024 135024
rect 62776 134984 65024 135012
rect 62776 134972 62782 134984
rect 65018 134972 65024 134984
rect 65076 134972 65082 135024
rect 135030 134904 135036 134956
rect 135088 134944 135094 134956
rect 136778 134944 136784 134956
rect 135088 134916 136784 134944
rect 135088 134904 135094 134916
rect 136778 134904 136784 134916
rect 136836 134904 136842 134956
rect 62810 134632 62816 134684
rect 62868 134672 62874 134684
rect 66306 134672 66312 134684
rect 62868 134644 66312 134672
rect 62868 134632 62874 134644
rect 66306 134632 66312 134644
rect 66364 134632 66370 134684
rect 100070 134632 100076 134684
rect 100128 134672 100134 134684
rect 102278 134672 102284 134684
rect 100128 134644 102284 134672
rect 100128 134632 100134 134644
rect 102278 134632 102284 134644
rect 102336 134632 102342 134684
rect 171830 134632 171836 134684
rect 171888 134672 171894 134684
rect 174222 134672 174228 134684
rect 171888 134644 174228 134672
rect 171888 134632 171894 134644
rect 174222 134632 174228 134644
rect 174280 134632 174286 134684
rect 135214 134496 135220 134548
rect 135272 134536 135278 134548
rect 136962 134536 136968 134548
rect 135272 134508 136968 134536
rect 135272 134496 135278 134508
rect 136962 134496 136968 134508
rect 137020 134496 137026 134548
rect 172658 134496 172664 134548
rect 172716 134536 172722 134548
rect 174314 134536 174320 134548
rect 172716 134508 174320 134536
rect 172716 134496 172722 134508
rect 174314 134496 174320 134508
rect 174372 134496 174378 134548
rect 62718 134428 62724 134480
rect 62776 134468 62782 134480
rect 66398 134468 66404 134480
rect 62776 134440 66404 134468
rect 62776 134428 62782 134440
rect 66398 134428 66404 134440
rect 66456 134428 66462 134480
rect 132641 134471 132699 134477
rect 132641 134437 132653 134471
rect 132687 134468 132699 134471
rect 132914 134468 132920 134480
rect 132687 134440 132920 134468
rect 132687 134437 132699 134440
rect 132641 134431 132699 134437
rect 132914 134428 132920 134440
rect 132972 134428 132978 134480
rect 135398 134428 135404 134480
rect 135456 134468 135462 134480
rect 136870 134468 136876 134480
rect 135456 134440 136876 134468
rect 135456 134428 135462 134440
rect 136870 134428 136876 134440
rect 136928 134428 136934 134480
rect 172198 133544 172204 133596
rect 172256 133584 172262 133596
rect 175326 133584 175332 133596
rect 172256 133556 175332 133584
rect 172256 133544 172262 133556
rect 175326 133544 175332 133556
rect 175384 133544 175390 133596
rect 100898 133136 100904 133188
rect 100956 133176 100962 133188
rect 102186 133176 102192 133188
rect 100956 133148 102192 133176
rect 100956 133136 100962 133148
rect 102186 133136 102192 133148
rect 102244 133136 102250 133188
rect 63546 133068 63552 133120
rect 63604 133108 63610 133120
rect 66398 133108 66404 133120
rect 63604 133080 66404 133108
rect 63604 133068 63610 133080
rect 66398 133068 66404 133080
rect 66456 133068 66462 133120
rect 135122 133068 135128 133120
rect 135180 133108 135186 133120
rect 136962 133108 136968 133120
rect 135180 133080 136968 133108
rect 135180 133068 135186 133080
rect 136962 133068 136968 133080
rect 137020 133068 137026 133120
rect 172658 133068 172664 133120
rect 172716 133108 172722 133120
rect 174866 133108 174872 133120
rect 172716 133080 174872 133108
rect 172716 133068 172722 133080
rect 174866 133068 174872 133080
rect 174924 133068 174930 133120
rect 63638 133000 63644 133052
rect 63696 133040 63702 133052
rect 65846 133040 65852 133052
rect 63696 133012 65852 133040
rect 63696 133000 63702 133012
rect 65846 133000 65852 133012
rect 65904 133000 65910 133052
rect 100070 133000 100076 133052
rect 100128 133040 100134 133052
rect 102094 133040 102100 133052
rect 100128 133012 102100 133040
rect 100128 133000 100134 133012
rect 102094 133000 102100 133012
rect 102152 133000 102158 133052
rect 135306 133000 135312 133052
rect 135364 133040 135370 133052
rect 136870 133040 136876 133052
rect 135364 133012 136876 133040
rect 135364 133000 135370 133012
rect 136870 133000 136876 133012
rect 136928 133000 136934 133052
rect 100990 132932 100996 132984
rect 101048 132972 101054 132984
rect 102370 132972 102376 132984
rect 101048 132944 102376 132972
rect 101048 132932 101054 132944
rect 102370 132932 102376 132944
rect 102428 132932 102434 132984
rect 172382 131912 172388 131964
rect 172440 131952 172446 131964
rect 175418 131952 175424 131964
rect 172440 131924 175424 131952
rect 172440 131912 172446 131924
rect 175418 131912 175424 131924
rect 175476 131912 175482 131964
rect 172658 131776 172664 131828
rect 172716 131816 172722 131828
rect 175142 131816 175148 131828
rect 172716 131788 175148 131816
rect 172716 131776 172722 131788
rect 175142 131776 175148 131788
rect 175200 131776 175206 131828
rect 63270 131708 63276 131760
rect 63328 131748 63334 131760
rect 65662 131748 65668 131760
rect 63328 131720 65668 131748
rect 63328 131708 63334 131720
rect 65662 131708 65668 131720
rect 65720 131708 65726 131760
rect 100898 131708 100904 131760
rect 100956 131748 100962 131760
rect 102002 131748 102008 131760
rect 100956 131720 102008 131748
rect 100956 131708 100962 131720
rect 102002 131708 102008 131720
rect 102060 131708 102066 131760
rect 134938 131708 134944 131760
rect 134996 131748 135002 131760
rect 136962 131748 136968 131760
rect 134996 131720 136968 131748
rect 134996 131708 135002 131720
rect 136962 131708 136968 131720
rect 137020 131708 137026 131760
rect 172014 131708 172020 131760
rect 172072 131748 172078 131760
rect 175234 131748 175240 131760
rect 172072 131720 175240 131748
rect 172072 131708 172078 131720
rect 175234 131708 175240 131720
rect 175292 131708 175298 131760
rect 63454 131640 63460 131692
rect 63512 131680 63518 131692
rect 66398 131680 66404 131692
rect 63512 131652 66404 131680
rect 63512 131640 63518 131652
rect 66398 131640 66404 131652
rect 66456 131640 66462 131692
rect 100438 131640 100444 131692
rect 100496 131680 100502 131692
rect 100496 131652 101036 131680
rect 100496 131640 100502 131652
rect 101008 131612 101036 131652
rect 135214 131640 135220 131692
rect 135272 131680 135278 131692
rect 136870 131680 136876 131692
rect 135272 131652 136876 131680
rect 135272 131640 135278 131652
rect 136870 131640 136876 131652
rect 136928 131640 136934 131692
rect 102370 131612 102376 131624
rect 101008 131584 102376 131612
rect 102370 131572 102376 131584
rect 102428 131572 102434 131624
rect 135306 131028 135312 131080
rect 135364 131068 135370 131080
rect 136778 131068 136784 131080
rect 135364 131040 136784 131068
rect 135364 131028 135370 131040
rect 136778 131028 136784 131040
rect 136836 131028 136842 131080
rect 62810 130756 62816 130808
rect 62868 130796 62874 130808
rect 65018 130796 65024 130808
rect 62868 130768 65024 130796
rect 62868 130756 62874 130768
rect 65018 130756 65024 130768
rect 65076 130756 65082 130808
rect 100438 130552 100444 130604
rect 100496 130592 100502 130604
rect 102278 130592 102284 130604
rect 100496 130564 102284 130592
rect 100496 130552 100502 130564
rect 102278 130552 102284 130564
rect 102336 130552 102342 130604
rect 172658 130552 172664 130604
rect 172716 130592 172722 130604
rect 174222 130592 174228 130604
rect 172716 130564 174228 130592
rect 172716 130552 172722 130564
rect 174222 130552 174228 130564
rect 174280 130552 174286 130604
rect 62626 130348 62632 130400
rect 62684 130388 62690 130400
rect 66398 130388 66404 130400
rect 62684 130360 66404 130388
rect 62684 130348 62690 130360
rect 66398 130348 66404 130360
rect 66456 130348 66462 130400
rect 100898 130348 100904 130400
rect 100956 130388 100962 130400
rect 102186 130388 102192 130400
rect 100956 130360 102192 130388
rect 100956 130348 100962 130360
rect 102186 130348 102192 130360
rect 102244 130348 102250 130400
rect 135030 130348 135036 130400
rect 135088 130388 135094 130400
rect 136962 130388 136968 130400
rect 135088 130360 136968 130388
rect 135088 130348 135094 130360
rect 136962 130348 136968 130360
rect 137020 130348 137026 130400
rect 62718 130280 62724 130332
rect 62776 130320 62782 130332
rect 66306 130320 66312 130332
rect 62776 130292 66312 130320
rect 62776 130280 62782 130292
rect 66306 130280 66312 130292
rect 66364 130280 66370 130332
rect 135398 130280 135404 130332
rect 135456 130320 135462 130332
rect 136870 130320 136876 130332
rect 135456 130292 136876 130320
rect 135456 130280 135462 130292
rect 136870 130280 136876 130292
rect 136928 130280 136934 130332
rect 172658 130280 172664 130332
rect 172716 130320 172722 130332
rect 174314 130320 174320 130332
rect 172716 130292 174320 130320
rect 172716 130280 172722 130292
rect 174314 130280 174320 130292
rect 174372 130280 174378 130332
rect 100990 130212 100996 130264
rect 101048 130252 101054 130264
rect 102370 130252 102376 130264
rect 101048 130224 102376 130252
rect 101048 130212 101054 130224
rect 102370 130212 102376 130224
rect 102428 130212 102434 130264
rect 171830 129328 171836 129380
rect 171888 129368 171894 129380
rect 174130 129368 174136 129380
rect 171888 129340 174136 129368
rect 171888 129328 171894 129340
rect 174130 129328 174136 129340
rect 174188 129328 174194 129380
rect 171830 129056 171836 129108
rect 171888 129096 171894 129108
rect 174498 129096 174504 129108
rect 171888 129068 174504 129096
rect 171888 129056 171894 129068
rect 174498 129056 174504 129068
rect 174556 129056 174562 129108
rect 62902 128988 62908 129040
rect 62960 129028 62966 129040
rect 66398 129028 66404 129040
rect 62960 129000 66404 129028
rect 62960 128988 62966 129000
rect 66398 128988 66404 129000
rect 66456 128988 66462 129040
rect 100898 128988 100904 129040
rect 100956 129028 100962 129040
rect 102002 129028 102008 129040
rect 100956 129000 102008 129028
rect 100956 128988 100962 129000
rect 102002 128988 102008 129000
rect 102060 128988 102066 129040
rect 135122 128988 135128 129040
rect 135180 129028 135186 129040
rect 136962 129028 136968 129040
rect 135180 129000 136968 129028
rect 135180 128988 135186 129000
rect 136962 128988 136968 129000
rect 137020 128988 137026 129040
rect 62810 128920 62816 128972
rect 62868 128960 62874 128972
rect 65478 128960 65484 128972
rect 62868 128932 65484 128960
rect 62868 128920 62874 128932
rect 65478 128920 65484 128932
rect 65536 128920 65542 128972
rect 100070 128920 100076 128972
rect 100128 128960 100134 128972
rect 101910 128960 101916 128972
rect 100128 128932 101916 128960
rect 100128 128920 100134 128932
rect 101910 128920 101916 128932
rect 101968 128920 101974 128972
rect 135306 128920 135312 128972
rect 135364 128960 135370 128972
rect 136870 128960 136876 128972
rect 135364 128932 136876 128960
rect 135364 128920 135370 128932
rect 136870 128920 136876 128932
rect 136928 128920 136934 128972
rect 100346 127832 100352 127884
rect 100404 127872 100410 127884
rect 102278 127872 102284 127884
rect 100404 127844 102284 127872
rect 100404 127832 100410 127844
rect 102278 127832 102284 127844
rect 102336 127832 102342 127884
rect 172566 127832 172572 127884
rect 172624 127872 172630 127884
rect 174222 127872 174228 127884
rect 172624 127844 174228 127872
rect 172624 127832 172630 127844
rect 174222 127832 174228 127844
rect 174280 127832 174286 127884
rect 100530 127560 100536 127612
rect 100588 127600 100594 127612
rect 102002 127600 102008 127612
rect 100588 127572 102008 127600
rect 100588 127560 100594 127572
rect 102002 127560 102008 127572
rect 102060 127560 102066 127612
rect 135214 127560 135220 127612
rect 135272 127600 135278 127612
rect 136870 127600 136876 127612
rect 135272 127572 136876 127600
rect 135272 127560 135278 127572
rect 136870 127560 136876 127572
rect 136928 127560 136934 127612
rect 171554 127560 171560 127612
rect 171612 127600 171618 127612
rect 174590 127600 174596 127612
rect 171612 127572 174596 127600
rect 171612 127560 171618 127572
rect 174590 127560 174596 127572
rect 174648 127560 174654 127612
rect 62626 127492 62632 127544
rect 62684 127532 62690 127544
rect 66398 127532 66404 127544
rect 62684 127504 66404 127532
rect 62684 127492 62690 127504
rect 66398 127492 66404 127504
rect 66456 127492 66462 127544
rect 222709 127535 222767 127541
rect 222709 127501 222721 127535
rect 222755 127532 222767 127535
rect 222798 127532 222804 127544
rect 222755 127504 222804 127532
rect 222755 127501 222767 127504
rect 222709 127495 222767 127501
rect 222798 127492 222804 127504
rect 222856 127492 222862 127544
rect 134662 127152 134668 127204
rect 134720 127192 134726 127204
rect 136778 127192 136784 127204
rect 134720 127164 136784 127192
rect 134720 127152 134726 127164
rect 136778 127152 136784 127164
rect 136836 127152 136842 127204
rect 62810 126880 62816 126932
rect 62868 126920 62874 126932
rect 65018 126920 65024 126932
rect 62868 126892 65024 126920
rect 62868 126880 62874 126892
rect 65018 126880 65024 126892
rect 65076 126880 65082 126932
rect 172198 126472 172204 126524
rect 172256 126512 172262 126524
rect 174314 126512 174320 126524
rect 172256 126484 174320 126512
rect 172256 126472 172262 126484
rect 174314 126472 174320 126484
rect 174372 126472 174378 126524
rect 100806 126268 100812 126320
rect 100864 126308 100870 126320
rect 102094 126308 102100 126320
rect 100864 126280 102100 126308
rect 100864 126268 100870 126280
rect 102094 126268 102100 126280
rect 102152 126268 102158 126320
rect 62718 126200 62724 126252
rect 62776 126240 62782 126252
rect 66306 126240 66312 126252
rect 62776 126212 66312 126240
rect 62776 126200 62782 126212
rect 66306 126200 66312 126212
rect 66364 126200 66370 126252
rect 100898 126200 100904 126252
rect 100956 126240 100962 126252
rect 102278 126240 102284 126252
rect 100956 126212 102284 126240
rect 100956 126200 100962 126212
rect 102278 126200 102284 126212
rect 102336 126200 102342 126252
rect 135030 126200 135036 126252
rect 135088 126240 135094 126252
rect 136962 126240 136968 126252
rect 135088 126212 136968 126240
rect 135088 126200 135094 126212
rect 136962 126200 136968 126212
rect 137020 126200 137026 126252
rect 172658 126200 172664 126252
rect 172716 126240 172722 126252
rect 174498 126240 174504 126252
rect 172716 126212 174504 126240
rect 172716 126200 172722 126212
rect 174498 126200 174504 126212
rect 174556 126200 174562 126252
rect 62902 126132 62908 126184
rect 62960 126172 62966 126184
rect 66398 126172 66404 126184
rect 62960 126144 66404 126172
rect 62960 126132 62966 126144
rect 66398 126132 66404 126144
rect 66456 126132 66462 126184
rect 100438 126132 100444 126184
rect 100496 126172 100502 126184
rect 100496 126144 101036 126172
rect 100496 126132 100502 126144
rect 101008 126104 101036 126144
rect 135306 126132 135312 126184
rect 135364 126172 135370 126184
rect 136870 126172 136876 126184
rect 135364 126144 136876 126172
rect 135364 126132 135370 126144
rect 136870 126132 136876 126144
rect 136928 126132 136934 126184
rect 172014 126132 172020 126184
rect 172072 126172 172078 126184
rect 174130 126172 174136 126184
rect 172072 126144 174136 126172
rect 172072 126132 172078 126144
rect 174130 126132 174136 126144
rect 174188 126132 174194 126184
rect 102370 126104 102376 126116
rect 101008 126076 102376 126104
rect 102370 126064 102376 126076
rect 102428 126064 102434 126116
rect 135398 125656 135404 125708
rect 135456 125696 135462 125708
rect 136778 125696 136784 125708
rect 135456 125668 136784 125696
rect 135456 125656 135462 125668
rect 136778 125656 136784 125668
rect 136836 125656 136842 125708
rect 62810 125520 62816 125572
rect 62868 125560 62874 125572
rect 65018 125560 65024 125572
rect 62868 125532 65024 125560
rect 62868 125520 62874 125532
rect 65018 125520 65024 125532
rect 65076 125520 65082 125572
rect 171830 125248 171836 125300
rect 171888 125288 171894 125300
rect 174222 125288 174228 125300
rect 171888 125260 174228 125288
rect 171888 125248 171894 125260
rect 174222 125248 174228 125260
rect 174280 125248 174286 125300
rect 100806 124840 100812 124892
rect 100864 124880 100870 124892
rect 102186 124880 102192 124892
rect 100864 124852 102192 124880
rect 100864 124840 100870 124852
rect 102186 124840 102192 124852
rect 102244 124840 102250 124892
rect 172198 124840 172204 124892
rect 172256 124880 172262 124892
rect 174590 124880 174596 124892
rect 172256 124852 174596 124880
rect 172256 124840 172262 124852
rect 174590 124840 174596 124852
rect 174648 124840 174654 124892
rect 62626 124772 62632 124824
rect 62684 124812 62690 124824
rect 66398 124812 66404 124824
rect 62684 124784 66404 124812
rect 62684 124772 62690 124784
rect 66398 124772 66404 124784
rect 66456 124772 66462 124824
rect 100898 124772 100904 124824
rect 100956 124812 100962 124824
rect 100956 124784 101036 124812
rect 100956 124772 100962 124784
rect 101008 124744 101036 124784
rect 135122 124772 135128 124824
rect 135180 124812 135186 124824
rect 136870 124812 136876 124824
rect 135180 124784 136876 124812
rect 135180 124772 135186 124784
rect 136870 124772 136876 124784
rect 136928 124772 136934 124824
rect 222706 124812 222712 124824
rect 222667 124784 222712 124812
rect 222706 124772 222712 124784
rect 222764 124772 222770 124824
rect 102370 124744 102376 124756
rect 101008 124716 102376 124744
rect 102370 124704 102376 124716
rect 102428 124704 102434 124756
rect 135214 124228 135220 124280
rect 135272 124268 135278 124280
rect 136778 124268 136784 124280
rect 135272 124240 136784 124268
rect 135272 124228 135278 124240
rect 136778 124228 136784 124240
rect 136836 124228 136842 124280
rect 62810 123752 62816 123804
rect 62868 123792 62874 123804
rect 65018 123792 65024 123804
rect 62868 123764 65024 123792
rect 62868 123752 62874 123764
rect 65018 123752 65024 123764
rect 65076 123752 65082 123804
rect 172566 123480 172572 123532
rect 172624 123520 172630 123532
rect 175326 123520 175332 123532
rect 172624 123492 175332 123520
rect 172624 123480 172630 123492
rect 175326 123480 175332 123492
rect 175384 123480 175390 123532
rect 63546 123344 63552 123396
rect 63604 123384 63610 123396
rect 66398 123384 66404 123396
rect 63604 123356 66404 123384
rect 63604 123344 63610 123356
rect 66398 123344 66404 123356
rect 66456 123344 66462 123396
rect 100254 123344 100260 123396
rect 100312 123384 100318 123396
rect 102278 123384 102284 123396
rect 100312 123356 102284 123384
rect 100312 123344 100318 123356
rect 102278 123344 102284 123356
rect 102336 123344 102342 123396
rect 135398 123344 135404 123396
rect 135456 123384 135462 123396
rect 136870 123384 136876 123396
rect 135456 123356 136876 123384
rect 135456 123344 135462 123356
rect 136870 123344 136876 123356
rect 136928 123344 136934 123396
rect 171830 123344 171836 123396
rect 171888 123384 171894 123396
rect 174130 123384 174136 123396
rect 171888 123356 174136 123384
rect 171888 123344 171894 123356
rect 174130 123344 174136 123356
rect 174188 123344 174194 123396
rect 135306 122868 135312 122920
rect 135364 122908 135370 122920
rect 136778 122908 136784 122920
rect 135364 122880 136784 122908
rect 135364 122868 135370 122880
rect 136778 122868 136784 122880
rect 136836 122868 136842 122920
rect 62810 122664 62816 122716
rect 62868 122704 62874 122716
rect 65018 122704 65024 122716
rect 62868 122676 65024 122704
rect 62868 122664 62874 122676
rect 65018 122664 65024 122676
rect 65076 122664 65082 122716
rect 171830 122392 171836 122444
rect 171888 122432 171894 122444
rect 175050 122432 175056 122444
rect 171888 122404 175056 122432
rect 171888 122392 171894 122404
rect 175050 122392 175056 122404
rect 175108 122392 175114 122444
rect 100162 122188 100168 122240
rect 100220 122228 100226 122240
rect 102278 122228 102284 122240
rect 100220 122200 102284 122228
rect 100220 122188 100226 122200
rect 102278 122188 102284 122200
rect 102336 122188 102342 122240
rect 100898 122120 100904 122172
rect 100956 122160 100962 122172
rect 102002 122160 102008 122172
rect 100956 122132 102008 122160
rect 100956 122120 100962 122132
rect 102002 122120 102008 122132
rect 102060 122120 102066 122172
rect 135122 122120 135128 122172
rect 135180 122160 135186 122172
rect 137054 122160 137060 122172
rect 135180 122132 137060 122160
rect 135180 122120 135186 122132
rect 137054 122120 137060 122132
rect 137112 122120 137118 122172
rect 172014 122120 172020 122172
rect 172072 122160 172078 122172
rect 175418 122160 175424 122172
rect 172072 122132 175424 122160
rect 172072 122120 172078 122132
rect 175418 122120 175424 122132
rect 175476 122120 175482 122172
rect 63454 122052 63460 122104
rect 63512 122092 63518 122104
rect 66306 122092 66312 122104
rect 63512 122064 66312 122092
rect 63512 122052 63518 122064
rect 66306 122052 66312 122064
rect 66364 122052 66370 122104
rect 135214 122052 135220 122104
rect 135272 122092 135278 122104
rect 136962 122092 136968 122104
rect 135272 122064 136968 122092
rect 135272 122052 135278 122064
rect 136962 122052 136968 122064
rect 137020 122052 137026 122104
rect 63638 121984 63644 122036
rect 63696 122024 63702 122036
rect 66398 122024 66404 122036
rect 63696 121996 66404 122024
rect 63696 121984 63702 121996
rect 66398 121984 66404 121996
rect 66456 121984 66462 122036
rect 100622 121984 100628 122036
rect 100680 122024 100686 122036
rect 102094 122024 102100 122036
rect 100680 121996 102100 122024
rect 100680 121984 100686 121996
rect 102094 121984 102100 121996
rect 102152 121984 102158 122036
rect 136870 122024 136876 122036
rect 135508 121996 136876 122024
rect 100990 121916 100996 121968
rect 101048 121956 101054 121968
rect 102370 121956 102376 121968
rect 101048 121928 102376 121956
rect 101048 121916 101054 121928
rect 102370 121916 102376 121928
rect 102428 121916 102434 121968
rect 135306 121916 135312 121968
rect 135364 121956 135370 121968
rect 135508 121956 135536 121996
rect 136870 121984 136876 121996
rect 136928 121984 136934 122036
rect 172658 121984 172664 122036
rect 172716 122024 172722 122036
rect 175142 122024 175148 122036
rect 172716 121996 175148 122024
rect 172716 121984 172722 121996
rect 175142 121984 175148 121996
rect 175200 121984 175206 122036
rect 135364 121928 135536 121956
rect 135364 121916 135370 121928
rect 62810 121440 62816 121492
rect 62868 121480 62874 121492
rect 65018 121480 65024 121492
rect 62868 121452 65024 121480
rect 62868 121440 62874 121452
rect 65018 121440 65024 121452
rect 65076 121440 65082 121492
rect 100898 120896 100904 120948
rect 100956 120936 100962 120948
rect 102186 120936 102192 120948
rect 100956 120908 102192 120936
rect 100956 120896 100962 120908
rect 102186 120896 102192 120908
rect 102244 120896 102250 120948
rect 172106 120896 172112 120948
rect 172164 120936 172170 120948
rect 174314 120936 174320 120948
rect 172164 120908 174320 120936
rect 172164 120896 172170 120908
rect 174314 120896 174320 120908
rect 174372 120896 174378 120948
rect 172658 120760 172664 120812
rect 172716 120800 172722 120812
rect 174222 120800 174228 120812
rect 172716 120772 174228 120800
rect 172716 120760 172722 120772
rect 174222 120760 174228 120772
rect 174280 120760 174286 120812
rect 100070 120624 100076 120676
rect 100128 120664 100134 120676
rect 100128 120636 101036 120664
rect 100128 120624 100134 120636
rect 101008 120596 101036 120636
rect 102370 120596 102376 120608
rect 101008 120568 102376 120596
rect 102370 120556 102376 120568
rect 102428 120556 102434 120608
rect 134846 120216 134852 120268
rect 134904 120256 134910 120268
rect 136778 120256 136784 120268
rect 134904 120228 136784 120256
rect 134904 120216 134910 120228
rect 136778 120216 136784 120228
rect 136836 120216 136842 120268
rect 62810 119944 62816 119996
rect 62868 119984 62874 119996
rect 65018 119984 65024 119996
rect 62868 119956 65024 119984
rect 62868 119944 62874 119956
rect 65018 119944 65024 119956
rect 65076 119944 65082 119996
rect 171830 119672 171836 119724
rect 171888 119712 171894 119724
rect 174130 119712 174136 119724
rect 171888 119684 174136 119712
rect 171888 119672 171894 119684
rect 174130 119672 174136 119684
rect 174188 119672 174194 119724
rect 171830 119400 171836 119452
rect 171888 119440 171894 119452
rect 174498 119440 174504 119452
rect 171888 119412 174504 119440
rect 171888 119400 171894 119412
rect 174498 119400 174504 119412
rect 174556 119400 174562 119452
rect 62902 119264 62908 119316
rect 62960 119304 62966 119316
rect 65478 119304 65484 119316
rect 62960 119276 65484 119304
rect 62960 119264 62966 119276
rect 65478 119264 65484 119276
rect 65536 119264 65542 119316
rect 100438 119264 100444 119316
rect 100496 119304 100502 119316
rect 102278 119304 102284 119316
rect 100496 119276 102284 119304
rect 100496 119264 100502 119276
rect 102278 119264 102284 119276
rect 102336 119264 102342 119316
rect 135214 119264 135220 119316
rect 135272 119304 135278 119316
rect 136870 119304 136876 119316
rect 135272 119276 136876 119304
rect 135272 119264 135278 119276
rect 136870 119264 136876 119276
rect 136928 119264 136934 119316
rect 62718 119128 62724 119180
rect 62776 119168 62782 119180
rect 66214 119168 66220 119180
rect 62776 119140 66220 119168
rect 62776 119128 62782 119140
rect 66214 119128 66220 119140
rect 66272 119128 66278 119180
rect 135306 119128 135312 119180
rect 135364 119168 135370 119180
rect 136962 119168 136968 119180
rect 135364 119140 136968 119168
rect 135364 119128 135370 119140
rect 136962 119128 136968 119140
rect 137020 119128 137026 119180
rect 62810 118720 62816 118772
rect 62868 118760 62874 118772
rect 65018 118760 65024 118772
rect 62868 118732 65024 118760
rect 62868 118720 62874 118732
rect 65018 118720 65024 118732
rect 65076 118720 65082 118772
rect 135306 118516 135312 118568
rect 135364 118556 135370 118568
rect 136778 118556 136784 118568
rect 135364 118528 136784 118556
rect 135364 118516 135370 118528
rect 136778 118516 136784 118528
rect 136836 118516 136842 118568
rect 171646 118176 171652 118228
rect 171704 118216 171710 118228
rect 173946 118216 173952 118228
rect 171704 118188 173952 118216
rect 171704 118176 171710 118188
rect 173946 118176 173952 118188
rect 174004 118176 174010 118228
rect 100622 118108 100628 118160
rect 100680 118148 100686 118160
rect 102278 118148 102284 118160
rect 100680 118120 102284 118148
rect 100680 118108 100686 118120
rect 102278 118108 102284 118120
rect 102336 118108 102342 118160
rect 172658 118040 172664 118092
rect 172716 118080 172722 118092
rect 174314 118080 174320 118092
rect 172716 118052 174320 118080
rect 172716 118040 172722 118052
rect 174314 118040 174320 118052
rect 174372 118040 174378 118092
rect 135122 117904 135128 117956
rect 135180 117944 135186 117956
rect 136870 117944 136876 117956
rect 135180 117916 136876 117944
rect 135180 117904 135186 117916
rect 136870 117904 136876 117916
rect 136928 117904 136934 117956
rect 62718 117836 62724 117888
rect 62776 117876 62782 117888
rect 66398 117876 66404 117888
rect 62776 117848 66404 117876
rect 62776 117836 62782 117848
rect 66398 117836 66404 117848
rect 66456 117836 66462 117888
rect 100254 117836 100260 117888
rect 100312 117876 100318 117888
rect 100312 117848 101036 117876
rect 100312 117836 100318 117848
rect 101008 117808 101036 117848
rect 132914 117836 132920 117888
rect 132972 117836 132978 117888
rect 136962 117876 136968 117888
rect 135508 117848 136968 117876
rect 102462 117808 102468 117820
rect 101008 117780 102468 117808
rect 102462 117768 102468 117780
rect 102520 117768 102526 117820
rect 132638 117808 132644 117820
rect 132599 117780 132644 117808
rect 132638 117768 132644 117780
rect 132696 117768 132702 117820
rect 100990 117700 100996 117752
rect 101048 117740 101054 117752
rect 102370 117740 102376 117752
rect 101048 117712 102376 117740
rect 101048 117700 101054 117712
rect 102370 117700 102376 117712
rect 102428 117700 102434 117752
rect 132638 117632 132644 117684
rect 132696 117672 132702 117684
rect 132932 117672 132960 117836
rect 134110 117768 134116 117820
rect 134168 117808 134174 117820
rect 135508 117808 135536 117848
rect 136962 117836 136968 117848
rect 137020 117836 137026 117888
rect 171830 117836 171836 117888
rect 171888 117876 171894 117888
rect 174038 117876 174044 117888
rect 171888 117848 174044 117876
rect 171888 117836 171894 117848
rect 174038 117836 174044 117848
rect 174096 117836 174102 117888
rect 134168 117780 135536 117808
rect 134168 117768 134174 117780
rect 132696 117644 132960 117672
rect 132696 117632 132702 117644
rect 62810 117292 62816 117344
rect 62868 117332 62874 117344
rect 65018 117332 65024 117344
rect 62868 117304 65024 117332
rect 62868 117292 62874 117304
rect 65018 117292 65024 117304
rect 65076 117292 65082 117344
rect 62810 117156 62816 117208
rect 62868 117196 62874 117208
rect 64926 117196 64932 117208
rect 62868 117168 64932 117196
rect 62868 117156 62874 117168
rect 64926 117156 64932 117168
rect 64984 117156 64990 117208
rect 134662 117156 134668 117208
rect 134720 117196 134726 117208
rect 136778 117196 136784 117208
rect 134720 117168 136784 117196
rect 134720 117156 134726 117168
rect 136778 117156 136784 117168
rect 136836 117156 136842 117208
rect 100254 116680 100260 116732
rect 100312 116720 100318 116732
rect 102186 116720 102192 116732
rect 100312 116692 102192 116720
rect 100312 116680 100318 116692
rect 102186 116680 102192 116692
rect 102244 116680 102250 116732
rect 172658 116544 172664 116596
rect 172716 116584 172722 116596
rect 174130 116584 174136 116596
rect 172716 116556 174136 116584
rect 172716 116544 172722 116556
rect 174130 116544 174136 116556
rect 174188 116544 174194 116596
rect 100898 116476 100904 116528
rect 100956 116516 100962 116528
rect 100956 116488 101036 116516
rect 100956 116476 100962 116488
rect 101008 116448 101036 116488
rect 135306 116476 135312 116528
rect 135364 116516 135370 116528
rect 136870 116516 136876 116528
rect 135364 116488 136876 116516
rect 135364 116476 135370 116488
rect 136870 116476 136876 116488
rect 136928 116476 136934 116528
rect 172566 116476 172572 116528
rect 172624 116516 172630 116528
rect 174222 116516 174228 116528
rect 172624 116488 174228 116516
rect 172624 116476 172630 116488
rect 174222 116476 174228 116488
rect 174280 116476 174286 116528
rect 102370 116448 102376 116460
rect 101008 116420 102376 116448
rect 102370 116408 102376 116420
rect 102428 116408 102434 116460
rect 100530 116340 100536 116392
rect 100588 116380 100594 116392
rect 102646 116380 102652 116392
rect 100588 116352 102652 116380
rect 100588 116340 100594 116352
rect 102646 116340 102652 116352
rect 102704 116340 102710 116392
rect 62810 115728 62816 115780
rect 62868 115768 62874 115780
rect 65018 115768 65024 115780
rect 62868 115740 65024 115768
rect 62868 115728 62874 115740
rect 65018 115728 65024 115740
rect 65076 115728 65082 115780
rect 134846 115592 134852 115644
rect 134904 115632 134910 115644
rect 136778 115632 136784 115644
rect 134904 115604 136784 115632
rect 134904 115592 134910 115604
rect 136778 115592 136784 115604
rect 136836 115592 136842 115644
rect 171830 115592 171836 115644
rect 171888 115632 171894 115644
rect 174038 115632 174044 115644
rect 171888 115604 174044 115632
rect 171888 115592 171894 115604
rect 174038 115592 174044 115604
rect 174096 115592 174102 115644
rect 100898 115456 100904 115508
rect 100956 115496 100962 115508
rect 102278 115496 102284 115508
rect 100956 115468 102284 115496
rect 100956 115456 100962 115468
rect 102278 115456 102284 115468
rect 102336 115456 102342 115508
rect 222614 115048 222620 115100
rect 222672 115088 222678 115100
rect 222982 115088 222988 115100
rect 222672 115060 222988 115088
rect 222672 115048 222678 115060
rect 222982 115048 222988 115060
rect 223040 115048 223046 115100
rect 62810 114844 62816 114896
rect 62868 114884 62874 114896
rect 66398 114884 66404 114896
rect 62868 114856 66404 114884
rect 62868 114844 62874 114856
rect 66398 114844 66404 114856
rect 66456 114844 66462 114896
rect 62810 114572 62816 114624
rect 62868 114612 62874 114624
rect 65018 114612 65024 114624
rect 62868 114584 65024 114612
rect 62868 114572 62874 114584
rect 65018 114572 65024 114584
rect 65076 114572 65082 114624
rect 134846 114436 134852 114488
rect 134904 114476 134910 114488
rect 136778 114476 136784 114488
rect 134904 114448 136784 114476
rect 134904 114436 134910 114448
rect 136778 114436 136784 114448
rect 136836 114436 136842 114488
rect 30426 114300 30432 114352
rect 30484 114340 30490 114352
rect 92710 114340 92716 114352
rect 30484 114312 92716 114340
rect 30484 114300 30490 114312
rect 92710 114300 92716 114312
rect 92768 114300 92774 114352
rect 113502 113620 113508 113672
rect 113560 113660 113566 113672
rect 114376 113660 114382 113672
rect 113560 113632 114382 113660
rect 113560 113620 113566 113632
rect 114376 113620 114382 113632
rect 114434 113620 114440 113672
rect 132086 113620 132092 113672
rect 132144 113660 132150 113672
rect 132641 113663 132699 113669
rect 132641 113660 132653 113663
rect 132144 113632 132653 113660
rect 132144 113620 132150 113632
rect 132641 113629 132653 113632
rect 132687 113660 132699 113663
rect 144874 113660 144880 113672
rect 132687 113632 144880 113660
rect 132687 113629 132699 113632
rect 132641 113623 132699 113629
rect 144874 113620 144880 113632
rect 144932 113660 144938 113672
rect 204674 113660 204680 113672
rect 144932 113632 204680 113660
rect 144932 113620 144938 113632
rect 204674 113620 204680 113632
rect 204732 113620 204738 113672
rect 154810 113552 154816 113604
rect 154868 113592 154874 113604
rect 207250 113592 207256 113604
rect 154868 113564 207256 113592
rect 154868 113552 154874 113564
rect 207250 113552 207256 113564
rect 207308 113552 207314 113604
rect 194646 113144 194652 113196
rect 194704 113184 194710 113196
rect 198234 113184 198240 113196
rect 194704 113156 198240 113184
rect 194704 113144 194710 113156
rect 198234 113144 198240 113156
rect 198292 113144 198298 113196
rect 189402 113076 189408 113128
rect 189460 113116 189466 113128
rect 190230 113116 190236 113128
rect 189460 113088 190236 113116
rect 189460 113076 189466 113088
rect 190230 113076 190236 113088
rect 190288 113076 190294 113128
rect 191334 113076 191340 113128
rect 191392 113116 191398 113128
rect 193082 113116 193088 113128
rect 191392 113088 193088 113116
rect 191392 113076 191398 113088
rect 193082 113076 193088 113088
rect 193140 113076 193146 113128
rect 193726 113076 193732 113128
rect 193784 113116 193790 113128
rect 196118 113116 196124 113128
rect 193784 113088 196124 113116
rect 193784 113076 193790 113088
rect 196118 113076 196124 113088
rect 196176 113076 196182 113128
rect 198510 113076 198516 113128
rect 198568 113116 198574 113128
rect 203386 113116 203392 113128
rect 198568 113088 203392 113116
rect 198568 113076 198574 113088
rect 203386 113076 203392 113088
rect 203444 113076 203450 113128
rect 195750 113008 195756 113060
rect 195808 113048 195814 113060
rect 199338 113048 199344 113060
rect 195808 113020 199344 113048
rect 195808 113008 195814 113020
rect 199338 113008 199344 113020
rect 199396 113008 199402 113060
rect 72010 112940 72016 112992
rect 72068 112980 72074 112992
rect 72838 112980 72844 112992
rect 72068 112952 72844 112980
rect 72068 112940 72074 112952
rect 72838 112940 72844 112952
rect 72896 112980 72902 112992
rect 103658 112980 103664 112992
rect 72896 112952 103664 112980
rect 72896 112940 72902 112952
rect 103658 112940 103664 112952
rect 103716 112940 103722 112992
rect 132638 112940 132644 112992
rect 132696 112980 132702 112992
rect 164838 112980 164844 112992
rect 132696 112952 164844 112980
rect 132696 112940 132702 112952
rect 164838 112940 164844 112952
rect 164896 112940 164902 112992
rect 198878 112940 198884 112992
rect 198936 112980 198942 112992
rect 203938 112980 203944 112992
rect 198936 112952 203944 112980
rect 198936 112940 198942 112952
rect 203938 112940 203944 112952
rect 203996 112940 204002 112992
rect 196118 112872 196124 112924
rect 196176 112912 196182 112924
rect 199982 112912 199988 112924
rect 196176 112884 199988 112912
rect 196176 112872 196182 112884
rect 199982 112872 199988 112884
rect 200040 112872 200046 112924
rect 81670 112736 81676 112788
rect 81728 112776 81734 112788
rect 82498 112776 82504 112788
rect 81728 112748 82504 112776
rect 81728 112736 81734 112748
rect 82498 112736 82504 112748
rect 82556 112736 82562 112788
rect 194554 112736 194560 112788
rect 194612 112776 194618 112788
rect 197682 112776 197688 112788
rect 194612 112748 197688 112776
rect 194612 112736 194618 112748
rect 197682 112736 197688 112748
rect 197740 112736 197746 112788
rect 197314 112600 197320 112652
rect 197372 112640 197378 112652
rect 201638 112640 201644 112652
rect 197372 112612 201644 112640
rect 197372 112600 197378 112612
rect 201638 112600 201644 112612
rect 201696 112600 201702 112652
rect 190506 112532 190512 112584
rect 190564 112572 190570 112584
rect 191978 112572 191984 112584
rect 190564 112544 191984 112572
rect 190564 112532 190570 112544
rect 191978 112532 191984 112544
rect 192036 112532 192042 112584
rect 192530 112532 192536 112584
rect 192588 112572 192594 112584
rect 194738 112572 194744 112584
rect 192588 112544 194744 112572
rect 192588 112532 192594 112544
rect 194738 112532 194744 112544
rect 194796 112532 194802 112584
rect 196486 112532 196492 112584
rect 196544 112572 196550 112584
rect 200534 112572 200540 112584
rect 196544 112544 200540 112572
rect 196544 112532 196550 112544
rect 200534 112532 200540 112544
rect 200592 112532 200598 112584
rect 190138 112464 190144 112516
rect 190196 112504 190202 112516
rect 191426 112504 191432 112516
rect 190196 112476 191432 112504
rect 190196 112464 190202 112476
rect 191426 112464 191432 112476
rect 191484 112464 191490 112516
rect 196946 112464 196952 112516
rect 197004 112504 197010 112516
rect 201086 112504 201092 112516
rect 197004 112476 201092 112504
rect 197004 112464 197010 112476
rect 201086 112464 201092 112476
rect 201144 112464 201150 112516
rect 189678 112396 189684 112448
rect 189736 112436 189742 112448
rect 190782 112436 190788 112448
rect 189736 112408 190788 112436
rect 189736 112396 189742 112408
rect 190782 112396 190788 112408
rect 190840 112396 190846 112448
rect 192898 112396 192904 112448
rect 192956 112436 192962 112448
rect 192956 112408 194416 112436
rect 192956 112396 192962 112408
rect 193174 112328 193180 112380
rect 193232 112368 193238 112380
rect 194186 112368 194192 112380
rect 193232 112340 194192 112368
rect 193232 112328 193238 112340
rect 194186 112328 194192 112340
rect 194244 112328 194250 112380
rect 103658 112260 103664 112312
rect 103716 112300 103722 112312
rect 109454 112300 109460 112312
rect 103716 112272 109460 112300
rect 103716 112260 103722 112272
rect 109454 112260 109460 112272
rect 109512 112300 109518 112312
rect 132086 112300 132092 112312
rect 109512 112272 132092 112300
rect 109512 112260 109518 112272
rect 132086 112260 132092 112272
rect 132144 112260 132150 112312
rect 194388 112300 194416 112408
rect 197498 112396 197504 112448
rect 197556 112436 197562 112448
rect 201638 112436 201644 112448
rect 197556 112408 201644 112436
rect 197556 112396 197562 112408
rect 201638 112396 201644 112408
rect 201696 112396 201702 112448
rect 198142 112328 198148 112380
rect 198200 112368 198206 112380
rect 202834 112368 202840 112380
rect 198200 112340 202840 112368
rect 198200 112328 198206 112340
rect 202834 112328 202840 112340
rect 202892 112328 202898 112380
rect 195382 112300 195388 112312
rect 194388 112272 195388 112300
rect 195382 112260 195388 112272
rect 195440 112260 195446 112312
rect 110006 112192 110012 112244
rect 110064 112232 110070 112244
rect 132638 112232 132644 112244
rect 110064 112204 132644 112232
rect 110064 112192 110070 112204
rect 132638 112192 132644 112204
rect 132696 112192 132702 112244
rect 194186 112192 194192 112244
rect 194244 112232 194250 112244
rect 195934 112232 195940 112244
rect 194244 112204 195940 112232
rect 194244 112192 194250 112204
rect 195934 112192 195940 112204
rect 195992 112192 195998 112244
rect 52598 112124 52604 112176
rect 52656 112164 52662 112176
rect 57014 112164 57020 112176
rect 52656 112136 57020 112164
rect 52656 112124 52662 112136
rect 57014 112124 57020 112136
rect 57072 112124 57078 112176
rect 81670 112124 81676 112176
rect 81728 112164 81734 112176
rect 110466 112164 110472 112176
rect 81728 112136 110472 112164
rect 81728 112124 81734 112136
rect 110466 112124 110472 112136
rect 110524 112124 110530 112176
rect 121046 112124 121052 112176
rect 121104 112164 121110 112176
rect 124726 112164 124732 112176
rect 121104 112136 124732 112164
rect 121104 112124 121110 112136
rect 124726 112124 124732 112136
rect 124784 112124 124790 112176
rect 51034 112056 51040 112108
rect 51092 112096 51098 112108
rect 54254 112096 54260 112108
rect 51092 112068 54260 112096
rect 51092 112056 51098 112068
rect 54254 112056 54260 112068
rect 54312 112056 54318 112108
rect 190598 112056 190604 112108
rect 190656 112096 190662 112108
rect 192254 112096 192260 112108
rect 190656 112068 192260 112096
rect 190656 112056 190662 112068
rect 192254 112056 192260 112068
rect 192312 112056 192318 112108
rect 53058 111988 53064 112040
rect 53116 112028 53122 112040
rect 57658 112028 57664 112040
rect 53116 112000 57664 112028
rect 53116 111988 53122 112000
rect 57658 111988 57664 112000
rect 57716 111988 57722 112040
rect 51862 111920 51868 111972
rect 51920 111960 51926 111972
rect 55634 111960 55640 111972
rect 51920 111932 55640 111960
rect 51920 111920 51926 111932
rect 55634 111920 55640 111932
rect 55692 111920 55698 111972
rect 122242 111920 122248 111972
rect 122300 111960 122306 111972
rect 126382 111960 126388 111972
rect 122300 111932 126388 111960
rect 122300 111920 122306 111932
rect 126382 111920 126388 111932
rect 126440 111920 126446 111972
rect 35210 111852 35216 111904
rect 35268 111892 35274 111904
rect 39810 111892 39816 111904
rect 35268 111864 39816 111892
rect 35268 111852 35274 111864
rect 39810 111852 39816 111864
rect 39868 111852 39874 111904
rect 52506 111852 52512 111904
rect 52564 111892 52570 111904
rect 56370 111892 56376 111904
rect 52564 111864 56376 111892
rect 52564 111852 52570 111864
rect 56370 111852 56376 111864
rect 56428 111852 56434 111904
rect 117826 111852 117832 111904
rect 117884 111892 117890 111904
rect 120310 111892 120316 111904
rect 117884 111864 120316 111892
rect 117884 111852 117890 111864
rect 120310 111852 120316 111864
rect 120368 111852 120374 111904
rect 123070 111892 123076 111904
rect 120420 111864 123076 111892
rect 53794 111784 53800 111836
rect 53852 111824 53858 111836
rect 59038 111824 59044 111836
rect 53852 111796 59044 111824
rect 53852 111784 53858 111796
rect 59038 111784 59044 111796
rect 59096 111784 59102 111836
rect 113042 111784 113048 111836
rect 113100 111824 113106 111836
rect 113778 111824 113784 111836
rect 113100 111796 113784 111824
rect 113100 111784 113106 111796
rect 113778 111784 113784 111796
rect 113836 111784 113842 111836
rect 119850 111784 119856 111836
rect 119908 111824 119914 111836
rect 120420 111824 120448 111864
rect 123070 111852 123076 111864
rect 123128 111852 123134 111904
rect 119908 111796 120448 111824
rect 119908 111784 119914 111796
rect 122702 111784 122708 111836
rect 122760 111824 122766 111836
rect 126934 111824 126940 111836
rect 122760 111796 126940 111824
rect 122760 111784 122766 111796
rect 126934 111784 126940 111796
rect 126992 111784 126998 111836
rect 34474 111716 34480 111768
rect 34532 111756 34538 111768
rect 39442 111756 39448 111768
rect 34532 111728 39448 111756
rect 34532 111716 34538 111728
rect 39442 111716 39448 111728
rect 39500 111716 39506 111768
rect 54254 111716 54260 111768
rect 54312 111756 54318 111768
rect 59774 111756 59780 111768
rect 54312 111728 59780 111756
rect 54312 111716 54318 111728
rect 59774 111716 59780 111728
rect 59832 111716 59838 111768
rect 120310 111716 120316 111768
rect 120368 111756 120374 111768
rect 123622 111756 123628 111768
rect 120368 111728 123628 111756
rect 120368 111716 120374 111728
rect 123622 111716 123628 111728
rect 123680 111716 123686 111768
rect 35854 111648 35860 111700
rect 35912 111688 35918 111700
rect 40270 111688 40276 111700
rect 35912 111660 40276 111688
rect 35912 111648 35918 111660
rect 40270 111648 40276 111660
rect 40328 111648 40334 111700
rect 53426 111648 53432 111700
rect 53484 111688 53490 111700
rect 58394 111688 58400 111700
rect 53484 111660 58400 111688
rect 53484 111648 53490 111660
rect 58394 111648 58400 111660
rect 58452 111648 58458 111700
rect 33830 111580 33836 111632
rect 33888 111620 33894 111632
rect 39074 111620 39080 111632
rect 33888 111592 39080 111620
rect 33888 111580 33894 111592
rect 39074 111580 39080 111592
rect 39132 111580 39138 111632
rect 54622 111580 54628 111632
rect 54680 111620 54686 111632
rect 60418 111620 60424 111632
rect 54680 111592 60424 111620
rect 54680 111580 54686 111592
rect 60418 111580 60424 111592
rect 60476 111580 60482 111632
rect 123070 111580 123076 111632
rect 123128 111620 123134 111632
rect 127486 111620 127492 111632
rect 123128 111592 127492 111620
rect 123128 111580 123134 111592
rect 127486 111580 127492 111592
rect 127544 111580 127550 111632
rect 37878 111512 37884 111564
rect 37936 111552 37942 111564
rect 41466 111552 41472 111564
rect 37936 111524 41472 111552
rect 37936 111512 37942 111524
rect 41466 111512 41472 111524
rect 41524 111512 41530 111564
rect 123438 111512 123444 111564
rect 123496 111552 123502 111564
rect 128038 111552 128044 111564
rect 123496 111524 128044 111552
rect 123496 111512 123502 111524
rect 128038 111512 128044 111524
rect 128096 111512 128102 111564
rect 39258 111444 39264 111496
rect 39316 111484 39322 111496
rect 42202 111484 42208 111496
rect 39316 111456 42208 111484
rect 39316 111444 39322 111456
rect 42202 111444 42208 111456
rect 42260 111444 42266 111496
rect 118654 111444 118660 111496
rect 118712 111484 118718 111496
rect 121414 111484 121420 111496
rect 118712 111456 121420 111484
rect 118712 111444 118718 111456
rect 121414 111444 121420 111456
rect 121472 111444 121478 111496
rect 124266 111444 124272 111496
rect 124324 111484 124330 111496
rect 129142 111484 129148 111496
rect 124324 111456 129148 111484
rect 124324 111444 124330 111456
rect 129142 111444 129148 111456
rect 129200 111444 129206 111496
rect 39994 111376 40000 111428
rect 40052 111416 40058 111428
rect 42294 111416 42300 111428
rect 40052 111388 42300 111416
rect 40052 111376 40058 111388
rect 42294 111376 42300 111388
rect 42352 111376 42358 111428
rect 48274 111376 48280 111428
rect 48332 111416 48338 111428
rect 49470 111416 49476 111428
rect 48332 111388 49476 111416
rect 48332 111376 48338 111388
rect 49470 111376 49476 111388
rect 49528 111376 49534 111428
rect 50666 111376 50672 111428
rect 50724 111416 50730 111428
rect 53610 111416 53616 111428
rect 50724 111388 53616 111416
rect 50724 111376 50730 111388
rect 53610 111376 53616 111388
rect 53668 111376 53674 111428
rect 114238 111376 114244 111428
rect 114296 111416 114302 111428
rect 115434 111416 115440 111428
rect 114296 111388 115440 111416
rect 114296 111376 114302 111388
rect 115434 111376 115440 111388
rect 115492 111376 115498 111428
rect 116630 111376 116636 111428
rect 116688 111416 116694 111428
rect 118746 111416 118752 111428
rect 116688 111388 118752 111416
rect 116688 111376 116694 111388
rect 118746 111376 118752 111388
rect 118804 111376 118810 111428
rect 121506 111376 121512 111428
rect 121564 111416 121570 111428
rect 125278 111416 125284 111428
rect 121564 111388 125284 111416
rect 121564 111376 121570 111388
rect 125278 111376 125284 111388
rect 125336 111376 125342 111428
rect 125830 111416 125836 111428
rect 125388 111388 125836 111416
rect 40638 111308 40644 111360
rect 40696 111348 40702 111360
rect 43030 111348 43036 111360
rect 40696 111320 43036 111348
rect 40696 111308 40702 111320
rect 43030 111308 43036 111320
rect 43088 111308 43094 111360
rect 43398 111308 43404 111360
rect 43456 111348 43462 111360
rect 44594 111348 44600 111360
rect 43456 111320 44600 111348
rect 43456 111308 43462 111320
rect 44594 111308 44600 111320
rect 44652 111308 44658 111360
rect 47814 111308 47820 111360
rect 47872 111348 47878 111360
rect 48826 111348 48832 111360
rect 47872 111320 48832 111348
rect 47872 111308 47878 111320
rect 48826 111308 48832 111320
rect 48884 111308 48890 111360
rect 49838 111308 49844 111360
rect 49896 111348 49902 111360
rect 52230 111348 52236 111360
rect 49896 111320 52236 111348
rect 49896 111308 49902 111320
rect 52230 111308 52236 111320
rect 52288 111308 52294 111360
rect 113870 111308 113876 111360
rect 113928 111348 113934 111360
rect 114882 111348 114888 111360
rect 113928 111320 114888 111348
rect 113928 111308 113934 111320
rect 114882 111308 114888 111320
rect 114940 111308 114946 111360
rect 116262 111308 116268 111360
rect 116320 111348 116326 111360
rect 118194 111348 118200 111360
rect 116320 111320 118200 111348
rect 116320 111308 116326 111320
rect 118194 111308 118200 111320
rect 118252 111308 118258 111360
rect 118286 111308 118292 111360
rect 118344 111348 118350 111360
rect 120862 111348 120868 111360
rect 118344 111320 120868 111348
rect 118344 111308 118350 111320
rect 120862 111308 120868 111320
rect 120920 111308 120926 111360
rect 121874 111308 121880 111360
rect 121932 111348 121938 111360
rect 125388 111348 125416 111388
rect 125830 111376 125836 111388
rect 125888 111376 125894 111428
rect 126290 111376 126296 111428
rect 126348 111416 126354 111428
rect 131902 111416 131908 111428
rect 126348 111388 131908 111416
rect 126348 111376 126354 111388
rect 131902 111376 131908 111388
rect 131960 111376 131966 111428
rect 182226 111376 182232 111428
rect 182284 111416 182290 111428
rect 183238 111416 183244 111428
rect 182284 111388 183244 111416
rect 182284 111376 182290 111388
rect 183238 111376 183244 111388
rect 183296 111376 183302 111428
rect 191978 111376 191984 111428
rect 192036 111416 192042 111428
rect 194278 111416 194284 111428
rect 192036 111388 194284 111416
rect 192036 111376 192042 111388
rect 194278 111376 194284 111388
rect 194336 111376 194342 111428
rect 195290 111376 195296 111428
rect 195348 111416 195354 111428
rect 198786 111416 198792 111428
rect 195348 111388 198792 111416
rect 195348 111376 195354 111388
rect 198786 111376 198792 111388
rect 198844 111376 198850 111428
rect 121932 111320 125416 111348
rect 121932 111308 121938 111320
rect 125462 111308 125468 111360
rect 125520 111348 125526 111360
rect 130798 111348 130804 111360
rect 125520 111320 130804 111348
rect 125520 111308 125526 111320
rect 130798 111308 130804 111320
rect 130856 111308 130862 111360
rect 182870 111308 182876 111360
rect 182928 111348 182934 111360
rect 183790 111348 183796 111360
rect 182928 111320 183796 111348
rect 182928 111308 182934 111320
rect 183790 111308 183796 111320
rect 183848 111308 183854 111360
rect 191702 111308 191708 111360
rect 191760 111348 191766 111360
rect 193634 111348 193640 111360
rect 191760 111320 193640 111348
rect 191760 111308 191766 111320
rect 193634 111308 193640 111320
rect 193692 111308 193698 111360
rect 194094 111308 194100 111360
rect 194152 111348 194158 111360
rect 197130 111348 197136 111360
rect 194152 111320 197136 111348
rect 194152 111308 194158 111320
rect 197130 111308 197136 111320
rect 197188 111308 197194 111360
rect 37234 111240 37240 111292
rect 37292 111280 37298 111292
rect 41006 111280 41012 111292
rect 37292 111252 41012 111280
rect 37292 111240 37298 111252
rect 41006 111240 41012 111252
rect 41064 111240 41070 111292
rect 48642 111240 48648 111292
rect 48700 111280 48706 111292
rect 50206 111280 50212 111292
rect 48700 111252 50212 111280
rect 48700 111240 48706 111252
rect 50206 111240 50212 111252
rect 50264 111240 50270 111292
rect 51402 111240 51408 111292
rect 51460 111280 51466 111292
rect 54990 111280 54996 111292
rect 51460 111252 54996 111280
rect 51460 111240 51466 111252
rect 54990 111240 54996 111252
rect 55048 111240 55054 111292
rect 114698 111240 114704 111292
rect 114756 111280 114762 111292
rect 115986 111280 115992 111292
rect 114756 111252 115992 111280
rect 114756 111240 114762 111252
rect 115986 111240 115992 111252
rect 116044 111240 116050 111292
rect 117458 111240 117464 111292
rect 117516 111280 117522 111292
rect 119758 111280 119764 111292
rect 117516 111252 119764 111280
rect 117516 111240 117522 111252
rect 119758 111240 119764 111252
rect 119816 111240 119822 111292
rect 120678 111240 120684 111292
rect 120736 111280 120742 111292
rect 124174 111280 124180 111292
rect 120736 111252 124180 111280
rect 120736 111240 120742 111252
rect 124174 111240 124180 111252
rect 124232 111240 124238 111292
rect 125094 111240 125100 111292
rect 125152 111280 125158 111292
rect 130246 111280 130252 111292
rect 125152 111252 130252 111280
rect 125152 111240 125158 111252
rect 130246 111240 130252 111252
rect 130304 111240 130310 111292
rect 36590 111172 36596 111224
rect 36648 111212 36654 111224
rect 40638 111212 40644 111224
rect 36648 111184 40644 111212
rect 36648 111172 36654 111184
rect 40638 111172 40644 111184
rect 40696 111172 40702 111224
rect 41282 111172 41288 111224
rect 41340 111212 41346 111224
rect 43398 111212 43404 111224
rect 41340 111184 43404 111212
rect 41340 111172 41346 111184
rect 43398 111172 43404 111184
rect 43456 111172 43462 111224
rect 44318 111172 44324 111224
rect 44376 111212 44382 111224
rect 45054 111212 45060 111224
rect 44376 111184 45060 111212
rect 44376 111172 44382 111184
rect 45054 111172 45060 111184
rect 45112 111172 45118 111224
rect 49470 111172 49476 111224
rect 49528 111212 49534 111224
rect 51586 111212 51592 111224
rect 49528 111184 51592 111212
rect 49528 111172 49534 111184
rect 51586 111172 51592 111184
rect 51644 111172 51650 111224
rect 115434 111172 115440 111224
rect 115492 111212 115498 111224
rect 117090 111212 117096 111224
rect 115492 111184 117096 111212
rect 115492 111172 115498 111184
rect 117090 111172 117096 111184
rect 117148 111172 117154 111224
rect 119482 111172 119488 111224
rect 119540 111212 119546 111224
rect 122518 111212 122524 111224
rect 119540 111184 122524 111212
rect 119540 111172 119546 111184
rect 122518 111172 122524 111184
rect 122576 111172 122582 111224
rect 124634 111172 124640 111224
rect 124692 111212 124698 111224
rect 129694 111212 129700 111224
rect 124692 111184 129700 111212
rect 124692 111172 124698 111184
rect 129694 111172 129700 111184
rect 129752 111172 129758 111224
rect 177442 111172 177448 111224
rect 177500 111212 177506 111224
rect 178270 111212 178276 111224
rect 177500 111184 178276 111212
rect 177500 111172 177506 111184
rect 178270 111172 178276 111184
rect 178328 111172 178334 111224
rect 42018 111104 42024 111156
rect 42076 111144 42082 111156
rect 43858 111144 43864 111156
rect 42076 111116 43864 111144
rect 42076 111104 42082 111116
rect 43858 111104 43864 111116
rect 43916 111104 43922 111156
rect 50206 111104 50212 111156
rect 50264 111144 50270 111156
rect 52966 111144 52972 111156
rect 50264 111116 52972 111144
rect 50264 111104 50270 111116
rect 52966 111104 52972 111116
rect 53024 111104 53030 111156
rect 105406 111104 105412 111156
rect 105464 111144 105470 111156
rect 107154 111144 107160 111156
rect 105464 111116 107160 111144
rect 105464 111104 105470 111116
rect 107154 111104 107160 111116
rect 107212 111104 107218 111156
rect 119114 111104 119120 111156
rect 119172 111144 119178 111156
rect 121966 111144 121972 111156
rect 119172 111116 121972 111144
rect 119172 111104 119178 111116
rect 121966 111104 121972 111116
rect 122024 111104 122030 111156
rect 123898 111104 123904 111156
rect 123956 111144 123962 111156
rect 128590 111144 128596 111156
rect 123956 111116 128596 111144
rect 123956 111104 123962 111116
rect 128590 111104 128596 111116
rect 128648 111104 128654 111156
rect 177074 111104 177080 111156
rect 177132 111144 177138 111156
rect 178822 111144 178828 111156
rect 177132 111116 178828 111144
rect 177132 111104 177138 111116
rect 178822 111104 178828 111116
rect 178880 111104 178886 111156
rect 38614 111036 38620 111088
rect 38672 111076 38678 111088
rect 41834 111076 41840 111088
rect 38672 111048 41840 111076
rect 38672 111036 38678 111048
rect 41834 111036 41840 111048
rect 41892 111036 41898 111088
rect 49010 111036 49016 111088
rect 49068 111076 49074 111088
rect 50850 111076 50856 111088
rect 49068 111048 50856 111076
rect 49068 111036 49074 111048
rect 50850 111036 50856 111048
rect 50908 111036 50914 111088
rect 105682 111036 105688 111088
rect 105740 111076 105746 111088
rect 107706 111076 107712 111088
rect 105740 111048 107712 111076
rect 105740 111036 105746 111048
rect 107706 111036 107712 111048
rect 107764 111036 107770 111088
rect 115894 111036 115900 111088
rect 115952 111076 115958 111088
rect 117642 111076 117648 111088
rect 115952 111048 117648 111076
rect 115952 111036 115958 111048
rect 117642 111036 117648 111048
rect 117700 111036 117706 111088
rect 126658 111036 126664 111088
rect 126716 111076 126722 111088
rect 132178 111076 132184 111088
rect 126716 111048 132184 111076
rect 126716 111036 126722 111048
rect 132178 111036 132184 111048
rect 132236 111036 132242 111088
rect 176982 111036 176988 111088
rect 177040 111076 177046 111088
rect 179374 111076 179380 111088
rect 177040 111048 179380 111076
rect 177040 111036 177046 111048
rect 179374 111036 179380 111048
rect 179432 111036 179438 111088
rect 42662 110968 42668 111020
rect 42720 111008 42726 111020
rect 44226 111008 44232 111020
rect 42720 110980 44232 111008
rect 42720 110968 42726 110980
rect 44226 110968 44232 110980
rect 44284 110968 44290 111020
rect 105222 110968 105228 111020
rect 105280 111008 105286 111020
rect 106602 111008 106608 111020
rect 105280 110980 106608 111008
rect 105280 110968 105286 110980
rect 106602 110968 106608 110980
rect 106660 110968 106666 111020
rect 108810 111008 108816 111020
rect 106712 110980 108816 111008
rect 105774 110900 105780 110952
rect 105832 110940 105838 110952
rect 106712 110940 106740 110980
rect 108810 110968 108816 110980
rect 108868 110968 108874 111020
rect 115066 110968 115072 111020
rect 115124 111008 115130 111020
rect 116538 111008 116544 111020
rect 115124 110980 116544 111008
rect 115124 110968 115130 110980
rect 116538 110968 116544 110980
rect 116596 110968 116602 111020
rect 117090 110968 117096 111020
rect 117148 111008 117154 111020
rect 119206 111008 119212 111020
rect 117148 110980 119212 111008
rect 117148 110968 117154 110980
rect 119206 110968 119212 110980
rect 119264 110968 119270 111020
rect 125830 110968 125836 111020
rect 125888 111008 125894 111020
rect 131350 111008 131356 111020
rect 125888 110980 131356 111008
rect 125888 110968 125894 110980
rect 131350 110968 131356 110980
rect 131408 110968 131414 111020
rect 177258 110968 177264 111020
rect 177316 111008 177322 111020
rect 180018 111008 180024 111020
rect 177316 110980 180024 111008
rect 177316 110968 177322 110980
rect 180018 110968 180024 110980
rect 180076 110968 180082 111020
rect 181674 110968 181680 111020
rect 181732 111008 181738 111020
rect 183100 111008 183106 111020
rect 181732 110980 183106 111008
rect 181732 110968 181738 110980
rect 183100 110968 183106 110980
rect 183158 110968 183164 111020
rect 183422 110968 183428 111020
rect 183480 111008 183486 111020
rect 184296 111008 184302 111020
rect 183480 110980 184302 111008
rect 183480 110968 183486 110980
rect 184296 110968 184302 110980
rect 184354 110968 184360 111020
rect 105832 110912 106740 110940
rect 105832 110900 105838 110912
rect 177718 110900 177724 110952
rect 177776 110940 177782 110952
rect 181122 110940 181128 110952
rect 177776 110912 181128 110940
rect 177776 110900 177782 110912
rect 181122 110900 181128 110912
rect 181180 110900 181186 110952
rect 222706 110220 222712 110272
rect 222764 110260 222770 110272
rect 222801 110263 222859 110269
rect 222801 110260 222813 110263
rect 222764 110232 222813 110260
rect 222764 110220 222770 110232
rect 222801 110229 222813 110232
rect 222847 110229 222859 110263
rect 222801 110223 222859 110229
rect 177166 109472 177172 109524
rect 177224 109512 177230 109524
rect 180570 109512 180576 109524
rect 177224 109484 180576 109512
rect 177224 109472 177230 109484
rect 180570 109472 180576 109484
rect 180628 109472 180634 109524
rect 105314 109132 105320 109184
rect 105372 109172 105378 109184
rect 108258 109172 108264 109184
rect 105372 109144 108264 109172
rect 105372 109132 105378 109144
rect 108258 109132 108264 109144
rect 108316 109132 108322 109184
rect 222798 107948 222804 107960
rect 222759 107920 222804 107948
rect 222798 107908 222804 107920
rect 222856 107908 222862 107960
rect 106418 107160 106424 107212
rect 106476 107200 106482 107212
rect 107890 107200 107896 107212
rect 106476 107172 107896 107200
rect 106476 107160 106482 107172
rect 107890 107160 107896 107172
rect 107948 107160 107954 107212
rect 177534 106820 177540 106872
rect 177592 106860 177598 106872
rect 179650 106860 179656 106872
rect 177592 106832 179656 106860
rect 177592 106820 177598 106832
rect 179650 106820 179656 106832
rect 179708 106820 179714 106872
rect 32634 104032 32640 104084
rect 32692 104072 32698 104084
rect 37418 104072 37424 104084
rect 32692 104044 37424 104072
rect 32692 104032 32698 104044
rect 37418 104032 37424 104044
rect 37476 104032 37482 104084
rect 56830 104032 56836 104084
rect 56888 104072 56894 104084
rect 59866 104072 59872 104084
rect 56888 104044 59872 104072
rect 56888 104032 56894 104044
rect 59866 104032 59872 104044
rect 59924 104032 59930 104084
rect 105774 104032 105780 104084
rect 105832 104072 105838 104084
rect 108442 104072 108448 104084
rect 105832 104044 108448 104072
rect 105832 104032 105838 104044
rect 108442 104032 108448 104044
rect 108500 104032 108506 104084
rect 177810 104032 177816 104084
rect 177868 104072 177874 104084
rect 179650 104072 179656 104084
rect 177868 104044 179656 104072
rect 177868 104032 177874 104044
rect 179650 104032 179656 104044
rect 179708 104032 179714 104084
rect 106326 101312 106332 101364
rect 106384 101352 106390 101364
rect 107890 101352 107896 101364
rect 106384 101324 107896 101352
rect 106384 101312 106390 101324
rect 107890 101312 107896 101324
rect 107948 101312 107954 101364
rect 177626 101312 177632 101364
rect 177684 101352 177690 101364
rect 179650 101352 179656 101364
rect 177684 101324 179656 101352
rect 177684 101312 177690 101324
rect 179650 101312 179656 101324
rect 179708 101312 179714 101364
rect 105958 101244 105964 101296
rect 106016 101284 106022 101296
rect 108534 101284 108540 101296
rect 106016 101256 108540 101284
rect 106016 101244 106022 101256
rect 108534 101244 108540 101256
rect 108592 101244 108598 101296
rect 176982 101244 176988 101296
rect 177040 101284 177046 101296
rect 180294 101284 180300 101296
rect 177040 101256 180300 101284
rect 177040 101244 177046 101256
rect 180294 101244 180300 101256
rect 180352 101244 180358 101296
rect 106418 99884 106424 99936
rect 106476 99924 106482 99936
rect 107890 99924 107896 99936
rect 106476 99896 107896 99924
rect 106476 99884 106482 99896
rect 107890 99884 107896 99896
rect 107948 99884 107954 99936
rect 177718 99884 177724 99936
rect 177776 99924 177782 99936
rect 179650 99924 179656 99936
rect 177776 99896 179656 99924
rect 177776 99884 177782 99896
rect 179650 99884 179656 99896
rect 179708 99884 179714 99936
rect 106234 97640 106240 97692
rect 106292 97680 106298 97692
rect 107890 97680 107896 97692
rect 106292 97652 107896 97680
rect 106292 97640 106298 97652
rect 107890 97640 107896 97652
rect 107948 97640 107954 97692
rect 177534 97164 177540 97216
rect 177592 97204 177598 97216
rect 179650 97204 179656 97216
rect 177592 97176 179656 97204
rect 177592 97164 177598 97176
rect 179650 97164 179656 97176
rect 179708 97164 179714 97216
rect 222982 97096 222988 97148
rect 223040 97136 223046 97148
rect 223534 97136 223540 97148
rect 223040 97108 223540 97136
rect 223040 97096 223046 97108
rect 223534 97096 223540 97108
rect 223592 97096 223598 97148
rect 132362 95776 132368 95788
rect 132323 95748 132368 95776
rect 132362 95736 132368 95748
rect 132420 95736 132426 95788
rect 106510 94784 106516 94836
rect 106568 94824 106574 94836
rect 108442 94824 108448 94836
rect 106568 94796 108448 94824
rect 106568 94784 106574 94796
rect 108442 94784 108448 94796
rect 108500 94784 108506 94836
rect 177442 94308 177448 94360
rect 177500 94348 177506 94360
rect 179558 94348 179564 94360
rect 177500 94320 179564 94348
rect 177500 94308 177506 94320
rect 179558 94308 179564 94320
rect 179616 94308 179622 94360
rect 222798 92540 222804 92592
rect 222856 92580 222862 92592
rect 223534 92580 223540 92592
rect 222856 92552 223540 92580
rect 222856 92540 222862 92552
rect 223534 92540 223540 92552
rect 223592 92540 223598 92592
rect 105866 91656 105872 91708
rect 105924 91696 105930 91708
rect 107798 91696 107804 91708
rect 105924 91668 107804 91696
rect 105924 91656 105930 91668
rect 107798 91656 107804 91668
rect 107856 91656 107862 91708
rect 177534 91656 177540 91708
rect 177592 91696 177598 91708
rect 179558 91696 179564 91708
rect 177592 91668 179564 91696
rect 177592 91656 177598 91668
rect 179558 91656 179564 91668
rect 179616 91656 179622 91708
rect 201086 91588 201092 91640
rect 201144 91628 201150 91640
rect 204490 91628 204496 91640
rect 201144 91600 204496 91628
rect 201144 91588 201150 91600
rect 204490 91588 204496 91600
rect 204548 91588 204554 91640
rect 28862 90228 28868 90280
rect 28920 90268 28926 90280
rect 36406 90268 36412 90280
rect 28920 90240 36412 90268
rect 28920 90228 28926 90240
rect 36406 90228 36412 90240
rect 36464 90228 36470 90280
rect 54809 90271 54867 90277
rect 54809 90237 54821 90271
rect 54855 90268 54867 90271
rect 59590 90268 59596 90280
rect 54855 90240 59596 90268
rect 54855 90237 54867 90240
rect 54809 90231 54867 90237
rect 59590 90228 59596 90240
rect 59648 90228 59654 90280
rect 105222 90228 105228 90280
rect 105280 90268 105286 90280
rect 107890 90268 107896 90280
rect 105280 90240 107896 90268
rect 105280 90228 105286 90240
rect 107890 90228 107896 90240
rect 107948 90228 107954 90280
rect 177350 90228 177356 90280
rect 177408 90268 177414 90280
rect 179650 90268 179656 90280
rect 177408 90240 179656 90268
rect 177408 90228 177414 90240
rect 179650 90228 179656 90240
rect 179708 90228 179714 90280
rect 105130 89208 105136 89260
rect 105188 89248 105194 89260
rect 107798 89248 107804 89260
rect 105188 89220 107804 89248
rect 105188 89208 105194 89220
rect 107798 89208 107804 89220
rect 107856 89208 107862 89260
rect 177350 89140 177356 89192
rect 177408 89180 177414 89192
rect 179558 89180 179564 89192
rect 177408 89152 179564 89180
rect 177408 89140 177414 89152
rect 179558 89140 179564 89152
rect 179616 89140 179622 89192
rect 132365 88775 132423 88781
rect 132365 88741 132377 88775
rect 132411 88772 132423 88775
rect 132546 88772 132552 88784
rect 132411 88744 132552 88772
rect 132411 88741 132423 88744
rect 132365 88735 132423 88741
rect 132546 88732 132552 88744
rect 132604 88732 132610 88784
rect 177350 88188 177356 88240
rect 177408 88228 177414 88240
rect 179466 88228 179472 88240
rect 177408 88200 179472 88228
rect 177408 88188 177414 88200
rect 179466 88188 179472 88200
rect 179524 88188 179530 88240
rect 105866 87712 105872 87764
rect 105924 87752 105930 87764
rect 107706 87752 107712 87764
rect 105924 87724 107712 87752
rect 105924 87712 105930 87724
rect 107706 87712 107712 87724
rect 107764 87712 107770 87764
rect 54806 86120 54812 86132
rect 54767 86092 54812 86120
rect 54806 86080 54812 86092
rect 54864 86080 54870 86132
rect 105590 86080 105596 86132
rect 105648 86120 105654 86132
rect 108718 86120 108724 86132
rect 105648 86092 108724 86120
rect 105648 86080 105654 86092
rect 108718 86080 108724 86092
rect 108776 86080 108782 86132
rect 178086 86080 178092 86132
rect 178144 86120 178150 86132
rect 180478 86120 180484 86132
rect 178144 86092 180484 86120
rect 178144 86080 178150 86092
rect 180478 86080 180484 86092
rect 180536 86080 180542 86132
rect 222798 84788 222804 84840
rect 222856 84828 222862 84840
rect 223534 84828 223540 84840
rect 222856 84800 223540 84828
rect 222856 84788 222862 84800
rect 223534 84788 223540 84800
rect 223592 84788 223598 84840
rect 106326 84720 106332 84772
rect 106384 84760 106390 84772
rect 108810 84760 108816 84772
rect 106384 84732 108816 84760
rect 106384 84720 106390 84732
rect 108810 84720 108816 84732
rect 108868 84720 108874 84772
rect 177534 84720 177540 84772
rect 177592 84760 177598 84772
rect 179650 84760 179656 84772
rect 177592 84732 179656 84760
rect 177592 84720 177598 84732
rect 179650 84720 179656 84732
rect 179708 84720 179714 84772
rect 178178 83632 178184 83684
rect 178236 83672 178242 83684
rect 180386 83672 180392 83684
rect 178236 83644 180392 83672
rect 178236 83632 178242 83644
rect 180386 83632 180392 83644
rect 180444 83632 180450 83684
rect 105590 83360 105596 83412
rect 105648 83400 105654 83412
rect 108626 83400 108632 83412
rect 105648 83372 108632 83400
rect 105648 83360 105654 83372
rect 108626 83360 108632 83372
rect 108684 83360 108690 83412
rect 105498 82000 105504 82052
rect 105556 82040 105562 82052
rect 108534 82040 108540 82052
rect 105556 82012 108540 82040
rect 105556 82000 105562 82012
rect 108534 82000 108540 82012
rect 108592 82000 108598 82052
rect 177718 82000 177724 82052
rect 177776 82040 177782 82052
rect 180294 82040 180300 82052
rect 177776 82012 180300 82040
rect 177776 82000 177782 82012
rect 180294 82000 180300 82012
rect 180352 82000 180358 82052
rect 106510 81932 106516 81984
rect 106568 81972 106574 81984
rect 107890 81972 107896 81984
rect 106568 81944 107896 81972
rect 106568 81932 106574 81944
rect 107890 81932 107896 81944
rect 107948 81932 107954 81984
rect 105222 80572 105228 80624
rect 105280 80612 105286 80624
rect 108074 80612 108080 80624
rect 105280 80584 108080 80612
rect 105280 80572 105286 80584
rect 108074 80572 108080 80584
rect 108132 80572 108138 80624
rect 177350 80572 177356 80624
rect 177408 80612 177414 80624
rect 180018 80612 180024 80624
rect 177408 80584 180024 80612
rect 177408 80572 177414 80584
rect 180018 80572 180024 80584
rect 180076 80572 180082 80624
rect 105130 79688 105136 79740
rect 105188 79728 105194 79740
rect 107522 79728 107528 79740
rect 105188 79700 107528 79728
rect 105188 79688 105194 79700
rect 107522 79688 107528 79700
rect 107580 79688 107586 79740
rect 132546 79280 132552 79332
rect 132604 79280 132610 79332
rect 54806 79252 54812 79264
rect 54767 79224 54812 79252
rect 54806 79212 54812 79224
rect 54864 79212 54870 79264
rect 132564 79196 132592 79280
rect 178178 79212 178184 79264
rect 178236 79252 178242 79264
rect 179374 79252 179380 79264
rect 178236 79224 179380 79252
rect 178236 79212 178242 79224
rect 179374 79212 179380 79224
rect 179432 79212 179438 79264
rect 132546 79144 132552 79196
rect 132604 79144 132610 79196
rect 30518 77784 30524 77836
rect 30576 77824 30582 77836
rect 37418 77824 37424 77836
rect 30576 77796 37424 77824
rect 30576 77784 30582 77796
rect 37418 77784 37424 77796
rect 37476 77784 37482 77836
rect 57474 77580 57480 77632
rect 57532 77620 57538 77632
rect 59590 77620 59596 77632
rect 57532 77592 59596 77620
rect 57532 77580 57538 77592
rect 59590 77580 59596 77592
rect 59648 77580 59654 77632
rect 54806 76464 54812 76476
rect 54767 76436 54812 76464
rect 54806 76424 54812 76436
rect 54864 76424 54870 76476
rect 222982 75064 222988 75116
rect 223040 75104 223046 75116
rect 223534 75104 223540 75116
rect 223040 75076 223540 75104
rect 223040 75064 223046 75076
rect 223534 75064 223540 75076
rect 223592 75064 223598 75116
rect 222798 73568 222804 73620
rect 222856 73608 222862 73620
rect 223074 73608 223080 73620
rect 222856 73580 223080 73608
rect 222856 73568 222862 73580
rect 223074 73568 223080 73580
rect 223132 73568 223138 73620
rect 103198 72344 103204 72396
rect 103256 72384 103262 72396
rect 108350 72384 108356 72396
rect 103256 72356 108356 72384
rect 103256 72344 103262 72356
rect 108350 72344 108356 72356
rect 108408 72344 108414 72396
rect 177350 72344 177356 72396
rect 177408 72384 177414 72396
rect 180570 72384 180576 72396
rect 177408 72356 180576 72384
rect 177408 72344 177414 72356
rect 180570 72344 180576 72356
rect 180628 72344 180634 72396
rect 178362 70848 178368 70900
rect 178420 70888 178426 70900
rect 181122 70888 181128 70900
rect 178420 70860 181128 70888
rect 178420 70848 178426 70860
rect 181122 70848 181128 70860
rect 181180 70848 181186 70900
rect 106510 70508 106516 70560
rect 106568 70548 106574 70560
rect 109270 70548 109276 70560
rect 106568 70520 109276 70548
rect 106568 70508 106574 70520
rect 109270 70508 109276 70520
rect 109328 70508 109334 70560
rect 90134 69760 90140 69812
rect 90192 69800 90198 69812
rect 96761 69803 96819 69809
rect 96761 69800 96773 69803
rect 90192 69772 96773 69800
rect 90192 69760 90198 69772
rect 96761 69769 96773 69772
rect 96807 69769 96819 69803
rect 96761 69763 96819 69769
rect 49381 69735 49439 69741
rect 49381 69701 49393 69735
rect 49427 69732 49439 69735
rect 54806 69732 54812 69744
rect 49427 69704 54812 69732
rect 49427 69701 49439 69704
rect 49381 69695 49439 69701
rect 54806 69692 54812 69704
rect 54864 69692 54870 69744
rect 59038 69596 59044 69608
rect 57216 69568 59044 69596
rect 22238 69488 22244 69540
rect 22296 69528 22302 69540
rect 28678 69528 28684 69540
rect 22296 69500 28684 69528
rect 22296 69488 22302 69500
rect 28678 69488 28684 69500
rect 28736 69488 28742 69540
rect 36038 69488 36044 69540
rect 36096 69528 36102 69540
rect 40270 69528 40276 69540
rect 36096 69500 40276 69528
rect 36096 69488 36102 69500
rect 40270 69488 40276 69500
rect 40328 69488 40334 69540
rect 53794 69488 53800 69540
rect 53852 69528 53858 69540
rect 57216 69528 57244 69568
rect 59038 69556 59044 69568
rect 59096 69556 59102 69608
rect 131626 69596 131632 69608
rect 131276 69568 131632 69596
rect 53852 69500 57244 69528
rect 53852 69488 53858 69500
rect 126290 69488 126296 69540
rect 126348 69528 126354 69540
rect 131276 69528 131304 69568
rect 131626 69556 131632 69568
rect 131684 69556 131690 69608
rect 203938 69596 203944 69608
rect 202116 69568 203944 69596
rect 126348 69500 131304 69528
rect 126348 69488 126354 69500
rect 198878 69488 198884 69540
rect 198936 69528 198942 69540
rect 202116 69528 202144 69568
rect 203938 69556 203944 69568
rect 203996 69556 204002 69608
rect 198936 69500 202144 69528
rect 198936 69488 198942 69500
rect 202190 69488 202196 69540
rect 202248 69528 202254 69540
rect 202248 69500 209964 69528
rect 202248 69488 202254 69500
rect 16626 69420 16632 69472
rect 16684 69460 16690 69472
rect 31898 69460 31904 69472
rect 16684 69432 31904 69460
rect 16684 69420 16690 69432
rect 31898 69420 31904 69432
rect 31956 69420 31962 69472
rect 35578 69420 35584 69472
rect 35636 69460 35642 69472
rect 39810 69460 39816 69472
rect 35636 69432 39816 69460
rect 35636 69420 35642 69432
rect 39810 69420 39816 69432
rect 39868 69420 39874 69472
rect 54254 69420 54260 69472
rect 54312 69460 54318 69472
rect 59406 69460 59412 69472
rect 54312 69432 59412 69460
rect 54312 69420 54318 69432
rect 59406 69420 59412 69432
rect 59464 69420 59470 69472
rect 198510 69420 198516 69472
rect 198568 69460 198574 69472
rect 202926 69460 202932 69472
rect 198568 69432 202932 69460
rect 198568 69420 198574 69432
rect 202926 69420 202932 69432
rect 202984 69420 202990 69472
rect 209936 69460 209964 69500
rect 210562 69460 210568 69472
rect 209936 69432 210568 69460
rect 210562 69420 210568 69432
rect 210620 69420 210626 69472
rect 34106 69352 34112 69404
rect 34164 69392 34170 69404
rect 39074 69392 39080 69404
rect 34164 69364 39080 69392
rect 34164 69352 34170 69364
rect 39074 69352 39080 69364
rect 39132 69352 39138 69404
rect 55358 69352 55364 69404
rect 55416 69392 55422 69404
rect 60142 69392 60148 69404
rect 55416 69364 60148 69392
rect 55416 69352 55422 69364
rect 60142 69352 60148 69364
rect 60200 69352 60206 69404
rect 196118 69352 196124 69404
rect 196176 69392 196182 69404
rect 199982 69392 199988 69404
rect 196176 69364 199988 69392
rect 196176 69352 196182 69364
rect 199982 69352 199988 69364
rect 200040 69352 200046 69404
rect 34658 69284 34664 69336
rect 34716 69324 34722 69336
rect 39442 69324 39448 69336
rect 34716 69296 39448 69324
rect 34716 69284 34722 69296
rect 39442 69284 39448 69296
rect 39500 69284 39506 69336
rect 53426 69284 53432 69336
rect 53484 69324 53490 69336
rect 58118 69324 58124 69336
rect 53484 69296 58124 69324
rect 53484 69284 53490 69296
rect 58118 69284 58124 69296
rect 58176 69284 58182 69336
rect 120310 69284 120316 69336
rect 120368 69324 120374 69336
rect 123070 69324 123076 69336
rect 120368 69296 123076 69324
rect 120368 69284 120374 69296
rect 123070 69284 123076 69296
rect 123128 69284 123134 69336
rect 200994 69284 201000 69336
rect 201052 69324 201058 69336
rect 215898 69324 215904 69336
rect 201052 69296 215904 69324
rect 201052 69284 201058 69296
rect 215898 69284 215904 69296
rect 215956 69284 215962 69336
rect 52230 69216 52236 69268
rect 52288 69256 52294 69268
rect 56370 69256 56376 69268
rect 52288 69228 56376 69256
rect 52288 69216 52294 69228
rect 56370 69216 56376 69228
rect 56428 69216 56434 69268
rect 125094 69216 125100 69268
rect 125152 69256 125158 69268
rect 129878 69256 129884 69268
rect 125152 69228 129884 69256
rect 125152 69216 125158 69228
rect 129878 69216 129884 69228
rect 129936 69216 129942 69268
rect 194094 69216 194100 69268
rect 194152 69256 194158 69268
rect 197130 69256 197136 69268
rect 194152 69228 197136 69256
rect 194152 69216 194158 69228
rect 197130 69216 197136 69228
rect 197188 69216 197194 69268
rect 197314 69216 197320 69268
rect 197372 69256 197378 69268
rect 201638 69256 201644 69268
rect 197372 69228 201644 69256
rect 197372 69216 197378 69228
rect 201638 69216 201644 69228
rect 201696 69216 201702 69268
rect 39994 69148 40000 69200
rect 40052 69188 40058 69200
rect 42662 69188 42668 69200
rect 40052 69160 42668 69188
rect 40052 69148 40058 69160
rect 42662 69148 42668 69160
rect 42720 69148 42726 69200
rect 51402 69148 51408 69200
rect 51460 69188 51466 69200
rect 54990 69188 54996 69200
rect 51460 69160 54996 69188
rect 51460 69148 51466 69160
rect 54990 69148 54996 69160
rect 55048 69148 55054 69200
rect 118286 69148 118292 69200
rect 118344 69188 118350 69200
rect 120310 69188 120316 69200
rect 118344 69160 120316 69188
rect 118344 69148 118350 69160
rect 120310 69148 120316 69160
rect 120368 69148 120374 69200
rect 125830 69148 125836 69200
rect 125888 69188 125894 69200
rect 131258 69188 131264 69200
rect 125888 69160 131264 69188
rect 125888 69148 125894 69160
rect 131258 69148 131264 69160
rect 131316 69148 131322 69200
rect 182226 69148 182232 69200
rect 182284 69188 182290 69200
rect 183238 69188 183244 69200
rect 182284 69160 183244 69188
rect 182284 69148 182290 69160
rect 183238 69148 183244 69160
rect 183296 69148 183302 69200
rect 192530 69148 192536 69200
rect 192588 69188 192594 69200
rect 194830 69188 194836 69200
rect 192588 69160 194836 69188
rect 192588 69148 192594 69160
rect 194830 69148 194836 69160
rect 194888 69148 194894 69200
rect 197406 69148 197412 69200
rect 197464 69188 197470 69200
rect 201822 69188 201828 69200
rect 197464 69160 201828 69188
rect 197464 69148 197470 69160
rect 201822 69148 201828 69160
rect 201880 69148 201886 69200
rect 36590 69080 36596 69132
rect 36648 69120 36654 69132
rect 40638 69120 40644 69132
rect 36648 69092 40644 69120
rect 36648 69080 36654 69092
rect 40638 69080 40644 69092
rect 40696 69080 40702 69132
rect 41282 69080 41288 69132
rect 41340 69120 41346 69132
rect 43398 69120 43404 69132
rect 41340 69092 43404 69120
rect 41340 69080 41346 69092
rect 43398 69080 43404 69092
rect 43456 69080 43462 69132
rect 49470 69080 49476 69132
rect 49528 69120 49534 69132
rect 51586 69120 51592 69132
rect 49528 69092 51592 69120
rect 49528 69080 49534 69092
rect 51586 69080 51592 69092
rect 51644 69080 51650 69132
rect 51862 69080 51868 69132
rect 51920 69120 51926 69132
rect 55634 69120 55640 69132
rect 51920 69092 55640 69120
rect 51920 69080 51926 69092
rect 55634 69080 55640 69092
rect 55692 69080 55698 69132
rect 117458 69080 117464 69132
rect 117516 69120 117522 69132
rect 119022 69120 119028 69132
rect 117516 69092 119028 69120
rect 117516 69080 117522 69092
rect 119022 69080 119028 69092
rect 119080 69080 119086 69132
rect 122702 69080 122708 69132
rect 122760 69120 122766 69132
rect 126474 69120 126480 69132
rect 122760 69092 126480 69120
rect 122760 69080 122766 69092
rect 126474 69080 126480 69092
rect 126532 69080 126538 69132
rect 126658 69080 126664 69132
rect 126716 69120 126722 69132
rect 132178 69120 132184 69132
rect 126716 69092 132184 69120
rect 126716 69080 126722 69092
rect 132178 69080 132184 69092
rect 132236 69080 132242 69132
rect 181674 69080 181680 69132
rect 181732 69120 181738 69132
rect 182778 69120 182784 69132
rect 181732 69092 182784 69120
rect 181732 69080 181738 69092
rect 182778 69080 182784 69092
rect 182836 69080 182842 69132
rect 189678 69080 189684 69132
rect 189736 69120 189742 69132
rect 190690 69120 190696 69132
rect 189736 69092 190696 69120
rect 189736 69080 189742 69092
rect 190690 69080 190696 69092
rect 190748 69080 190754 69132
rect 191794 69080 191800 69132
rect 191852 69120 191858 69132
rect 194278 69120 194284 69132
rect 191852 69092 194284 69120
rect 191852 69080 191858 69092
rect 194278 69080 194284 69092
rect 194336 69080 194342 69132
rect 194554 69080 194560 69132
rect 194612 69120 194618 69132
rect 197682 69120 197688 69132
rect 194612 69092 197688 69120
rect 194612 69080 194618 69092
rect 197682 69080 197688 69092
rect 197740 69080 197746 69132
rect 198142 69080 198148 69132
rect 198200 69120 198206 69132
rect 202834 69120 202840 69132
rect 198200 69092 202840 69120
rect 198200 69080 198206 69092
rect 202834 69080 202840 69092
rect 202892 69080 202898 69132
rect 37234 69012 37240 69064
rect 37292 69052 37298 69064
rect 41006 69052 41012 69064
rect 37292 69024 41012 69052
rect 37292 69012 37298 69024
rect 41006 69012 41012 69024
rect 41064 69012 41070 69064
rect 42662 69012 42668 69064
rect 42720 69052 42726 69064
rect 44226 69052 44232 69064
rect 42720 69024 44232 69052
rect 42720 69012 42726 69024
rect 44226 69012 44232 69024
rect 44284 69012 44290 69064
rect 53058 69012 53064 69064
rect 53116 69052 53122 69064
rect 57658 69052 57664 69064
rect 53116 69024 57664 69052
rect 53116 69012 53122 69024
rect 57658 69012 57664 69024
rect 57716 69012 57722 69064
rect 62718 69012 62724 69064
rect 62776 69052 62782 69064
rect 68974 69052 68980 69064
rect 62776 69024 68980 69052
rect 62776 69012 62782 69024
rect 68974 69012 68980 69024
rect 69032 69012 69038 69064
rect 92342 69012 92348 69064
rect 92400 69052 92406 69064
rect 97034 69052 97040 69064
rect 92400 69024 97040 69052
rect 92400 69012 92406 69024
rect 97034 69012 97040 69024
rect 97092 69012 97098 69064
rect 118654 69012 118660 69064
rect 118712 69052 118718 69064
rect 120586 69052 120592 69064
rect 118712 69024 120592 69052
rect 118712 69012 118718 69024
rect 120586 69012 120592 69024
rect 120644 69012 120650 69064
rect 123714 69012 123720 69064
rect 123772 69052 123778 69064
rect 127578 69052 127584 69064
rect 123772 69024 127584 69052
rect 123772 69012 123778 69024
rect 127578 69012 127584 69024
rect 127636 69012 127642 69064
rect 192898 69012 192904 69064
rect 192956 69052 192962 69064
rect 195382 69052 195388 69064
rect 192956 69024 195388 69052
rect 192956 69012 192962 69024
rect 195382 69012 195388 69024
rect 195440 69012 195446 69064
rect 196946 69012 196952 69064
rect 197004 69052 197010 69064
rect 201086 69052 201092 69064
rect 197004 69024 201092 69052
rect 197004 69012 197010 69024
rect 201086 69012 201092 69024
rect 201144 69012 201150 69064
rect 40638 68944 40644 68996
rect 40696 68984 40702 68996
rect 43030 68984 43036 68996
rect 40696 68956 43036 68984
rect 40696 68944 40702 68956
rect 43030 68944 43036 68956
rect 43088 68944 43094 68996
rect 43398 68944 43404 68996
rect 43456 68984 43462 68996
rect 44594 68984 44600 68996
rect 43456 68956 44600 68984
rect 43456 68944 43462 68956
rect 44594 68944 44600 68956
rect 44652 68944 44658 68996
rect 47814 68944 47820 68996
rect 47872 68984 47878 68996
rect 48550 68984 48556 68996
rect 47872 68956 48556 68984
rect 47872 68944 47878 68956
rect 48550 68944 48556 68956
rect 48608 68944 48614 68996
rect 48642 68944 48648 68996
rect 48700 68984 48706 68996
rect 49930 68984 49936 68996
rect 48700 68956 49936 68984
rect 48700 68944 48706 68956
rect 49930 68944 49936 68956
rect 49988 68944 49994 68996
rect 50666 68944 50672 68996
rect 50724 68984 50730 68996
rect 53610 68984 53616 68996
rect 50724 68956 53616 68984
rect 50724 68944 50730 68956
rect 53610 68944 53616 68956
rect 53668 68944 53674 68996
rect 54622 68944 54628 68996
rect 54680 68984 54686 68996
rect 55358 68984 55364 68996
rect 54680 68956 55364 68984
rect 54680 68944 54686 68956
rect 55358 68944 55364 68956
rect 55416 68944 55422 68996
rect 88938 68944 88944 68996
rect 88996 68984 89002 68996
rect 96850 68984 96856 68996
rect 88996 68956 96856 68984
rect 88996 68944 89002 68956
rect 96850 68944 96856 68956
rect 96908 68944 96914 68996
rect 125462 68944 125468 68996
rect 125520 68984 125526 68996
rect 130430 68984 130436 68996
rect 125520 68956 130436 68984
rect 125520 68944 125526 68956
rect 130430 68944 130436 68956
rect 130488 68944 130494 68996
rect 158766 68944 158772 68996
rect 158824 68984 158830 68996
rect 165114 68984 165120 68996
rect 158824 68956 165120 68984
rect 158824 68944 158830 68956
rect 165114 68944 165120 68956
rect 165172 68944 165178 68996
rect 193358 68944 193364 68996
rect 193416 68984 193422 68996
rect 195934 68984 195940 68996
rect 193416 68956 195940 68984
rect 193416 68944 193422 68956
rect 195934 68944 195940 68956
rect 195992 68944 195998 68996
rect 196486 68944 196492 68996
rect 196544 68984 196550 68996
rect 200534 68984 200540 68996
rect 196544 68956 200540 68984
rect 196544 68944 196550 68956
rect 200534 68944 200540 68956
rect 200592 68944 200598 68996
rect 42018 68876 42024 68928
rect 42076 68916 42082 68928
rect 43858 68916 43864 68928
rect 42076 68888 43864 68916
rect 42076 68876 42082 68888
rect 43858 68876 43864 68888
rect 43916 68876 43922 68928
rect 52598 68876 52604 68928
rect 52656 68916 52662 68928
rect 56738 68916 56744 68928
rect 52656 68888 56744 68916
rect 52656 68876 52662 68888
rect 56738 68876 56744 68888
rect 56796 68876 56802 68928
rect 62902 68876 62908 68928
rect 62960 68916 62966 68928
rect 67870 68916 67876 68928
rect 62960 68888 67876 68916
rect 62960 68876 62966 68888
rect 67870 68876 67876 68888
rect 67928 68876 67934 68928
rect 83418 68876 83424 68928
rect 83476 68916 83482 68928
rect 87190 68916 87196 68928
rect 83476 68888 87196 68916
rect 83476 68876 83482 68888
rect 87190 68876 87196 68888
rect 87248 68876 87254 68928
rect 87834 68876 87840 68928
rect 87892 68916 87898 68928
rect 94734 68916 94740 68928
rect 87892 68888 94740 68916
rect 87892 68876 87898 68888
rect 94734 68876 94740 68888
rect 94792 68876 94798 68928
rect 124266 68876 124272 68928
rect 124324 68916 124330 68928
rect 128682 68916 128688 68928
rect 124324 68888 128688 68916
rect 124324 68876 124330 68888
rect 128682 68876 128688 68888
rect 128740 68876 128746 68928
rect 151038 68876 151044 68928
rect 151096 68916 151102 68928
rect 152050 68916 152056 68928
rect 151096 68888 152056 68916
rect 151096 68876 151102 68888
rect 152050 68876 152056 68888
rect 152108 68876 152114 68928
rect 159870 68876 159876 68928
rect 159928 68916 159934 68928
rect 167046 68916 167052 68928
rect 159928 68888 167052 68916
rect 159928 68876 159934 68888
rect 167046 68876 167052 68888
rect 167104 68876 167110 68928
rect 168794 68876 168800 68928
rect 168852 68916 168858 68928
rect 173854 68916 173860 68928
rect 168852 68888 173860 68916
rect 168852 68876 168858 68888
rect 173854 68876 173860 68888
rect 173912 68876 173918 68928
rect 190598 68876 190604 68928
rect 190656 68916 190662 68928
rect 192530 68916 192536 68928
rect 190656 68888 192536 68916
rect 190656 68876 190662 68888
rect 192530 68876 192536 68888
rect 192588 68876 192594 68928
rect 195750 68876 195756 68928
rect 195808 68916 195814 68928
rect 199338 68916 199344 68928
rect 195808 68888 199344 68916
rect 195808 68876 195814 68888
rect 199338 68876 199344 68888
rect 199396 68876 199402 68928
rect 31898 68808 31904 68860
rect 31956 68848 31962 68860
rect 36041 68851 36099 68857
rect 36041 68848 36053 68851
rect 31956 68820 36053 68848
rect 31956 68808 31962 68820
rect 36041 68817 36053 68820
rect 36087 68817 36099 68851
rect 36041 68811 36099 68817
rect 39258 68808 39264 68860
rect 39316 68848 39322 68860
rect 42202 68848 42208 68860
rect 39316 68820 42208 68848
rect 39316 68808 39322 68820
rect 42202 68808 42208 68820
rect 42260 68808 42266 68860
rect 51034 68808 51040 68860
rect 51092 68848 51098 68860
rect 54254 68848 54260 68860
rect 51092 68820 54260 68848
rect 51092 68808 51098 68820
rect 54254 68808 54260 68820
rect 54312 68808 54318 68860
rect 62810 68808 62816 68860
rect 62868 68848 62874 68860
rect 70078 68848 70084 68860
rect 62868 68820 70084 68848
rect 62868 68808 62874 68820
rect 70078 68808 70084 68820
rect 70136 68808 70142 68860
rect 82314 68808 82320 68860
rect 82372 68848 82378 68860
rect 85350 68848 85356 68860
rect 82372 68820 85356 68848
rect 82372 68808 82378 68820
rect 85350 68808 85356 68820
rect 85408 68808 85414 68860
rect 93446 68808 93452 68860
rect 93504 68848 93510 68860
rect 102830 68848 102836 68860
rect 93504 68820 102836 68848
rect 93504 68808 93510 68820
rect 102830 68808 102836 68820
rect 102888 68808 102894 68860
rect 122242 68808 122248 68860
rect 122300 68848 122306 68860
rect 125830 68848 125836 68860
rect 122300 68820 125836 68848
rect 122300 68808 122306 68820
rect 125830 68808 125836 68820
rect 125888 68808 125894 68860
rect 140826 68808 140832 68860
rect 140884 68848 140890 68860
rect 144322 68848 144328 68860
rect 140884 68820 144328 68848
rect 140884 68808 140890 68820
rect 144322 68808 144328 68820
rect 144380 68808 144386 68860
rect 160974 68808 160980 68860
rect 161032 68848 161038 68860
rect 168886 68848 168892 68860
rect 161032 68820 168892 68848
rect 161032 68808 161038 68820
rect 168886 68808 168892 68820
rect 168944 68808 168950 68860
rect 169898 68808 169904 68860
rect 169956 68848 169962 68860
rect 173946 68848 173952 68860
rect 169956 68820 173952 68848
rect 169956 68808 169962 68820
rect 173946 68808 173952 68820
rect 174004 68808 174010 68860
rect 193726 68808 193732 68860
rect 193784 68848 193790 68860
rect 196486 68848 196492 68860
rect 193784 68820 196492 68848
rect 193784 68808 193790 68820
rect 196486 68808 196492 68820
rect 196544 68808 196550 68860
rect 205134 68808 205140 68860
rect 205192 68848 205198 68860
rect 221234 68848 221240 68860
rect 205192 68820 221240 68848
rect 205192 68808 205198 68820
rect 221234 68808 221240 68820
rect 221292 68808 221298 68860
rect 27574 68740 27580 68792
rect 27632 68780 27638 68792
rect 49381 68783 49439 68789
rect 49381 68780 49393 68783
rect 27632 68752 49393 68780
rect 27632 68740 27638 68752
rect 49381 68749 49393 68752
rect 49427 68749 49439 68783
rect 49381 68743 49439 68749
rect 50206 68740 50212 68792
rect 50264 68780 50270 68792
rect 52966 68780 52972 68792
rect 50264 68752 52972 68780
rect 50264 68740 50270 68752
rect 52966 68740 52972 68752
rect 53024 68740 53030 68792
rect 121874 68740 121880 68792
rect 121932 68780 121938 68792
rect 125186 68780 125192 68792
rect 121932 68752 125192 68780
rect 121932 68740 121938 68752
rect 125186 68740 125192 68752
rect 125244 68740 125250 68792
rect 195290 68740 195296 68792
rect 195348 68780 195354 68792
rect 198786 68780 198792 68792
rect 195348 68752 198792 68780
rect 195348 68740 195354 68752
rect 198786 68740 198792 68752
rect 198844 68740 198850 68792
rect 36041 68715 36099 68721
rect 36041 68681 36053 68715
rect 36087 68712 36099 68715
rect 96761 68715 96819 68721
rect 36087 68684 45836 68712
rect 36087 68681 36099 68684
rect 36041 68675 36099 68681
rect 37878 68536 37884 68588
rect 37936 68576 37942 68588
rect 41466 68576 41472 68588
rect 37936 68548 41472 68576
rect 37936 68536 37942 68548
rect 41466 68536 41472 68548
rect 41524 68536 41530 68588
rect 45808 68576 45836 68684
rect 96761 68681 96773 68715
rect 96807 68681 96819 68715
rect 96761 68675 96819 68681
rect 96776 68644 96804 68675
rect 102278 68672 102284 68724
rect 102336 68712 102342 68724
rect 174314 68712 174320 68724
rect 102336 68684 174320 68712
rect 102336 68672 102342 68684
rect 174314 68672 174320 68684
rect 174372 68672 174378 68724
rect 99521 68647 99579 68653
rect 99521 68644 99533 68647
rect 96776 68616 99533 68644
rect 99521 68613 99533 68616
rect 99567 68613 99579 68647
rect 99521 68607 99579 68613
rect 101174 68604 101180 68656
rect 101232 68644 101238 68656
rect 173210 68644 173216 68656
rect 101232 68616 173216 68644
rect 101232 68604 101238 68616
rect 173210 68604 173216 68616
rect 173268 68604 173274 68656
rect 194646 68604 194652 68656
rect 194704 68644 194710 68656
rect 198234 68644 198240 68656
rect 194704 68616 198240 68644
rect 194704 68604 194710 68616
rect 198234 68604 198240 68616
rect 198292 68604 198298 68656
rect 57474 68576 57480 68588
rect 45808 68548 57480 68576
rect 57474 68536 57480 68548
rect 57532 68536 57538 68588
rect 120678 68536 120684 68588
rect 120736 68576 120742 68588
rect 123438 68576 123444 68588
rect 120736 68548 123444 68576
rect 120736 68536 120742 68548
rect 123438 68536 123444 68548
rect 123496 68536 123502 68588
rect 125002 68536 125008 68588
rect 125060 68576 125066 68588
rect 129326 68576 129332 68588
rect 125060 68548 129332 68576
rect 125060 68536 125066 68548
rect 129326 68536 129332 68548
rect 129384 68536 129390 68588
rect 191702 68536 191708 68588
rect 191760 68576 191766 68588
rect 193634 68576 193640 68588
rect 191760 68548 193640 68576
rect 191760 68536 191766 68548
rect 193634 68536 193640 68548
rect 193692 68536 193698 68588
rect 38614 68468 38620 68520
rect 38672 68508 38678 68520
rect 41834 68508 41840 68520
rect 38672 68480 41840 68508
rect 38672 68468 38678 68480
rect 41834 68468 41840 68480
rect 41892 68468 41898 68520
rect 99613 68511 99671 68517
rect 99613 68477 99625 68511
rect 99659 68508 99671 68511
rect 110009 68511 110067 68517
rect 110009 68508 110021 68511
rect 99659 68480 110021 68508
rect 99659 68477 99671 68480
rect 99613 68471 99671 68477
rect 110009 68477 110021 68480
rect 110055 68477 110067 68511
rect 110009 68471 110067 68477
rect 110558 68468 110564 68520
rect 110616 68508 110622 68520
rect 111478 68508 111484 68520
rect 110616 68480 111484 68508
rect 110616 68468 110622 68480
rect 111478 68468 111484 68480
rect 111536 68468 111542 68520
rect 116630 68468 116636 68520
rect 116688 68508 116694 68520
rect 117642 68508 117648 68520
rect 116688 68480 117648 68508
rect 116688 68468 116694 68480
rect 117642 68468 117648 68480
rect 117700 68468 117706 68520
rect 119482 68468 119488 68520
rect 119540 68508 119546 68520
rect 121690 68508 121696 68520
rect 119540 68480 121696 68508
rect 119540 68468 119546 68480
rect 121690 68468 121696 68480
rect 121748 68468 121754 68520
rect 123898 68468 123904 68520
rect 123956 68508 123962 68520
rect 128130 68508 128136 68520
rect 123956 68480 128136 68508
rect 123956 68468 123962 68480
rect 128130 68468 128136 68480
rect 128188 68468 128194 68520
rect 49838 68400 49844 68452
rect 49896 68440 49902 68452
rect 52230 68440 52236 68452
rect 49896 68412 52236 68440
rect 49896 68400 49902 68412
rect 52230 68400 52236 68412
rect 52288 68400 52294 68452
rect 74586 68400 74592 68452
rect 74644 68440 74650 68452
rect 75598 68440 75604 68452
rect 74644 68412 75604 68440
rect 74644 68400 74650 68412
rect 75598 68400 75604 68412
rect 75656 68400 75662 68452
rect 94550 68400 94556 68452
rect 94608 68440 94614 68452
rect 102738 68440 102744 68452
rect 94608 68412 102744 68440
rect 94608 68400 94614 68412
rect 102738 68400 102744 68412
rect 102796 68400 102802 68452
rect 110098 68400 110104 68452
rect 110156 68440 110162 68452
rect 111110 68440 111116 68452
rect 110156 68412 111116 68440
rect 110156 68400 110162 68412
rect 111110 68400 111116 68412
rect 111168 68400 111174 68452
rect 116262 68400 116268 68452
rect 116320 68440 116326 68452
rect 117090 68440 117096 68452
rect 116320 68412 117096 68440
rect 116320 68400 116326 68412
rect 117090 68400 117096 68412
rect 117148 68400 117154 68452
rect 182870 68400 182876 68452
rect 182928 68440 182934 68452
rect 183606 68440 183612 68452
rect 182928 68412 183612 68440
rect 182928 68400 182934 68412
rect 183606 68400 183612 68412
rect 183664 68400 183670 68452
rect 86730 68332 86736 68384
rect 86788 68372 86794 68384
rect 92802 68372 92808 68384
rect 86788 68344 92808 68372
rect 86788 68332 86794 68344
rect 92802 68332 92808 68344
rect 92860 68332 92866 68384
rect 97862 68332 97868 68384
rect 97920 68372 97926 68384
rect 102554 68372 102560 68384
rect 97920 68344 102560 68372
rect 97920 68332 97926 68344
rect 102554 68332 102560 68344
rect 102612 68332 102618 68384
rect 110193 68375 110251 68381
rect 110193 68341 110205 68375
rect 110239 68372 110251 68375
rect 116173 68375 116231 68381
rect 116173 68372 116185 68375
rect 110239 68344 116185 68372
rect 110239 68341 110251 68344
rect 110193 68335 110251 68341
rect 116173 68341 116185 68344
rect 116219 68341 116231 68375
rect 116173 68335 116231 68341
rect 119850 68332 119856 68384
rect 119908 68372 119914 68384
rect 122334 68372 122340 68384
rect 119908 68344 122340 68372
rect 119908 68332 119914 68344
rect 122334 68332 122340 68344
rect 122392 68332 122398 68384
rect 123346 68332 123352 68384
rect 123404 68372 123410 68384
rect 127302 68372 127308 68384
rect 123404 68344 127308 68372
rect 123404 68332 123410 68344
rect 127302 68332 127308 68344
rect 127360 68332 127366 68384
rect 155454 68332 155460 68384
rect 155512 68372 155518 68384
rect 159502 68372 159508 68384
rect 155512 68344 159508 68372
rect 155512 68332 155518 68344
rect 159502 68332 159508 68344
rect 159560 68332 159566 68384
rect 62994 68264 63000 68316
rect 63052 68304 63058 68316
rect 64558 68304 64564 68316
rect 63052 68276 64564 68304
rect 63052 68264 63058 68276
rect 64558 68264 64564 68276
rect 64616 68264 64622 68316
rect 70814 68304 70820 68316
rect 69084 68276 70820 68304
rect 62350 68196 62356 68248
rect 62408 68236 62414 68248
rect 63454 68236 63460 68248
rect 62408 68208 63460 68236
rect 62408 68196 62414 68208
rect 63454 68196 63460 68208
rect 63512 68196 63518 68248
rect 63362 68128 63368 68180
rect 63420 68168 63426 68180
rect 69084 68168 69112 68276
rect 70814 68264 70820 68276
rect 70872 68264 70878 68316
rect 70998 68264 71004 68316
rect 71056 68304 71062 68316
rect 73390 68304 73396 68316
rect 71056 68276 73396 68304
rect 71056 68264 71062 68276
rect 73390 68264 73396 68276
rect 73448 68264 73454 68316
rect 81210 68264 81216 68316
rect 81268 68304 81274 68316
rect 83510 68304 83516 68316
rect 81268 68276 83516 68304
rect 81268 68264 81274 68276
rect 83510 68264 83516 68276
rect 83568 68264 83574 68316
rect 85626 68264 85632 68316
rect 85684 68304 85690 68316
rect 90962 68304 90968 68316
rect 85684 68276 90968 68304
rect 85684 68264 85690 68276
rect 90962 68264 90968 68276
rect 91020 68264 91026 68316
rect 95654 68264 95660 68316
rect 95712 68304 95718 68316
rect 102646 68304 102652 68316
rect 95712 68276 102652 68304
rect 95712 68264 95718 68276
rect 102646 68264 102652 68276
rect 102704 68264 102710 68316
rect 121506 68264 121512 68316
rect 121564 68304 121570 68316
rect 124634 68304 124640 68316
rect 121564 68276 124640 68304
rect 121564 68264 121570 68276
rect 124634 68264 124640 68276
rect 124692 68264 124698 68316
rect 124729 68307 124787 68313
rect 124729 68273 124741 68307
rect 124775 68304 124787 68307
rect 132546 68304 132552 68316
rect 124775 68276 132552 68304
rect 124775 68273 124787 68276
rect 124729 68267 124787 68273
rect 132546 68264 132552 68276
rect 132604 68264 132610 68316
rect 144506 68264 144512 68316
rect 144564 68304 144570 68316
rect 146530 68304 146536 68316
rect 144564 68276 146536 68304
rect 144564 68264 144570 68276
rect 146530 68264 146536 68276
rect 146588 68264 146594 68316
rect 153246 68264 153252 68316
rect 153304 68304 153310 68316
rect 155822 68304 155828 68316
rect 153304 68276 155828 68304
rect 153304 68264 153310 68276
rect 155822 68264 155828 68276
rect 155880 68264 155886 68316
rect 156558 68264 156564 68316
rect 156616 68304 156622 68316
rect 161434 68304 161440 68316
rect 156616 68276 161440 68304
rect 156616 68264 156622 68276
rect 161434 68264 161440 68276
rect 161492 68264 161498 68316
rect 163274 68304 163280 68316
rect 161636 68276 163280 68304
rect 69158 68196 69164 68248
rect 69216 68236 69222 68248
rect 72286 68236 72292 68248
rect 69216 68208 72292 68236
rect 69216 68196 69222 68208
rect 72286 68196 72292 68208
rect 72344 68196 72350 68248
rect 72838 68196 72844 68248
rect 72896 68236 72902 68248
rect 74494 68236 74500 68248
rect 72896 68208 74500 68236
rect 72896 68196 72902 68208
rect 74494 68196 74500 68208
rect 74552 68196 74558 68248
rect 80106 68196 80112 68248
rect 80164 68236 80170 68248
rect 81670 68236 81676 68248
rect 80164 68208 81676 68236
rect 80164 68196 80170 68208
rect 81670 68196 81676 68208
rect 81728 68196 81734 68248
rect 84522 68196 84528 68248
rect 84580 68236 84586 68248
rect 89122 68236 89128 68248
rect 84580 68208 89128 68236
rect 84580 68196 84586 68208
rect 89122 68196 89128 68208
rect 89180 68196 89186 68248
rect 98966 68196 98972 68248
rect 99024 68236 99030 68248
rect 100346 68236 100352 68248
rect 99024 68208 100352 68236
rect 99024 68196 99030 68208
rect 100346 68196 100352 68208
rect 100404 68196 100410 68248
rect 121046 68196 121052 68248
rect 121104 68236 121110 68248
rect 124450 68236 124456 68248
rect 121104 68208 124456 68236
rect 121104 68196 121110 68208
rect 124450 68196 124456 68208
rect 124508 68196 124514 68248
rect 134478 68196 134484 68248
rect 134536 68236 134542 68248
rect 136594 68236 136600 68248
rect 134536 68208 136600 68236
rect 134536 68196 134542 68208
rect 136594 68196 136600 68208
rect 136652 68196 136658 68248
rect 142666 68196 142672 68248
rect 142724 68236 142730 68248
rect 145426 68236 145432 68248
rect 142724 68208 145432 68236
rect 142724 68196 142730 68208
rect 145426 68196 145432 68208
rect 145484 68196 145490 68248
rect 146438 68196 146444 68248
rect 146496 68236 146502 68248
rect 147634 68236 147640 68248
rect 146496 68208 147640 68236
rect 146496 68196 146502 68208
rect 147634 68196 147640 68208
rect 147692 68196 147698 68248
rect 152142 68196 152148 68248
rect 152200 68236 152206 68248
rect 153890 68236 153896 68248
rect 152200 68208 153896 68236
rect 152200 68196 152206 68208
rect 153890 68196 153896 68208
rect 153948 68196 153954 68248
rect 154350 68196 154356 68248
rect 154408 68236 154414 68248
rect 157662 68236 157668 68248
rect 154408 68208 157668 68236
rect 154408 68196 154414 68208
rect 157662 68196 157668 68208
rect 157720 68196 157726 68248
rect 157938 68196 157944 68248
rect 157996 68236 158002 68248
rect 161636 68236 161664 68276
rect 163274 68264 163280 68276
rect 163332 68264 163338 68316
rect 165482 68264 165488 68316
rect 165540 68304 165546 68316
rect 167138 68304 167144 68316
rect 165540 68276 167144 68304
rect 165540 68264 165546 68276
rect 167138 68264 167144 68276
rect 167196 68264 167202 68316
rect 167690 68264 167696 68316
rect 167748 68304 167754 68316
rect 169530 68304 169536 68316
rect 167748 68276 169536 68304
rect 167748 68264 167754 68276
rect 169530 68264 169536 68276
rect 169588 68264 169594 68316
rect 171002 68264 171008 68316
rect 171060 68304 171066 68316
rect 174038 68304 174044 68316
rect 171060 68276 174044 68304
rect 171060 68264 171066 68276
rect 174038 68264 174044 68276
rect 174096 68264 174102 68316
rect 157996 68208 161664 68236
rect 157996 68196 158002 68208
rect 164378 68196 164384 68248
rect 164436 68236 164442 68248
rect 169254 68236 169260 68248
rect 164436 68208 169260 68236
rect 164436 68196 164442 68208
rect 169254 68196 169260 68208
rect 169312 68196 169318 68248
rect 172106 68196 172112 68248
rect 172164 68236 172170 68248
rect 172164 68208 174084 68236
rect 172164 68196 172170 68208
rect 63420 68140 69112 68168
rect 63420 68128 63426 68140
rect 135306 68128 135312 68180
rect 135364 68168 135370 68180
rect 143218 68168 143224 68180
rect 135364 68140 143224 68168
rect 135364 68128 135370 68140
rect 143218 68128 143224 68140
rect 143276 68128 143282 68180
rect 174056 68168 174084 68208
rect 174682 68168 174688 68180
rect 174056 68140 174688 68168
rect 174682 68128 174688 68140
rect 174740 68128 174746 68180
rect 100070 68060 100076 68112
rect 100128 68100 100134 68112
rect 102462 68100 102468 68112
rect 100128 68072 102468 68100
rect 100128 68060 100134 68072
rect 102462 68060 102468 68072
rect 102520 68060 102526 68112
rect 116173 68103 116231 68109
rect 116173 68069 116185 68103
rect 116219 68100 116231 68103
rect 124729 68103 124787 68109
rect 124729 68100 124741 68103
rect 116219 68072 124741 68100
rect 116219 68069 116231 68072
rect 116173 68063 116231 68069
rect 124729 68069 124741 68072
rect 124775 68069 124787 68103
rect 124729 68063 124787 68069
rect 135030 68060 135036 68112
rect 135088 68100 135094 68112
rect 142114 68100 142120 68112
rect 135088 68072 142120 68100
rect 135088 68060 135094 68072
rect 142114 68060 142120 68072
rect 142172 68060 142178 68112
rect 100346 67516 100352 67568
rect 100404 67556 100410 67568
rect 102370 67556 102376 67568
rect 100404 67528 102376 67556
rect 100404 67516 100410 67528
rect 102370 67516 102376 67528
rect 102428 67516 102434 67568
rect 134662 66700 134668 66752
rect 134720 66740 134726 66752
rect 139538 66740 139544 66752
rect 134720 66712 139544 66740
rect 134720 66700 134726 66712
rect 139538 66700 139544 66712
rect 139596 66700 139602 66752
rect 135306 66428 135312 66480
rect 135364 66468 135370 66480
rect 141010 66468 141016 66480
rect 135364 66440 141016 66468
rect 135364 66428 135370 66440
rect 141010 66428 141016 66440
rect 141068 66428 141074 66480
rect 96758 65952 96764 66004
rect 96816 65992 96822 66004
rect 102370 65992 102376 66004
rect 96816 65964 102376 65992
rect 96816 65952 96822 65964
rect 102370 65952 102376 65964
rect 102428 65952 102434 66004
rect 63270 65544 63276 65596
rect 63328 65584 63334 65596
rect 66398 65584 66404 65596
rect 63328 65556 66404 65584
rect 63328 65544 63334 65556
rect 66398 65544 66404 65556
rect 66456 65544 66462 65596
rect 166586 65544 166592 65596
rect 166644 65544 166650 65596
rect 167138 65544 167144 65596
rect 167196 65544 167202 65596
rect 100898 65408 100904 65460
rect 100956 65448 100962 65460
rect 102554 65448 102560 65460
rect 100956 65420 102560 65448
rect 100956 65408 100962 65420
rect 102554 65408 102560 65420
rect 102612 65408 102618 65460
rect 134662 65408 134668 65460
rect 134720 65448 134726 65460
rect 136870 65448 136876 65460
rect 134720 65420 136876 65448
rect 134720 65408 134726 65420
rect 136870 65408 136876 65420
rect 136928 65408 136934 65460
rect 62810 65340 62816 65392
rect 62868 65380 62874 65392
rect 66306 65380 66312 65392
rect 62868 65352 66312 65380
rect 62868 65340 62874 65352
rect 66306 65340 66312 65352
rect 66364 65340 66370 65392
rect 135030 65340 135036 65392
rect 135088 65380 135094 65392
rect 137698 65380 137704 65392
rect 135088 65352 137704 65380
rect 135088 65340 135094 65352
rect 137698 65340 137704 65352
rect 137756 65340 137762 65392
rect 62718 65272 62724 65324
rect 62776 65312 62782 65324
rect 65662 65312 65668 65324
rect 62776 65284 65668 65312
rect 62776 65272 62782 65284
rect 65662 65272 65668 65284
rect 65720 65272 65726 65324
rect 166604 65312 166632 65544
rect 167156 65380 167184 65544
rect 174222 65380 174228 65392
rect 167156 65352 174228 65380
rect 174222 65340 174228 65352
rect 174280 65340 174286 65392
rect 174130 65312 174136 65324
rect 166604 65284 174136 65312
rect 174130 65272 174136 65284
rect 174188 65272 174194 65324
rect 135306 65204 135312 65256
rect 135364 65244 135370 65256
rect 138158 65244 138164 65256
rect 135364 65216 138164 65244
rect 135364 65204 135370 65216
rect 138158 65204 138164 65216
rect 138216 65204 138222 65256
rect 63546 64320 63552 64372
rect 63604 64360 63610 64372
rect 66398 64360 66404 64372
rect 63604 64332 66404 64360
rect 63604 64320 63610 64332
rect 66398 64320 66404 64332
rect 66456 64320 66462 64372
rect 100622 64320 100628 64372
rect 100680 64360 100686 64372
rect 102462 64360 102468 64372
rect 100680 64332 102468 64360
rect 100680 64320 100686 64332
rect 102462 64320 102468 64332
rect 102520 64320 102526 64372
rect 63454 64184 63460 64236
rect 63512 64224 63518 64236
rect 66398 64224 66404 64236
rect 63512 64196 66404 64224
rect 63512 64184 63518 64196
rect 66398 64184 66404 64196
rect 66456 64184 66462 64236
rect 135398 64116 135404 64168
rect 135456 64156 135462 64168
rect 136962 64156 136968 64168
rect 135456 64128 136968 64156
rect 135456 64116 135462 64128
rect 136962 64116 136968 64128
rect 137020 64116 137026 64168
rect 100898 64048 100904 64100
rect 100956 64088 100962 64100
rect 102646 64088 102652 64100
rect 100956 64060 102652 64088
rect 100956 64048 100962 64060
rect 102646 64048 102652 64060
rect 102704 64048 102710 64100
rect 135030 64048 135036 64100
rect 135088 64088 135094 64100
rect 136870 64088 136876 64100
rect 135088 64060 136876 64088
rect 135088 64048 135094 64060
rect 136870 64048 136876 64060
rect 136928 64048 136934 64100
rect 169254 63980 169260 64032
rect 169312 64020 169318 64032
rect 174130 64020 174136 64032
rect 169312 63992 174136 64020
rect 169312 63980 169318 63992
rect 174130 63980 174136 63992
rect 174188 63980 174194 64032
rect 97034 63776 97040 63828
rect 97092 63816 97098 63828
rect 102370 63816 102376 63828
rect 97092 63788 102376 63816
rect 97092 63776 97098 63788
rect 102370 63776 102376 63788
rect 102428 63776 102434 63828
rect 171830 63708 171836 63760
rect 171888 63748 171894 63760
rect 174222 63748 174228 63760
rect 171888 63720 174228 63748
rect 171888 63708 171894 63720
rect 174222 63708 174228 63720
rect 174280 63708 174286 63760
rect 172014 63232 172020 63284
rect 172072 63272 172078 63284
rect 173854 63272 173860 63284
rect 172072 63244 173860 63272
rect 172072 63232 172078 63244
rect 173854 63232 173860 63244
rect 173912 63232 173918 63284
rect 62810 62960 62816 63012
rect 62868 63000 62874 63012
rect 66398 63000 66404 63012
rect 62868 62972 66404 63000
rect 62868 62960 62874 62972
rect 66398 62960 66404 62972
rect 66456 62960 66462 63012
rect 100438 62960 100444 63012
rect 100496 63000 100502 63012
rect 102370 63000 102376 63012
rect 100496 62972 102376 63000
rect 100496 62960 100502 62972
rect 102370 62960 102376 62972
rect 102428 62960 102434 63012
rect 63178 62688 63184 62740
rect 63236 62728 63242 62740
rect 66306 62728 66312 62740
rect 63236 62700 66312 62728
rect 63236 62688 63242 62700
rect 66306 62688 66312 62700
rect 66364 62688 66370 62740
rect 100898 62688 100904 62740
rect 100956 62728 100962 62740
rect 102554 62728 102560 62740
rect 100956 62700 102560 62728
rect 100956 62688 100962 62700
rect 102554 62688 102560 62700
rect 102612 62688 102618 62740
rect 134478 62688 134484 62740
rect 134536 62728 134542 62740
rect 136962 62728 136968 62740
rect 134536 62700 136968 62728
rect 134536 62688 134542 62700
rect 136962 62688 136968 62700
rect 137020 62688 137026 62740
rect 13314 62620 13320 62672
rect 13372 62660 13378 62672
rect 29230 62660 29236 62672
rect 13372 62632 29236 62660
rect 13372 62620 13378 62632
rect 29230 62620 29236 62632
rect 29288 62620 29294 62672
rect 135306 62620 135312 62672
rect 135364 62660 135370 62672
rect 136870 62660 136876 62672
rect 135364 62632 136876 62660
rect 135364 62620 135370 62632
rect 136870 62620 136876 62632
rect 136928 62620 136934 62672
rect 171646 62552 171652 62604
rect 171704 62592 171710 62604
rect 174314 62592 174320 62604
rect 171704 62564 174320 62592
rect 171704 62552 171710 62564
rect 174314 62552 174320 62564
rect 174372 62552 174378 62604
rect 171738 62484 171744 62536
rect 171796 62524 171802 62536
rect 174130 62524 174136 62536
rect 171796 62496 174136 62524
rect 171796 62484 171802 62496
rect 174130 62484 174136 62496
rect 174188 62484 174194 62536
rect 171646 62008 171652 62060
rect 171704 62048 171710 62060
rect 174038 62048 174044 62060
rect 171704 62020 174044 62048
rect 171704 62008 171710 62020
rect 174038 62008 174044 62020
rect 174096 62008 174102 62060
rect 62718 61736 62724 61788
rect 62776 61776 62782 61788
rect 66398 61776 66404 61788
rect 62776 61748 66404 61776
rect 62776 61736 62782 61748
rect 66398 61736 66404 61748
rect 66456 61736 66462 61788
rect 63730 61464 63736 61516
rect 63788 61504 63794 61516
rect 66306 61504 66312 61516
rect 63788 61476 66312 61504
rect 63788 61464 63794 61476
rect 66306 61464 66312 61476
rect 66364 61464 66370 61516
rect 100898 61328 100904 61380
rect 100956 61368 100962 61380
rect 102738 61368 102744 61380
rect 100956 61340 102744 61368
rect 100956 61328 100962 61340
rect 102738 61328 102744 61340
rect 102796 61328 102802 61380
rect 172658 61328 172664 61380
rect 172716 61368 172722 61380
rect 173946 61368 173952 61380
rect 172716 61340 173952 61368
rect 172716 61328 172722 61340
rect 173946 61328 173952 61340
rect 174004 61328 174010 61380
rect 100254 61260 100260 61312
rect 100312 61300 100318 61312
rect 102462 61300 102468 61312
rect 100312 61272 102468 61300
rect 100312 61260 100318 61272
rect 102462 61260 102468 61272
rect 102520 61260 102526 61312
rect 135214 61260 135220 61312
rect 135272 61300 135278 61312
rect 136870 61300 136876 61312
rect 135272 61272 136876 61300
rect 135272 61260 135278 61272
rect 136870 61260 136876 61272
rect 136928 61260 136934 61312
rect 172750 61192 172756 61244
rect 172808 61232 172814 61244
rect 174130 61232 174136 61244
rect 172808 61204 174136 61232
rect 172808 61192 172814 61204
rect 174130 61192 174136 61204
rect 174188 61192 174194 61244
rect 134846 60920 134852 60972
rect 134904 60960 134910 60972
rect 136778 60960 136784 60972
rect 134904 60932 136784 60960
rect 134904 60920 134910 60932
rect 136778 60920 136784 60932
rect 136836 60920 136842 60972
rect 100622 60308 100628 60360
rect 100680 60348 100686 60360
rect 102646 60348 102652 60360
rect 100680 60320 102652 60348
rect 100680 60308 100686 60320
rect 102646 60308 102652 60320
rect 102704 60308 102710 60360
rect 100898 60172 100904 60224
rect 100956 60212 100962 60224
rect 102370 60212 102376 60224
rect 100956 60184 102376 60212
rect 100956 60172 100962 60184
rect 102370 60172 102376 60184
rect 102428 60172 102434 60224
rect 62626 60104 62632 60156
rect 62684 60144 62690 60156
rect 66398 60144 66404 60156
rect 62684 60116 66404 60144
rect 62684 60104 62690 60116
rect 66398 60104 66404 60116
rect 66456 60104 66462 60156
rect 134478 60036 134484 60088
rect 134536 60076 134542 60088
rect 136962 60076 136968 60088
rect 134536 60048 136968 60076
rect 134536 60036 134542 60048
rect 136962 60036 136968 60048
rect 137020 60036 137026 60088
rect 62810 59968 62816 60020
rect 62868 60008 62874 60020
rect 66306 60008 66312 60020
rect 62868 59980 66312 60008
rect 62868 59968 62874 59980
rect 66306 59968 66312 59980
rect 66364 59968 66370 60020
rect 99702 59968 99708 60020
rect 99760 60008 99766 60020
rect 102554 60008 102560 60020
rect 99760 59980 102560 60008
rect 99760 59968 99766 59980
rect 102554 59968 102560 59980
rect 102612 59968 102618 60020
rect 172658 59968 172664 60020
rect 172716 60008 172722 60020
rect 173762 60008 173768 60020
rect 172716 59980 173768 60008
rect 172716 59968 172722 59980
rect 173762 59968 173768 59980
rect 173820 59968 173826 60020
rect 63730 59900 63736 59952
rect 63788 59940 63794 59952
rect 66214 59940 66220 59952
rect 63788 59912 66220 59940
rect 63788 59900 63794 59912
rect 66214 59900 66220 59912
rect 66272 59900 66278 59952
rect 135398 59900 135404 59952
rect 135456 59940 135462 59952
rect 136870 59940 136876 59952
rect 135456 59912 136876 59940
rect 135456 59900 135462 59912
rect 136870 59900 136876 59912
rect 136928 59900 136934 59952
rect 172198 59900 172204 59952
rect 172256 59940 172262 59952
rect 174038 59940 174044 59952
rect 172256 59912 174044 59940
rect 172256 59900 172262 59912
rect 174038 59900 174044 59912
rect 174096 59900 174102 59952
rect 134386 59832 134392 59884
rect 134444 59872 134450 59884
rect 136778 59872 136784 59884
rect 134444 59844 136784 59872
rect 134444 59832 134450 59844
rect 136778 59832 136784 59844
rect 136836 59832 136842 59884
rect 172658 58812 172664 58864
rect 172716 58852 172722 58864
rect 174038 58852 174044 58864
rect 172716 58824 174044 58852
rect 172716 58812 172722 58824
rect 174038 58812 174044 58824
rect 174096 58812 174102 58864
rect 100622 58744 100628 58796
rect 100680 58784 100686 58796
rect 102462 58784 102468 58796
rect 100680 58756 102468 58784
rect 100680 58744 100686 58756
rect 102462 58744 102468 58756
rect 102520 58744 102526 58796
rect 62902 58608 62908 58660
rect 62960 58648 62966 58660
rect 66398 58648 66404 58660
rect 62960 58620 66404 58648
rect 62960 58608 62966 58620
rect 66398 58608 66404 58620
rect 66456 58608 66462 58660
rect 100622 58608 100628 58660
rect 100680 58648 100686 58660
rect 102646 58648 102652 58660
rect 100680 58620 102652 58648
rect 100680 58608 100686 58620
rect 102646 58608 102652 58620
rect 102704 58608 102710 58660
rect 172658 58608 172664 58660
rect 172716 58648 172722 58660
rect 173854 58648 173860 58660
rect 172716 58620 173860 58648
rect 172716 58608 172722 58620
rect 173854 58608 173860 58620
rect 173912 58608 173918 58660
rect 63546 58540 63552 58592
rect 63604 58580 63610 58592
rect 66306 58580 66312 58592
rect 63604 58552 66312 58580
rect 63604 58540 63610 58552
rect 66306 58540 66312 58552
rect 66364 58540 66370 58592
rect 135214 58540 135220 58592
rect 135272 58580 135278 58592
rect 136870 58580 136876 58592
rect 135272 58552 136876 58580
rect 135272 58540 135278 58552
rect 136870 58540 136876 58552
rect 136928 58540 136934 58592
rect 172750 58472 172756 58524
rect 172808 58512 172814 58524
rect 174130 58512 174136 58524
rect 172808 58484 174136 58512
rect 172808 58472 172814 58484
rect 174130 58472 174136 58484
rect 174188 58472 174194 58524
rect 135030 58404 135036 58456
rect 135088 58444 135094 58456
rect 136778 58444 136784 58456
rect 135088 58416 136784 58444
rect 135088 58404 135094 58416
rect 136778 58404 136784 58416
rect 136836 58404 136842 58456
rect 62810 57384 62816 57436
rect 62868 57424 62874 57436
rect 66398 57424 66404 57436
rect 62868 57396 66404 57424
rect 62868 57384 62874 57396
rect 66398 57384 66404 57396
rect 66456 57384 66462 57436
rect 100622 57384 100628 57436
rect 100680 57424 100686 57436
rect 102370 57424 102376 57436
rect 100680 57396 102376 57424
rect 100680 57384 100686 57396
rect 102370 57384 102376 57396
rect 102428 57384 102434 57436
rect 172658 57248 172664 57300
rect 172716 57288 172722 57300
rect 173946 57288 173952 57300
rect 172716 57260 173952 57288
rect 172716 57248 172722 57260
rect 173946 57248 173952 57260
rect 174004 57248 174010 57300
rect 100622 57180 100628 57232
rect 100680 57220 100686 57232
rect 102462 57220 102468 57232
rect 100680 57192 102468 57220
rect 100680 57180 100686 57192
rect 102462 57180 102468 57192
rect 102520 57180 102526 57232
rect 135398 57180 135404 57232
rect 135456 57220 135462 57232
rect 136962 57220 136968 57232
rect 135456 57192 136968 57220
rect 135456 57180 135462 57192
rect 136962 57180 136968 57192
rect 137020 57180 137026 57232
rect 172566 57180 172572 57232
rect 172624 57220 172630 57232
rect 173762 57220 173768 57232
rect 172624 57192 173768 57220
rect 172624 57180 172630 57192
rect 173762 57180 173768 57192
rect 173820 57180 173826 57232
rect 62718 57112 62724 57164
rect 62776 57152 62782 57164
rect 66398 57152 66404 57164
rect 62776 57124 66404 57152
rect 62776 57112 62782 57124
rect 66398 57112 66404 57124
rect 66456 57112 66462 57164
rect 100530 57112 100536 57164
rect 100588 57152 100594 57164
rect 102554 57152 102560 57164
rect 100588 57124 102560 57152
rect 100588 57112 100594 57124
rect 102554 57112 102560 57124
rect 102612 57112 102618 57164
rect 135306 57112 135312 57164
rect 135364 57152 135370 57164
rect 136870 57152 136876 57164
rect 135364 57124 136876 57152
rect 135364 57112 135370 57124
rect 136870 57112 136876 57124
rect 136928 57112 136934 57164
rect 172106 57112 172112 57164
rect 172164 57152 172170 57164
rect 174038 57152 174044 57164
rect 172164 57124 174044 57152
rect 172164 57112 172170 57124
rect 174038 57112 174044 57124
rect 174096 57112 174102 57164
rect 134570 57044 134576 57096
rect 134628 57084 134634 57096
rect 136778 57084 136784 57096
rect 134628 57056 136784 57084
rect 134628 57044 134634 57056
rect 136778 57044 136784 57056
rect 136836 57044 136842 57096
rect 62626 56976 62632 57028
rect 62684 57016 62690 57028
rect 65018 57016 65024 57028
rect 62684 56988 65024 57016
rect 62684 56976 62690 56988
rect 65018 56976 65024 56988
rect 65076 56976 65082 57028
rect 172658 56024 172664 56076
rect 172716 56064 172722 56076
rect 174038 56064 174044 56076
rect 172716 56036 174044 56064
rect 172716 56024 172722 56036
rect 174038 56024 174044 56036
rect 174096 56024 174102 56076
rect 63270 55888 63276 55940
rect 63328 55928 63334 55940
rect 66398 55928 66404 55940
rect 63328 55900 66404 55928
rect 63328 55888 63334 55900
rect 66398 55888 66404 55900
rect 66456 55888 66462 55940
rect 100622 55888 100628 55940
rect 100680 55928 100686 55940
rect 102370 55928 102376 55940
rect 100680 55900 102376 55928
rect 100680 55888 100686 55900
rect 102370 55888 102376 55900
rect 102428 55888 102434 55940
rect 63546 55752 63552 55804
rect 63604 55792 63610 55804
rect 66306 55792 66312 55804
rect 63604 55764 66312 55792
rect 63604 55752 63610 55764
rect 66306 55752 66312 55764
rect 66364 55752 66370 55804
rect 100898 55752 100904 55804
rect 100956 55792 100962 55804
rect 102646 55792 102652 55804
rect 100956 55764 102652 55792
rect 100956 55752 100962 55764
rect 102646 55752 102652 55764
rect 102704 55752 102710 55804
rect 134294 55752 134300 55804
rect 134352 55792 134358 55804
rect 136870 55792 136876 55804
rect 134352 55764 136876 55792
rect 134352 55752 134358 55764
rect 136870 55752 136876 55764
rect 136928 55752 136934 55804
rect 135030 55412 135036 55464
rect 135088 55452 135094 55464
rect 136778 55452 136784 55464
rect 135088 55424 136784 55452
rect 135088 55412 135094 55424
rect 136778 55412 136784 55424
rect 136836 55412 136842 55464
rect 100622 54800 100628 54852
rect 100680 54840 100686 54852
rect 102462 54840 102468 54852
rect 100680 54812 102468 54840
rect 100680 54800 100686 54812
rect 102462 54800 102468 54812
rect 102520 54800 102526 54852
rect 63362 54664 63368 54716
rect 63420 54704 63426 54716
rect 66398 54704 66404 54716
rect 63420 54676 66404 54704
rect 63420 54664 63426 54676
rect 66398 54664 66404 54676
rect 66456 54664 66462 54716
rect 100806 54528 100812 54580
rect 100864 54568 100870 54580
rect 102554 54568 102560 54580
rect 100864 54540 102560 54568
rect 100864 54528 100870 54540
rect 102554 54528 102560 54540
rect 102612 54528 102618 54580
rect 134202 54528 134208 54580
rect 134260 54568 134266 54580
rect 137146 54568 137152 54580
rect 134260 54540 137152 54568
rect 134260 54528 134266 54540
rect 137146 54528 137152 54540
rect 137204 54528 137210 54580
rect 63454 54392 63460 54444
rect 63512 54432 63518 54444
rect 66306 54432 66312 54444
rect 63512 54404 66312 54432
rect 63512 54392 63518 54404
rect 66306 54392 66312 54404
rect 66364 54392 66370 54444
rect 171738 54392 171744 54444
rect 171796 54432 171802 54444
rect 171796 54404 172796 54432
rect 171796 54392 171802 54404
rect 172768 54364 172796 54404
rect 174222 54364 174228 54376
rect 172768 54336 174228 54364
rect 174222 54324 174228 54336
rect 174280 54324 174286 54376
rect 172934 54052 172940 54104
rect 172992 54092 172998 54104
rect 174130 54092 174136 54104
rect 172992 54064 174136 54092
rect 172992 54052 172998 54064
rect 174130 54052 174136 54064
rect 174188 54052 174194 54104
rect 135122 53916 135128 53968
rect 135180 53956 135186 53968
rect 136778 53956 136784 53968
rect 135180 53928 136784 53956
rect 135180 53916 135186 53928
rect 136778 53916 136784 53928
rect 136836 53916 136842 53968
rect 62810 53304 62816 53356
rect 62868 53344 62874 53356
rect 66398 53344 66404 53356
rect 62868 53316 66404 53344
rect 62868 53304 62874 53316
rect 66398 53304 66404 53316
rect 66456 53304 66462 53356
rect 100622 53236 100628 53288
rect 100680 53276 100686 53288
rect 102738 53276 102744 53288
rect 100680 53248 102744 53276
rect 100680 53236 100686 53248
rect 102738 53236 102744 53248
rect 102796 53236 102802 53288
rect 172566 53168 172572 53220
rect 172624 53208 172630 53220
rect 174038 53208 174044 53220
rect 172624 53180 174044 53208
rect 172624 53168 172630 53180
rect 174038 53168 174044 53180
rect 174096 53168 174102 53220
rect 100622 53032 100628 53084
rect 100680 53072 100686 53084
rect 102370 53072 102376 53084
rect 100680 53044 102376 53072
rect 100680 53032 100686 53044
rect 102370 53032 102376 53044
rect 102428 53032 102434 53084
rect 172658 53032 172664 53084
rect 172716 53072 172722 53084
rect 173854 53072 173860 53084
rect 172716 53044 173860 53072
rect 172716 53032 172722 53044
rect 173854 53032 173860 53044
rect 173912 53032 173918 53084
rect 63730 52964 63736 53016
rect 63788 53004 63794 53016
rect 66306 53004 66312 53016
rect 63788 52976 66312 53004
rect 63788 52964 63794 52976
rect 66306 52964 66312 52976
rect 66364 52964 66370 53016
rect 135398 52964 135404 53016
rect 135456 53004 135462 53016
rect 136870 53004 136876 53016
rect 135456 52976 136876 53004
rect 135456 52964 135462 52976
rect 136870 52964 136876 52976
rect 136928 52964 136934 53016
rect 172842 52896 172848 52948
rect 172900 52936 172906 52948
rect 174130 52936 174136 52948
rect 172900 52908 174136 52936
rect 172900 52896 172906 52908
rect 174130 52896 174136 52908
rect 174188 52896 174194 52948
rect 135030 52828 135036 52880
rect 135088 52868 135094 52880
rect 136778 52868 136784 52880
rect 135088 52840 136784 52868
rect 135088 52828 135094 52840
rect 136778 52828 136784 52840
rect 136836 52828 136842 52880
rect 100622 52216 100628 52268
rect 100680 52256 100686 52268
rect 102646 52256 102652 52268
rect 100680 52228 102652 52256
rect 100680 52216 100686 52228
rect 102646 52216 102652 52228
rect 102704 52216 102710 52268
rect 62902 52080 62908 52132
rect 62960 52120 62966 52132
rect 66398 52120 66404 52132
rect 62960 52092 66404 52120
rect 62960 52080 62966 52092
rect 66398 52080 66404 52092
rect 66456 52080 66462 52132
rect 172658 51808 172664 51860
rect 172716 51848 172722 51860
rect 173946 51848 173952 51860
rect 172716 51820 173952 51848
rect 172716 51808 172722 51820
rect 173946 51808 173952 51820
rect 174004 51808 174010 51860
rect 62718 51672 62724 51724
rect 62776 51712 62782 51724
rect 66398 51712 66404 51724
rect 62776 51684 66404 51712
rect 62776 51672 62782 51684
rect 66398 51672 66404 51684
rect 66456 51672 66462 51724
rect 100622 51672 100628 51724
rect 100680 51712 100686 51724
rect 102462 51712 102468 51724
rect 100680 51684 102468 51712
rect 100680 51672 100686 51684
rect 102462 51672 102468 51684
rect 102520 51672 102526 51724
rect 172658 51672 172664 51724
rect 172716 51712 172722 51724
rect 173762 51712 173768 51724
rect 172716 51684 173768 51712
rect 172716 51672 172722 51684
rect 173762 51672 173768 51684
rect 173820 51672 173826 51724
rect 63730 51604 63736 51656
rect 63788 51644 63794 51656
rect 65662 51644 65668 51656
rect 63788 51616 65668 51644
rect 63788 51604 63794 51616
rect 65662 51604 65668 51616
rect 65720 51604 65726 51656
rect 100530 51604 100536 51656
rect 100588 51644 100594 51656
rect 102554 51644 102560 51656
rect 100588 51616 102560 51644
rect 100588 51604 100594 51616
rect 102554 51604 102560 51616
rect 102612 51604 102618 51656
rect 135306 51604 135312 51656
rect 135364 51644 135370 51656
rect 136870 51644 136876 51656
rect 135364 51616 136876 51644
rect 135364 51604 135370 51616
rect 136870 51604 136876 51616
rect 136928 51604 136934 51656
rect 172014 51604 172020 51656
rect 172072 51644 172078 51656
rect 174038 51644 174044 51656
rect 172072 51616 174044 51644
rect 172072 51604 172078 51616
rect 174038 51604 174044 51616
rect 174096 51604 174102 51656
rect 135030 51332 135036 51384
rect 135088 51372 135094 51384
rect 136778 51372 136784 51384
rect 135088 51344 136784 51372
rect 135088 51332 135094 51344
rect 136778 51332 136784 51344
rect 136836 51332 136842 51384
rect 135398 51060 135404 51112
rect 135456 51100 135462 51112
rect 136686 51100 136692 51112
rect 135456 51072 136692 51100
rect 135456 51060 135462 51072
rect 136686 51060 136692 51072
rect 136744 51060 136750 51112
rect 63822 50584 63828 50636
rect 63880 50624 63886 50636
rect 66398 50624 66404 50636
rect 63880 50596 66404 50624
rect 63880 50584 63886 50596
rect 66398 50584 66404 50596
rect 66456 50584 66462 50636
rect 171646 50584 171652 50636
rect 171704 50624 171710 50636
rect 174038 50624 174044 50636
rect 171704 50596 174044 50624
rect 171704 50584 171710 50596
rect 174038 50584 174044 50596
rect 174096 50584 174102 50636
rect 62810 50448 62816 50500
rect 62868 50488 62874 50500
rect 66398 50488 66404 50500
rect 62868 50460 66404 50488
rect 62868 50448 62874 50460
rect 66398 50448 66404 50460
rect 66456 50448 66462 50500
rect 100622 50448 100628 50500
rect 100680 50488 100686 50500
rect 102646 50488 102652 50500
rect 100680 50460 102652 50488
rect 100680 50448 100686 50460
rect 102646 50448 102652 50460
rect 102704 50448 102710 50500
rect 100622 50312 100628 50364
rect 100680 50352 100686 50364
rect 102370 50352 102376 50364
rect 100680 50324 102376 50352
rect 100680 50312 100686 50324
rect 102370 50312 102376 50324
rect 102428 50312 102434 50364
rect 135398 50244 135404 50296
rect 135456 50284 135462 50296
rect 136870 50284 136876 50296
rect 135456 50256 136876 50284
rect 135456 50244 135462 50256
rect 136870 50244 136876 50256
rect 136928 50244 136934 50296
rect 134846 50176 134852 50228
rect 134904 50216 134910 50228
rect 136778 50216 136784 50228
rect 134904 50188 136784 50216
rect 134904 50176 134910 50188
rect 136778 50176 136784 50188
rect 136836 50176 136842 50228
rect 100622 49224 100628 49276
rect 100680 49264 100686 49276
rect 102462 49264 102468 49276
rect 100680 49236 102468 49264
rect 100680 49224 100686 49236
rect 102462 49224 102468 49236
rect 102520 49224 102526 49276
rect 63730 48952 63736 49004
rect 63788 48992 63794 49004
rect 65478 48992 65484 49004
rect 63788 48964 65484 48992
rect 63788 48952 63794 48964
rect 65478 48952 65484 48964
rect 65536 48952 65542 49004
rect 100622 48952 100628 49004
rect 100680 48992 100686 49004
rect 102554 48992 102560 49004
rect 100680 48964 102560 48992
rect 100680 48952 100686 48964
rect 102554 48952 102560 48964
rect 102612 48952 102618 49004
rect 172658 48952 172664 49004
rect 172716 48992 172722 49004
rect 173946 48992 173952 49004
rect 172716 48964 173952 48992
rect 172716 48952 172722 48964
rect 173946 48952 173952 48964
rect 174004 48952 174010 49004
rect 62902 48884 62908 48936
rect 62960 48924 62966 48936
rect 66398 48924 66404 48936
rect 62960 48896 66404 48924
rect 62960 48884 62966 48896
rect 66398 48884 66404 48896
rect 66456 48884 66462 48936
rect 136870 48924 136876 48936
rect 135508 48896 136876 48924
rect 135306 48816 135312 48868
rect 135364 48856 135370 48868
rect 135508 48856 135536 48896
rect 136870 48884 136876 48896
rect 136928 48884 136934 48936
rect 171830 48884 171836 48936
rect 171888 48924 171894 48936
rect 174038 48924 174044 48936
rect 171888 48896 174044 48924
rect 171888 48884 171894 48896
rect 174038 48884 174044 48896
rect 174096 48884 174102 48936
rect 135364 48828 135536 48856
rect 135364 48816 135370 48828
rect 172750 48816 172756 48868
rect 172808 48856 172814 48868
rect 174130 48856 174136 48868
rect 172808 48828 174136 48856
rect 172808 48816 172814 48828
rect 174130 48816 174136 48828
rect 174188 48816 174194 48868
rect 134754 48408 134760 48460
rect 134812 48448 134818 48460
rect 136778 48448 136784 48460
rect 134812 48420 136784 48448
rect 134812 48408 134818 48420
rect 136778 48408 136784 48420
rect 136836 48408 136842 48460
rect 100622 47864 100628 47916
rect 100680 47904 100686 47916
rect 102646 47904 102652 47916
rect 100680 47876 102652 47904
rect 100680 47864 100686 47876
rect 102646 47864 102652 47876
rect 102704 47864 102710 47916
rect 100622 47592 100628 47644
rect 100680 47632 100686 47644
rect 102370 47632 102376 47644
rect 100680 47604 102376 47632
rect 100680 47592 100686 47604
rect 102370 47592 102376 47604
rect 102428 47592 102434 47644
rect 172106 47592 172112 47644
rect 172164 47632 172170 47644
rect 174038 47632 174044 47644
rect 172164 47604 174044 47632
rect 172164 47592 172170 47604
rect 174038 47592 174044 47604
rect 174096 47592 174102 47644
rect 172566 47524 172572 47576
rect 172624 47564 172630 47576
rect 173854 47564 173860 47576
rect 172624 47536 173860 47564
rect 172624 47524 172630 47536
rect 173854 47524 173860 47536
rect 173912 47524 173918 47576
rect 62810 47456 62816 47508
rect 62868 47496 62874 47508
rect 66398 47496 66404 47508
rect 62868 47468 66404 47496
rect 62868 47456 62874 47468
rect 66398 47456 66404 47468
rect 66456 47456 66462 47508
rect 100622 47456 100628 47508
rect 100680 47496 100686 47508
rect 102462 47496 102468 47508
rect 100680 47468 102468 47496
rect 100680 47456 100686 47468
rect 102462 47456 102468 47468
rect 102520 47456 102526 47508
rect 135398 47456 135404 47508
rect 135456 47496 135462 47508
rect 136870 47496 136876 47508
rect 135456 47468 136876 47496
rect 135456 47456 135462 47468
rect 136870 47456 136876 47468
rect 136928 47456 136934 47508
rect 172658 47456 172664 47508
rect 172716 47496 172722 47508
rect 172716 47468 172796 47496
rect 172716 47456 172722 47468
rect 172768 47428 172796 47468
rect 174222 47428 174228 47440
rect 172768 47400 174228 47428
rect 174222 47388 174228 47400
rect 174280 47388 174286 47440
rect 134846 47320 134852 47372
rect 134904 47360 134910 47372
rect 136778 47360 136784 47372
rect 134904 47332 136784 47360
rect 134904 47320 134910 47332
rect 136778 47320 136784 47332
rect 136836 47320 136842 47372
rect 62718 47184 62724 47236
rect 62776 47224 62782 47236
rect 65018 47224 65024 47236
rect 62776 47196 65024 47224
rect 62776 47184 62782 47196
rect 65018 47184 65024 47196
rect 65076 47184 65082 47236
rect 62902 47116 62908 47168
rect 62960 47156 62966 47168
rect 64926 47156 64932 47168
rect 62960 47128 64932 47156
rect 62960 47116 62966 47128
rect 64926 47116 64932 47128
rect 64984 47116 64990 47168
rect 135306 47116 135312 47168
rect 135364 47156 135370 47168
rect 136686 47156 136692 47168
rect 135364 47128 136692 47156
rect 135364 47116 135370 47128
rect 136686 47116 136692 47128
rect 136744 47116 136750 47168
rect 63730 46368 63736 46420
rect 63788 46408 63794 46420
rect 66398 46408 66404 46420
rect 63788 46380 66404 46408
rect 63788 46368 63794 46380
rect 66398 46368 66404 46380
rect 66456 46368 66462 46420
rect 172658 46368 172664 46420
rect 172716 46408 172722 46420
rect 174038 46408 174044 46420
rect 172716 46380 174044 46408
rect 172716 46368 172722 46380
rect 174038 46368 174044 46380
rect 174096 46368 174102 46420
rect 100622 46232 100628 46284
rect 100680 46272 100686 46284
rect 102554 46272 102560 46284
rect 100680 46244 102560 46272
rect 100680 46232 100686 46244
rect 102554 46232 102560 46244
rect 102612 46232 102618 46284
rect 100898 46096 100904 46148
rect 100956 46136 100962 46148
rect 102370 46136 102376 46148
rect 100956 46108 102376 46136
rect 100956 46096 100962 46108
rect 102370 46096 102376 46108
rect 102428 46096 102434 46148
rect 134662 46028 134668 46080
rect 134720 46068 134726 46080
rect 136778 46068 136784 46080
rect 134720 46040 136784 46068
rect 134720 46028 134726 46040
rect 136778 46028 136784 46040
rect 136836 46028 136842 46080
rect 100530 45212 100536 45264
rect 100588 45252 100594 45264
rect 102462 45252 102468 45264
rect 100588 45224 102468 45252
rect 100588 45212 100594 45224
rect 102462 45212 102468 45224
rect 102520 45212 102526 45264
rect 99978 44940 99984 44992
rect 100036 44980 100042 44992
rect 102554 44980 102560 44992
rect 100036 44952 102560 44980
rect 100036 44940 100042 44952
rect 102554 44940 102560 44952
rect 102612 44940 102618 44992
rect 63730 44804 63736 44856
rect 63788 44844 63794 44856
rect 66398 44844 66404 44856
rect 63788 44816 66404 44844
rect 63788 44804 63794 44816
rect 66398 44804 66404 44816
rect 66456 44804 66462 44856
rect 63638 44736 63644 44788
rect 63696 44776 63702 44788
rect 65662 44776 65668 44788
rect 63696 44748 65668 44776
rect 63696 44736 63702 44748
rect 65662 44736 65668 44748
rect 65720 44736 65726 44788
rect 171830 44736 171836 44788
rect 171888 44776 171894 44788
rect 171888 44748 172796 44776
rect 171888 44736 171894 44748
rect 62810 44668 62816 44720
rect 62868 44708 62874 44720
rect 65294 44708 65300 44720
rect 62868 44680 65300 44708
rect 62868 44668 62874 44680
rect 65294 44668 65300 44680
rect 65352 44668 65358 44720
rect 135030 44668 135036 44720
rect 135088 44708 135094 44720
rect 137514 44708 137520 44720
rect 135088 44680 137520 44708
rect 135088 44668 135094 44680
rect 137514 44668 137520 44680
rect 137572 44668 137578 44720
rect 172768 44640 172796 44748
rect 172842 44668 172848 44720
rect 172900 44708 172906 44720
rect 174130 44708 174136 44720
rect 172900 44680 174136 44708
rect 172900 44668 172906 44680
rect 174130 44668 174136 44680
rect 174188 44668 174194 44720
rect 174682 44640 174688 44652
rect 172768 44612 174688 44640
rect 174682 44600 174688 44612
rect 174740 44600 174746 44652
rect 135398 44396 135404 44448
rect 135456 44436 135462 44448
rect 136686 44436 136692 44448
rect 135456 44408 136692 44436
rect 135456 44396 135462 44408
rect 136686 44396 136692 44408
rect 136744 44396 136750 44448
rect 135030 44260 135036 44312
rect 135088 44300 135094 44312
rect 136778 44300 136784 44312
rect 135088 44272 136784 44300
rect 135088 44260 135094 44272
rect 136778 44260 136784 44272
rect 136836 44260 136842 44312
rect 172750 44260 172756 44312
rect 172808 44300 172814 44312
rect 174498 44300 174504 44312
rect 172808 44272 174504 44300
rect 172808 44260 172814 44272
rect 174498 44260 174504 44272
rect 174556 44260 174562 44312
rect 99886 44056 99892 44108
rect 99944 44096 99950 44108
rect 102278 44096 102284 44108
rect 99944 44068 102284 44096
rect 99944 44056 99950 44068
rect 102278 44056 102284 44068
rect 102336 44056 102342 44108
rect 63914 43512 63920 43564
rect 63972 43552 63978 43564
rect 66398 43552 66404 43564
rect 63972 43524 66404 43552
rect 63972 43512 63978 43524
rect 66398 43512 66404 43524
rect 66456 43512 66462 43564
rect 171830 43512 171836 43564
rect 171888 43552 171894 43564
rect 174038 43552 174044 43564
rect 171888 43524 174044 43552
rect 171888 43512 171894 43524
rect 174038 43512 174044 43524
rect 174096 43512 174102 43564
rect 63730 43308 63736 43360
rect 63788 43348 63794 43360
rect 65294 43348 65300 43360
rect 63788 43320 65300 43348
rect 63788 43308 63794 43320
rect 65294 43308 65300 43320
rect 65352 43308 65358 43360
rect 100622 43308 100628 43360
rect 100680 43348 100686 43360
rect 136870 43348 136876 43360
rect 100680 43320 101036 43348
rect 100680 43308 100686 43320
rect 101008 43280 101036 43320
rect 135508 43320 136876 43348
rect 102370 43280 102376 43292
rect 101008 43252 102376 43280
rect 102370 43240 102376 43252
rect 102428 43240 102434 43292
rect 134938 43240 134944 43292
rect 134996 43280 135002 43292
rect 135508 43280 135536 43320
rect 136870 43308 136876 43320
rect 136928 43308 136934 43360
rect 172658 43308 172664 43360
rect 172716 43348 172722 43360
rect 172716 43320 172796 43348
rect 172716 43308 172722 43320
rect 134996 43252 135536 43280
rect 172768 43280 172796 43320
rect 174222 43280 174228 43292
rect 172768 43252 174228 43280
rect 134996 43240 135002 43252
rect 174222 43240 174228 43252
rect 174280 43240 174286 43292
rect 135398 43036 135404 43088
rect 135456 43076 135462 43088
rect 136778 43076 136784 43088
rect 135456 43048 136784 43076
rect 135456 43036 135462 43048
rect 136778 43036 136784 43048
rect 136836 43036 136842 43088
rect 63822 42832 63828 42884
rect 63880 42872 63886 42884
rect 66398 42872 66404 42884
rect 63880 42844 66404 42872
rect 63880 42832 63886 42844
rect 66398 42832 66404 42844
rect 66456 42832 66462 42884
rect 100622 42628 100628 42680
rect 100680 42668 100686 42680
rect 102554 42668 102560 42680
rect 100680 42640 102560 42668
rect 100680 42628 100686 42640
rect 102554 42628 102560 42640
rect 102612 42628 102618 42680
rect 172382 42288 172388 42340
rect 172440 42328 172446 42340
rect 173946 42328 173952 42340
rect 172440 42300 173952 42328
rect 172440 42288 172446 42300
rect 173946 42288 173952 42300
rect 174004 42288 174010 42340
rect 100622 42152 100628 42204
rect 100680 42192 100686 42204
rect 102462 42192 102468 42204
rect 100680 42164 102468 42192
rect 100680 42152 100686 42164
rect 102462 42152 102468 42164
rect 102520 42152 102526 42204
rect 100622 42016 100628 42068
rect 100680 42056 100686 42068
rect 102370 42056 102376 42068
rect 100680 42028 102376 42056
rect 100680 42016 100686 42028
rect 102370 42016 102376 42028
rect 102428 42016 102434 42068
rect 172658 42016 172664 42068
rect 172716 42056 172722 42068
rect 174038 42056 174044 42068
rect 172716 42028 174044 42056
rect 172716 42016 172722 42028
rect 174038 42016 174044 42028
rect 174096 42016 174102 42068
rect 63730 41948 63736 42000
rect 63788 41988 63794 42000
rect 66398 41988 66404 42000
rect 63788 41960 66404 41988
rect 63788 41948 63794 41960
rect 66398 41948 66404 41960
rect 66456 41948 66462 42000
rect 136870 41988 136876 42000
rect 135508 41960 136876 41988
rect 135398 41880 135404 41932
rect 135456 41920 135462 41932
rect 135508 41920 135536 41960
rect 136870 41948 136876 41960
rect 136928 41948 136934 42000
rect 172566 41948 172572 42000
rect 172624 41988 172630 42000
rect 172624 41960 172888 41988
rect 172624 41948 172630 41960
rect 135456 41892 135536 41920
rect 172860 41920 172888 41960
rect 174130 41920 174136 41932
rect 172860 41892 174136 41920
rect 135456 41880 135462 41892
rect 174130 41880 174136 41892
rect 174188 41880 174194 41932
rect 135306 41812 135312 41864
rect 135364 41852 135370 41864
rect 136686 41852 136692 41864
rect 135364 41824 136692 41852
rect 135364 41812 135370 41824
rect 136686 41812 136692 41824
rect 136744 41812 136750 41864
rect 134846 41472 134852 41524
rect 134904 41512 134910 41524
rect 136778 41512 136784 41524
rect 134904 41484 136784 41512
rect 134904 41472 134910 41484
rect 136778 41472 136784 41484
rect 136836 41472 136842 41524
rect 62810 40520 62816 40572
rect 62868 40560 62874 40572
rect 65294 40560 65300 40572
rect 62868 40532 65300 40560
rect 62868 40520 62874 40532
rect 65294 40520 65300 40532
rect 65352 40520 65358 40572
rect 71918 39908 71924 39960
rect 71976 39948 71982 39960
rect 82498 39948 82504 39960
rect 71976 39920 82504 39948
rect 71976 39908 71982 39920
rect 82498 39908 82504 39920
rect 82556 39908 82562 39960
rect 143586 39908 143592 39960
rect 143644 39948 143650 39960
rect 154810 39948 154816 39960
rect 143644 39920 154816 39948
rect 143644 39908 143650 39920
rect 154810 39908 154816 39920
rect 154868 39908 154874 39960
rect 66306 39840 66312 39892
rect 66364 39880 66370 39892
rect 86270 39880 86276 39892
rect 66364 39852 86276 39880
rect 66364 39840 66370 39852
rect 86270 39840 86276 39852
rect 86328 39840 86334 39892
rect 138066 39840 138072 39892
rect 138124 39880 138130 39892
rect 158582 39880 158588 39892
rect 138124 39852 158588 39880
rect 138124 39840 138130 39852
rect 158582 39840 158588 39852
rect 158640 39840 158646 39892
rect 62810 39160 62816 39212
rect 62868 39200 62874 39212
rect 72562 39200 72568 39212
rect 62868 39172 72568 39200
rect 62868 39160 62874 39172
rect 72562 39160 72568 39172
rect 72620 39160 72626 39212
rect 93170 39160 93176 39212
rect 93228 39200 93234 39212
rect 102370 39200 102376 39212
rect 93228 39172 102376 39200
rect 93228 39160 93234 39172
rect 102370 39160 102376 39172
rect 102428 39160 102434 39212
rect 134478 39160 134484 39212
rect 134536 39200 134542 39212
rect 144874 39200 144880 39212
rect 134536 39172 144880 39200
rect 134536 39160 134542 39172
rect 144874 39160 144880 39172
rect 144932 39160 144938 39212
rect 164838 39160 164844 39212
rect 164896 39200 164902 39212
rect 174130 39200 174136 39212
rect 164896 39172 174136 39200
rect 164896 39160 164902 39172
rect 174130 39160 174136 39172
rect 174188 39160 174194 39212
rect 79370 37732 79376 37784
rect 79428 37772 79434 37784
rect 127762 37772 127768 37784
rect 79428 37744 127768 37772
rect 79428 37732 79434 37744
rect 127762 37732 127768 37744
rect 127820 37732 127826 37784
rect 151038 37732 151044 37784
rect 151096 37772 151102 37784
rect 200074 37772 200080 37784
rect 151096 37744 200080 37772
rect 151096 37732 151102 37744
rect 200074 37732 200080 37744
rect 200132 37732 200138 37784
rect 222522 37772 222528 37784
rect 222483 37744 222528 37772
rect 222522 37732 222528 37744
rect 222580 37732 222586 37784
rect 190782 37664 190788 37716
rect 190840 37704 190846 37716
rect 205134 37704 205140 37716
rect 190840 37676 205140 37704
rect 190840 37664 190846 37676
rect 205134 37664 205140 37676
rect 205192 37664 205198 37716
rect 30518 33584 30524 33636
rect 30576 33624 30582 33636
rect 66214 33624 66220 33636
rect 30576 33596 66220 33624
rect 30576 33584 30582 33596
rect 66214 33584 66220 33596
rect 66272 33584 66278 33636
rect 118838 33584 118844 33636
rect 118896 33624 118902 33636
rect 136870 33624 136876 33636
rect 118896 33596 136876 33624
rect 118896 33584 118902 33596
rect 136870 33584 136876 33596
rect 136928 33584 136934 33636
rect 222525 28187 222583 28193
rect 222525 28153 222537 28187
rect 222571 28184 222583 28187
rect 222706 28184 222712 28196
rect 222571 28156 222712 28184
rect 222571 28153 222583 28156
rect 222525 28147 222583 28153
rect 222706 28144 222712 28156
rect 222764 28144 222770 28196
rect 77990 12572 77996 12624
rect 78048 12612 78054 12624
rect 79048 12612 79054 12624
rect 78048 12584 79054 12612
rect 78048 12572 78054 12584
rect 79048 12572 79054 12584
rect 79106 12572 79112 12624
rect 86914 11688 86920 11740
rect 86972 11728 86978 11740
rect 132546 11728 132552 11740
rect 86972 11700 132552 11728
rect 86972 11688 86978 11700
rect 132546 11688 132552 11700
rect 132604 11688 132610 11740
rect 166034 11688 166040 11740
rect 166092 11728 166098 11740
rect 214242 11728 214248 11740
rect 166092 11700 214248 11728
rect 166092 11688 166098 11700
rect 214242 11688 214248 11700
rect 214300 11688 214306 11740
rect 93998 11620 94004 11672
rect 94056 11660 94062 11672
rect 187010 11660 187016 11672
rect 94056 11632 187016 11660
rect 94056 11620 94062 11632
rect 187010 11620 187016 11632
rect 187068 11620 187074 11672
rect 23526 10940 23532 10992
rect 23584 10980 23590 10992
rect 71274 10980 71280 10992
rect 23584 10952 71280 10980
rect 23584 10940 23590 10952
rect 71274 10940 71280 10952
rect 71332 10940 71338 10992
rect 105222 10940 105228 10992
rect 105280 10980 105286 10992
rect 151038 10980 151044 10992
rect 105280 10952 151044 10980
rect 105280 10940 105286 10952
rect 151038 10940 151044 10952
rect 151096 10940 151102 10992
rect 50758 10872 50764 10924
rect 50816 10912 50822 10924
rect 143586 10912 143592 10924
rect 50816 10884 143592 10912
rect 50816 10872 50822 10884
rect 143586 10872 143592 10884
rect 143644 10872 143650 10924
rect 158582 10396 158588 10448
rect 158640 10436 158646 10448
rect 159778 10436 159784 10448
rect 158640 10408 159784 10436
rect 158640 10396 158646 10408
rect 159778 10396 159784 10408
rect 159836 10396 159842 10448
<< via1 >>
rect 23532 244860 23584 244912
rect 70544 244860 70596 244912
rect 105228 244860 105280 244912
rect 149664 244860 149716 244912
rect 50764 244792 50816 244844
rect 142396 244792 142448 244844
rect 157484 244792 157536 244844
rect 159784 244792 159836 244844
rect 85632 242412 85684 242464
rect 132552 242140 132604 242192
rect 165304 242140 165356 242192
rect 214248 242140 214300 242192
rect 93360 242072 93412 242124
rect 187016 242072 187068 242124
rect 167788 229764 167840 229816
rect 168524 229764 168576 229816
rect 207256 223372 207308 223424
rect 223080 223372 223132 223424
rect 170088 222760 170140 222812
rect 207256 222760 207308 222812
rect 71280 217932 71332 217984
rect 143684 217932 143736 217984
rect 170088 217932 170140 217984
rect 46532 217864 46584 217916
rect 98236 217864 98288 217916
rect 98420 217864 98472 217916
rect 109276 217864 109328 217916
rect 118844 217864 118896 217916
rect 169996 217864 170048 217916
rect 109276 217252 109328 217304
rect 143684 217252 143736 217304
rect 37240 217184 37292 217236
rect 71280 217184 71332 217236
rect 79376 217184 79428 217236
rect 127768 217184 127820 217236
rect 81768 216572 81820 216624
rect 94004 216572 94056 216624
rect 158588 216572 158640 216624
rect 167236 216572 167288 216624
rect 91796 216504 91848 216556
rect 102376 216504 102428 216556
rect 164108 216504 164160 216556
rect 174228 216504 174280 216556
rect 86920 216436 86972 216488
rect 98328 216436 98380 216488
rect 154080 216436 154132 216488
rect 166040 216436 166092 216488
rect 62540 215756 62592 215808
rect 71832 215756 71884 215808
rect 135404 215756 135456 215808
rect 143776 215756 143828 215808
rect 100996 214600 101048 214652
rect 102376 214600 102428 214652
rect 62632 214464 62684 214516
rect 65024 214464 65076 214516
rect 135404 214464 135456 214516
rect 136784 214464 136836 214516
rect 171836 213988 171888 214040
rect 174044 213988 174096 214040
rect 100996 213308 101048 213360
rect 102376 213308 102428 213360
rect 135036 213308 135088 213360
rect 136784 213308 136836 213360
rect 62540 213240 62592 213292
rect 65024 213240 65076 213292
rect 63736 213036 63788 213088
rect 66220 213036 66272 213088
rect 100536 213036 100588 213088
rect 102468 213104 102520 213156
rect 135404 213104 135456 213156
rect 136876 213036 136928 213088
rect 172664 213036 172716 213088
rect 174228 213104 174280 213156
rect 171744 212968 171796 213020
rect 174044 212968 174096 213020
rect 101088 212220 101140 212272
rect 102376 212220 102428 212272
rect 134668 212084 134720 212136
rect 136968 212084 137020 212136
rect 100996 211880 101048 211932
rect 102376 211880 102428 211932
rect 62632 211744 62684 211796
rect 65024 211744 65076 211796
rect 134300 211744 134352 211796
rect 136876 211744 136928 211796
rect 62356 211676 62408 211728
rect 64932 211676 64984 211728
rect 172664 211608 172716 211660
rect 174228 211676 174280 211728
rect 172572 211404 172624 211456
rect 174044 211404 174096 211456
rect 62632 211064 62684 211116
rect 65484 211064 65536 211116
rect 171836 210724 171888 210776
rect 174136 210724 174188 210776
rect 62632 210384 62684 210436
rect 65024 210384 65076 210436
rect 207900 210316 207952 210368
rect 223540 210316 223592 210368
rect 171928 209636 171980 209688
rect 174136 209636 174188 209688
rect 62632 209500 62684 209552
rect 65484 209500 65536 209552
rect 62724 209024 62776 209076
rect 65024 209024 65076 209076
rect 135312 209024 135364 209076
rect 137704 209024 137756 209076
rect 171468 208888 171520 208940
rect 174596 208956 174648 209008
rect 62540 208072 62592 208124
rect 65668 208072 65720 208124
rect 135404 207664 135456 207716
rect 136876 207664 136928 207716
rect 172572 207324 172624 207376
rect 174044 207324 174096 207376
rect 62632 206848 62684 206900
rect 65668 206848 65720 206900
rect 172664 202224 172716 202276
rect 174228 202224 174280 202276
rect 62632 201884 62684 201936
rect 65024 201884 65076 201936
rect 172664 200728 172716 200780
rect 174136 200728 174188 200780
rect 100904 200660 100956 200712
rect 102376 200660 102428 200712
rect 135404 200456 135456 200508
rect 136784 200456 136836 200508
rect 62632 200388 62684 200440
rect 65024 200388 65076 200440
rect 171652 199368 171704 199420
rect 175240 199368 175292 199420
rect 100904 199300 100956 199352
rect 102376 199300 102428 199352
rect 134760 199096 134812 199148
rect 136784 199096 136836 199148
rect 62356 199028 62408 199080
rect 65024 199028 65076 199080
rect 172664 198144 172716 198196
rect 174136 198144 174188 198196
rect 100812 198008 100864 198060
rect 102376 198008 102428 198060
rect 172664 198008 172716 198060
rect 174228 198008 174280 198060
rect 62540 197804 62592 197856
rect 65668 197872 65720 197924
rect 100904 197872 100956 197924
rect 102468 197872 102520 197924
rect 62632 197736 62684 197788
rect 65024 197736 65076 197788
rect 135404 197736 135456 197788
rect 136784 197736 136836 197788
rect 135404 197396 135456 197448
rect 136692 197396 136744 197448
rect 172572 196784 172624 196836
rect 174136 196784 174188 196836
rect 100720 196648 100772 196700
rect 102376 196648 102428 196700
rect 62632 196444 62684 196496
rect 66220 196512 66272 196564
rect 100904 196512 100956 196564
rect 102468 196512 102520 196564
rect 172664 196512 172716 196564
rect 174228 196512 174280 196564
rect 135404 196376 135456 196428
rect 136784 196376 136836 196428
rect 62540 196308 62592 196360
rect 65024 196308 65076 196360
rect 135404 196172 135456 196224
rect 136692 196172 136744 196224
rect 100904 195424 100956 195476
rect 102560 195424 102612 195476
rect 172664 195288 172716 195340
rect 174136 195288 174188 195340
rect 172388 195220 172440 195272
rect 174228 195220 174280 195272
rect 62540 195084 62592 195136
rect 66404 195152 66456 195204
rect 100904 195152 100956 195204
rect 102376 195152 102428 195204
rect 135404 195084 135456 195136
rect 136876 195152 136928 195204
rect 62632 195016 62684 195068
rect 65024 195016 65076 195068
rect 135404 194812 135456 194864
rect 136784 194812 136836 194864
rect 100628 194336 100680 194388
rect 102468 194336 102520 194388
rect 171744 193928 171796 193980
rect 174136 193928 174188 193980
rect 172664 193860 172716 193912
rect 174228 193860 174280 193912
rect 100628 193792 100680 193844
rect 102376 193792 102428 193844
rect 62632 193656 62684 193708
rect 66404 193724 66456 193776
rect 135404 193656 135456 193708
rect 136784 193656 136836 193708
rect 62540 193588 62592 193640
rect 65024 193588 65076 193640
rect 135404 193452 135456 193504
rect 136692 193452 136744 193504
rect 99892 192908 99944 192960
rect 102468 192908 102520 192960
rect 172664 192704 172716 192756
rect 174228 192704 174280 192756
rect 172020 192636 172072 192688
rect 174136 192636 174188 192688
rect 171652 192568 171704 192620
rect 174320 192568 174372 192620
rect 62632 192432 62684 192484
rect 65668 192432 65720 192484
rect 100628 192432 100680 192484
rect 102376 192432 102428 192484
rect 100536 192364 100588 192416
rect 102652 192364 102704 192416
rect 135312 192364 135364 192416
rect 136876 192364 136928 192416
rect 135404 192296 135456 192348
rect 136784 192296 136836 192348
rect 62540 192228 62592 192280
rect 64932 192228 64984 192280
rect 135220 192092 135272 192144
rect 136692 192092 136744 192144
rect 62356 191616 62408 191668
rect 65024 191616 65076 191668
rect 100628 191208 100680 191260
rect 102284 191208 102336 191260
rect 172664 191208 172716 191260
rect 174044 191208 174096 191260
rect 171836 191072 171888 191124
rect 175332 191072 175384 191124
rect 100904 191004 100956 191056
rect 102560 191004 102612 191056
rect 134208 191004 134260 191056
rect 137152 191004 137204 191056
rect 62356 190800 62408 190852
rect 65024 190800 65076 190852
rect 135404 190732 135456 190784
rect 136784 190732 136836 190784
rect 100444 190120 100496 190172
rect 102376 190120 102428 190172
rect 171652 189916 171704 189968
rect 174412 189916 174464 189968
rect 99984 189848 100036 189900
rect 102468 189848 102520 189900
rect 171836 189712 171888 189764
rect 175424 189712 175476 189764
rect 63644 189644 63696 189696
rect 66404 189644 66456 189696
rect 62632 189508 62684 189560
rect 65208 189508 65260 189560
rect 134760 189236 134812 189288
rect 136784 189236 136836 189288
rect 62632 189032 62684 189084
rect 65024 189032 65076 189084
rect 134944 188148 134996 188200
rect 137244 188148 137296 188200
rect 116452 187604 116504 187656
rect 117418 187604 117470 187656
rect 183980 186856 184032 186908
rect 184440 186856 184492 186908
rect 188488 186856 188540 186908
rect 189132 186856 189184 186908
rect 36320 185428 36372 185480
rect 40644 185428 40696 185480
rect 41012 185428 41064 185480
rect 43404 185428 43456 185480
rect 43772 185428 43824 185480
rect 44692 185428 44744 185480
rect 49016 185428 49068 185480
rect 50580 185428 50632 185480
rect 50672 185428 50724 185480
rect 53340 185428 53392 185480
rect 53432 185428 53484 185480
rect 58124 185428 58176 185480
rect 110104 185428 110156 185480
rect 111116 185428 111168 185480
rect 117556 185428 117608 185480
rect 118936 185428 118988 185480
rect 120224 185428 120276 185480
rect 122340 185428 122392 185480
rect 122432 185428 122484 185480
rect 123444 185428 123496 185480
rect 124180 185428 124232 185480
rect 128136 185428 128188 185480
rect 182232 185428 182284 185480
rect 183244 185428 183296 185480
rect 188120 185428 188172 185480
rect 188580 185428 188632 185480
rect 190604 185428 190656 185480
rect 192536 185428 192588 185480
rect 192904 185428 192956 185480
rect 195388 185428 195440 185480
rect 197320 185428 197372 185480
rect 201644 185428 201696 185480
rect 40368 185360 40420 185412
rect 43036 185360 43088 185412
rect 43128 185360 43180 185412
rect 44600 185360 44652 185412
rect 49844 185360 49896 185412
rect 51960 185360 52012 185412
rect 110748 185360 110800 185412
rect 111484 185360 111536 185412
rect 118568 185360 118620 185412
rect 120316 185360 120368 185412
rect 124548 185360 124600 185412
rect 128688 185360 128740 185412
rect 191708 185360 191760 185412
rect 193640 185360 193692 185412
rect 194100 185360 194152 185412
rect 197136 185360 197188 185412
rect 37608 185292 37660 185344
rect 41472 185292 41524 185344
rect 41748 185292 41800 185344
rect 43864 185292 43916 185344
rect 52236 185292 52288 185344
rect 56100 185292 56152 185344
rect 123812 185292 123864 185344
rect 127584 185292 127636 185344
rect 176896 185292 176948 185344
rect 177724 185292 177776 185344
rect 192536 185292 192588 185344
rect 194836 185292 194888 185344
rect 195756 185292 195808 185344
rect 199344 185292 199396 185344
rect 39724 185224 39776 185276
rect 42668 185224 42720 185276
rect 49476 185224 49528 185276
rect 51316 185224 51368 185276
rect 53064 185224 53116 185276
rect 57388 185224 57440 185276
rect 105596 185224 105648 185276
rect 109276 185224 109328 185276
rect 118936 185224 118988 185276
rect 120592 185224 120644 185276
rect 123352 185224 123404 185276
rect 127308 185224 127360 185276
rect 193364 185224 193416 185276
rect 195940 185224 195992 185276
rect 196124 185224 196176 185276
rect 199988 185224 200040 185276
rect 36964 185156 37016 185208
rect 41012 185156 41064 185208
rect 50212 185156 50264 185208
rect 52696 185156 52748 185208
rect 122616 185156 122668 185208
rect 125836 185156 125888 185208
rect 177724 185156 177776 185208
rect 181128 185156 181180 185208
rect 194560 185156 194612 185208
rect 197688 185156 197740 185208
rect 34940 185088 34992 185140
rect 39540 185088 39592 185140
rect 42392 185088 42444 185140
rect 44232 185088 44284 185140
rect 52604 185088 52656 185140
rect 56744 185088 56796 185140
rect 122984 185088 123036 185140
rect 126388 185088 126440 185140
rect 190420 185088 190472 185140
rect 191984 185088 192036 185140
rect 193732 185088 193784 185140
rect 196492 185088 196544 185140
rect 38988 185020 39040 185072
rect 42208 185020 42260 185072
rect 48648 185020 48700 185072
rect 49936 185020 49988 185072
rect 51040 185020 51092 185072
rect 53984 185020 54036 185072
rect 121328 185020 121380 185072
rect 124456 185020 124508 185072
rect 194652 185020 194704 185072
rect 198240 185020 198292 185072
rect 38344 184952 38396 185004
rect 41840 184952 41892 185004
rect 51408 184952 51460 185004
rect 54720 184952 54772 185004
rect 121788 184952 121840 185004
rect 124640 184952 124692 185004
rect 181680 184952 181732 185004
rect 183106 184952 183158 185004
rect 183428 184952 183480 185004
rect 184302 184952 184354 185004
rect 188626 184952 188678 185004
rect 189684 184952 189736 185004
rect 189822 184952 189874 185004
rect 191432 184952 191484 185004
rect 191846 184952 191898 185004
rect 194284 184952 194336 185004
rect 197826 184952 197878 185004
rect 202840 184952 202892 185004
rect 51868 184884 51920 184936
rect 55364 184884 55416 184936
rect 122156 184884 122208 184936
rect 125192 184884 125244 184936
rect 182876 184884 182928 184936
rect 183842 184884 183894 184936
rect 189086 184884 189138 184936
rect 190236 184884 190288 184936
rect 191110 184884 191162 184936
rect 193088 184884 193140 184936
rect 196630 184884 196682 184936
rect 201092 184884 201144 184936
rect 189684 184816 189736 184868
rect 190788 184816 190840 184868
rect 196492 184816 196544 184868
rect 200540 184816 200592 184868
rect 195296 184748 195348 184800
rect 198792 184748 198844 184800
rect 35584 184408 35636 184460
rect 38160 184408 38212 184460
rect 39264 184408 39316 184460
rect 53984 184408 54036 184460
rect 54536 184408 54588 184460
rect 34204 184272 34256 184324
rect 33560 184068 33612 184120
rect 38896 184068 38948 184120
rect 106056 184340 106108 184392
rect 107160 184340 107212 184392
rect 176988 184340 177040 184392
rect 179380 184340 179432 184392
rect 59504 184204 59556 184256
rect 177632 184136 177684 184188
rect 178276 184136 178328 184188
rect 58768 184068 58820 184120
rect 105964 184068 106016 184120
rect 106608 184068 106660 184120
rect 106148 184000 106200 184052
rect 108356 184068 108408 184120
rect 177816 184068 177868 184120
rect 178828 184068 178880 184120
rect 177356 184000 177408 184052
rect 180576 184068 180628 184120
rect 105596 182368 105648 182420
rect 107896 182368 107948 182420
rect 177172 182164 177224 182216
rect 180024 182164 180076 182216
rect 105412 180328 105464 180380
rect 108080 180328 108132 180380
rect 178092 180328 178144 180380
rect 179656 180328 179708 180380
rect 106332 178560 106384 178612
rect 107896 178560 107948 178612
rect 177816 178560 177868 178612
rect 179656 178560 179708 178612
rect 32640 177200 32692 177252
rect 37424 177200 37476 177252
rect 106424 175840 106476 175892
rect 107896 175840 107948 175892
rect 177724 175840 177776 175892
rect 179656 175840 179708 175892
rect 57388 175772 57440 175824
rect 59596 175772 59648 175824
rect 177172 175568 177224 175620
rect 180300 175568 180352 175620
rect 106148 175364 106200 175416
rect 108540 175364 108592 175416
rect 105964 173052 106016 173104
rect 107896 173052 107948 173104
rect 177540 173052 177592 173104
rect 179656 173052 179708 173104
rect 105688 171692 105740 171744
rect 108080 171692 108132 171744
rect 178184 171692 178236 171744
rect 179656 171692 179708 171744
rect 222804 169108 222856 169160
rect 223540 169108 223592 169160
rect 201092 166116 201144 166168
rect 204496 166116 204548 166168
rect 177172 165300 177224 165352
rect 179564 165300 179616 165352
rect 105228 165232 105280 165284
rect 107804 165232 107856 165284
rect 28868 164756 28920 164808
rect 37424 164756 37476 164808
rect 54812 164756 54864 164808
rect 59596 164756 59648 164808
rect 177540 163600 177592 163652
rect 179564 163600 179616 163652
rect 105596 163464 105648 163516
rect 107436 163464 107488 163516
rect 105780 163396 105832 163448
rect 107804 163396 107856 163448
rect 176988 163396 177040 163448
rect 179196 163396 179248 163448
rect 105688 162036 105740 162088
rect 107804 162036 107856 162088
rect 176988 162036 177040 162088
rect 179564 162036 179616 162088
rect 105228 161016 105280 161068
rect 107712 161016 107764 161068
rect 177540 160880 177592 160932
rect 179472 160880 179524 160932
rect 105596 159520 105648 159572
rect 107620 159520 107672 159572
rect 177356 159248 177408 159300
rect 179380 159248 179432 159300
rect 105780 158296 105832 158348
rect 108724 158296 108776 158348
rect 177632 157956 177684 158008
rect 180484 157956 180536 158008
rect 106148 157888 106200 157940
rect 108632 157888 108684 157940
rect 178184 157888 178236 157940
rect 180392 157888 180444 157940
rect 222804 156868 222856 156920
rect 223540 156868 223592 156920
rect 106148 156664 106200 156716
rect 108540 156664 108592 156716
rect 177356 156460 177408 156512
rect 180300 156460 180352 156512
rect 105780 155304 105832 155356
rect 107896 155304 107948 155356
rect 178092 155100 178144 155152
rect 179656 155100 179708 155152
rect 57480 151496 57532 151548
rect 59596 151496 59648 151548
rect 200540 151496 200592 151548
rect 207348 151496 207400 151548
rect 105964 147008 106016 147060
rect 108356 147008 108408 147060
rect 177356 146872 177408 146924
rect 180576 146872 180628 146924
rect 178276 146124 178328 146176
rect 179012 146124 179064 146176
rect 22244 145172 22296 145224
rect 28684 145172 28736 145224
rect 207348 145172 207400 145224
rect 210016 145172 210068 145224
rect 210292 145172 210344 145224
rect 178368 145104 178420 145156
rect 181128 145104 181180 145156
rect 106700 144832 106752 144884
rect 109276 144832 109328 144884
rect 191846 144696 191898 144748
rect 194284 144696 194336 144748
rect 191478 144628 191530 144680
rect 193640 144628 193692 144680
rect 197826 144628 197878 144680
rect 202840 144628 202892 144680
rect 135496 144424 135548 144476
rect 136324 144424 136376 144476
rect 125836 144220 125888 144272
rect 131448 144220 131500 144272
rect 190604 144220 190656 144272
rect 192536 144220 192588 144272
rect 198884 144220 198936 144272
rect 203944 144220 203996 144272
rect 40644 144152 40696 144204
rect 43036 144152 43088 144204
rect 54260 144152 54312 144204
rect 59780 144152 59832 144204
rect 120224 144152 120276 144204
rect 122340 144152 122392 144204
rect 126664 144152 126716 144204
rect 132184 144152 132236 144204
rect 198516 144152 198568 144204
rect 203392 144152 203444 144204
rect 41288 144084 41340 144136
rect 43404 144084 43456 144136
rect 54628 144084 54680 144136
rect 60424 144084 60476 144136
rect 105228 144084 105280 144136
rect 105964 144084 106016 144136
rect 106516 144084 106568 144136
rect 107160 144084 107212 144136
rect 118936 144084 118988 144136
rect 120592 144084 120644 144136
rect 126296 144084 126348 144136
rect 131632 144084 131684 144136
rect 132644 144084 132696 144136
rect 174136 144084 174188 144136
rect 197504 144084 197556 144136
rect 202196 144084 202248 144136
rect 132644 143447 132696 143456
rect 132644 143413 132653 143447
rect 132653 143413 132687 143447
rect 132687 143413 132696 143447
rect 132644 143404 132696 143413
rect 34112 142656 34164 142708
rect 39080 142656 39132 142708
rect 39264 142656 39316 142708
rect 42208 142656 42260 142708
rect 43404 142656 43456 142708
rect 44600 142656 44652 142708
rect 48280 142656 48332 142708
rect 49476 142656 49528 142708
rect 51040 142656 51092 142708
rect 53800 142656 53852 142708
rect 58676 142656 58728 142708
rect 62816 142656 62868 142708
rect 16724 142588 16776 142640
rect 31904 142588 31956 142640
rect 34664 142588 34716 142640
rect 39448 142588 39500 142640
rect 42668 142588 42720 142640
rect 44232 142588 44284 142640
rect 47820 142588 47872 142640
rect 48832 142588 48884 142640
rect 49752 142588 49804 142640
rect 51592 142588 51644 142640
rect 53064 142588 53116 142640
rect 57664 142588 57716 142640
rect 37240 142520 37292 142572
rect 41012 142520 41064 142572
rect 50212 142520 50264 142572
rect 52972 142520 53024 142572
rect 53432 142520 53484 142572
rect 58124 142520 58176 142572
rect 66496 142656 66548 142708
rect 67876 142656 67928 142708
rect 72844 142656 72896 142708
rect 74500 142656 74552 142708
rect 74776 142656 74828 142708
rect 75604 142656 75656 142708
rect 80112 142656 80164 142708
rect 81676 142656 81728 142708
rect 84528 142656 84580 142708
rect 89128 142656 89180 142708
rect 95476 142656 95528 142708
rect 96764 142656 96816 142708
rect 110104 142656 110156 142708
rect 111116 142656 111168 142708
rect 120684 142656 120736 142708
rect 123444 142656 123496 142708
rect 125468 142656 125520 142708
rect 130436 142656 130488 142708
rect 153252 142656 153304 142708
rect 155828 142656 155880 142708
rect 156564 142656 156616 142708
rect 161440 142656 161492 142708
rect 182232 142656 182284 142708
rect 183244 142656 183296 142708
rect 189684 142656 189736 142708
rect 190788 142656 190840 142708
rect 191340 142656 191392 142708
rect 193088 142656 193140 142708
rect 196492 142656 196544 142708
rect 200540 142656 200592 142708
rect 201000 142656 201052 142708
rect 215904 142656 215956 142708
rect 81216 142588 81268 142640
rect 83516 142588 83568 142640
rect 86736 142588 86788 142640
rect 92808 142588 92860 142640
rect 119120 142588 119172 142640
rect 121144 142588 121196 142640
rect 123904 142588 123956 142640
rect 128136 142588 128188 142640
rect 154356 142588 154408 142640
rect 157668 142588 157720 142640
rect 163280 142588 163332 142640
rect 174412 142588 174464 142640
rect 189316 142588 189368 142640
rect 190236 142588 190288 142640
rect 190512 142588 190564 142640
rect 191984 142588 192036 142640
rect 194100 142588 194152 142640
rect 197136 142588 197188 142640
rect 71188 142520 71240 142572
rect 121052 142520 121104 142572
rect 124456 142520 124508 142572
rect 124640 142520 124692 142572
rect 129332 142520 129384 142572
rect 134116 142520 134168 142572
rect 143224 142520 143276 142572
rect 155460 142520 155512 142572
rect 159508 142520 159560 142572
rect 181680 142520 181732 142572
rect 182784 142520 182836 142572
rect 193732 142520 193784 142572
rect 196492 142520 196544 142572
rect 27580 142452 27632 142504
rect 36596 142384 36648 142436
rect 40368 142384 40420 142436
rect 48648 142384 48700 142436
rect 50212 142384 50264 142436
rect 50672 142452 50724 142504
rect 53616 142452 53668 142504
rect 54260 142452 54312 142504
rect 102284 142452 102336 142504
rect 174320 142452 174372 142504
rect 194560 142452 194612 142504
rect 197688 142452 197740 142504
rect 52236 142384 52288 142436
rect 56100 142384 56152 142436
rect 69164 142384 69216 142436
rect 72292 142384 72344 142436
rect 85632 142384 85684 142436
rect 90968 142384 91020 142436
rect 117464 142384 117516 142436
rect 118844 142384 118896 142436
rect 119488 142384 119540 142436
rect 121696 142384 121748 142436
rect 124272 142384 124324 142436
rect 128688 142384 128740 142436
rect 159876 142384 159928 142436
rect 167052 142384 167104 142436
rect 192904 142384 192956 142436
rect 195388 142384 195440 142436
rect 195756 142384 195808 142436
rect 199068 142384 199120 142436
rect 51868 142316 51920 142368
rect 55364 142316 55416 142368
rect 98972 142316 99024 142368
rect 102284 142316 102336 142368
rect 123720 142316 123772 142368
rect 127584 142316 127636 142368
rect 160980 142316 161032 142368
rect 168892 142316 168944 142368
rect 192444 142316 192496 142368
rect 194836 142316 194888 142368
rect 196952 142316 197004 142368
rect 201092 142316 201144 142368
rect 31904 142248 31956 142300
rect 40000 142248 40052 142300
rect 42300 142248 42352 142300
rect 38620 142180 38672 142232
rect 41840 142180 41892 142232
rect 37884 142112 37936 142164
rect 41472 142112 41524 142164
rect 42024 142112 42076 142164
rect 43864 142112 43916 142164
rect 51408 142248 51460 142300
rect 54996 142248 55048 142300
rect 62356 142248 62408 142300
rect 63460 142248 63512 142300
rect 116636 142248 116688 142300
rect 117648 142248 117700 142300
rect 120316 142248 120368 142300
rect 123076 142248 123128 142300
rect 125100 142248 125152 142300
rect 129884 142248 129936 142300
rect 167696 142248 167748 142300
rect 174320 142248 174372 142300
rect 182876 142248 182928 142300
rect 183612 142248 183664 142300
rect 193364 142248 193416 142300
rect 195940 142248 195992 142300
rect 197320 142248 197372 142300
rect 201644 142248 201696 142300
rect 49016 142180 49068 142232
rect 50856 142180 50908 142232
rect 49844 142044 49896 142096
rect 52236 142180 52288 142232
rect 121512 142180 121564 142232
rect 124640 142180 124692 142232
rect 134484 142180 134536 142232
rect 135496 142180 135548 142232
rect 142672 142180 142724 142232
rect 145432 142180 145484 142232
rect 172112 142180 172164 142232
rect 175240 142180 175292 142232
rect 196124 142180 196176 142232
rect 199620 142180 199672 142232
rect 54904 142112 54956 142164
rect 63460 142112 63512 142164
rect 64564 142112 64616 142164
rect 87840 142112 87892 142164
rect 94740 142112 94792 142164
rect 117096 142112 117148 142164
rect 118200 142112 118252 142164
rect 118292 142112 118344 142164
rect 119948 142112 120000 142164
rect 123352 142112 123404 142164
rect 126940 142112 126992 142164
rect 158772 142112 158824 142164
rect 165120 142112 165172 142164
rect 166592 142112 166644 142164
rect 175424 142112 175476 142164
rect 194652 142112 194704 142164
rect 198240 142112 198292 142164
rect 57480 142044 57532 142096
rect 134576 142044 134628 142096
rect 135588 142044 135640 142096
rect 165488 142044 165540 142096
rect 175148 142044 175200 142096
rect 195296 142044 195348 142096
rect 198792 142044 198844 142096
rect 222528 142044 222580 142096
rect 222804 142044 222856 142096
rect 52604 141976 52656 142028
rect 57020 141976 57072 142028
rect 83424 141976 83476 142028
rect 87288 141976 87340 142028
rect 88944 141976 88996 142028
rect 96856 141976 96908 142028
rect 100076 141976 100128 142028
rect 103112 141976 103164 142028
rect 110426 141976 110478 142028
rect 111484 141976 111536 142028
rect 113278 141976 113330 142028
rect 113508 141976 113560 142028
rect 116268 141976 116320 142028
rect 117418 141976 117470 142028
rect 117832 141976 117884 142028
rect 119718 141976 119770 142028
rect 121880 141976 121932 142028
rect 125514 141976 125566 142028
rect 134300 141976 134352 142028
rect 136876 141976 136928 142028
rect 168800 141976 168852 142028
rect 172848 141976 172900 142028
rect 190144 141976 190196 142028
rect 191432 141976 191484 142028
rect 207992 141976 208044 142028
rect 221240 141976 221292 142028
rect 101180 141908 101232 141960
rect 173216 141908 173268 141960
rect 207900 141908 207952 141960
rect 210016 141908 210068 141960
rect 222528 141908 222580 141960
rect 223540 141908 223592 141960
rect 71004 141840 71056 141892
rect 73396 141840 73448 141892
rect 132368 141840 132420 141892
rect 122892 141772 122944 141824
rect 126388 141772 126440 141824
rect 35584 141704 35636 141756
rect 39816 141704 39868 141756
rect 122248 141704 122300 141756
rect 125836 141704 125888 141756
rect 35952 141636 36004 141688
rect 40184 141636 40236 141688
rect 82320 141500 82372 141552
rect 85356 141500 85408 141552
rect 152148 141772 152200 141824
rect 153896 141772 153948 141824
rect 144512 141636 144564 141688
rect 146536 141636 146588 141688
rect 157944 141568 157996 141620
rect 163280 141568 163332 141620
rect 146444 141500 146496 141552
rect 147640 141500 147692 141552
rect 151044 141500 151096 141552
rect 152056 141500 152108 141552
rect 169904 141364 169956 141416
rect 90140 141296 90192 141348
rect 92348 141296 92400 141348
rect 93452 141296 93504 141348
rect 97868 141296 97920 141348
rect 62816 141228 62868 141280
rect 69256 141228 69308 141280
rect 62724 141160 62776 141212
rect 68060 141160 68112 141212
rect 132644 141296 132696 141348
rect 140832 141296 140884 141348
rect 144328 141296 144380 141348
rect 164384 141296 164436 141348
rect 171008 141296 171060 141348
rect 102376 141160 102428 141212
rect 174228 141228 174280 141280
rect 174780 141160 174832 141212
rect 135404 141092 135456 141144
rect 141108 141092 141160 141144
rect 135404 140684 135456 140736
rect 141016 140684 141068 140736
rect 62816 139868 62868 139920
rect 66496 139868 66548 139920
rect 95476 139868 95528 139920
rect 102376 139868 102428 139920
rect 172848 139868 172900 139920
rect 174964 139868 175016 139920
rect 95568 139800 95620 139852
rect 102468 139800 102520 139852
rect 135404 139800 135456 139852
rect 139544 139800 139596 139852
rect 62724 139732 62776 139784
rect 65116 139732 65168 139784
rect 94096 139732 94148 139784
rect 102560 139732 102612 139784
rect 62816 139596 62868 139648
rect 66588 139596 66640 139648
rect 135404 139460 135456 139512
rect 138256 139460 138308 139512
rect 172480 138712 172532 138764
rect 174228 138712 174280 138764
rect 62908 138644 62960 138696
rect 66404 138644 66456 138696
rect 135128 138644 135180 138696
rect 136968 138644 137020 138696
rect 172664 138644 172716 138696
rect 174320 138644 174372 138696
rect 62816 138576 62868 138628
rect 66220 138576 66272 138628
rect 135404 138576 135456 138628
rect 136876 138576 136928 138628
rect 102376 138508 102428 138560
rect 102468 138440 102520 138492
rect 174136 138440 174188 138492
rect 100996 138372 101048 138424
rect 62724 137216 62776 137268
rect 66220 137216 66272 137268
rect 135220 137216 135272 137268
rect 136968 137216 137020 137268
rect 172664 137216 172716 137268
rect 174044 137216 174096 137268
rect 62632 137148 62684 137200
rect 66404 137148 66456 137200
rect 135312 137148 135364 137200
rect 136876 137148 136928 137200
rect 172204 137148 172256 137200
rect 173952 137148 174004 137200
rect 100628 137012 100680 137064
rect 102836 137012 102888 137064
rect 100536 136672 100588 136724
rect 102468 136672 102520 136724
rect 172572 136128 172624 136180
rect 174136 136128 174188 136180
rect 100628 135992 100680 136044
rect 102192 135992 102244 136044
rect 172664 135992 172716 136044
rect 174504 135992 174556 136044
rect 62908 135856 62960 135908
rect 66036 135856 66088 135908
rect 100904 135856 100956 135908
rect 102100 135856 102152 135908
rect 134944 135856 134996 135908
rect 136968 135856 137020 135908
rect 63000 135788 63052 135840
rect 66404 135788 66456 135840
rect 135128 135788 135180 135840
rect 136876 135788 136928 135840
rect 172020 135788 172072 135840
rect 174320 135788 174372 135840
rect 100720 135720 100772 135772
rect 102376 135720 102428 135772
rect 100996 135652 101048 135704
rect 102468 135652 102520 135704
rect 100352 135584 100404 135636
rect 102652 135584 102704 135636
rect 62724 134972 62776 135024
rect 65024 134972 65076 135024
rect 135036 134904 135088 134956
rect 136784 134904 136836 134956
rect 62816 134632 62868 134684
rect 66312 134632 66364 134684
rect 100076 134632 100128 134684
rect 102284 134632 102336 134684
rect 171836 134632 171888 134684
rect 174228 134632 174280 134684
rect 135220 134496 135272 134548
rect 136968 134496 137020 134548
rect 172664 134496 172716 134548
rect 174320 134496 174372 134548
rect 62724 134428 62776 134480
rect 66404 134428 66456 134480
rect 132920 134428 132972 134480
rect 135404 134428 135456 134480
rect 136876 134428 136928 134480
rect 172204 133544 172256 133596
rect 175332 133544 175384 133596
rect 100904 133136 100956 133188
rect 102192 133136 102244 133188
rect 63552 133068 63604 133120
rect 66404 133068 66456 133120
rect 135128 133068 135180 133120
rect 136968 133068 137020 133120
rect 172664 133068 172716 133120
rect 174872 133068 174924 133120
rect 63644 133000 63696 133052
rect 65852 133000 65904 133052
rect 100076 133000 100128 133052
rect 102100 133000 102152 133052
rect 135312 133000 135364 133052
rect 136876 133000 136928 133052
rect 100996 132932 101048 132984
rect 102376 132932 102428 132984
rect 172388 131912 172440 131964
rect 175424 131912 175476 131964
rect 172664 131776 172716 131828
rect 175148 131776 175200 131828
rect 63276 131708 63328 131760
rect 65668 131708 65720 131760
rect 100904 131708 100956 131760
rect 102008 131708 102060 131760
rect 134944 131708 134996 131760
rect 136968 131708 137020 131760
rect 172020 131708 172072 131760
rect 175240 131708 175292 131760
rect 63460 131640 63512 131692
rect 66404 131640 66456 131692
rect 100444 131640 100496 131692
rect 135220 131640 135272 131692
rect 136876 131640 136928 131692
rect 102376 131572 102428 131624
rect 135312 131028 135364 131080
rect 136784 131028 136836 131080
rect 62816 130756 62868 130808
rect 65024 130756 65076 130808
rect 100444 130552 100496 130604
rect 102284 130552 102336 130604
rect 172664 130552 172716 130604
rect 174228 130552 174280 130604
rect 62632 130348 62684 130400
rect 66404 130348 66456 130400
rect 100904 130348 100956 130400
rect 102192 130348 102244 130400
rect 135036 130348 135088 130400
rect 136968 130348 137020 130400
rect 62724 130280 62776 130332
rect 66312 130280 66364 130332
rect 135404 130280 135456 130332
rect 136876 130280 136928 130332
rect 172664 130280 172716 130332
rect 174320 130280 174372 130332
rect 100996 130212 101048 130264
rect 102376 130212 102428 130264
rect 171836 129328 171888 129380
rect 174136 129328 174188 129380
rect 171836 129056 171888 129108
rect 174504 129056 174556 129108
rect 62908 128988 62960 129040
rect 66404 128988 66456 129040
rect 100904 128988 100956 129040
rect 102008 128988 102060 129040
rect 135128 128988 135180 129040
rect 136968 128988 137020 129040
rect 62816 128920 62868 128972
rect 65484 128920 65536 128972
rect 100076 128920 100128 128972
rect 101916 128920 101968 128972
rect 135312 128920 135364 128972
rect 136876 128920 136928 128972
rect 100352 127832 100404 127884
rect 102284 127832 102336 127884
rect 172572 127832 172624 127884
rect 174228 127832 174280 127884
rect 100536 127560 100588 127612
rect 102008 127560 102060 127612
rect 135220 127560 135272 127612
rect 136876 127560 136928 127612
rect 171560 127560 171612 127612
rect 174596 127560 174648 127612
rect 62632 127492 62684 127544
rect 66404 127492 66456 127544
rect 222804 127492 222856 127544
rect 134668 127152 134720 127204
rect 136784 127152 136836 127204
rect 62816 126880 62868 126932
rect 65024 126880 65076 126932
rect 172204 126472 172256 126524
rect 174320 126472 174372 126524
rect 100812 126268 100864 126320
rect 102100 126268 102152 126320
rect 62724 126200 62776 126252
rect 66312 126200 66364 126252
rect 100904 126200 100956 126252
rect 102284 126200 102336 126252
rect 135036 126200 135088 126252
rect 136968 126200 137020 126252
rect 172664 126200 172716 126252
rect 174504 126200 174556 126252
rect 62908 126132 62960 126184
rect 66404 126132 66456 126184
rect 100444 126132 100496 126184
rect 135312 126132 135364 126184
rect 136876 126132 136928 126184
rect 172020 126132 172072 126184
rect 174136 126132 174188 126184
rect 102376 126064 102428 126116
rect 135404 125656 135456 125708
rect 136784 125656 136836 125708
rect 62816 125520 62868 125572
rect 65024 125520 65076 125572
rect 171836 125248 171888 125300
rect 174228 125248 174280 125300
rect 100812 124840 100864 124892
rect 102192 124840 102244 124892
rect 172204 124840 172256 124892
rect 174596 124840 174648 124892
rect 62632 124772 62684 124824
rect 66404 124772 66456 124824
rect 100904 124772 100956 124824
rect 135128 124772 135180 124824
rect 136876 124772 136928 124824
rect 222712 124815 222764 124824
rect 222712 124781 222721 124815
rect 222721 124781 222755 124815
rect 222755 124781 222764 124815
rect 222712 124772 222764 124781
rect 102376 124704 102428 124756
rect 135220 124228 135272 124280
rect 136784 124228 136836 124280
rect 62816 123752 62868 123804
rect 65024 123752 65076 123804
rect 172572 123480 172624 123532
rect 175332 123480 175384 123532
rect 63552 123344 63604 123396
rect 66404 123344 66456 123396
rect 100260 123344 100312 123396
rect 102284 123344 102336 123396
rect 135404 123344 135456 123396
rect 136876 123344 136928 123396
rect 171836 123344 171888 123396
rect 174136 123344 174188 123396
rect 135312 122868 135364 122920
rect 136784 122868 136836 122920
rect 62816 122664 62868 122716
rect 65024 122664 65076 122716
rect 171836 122392 171888 122444
rect 175056 122392 175108 122444
rect 100168 122188 100220 122240
rect 102284 122188 102336 122240
rect 100904 122120 100956 122172
rect 102008 122120 102060 122172
rect 135128 122120 135180 122172
rect 137060 122120 137112 122172
rect 172020 122120 172072 122172
rect 175424 122120 175476 122172
rect 63460 122052 63512 122104
rect 66312 122052 66364 122104
rect 135220 122052 135272 122104
rect 136968 122052 137020 122104
rect 63644 121984 63696 122036
rect 66404 121984 66456 122036
rect 100628 121984 100680 122036
rect 102100 121984 102152 122036
rect 100996 121916 101048 121968
rect 102376 121916 102428 121968
rect 135312 121916 135364 121968
rect 136876 121984 136928 122036
rect 172664 121984 172716 122036
rect 175148 121984 175200 122036
rect 62816 121440 62868 121492
rect 65024 121440 65076 121492
rect 100904 120896 100956 120948
rect 102192 120896 102244 120948
rect 172112 120896 172164 120948
rect 174320 120896 174372 120948
rect 172664 120760 172716 120812
rect 174228 120760 174280 120812
rect 100076 120624 100128 120676
rect 102376 120556 102428 120608
rect 134852 120216 134904 120268
rect 136784 120216 136836 120268
rect 62816 119944 62868 119996
rect 65024 119944 65076 119996
rect 171836 119672 171888 119724
rect 174136 119672 174188 119724
rect 171836 119400 171888 119452
rect 174504 119400 174556 119452
rect 62908 119264 62960 119316
rect 65484 119264 65536 119316
rect 100444 119264 100496 119316
rect 102284 119264 102336 119316
rect 135220 119264 135272 119316
rect 136876 119264 136928 119316
rect 62724 119128 62776 119180
rect 66220 119128 66272 119180
rect 135312 119128 135364 119180
rect 136968 119128 137020 119180
rect 62816 118720 62868 118772
rect 65024 118720 65076 118772
rect 135312 118516 135364 118568
rect 136784 118516 136836 118568
rect 171652 118176 171704 118228
rect 173952 118176 174004 118228
rect 100628 118108 100680 118160
rect 102284 118108 102336 118160
rect 172664 118040 172716 118092
rect 174320 118040 174372 118092
rect 135128 117904 135180 117956
rect 136876 117904 136928 117956
rect 62724 117836 62776 117888
rect 66404 117836 66456 117888
rect 100260 117836 100312 117888
rect 132920 117836 132972 117888
rect 102468 117768 102520 117820
rect 132644 117811 132696 117820
rect 132644 117777 132653 117811
rect 132653 117777 132687 117811
rect 132687 117777 132696 117811
rect 132644 117768 132696 117777
rect 100996 117700 101048 117752
rect 102376 117700 102428 117752
rect 132644 117632 132696 117684
rect 134116 117768 134168 117820
rect 136968 117836 137020 117888
rect 171836 117836 171888 117888
rect 174044 117836 174096 117888
rect 62816 117292 62868 117344
rect 65024 117292 65076 117344
rect 62816 117156 62868 117208
rect 64932 117156 64984 117208
rect 134668 117156 134720 117208
rect 136784 117156 136836 117208
rect 100260 116680 100312 116732
rect 102192 116680 102244 116732
rect 172664 116544 172716 116596
rect 174136 116544 174188 116596
rect 100904 116476 100956 116528
rect 135312 116476 135364 116528
rect 136876 116476 136928 116528
rect 172572 116476 172624 116528
rect 174228 116476 174280 116528
rect 102376 116408 102428 116460
rect 100536 116340 100588 116392
rect 102652 116340 102704 116392
rect 62816 115728 62868 115780
rect 65024 115728 65076 115780
rect 134852 115592 134904 115644
rect 136784 115592 136836 115644
rect 171836 115592 171888 115644
rect 174044 115592 174096 115644
rect 100904 115456 100956 115508
rect 102284 115456 102336 115508
rect 222620 115048 222672 115100
rect 222988 115048 223040 115100
rect 62816 114844 62868 114896
rect 66404 114844 66456 114896
rect 62816 114572 62868 114624
rect 65024 114572 65076 114624
rect 134852 114436 134904 114488
rect 136784 114436 136836 114488
rect 30432 114300 30484 114352
rect 92716 114300 92768 114352
rect 113508 113620 113560 113672
rect 114382 113620 114434 113672
rect 132092 113620 132144 113672
rect 144880 113620 144932 113672
rect 204680 113620 204732 113672
rect 154816 113552 154868 113604
rect 207256 113552 207308 113604
rect 194652 113144 194704 113196
rect 198240 113144 198292 113196
rect 189408 113076 189460 113128
rect 190236 113076 190288 113128
rect 191340 113076 191392 113128
rect 193088 113076 193140 113128
rect 193732 113076 193784 113128
rect 196124 113076 196176 113128
rect 198516 113076 198568 113128
rect 203392 113076 203444 113128
rect 195756 113008 195808 113060
rect 199344 113008 199396 113060
rect 72016 112940 72068 112992
rect 72844 112940 72896 112992
rect 103664 112940 103716 112992
rect 132644 112940 132696 112992
rect 164844 112940 164896 112992
rect 198884 112940 198936 112992
rect 203944 112940 203996 112992
rect 196124 112872 196176 112924
rect 199988 112872 200040 112924
rect 81676 112736 81728 112788
rect 82504 112736 82556 112788
rect 194560 112736 194612 112788
rect 197688 112736 197740 112788
rect 197320 112600 197372 112652
rect 201644 112600 201696 112652
rect 190512 112532 190564 112584
rect 191984 112532 192036 112584
rect 192536 112532 192588 112584
rect 194744 112532 194796 112584
rect 196492 112532 196544 112584
rect 200540 112532 200592 112584
rect 190144 112464 190196 112516
rect 191432 112464 191484 112516
rect 196952 112464 197004 112516
rect 201092 112464 201144 112516
rect 189684 112396 189736 112448
rect 190788 112396 190840 112448
rect 192904 112396 192956 112448
rect 193180 112328 193232 112380
rect 194192 112328 194244 112380
rect 103664 112260 103716 112312
rect 109460 112260 109512 112312
rect 132092 112260 132144 112312
rect 197504 112396 197556 112448
rect 201644 112396 201696 112448
rect 198148 112328 198200 112380
rect 202840 112328 202892 112380
rect 195388 112260 195440 112312
rect 110012 112192 110064 112244
rect 132644 112192 132696 112244
rect 194192 112192 194244 112244
rect 195940 112192 195992 112244
rect 52604 112124 52656 112176
rect 57020 112124 57072 112176
rect 81676 112124 81728 112176
rect 110472 112124 110524 112176
rect 121052 112124 121104 112176
rect 124732 112124 124784 112176
rect 51040 112056 51092 112108
rect 54260 112056 54312 112108
rect 190604 112056 190656 112108
rect 192260 112056 192312 112108
rect 53064 111988 53116 112040
rect 57664 111988 57716 112040
rect 51868 111920 51920 111972
rect 55640 111920 55692 111972
rect 122248 111920 122300 111972
rect 126388 111920 126440 111972
rect 35216 111852 35268 111904
rect 39816 111852 39868 111904
rect 52512 111852 52564 111904
rect 56376 111852 56428 111904
rect 117832 111852 117884 111904
rect 120316 111852 120368 111904
rect 53800 111784 53852 111836
rect 59044 111784 59096 111836
rect 113048 111784 113100 111836
rect 113784 111784 113836 111836
rect 119856 111784 119908 111836
rect 123076 111852 123128 111904
rect 122708 111784 122760 111836
rect 126940 111784 126992 111836
rect 34480 111716 34532 111768
rect 39448 111716 39500 111768
rect 54260 111716 54312 111768
rect 59780 111716 59832 111768
rect 120316 111716 120368 111768
rect 123628 111716 123680 111768
rect 35860 111648 35912 111700
rect 40276 111648 40328 111700
rect 53432 111648 53484 111700
rect 58400 111648 58452 111700
rect 33836 111580 33888 111632
rect 39080 111580 39132 111632
rect 54628 111580 54680 111632
rect 60424 111580 60476 111632
rect 123076 111580 123128 111632
rect 127492 111580 127544 111632
rect 37884 111512 37936 111564
rect 41472 111512 41524 111564
rect 123444 111512 123496 111564
rect 128044 111512 128096 111564
rect 39264 111444 39316 111496
rect 42208 111444 42260 111496
rect 118660 111444 118712 111496
rect 121420 111444 121472 111496
rect 124272 111444 124324 111496
rect 129148 111444 129200 111496
rect 40000 111376 40052 111428
rect 42300 111376 42352 111428
rect 48280 111376 48332 111428
rect 49476 111376 49528 111428
rect 50672 111376 50724 111428
rect 53616 111376 53668 111428
rect 114244 111376 114296 111428
rect 115440 111376 115492 111428
rect 116636 111376 116688 111428
rect 118752 111376 118804 111428
rect 121512 111376 121564 111428
rect 125284 111376 125336 111428
rect 40644 111308 40696 111360
rect 43036 111308 43088 111360
rect 43404 111308 43456 111360
rect 44600 111308 44652 111360
rect 47820 111308 47872 111360
rect 48832 111308 48884 111360
rect 49844 111308 49896 111360
rect 52236 111308 52288 111360
rect 113876 111308 113928 111360
rect 114888 111308 114940 111360
rect 116268 111308 116320 111360
rect 118200 111308 118252 111360
rect 118292 111308 118344 111360
rect 120868 111308 120920 111360
rect 121880 111308 121932 111360
rect 125836 111376 125888 111428
rect 126296 111376 126348 111428
rect 131908 111376 131960 111428
rect 182232 111376 182284 111428
rect 183244 111376 183296 111428
rect 191984 111376 192036 111428
rect 194284 111376 194336 111428
rect 195296 111376 195348 111428
rect 198792 111376 198844 111428
rect 125468 111308 125520 111360
rect 130804 111308 130856 111360
rect 182876 111308 182928 111360
rect 183796 111308 183848 111360
rect 191708 111308 191760 111360
rect 193640 111308 193692 111360
rect 194100 111308 194152 111360
rect 197136 111308 197188 111360
rect 37240 111240 37292 111292
rect 41012 111240 41064 111292
rect 48648 111240 48700 111292
rect 50212 111240 50264 111292
rect 51408 111240 51460 111292
rect 54996 111240 55048 111292
rect 114704 111240 114756 111292
rect 115992 111240 116044 111292
rect 117464 111240 117516 111292
rect 119764 111240 119816 111292
rect 120684 111240 120736 111292
rect 124180 111240 124232 111292
rect 125100 111240 125152 111292
rect 130252 111240 130304 111292
rect 36596 111172 36648 111224
rect 40644 111172 40696 111224
rect 41288 111172 41340 111224
rect 43404 111172 43456 111224
rect 44324 111172 44376 111224
rect 45060 111172 45112 111224
rect 49476 111172 49528 111224
rect 51592 111172 51644 111224
rect 115440 111172 115492 111224
rect 117096 111172 117148 111224
rect 119488 111172 119540 111224
rect 122524 111172 122576 111224
rect 124640 111172 124692 111224
rect 129700 111172 129752 111224
rect 177448 111172 177500 111224
rect 178276 111172 178328 111224
rect 42024 111104 42076 111156
rect 43864 111104 43916 111156
rect 50212 111104 50264 111156
rect 52972 111104 53024 111156
rect 105412 111104 105464 111156
rect 107160 111104 107212 111156
rect 119120 111104 119172 111156
rect 121972 111104 122024 111156
rect 123904 111104 123956 111156
rect 128596 111104 128648 111156
rect 177080 111104 177132 111156
rect 178828 111104 178880 111156
rect 38620 111036 38672 111088
rect 41840 111036 41892 111088
rect 49016 111036 49068 111088
rect 50856 111036 50908 111088
rect 105688 111036 105740 111088
rect 107712 111036 107764 111088
rect 115900 111036 115952 111088
rect 117648 111036 117700 111088
rect 126664 111036 126716 111088
rect 132184 111036 132236 111088
rect 176988 111036 177040 111088
rect 179380 111036 179432 111088
rect 42668 110968 42720 111020
rect 44232 110968 44284 111020
rect 105228 110968 105280 111020
rect 106608 110968 106660 111020
rect 105780 110900 105832 110952
rect 108816 110968 108868 111020
rect 115072 110968 115124 111020
rect 116544 110968 116596 111020
rect 117096 110968 117148 111020
rect 119212 110968 119264 111020
rect 125836 110968 125888 111020
rect 131356 110968 131408 111020
rect 177264 110968 177316 111020
rect 180024 110968 180076 111020
rect 181680 110968 181732 111020
rect 183106 110968 183158 111020
rect 183428 110968 183480 111020
rect 184302 110968 184354 111020
rect 177724 110900 177776 110952
rect 181128 110900 181180 110952
rect 222712 110220 222764 110272
rect 177172 109472 177224 109524
rect 180576 109472 180628 109524
rect 105320 109132 105372 109184
rect 108264 109132 108316 109184
rect 222804 107951 222856 107960
rect 222804 107917 222813 107951
rect 222813 107917 222847 107951
rect 222847 107917 222856 107951
rect 222804 107908 222856 107917
rect 106424 107160 106476 107212
rect 107896 107160 107948 107212
rect 177540 106820 177592 106872
rect 179656 106820 179708 106872
rect 32640 104032 32692 104084
rect 37424 104032 37476 104084
rect 56836 104032 56888 104084
rect 59872 104032 59924 104084
rect 105780 104032 105832 104084
rect 108448 104032 108500 104084
rect 177816 104032 177868 104084
rect 179656 104032 179708 104084
rect 106332 101312 106384 101364
rect 107896 101312 107948 101364
rect 177632 101312 177684 101364
rect 179656 101312 179708 101364
rect 105964 101244 106016 101296
rect 108540 101244 108592 101296
rect 176988 101244 177040 101296
rect 180300 101244 180352 101296
rect 106424 99884 106476 99936
rect 107896 99884 107948 99936
rect 177724 99884 177776 99936
rect 179656 99884 179708 99936
rect 106240 97640 106292 97692
rect 107896 97640 107948 97692
rect 177540 97164 177592 97216
rect 179656 97164 179708 97216
rect 222988 97096 223040 97148
rect 223540 97096 223592 97148
rect 132368 95779 132420 95788
rect 132368 95745 132377 95779
rect 132377 95745 132411 95779
rect 132411 95745 132420 95779
rect 132368 95736 132420 95745
rect 106516 94784 106568 94836
rect 108448 94784 108500 94836
rect 177448 94308 177500 94360
rect 179564 94308 179616 94360
rect 222804 92540 222856 92592
rect 223540 92540 223592 92592
rect 105872 91656 105924 91708
rect 107804 91656 107856 91708
rect 177540 91656 177592 91708
rect 179564 91656 179616 91708
rect 201092 91588 201144 91640
rect 204496 91588 204548 91640
rect 28868 90228 28920 90280
rect 36412 90228 36464 90280
rect 59596 90228 59648 90280
rect 105228 90228 105280 90280
rect 107896 90228 107948 90280
rect 177356 90228 177408 90280
rect 179656 90228 179708 90280
rect 105136 89208 105188 89260
rect 107804 89208 107856 89260
rect 177356 89140 177408 89192
rect 179564 89140 179616 89192
rect 132552 88732 132604 88784
rect 177356 88188 177408 88240
rect 179472 88188 179524 88240
rect 105872 87712 105924 87764
rect 107712 87712 107764 87764
rect 54812 86123 54864 86132
rect 54812 86089 54821 86123
rect 54821 86089 54855 86123
rect 54855 86089 54864 86123
rect 54812 86080 54864 86089
rect 105596 86080 105648 86132
rect 108724 86080 108776 86132
rect 178092 86080 178144 86132
rect 180484 86080 180536 86132
rect 222804 84788 222856 84840
rect 223540 84788 223592 84840
rect 106332 84720 106384 84772
rect 108816 84720 108868 84772
rect 177540 84720 177592 84772
rect 179656 84720 179708 84772
rect 178184 83632 178236 83684
rect 180392 83632 180444 83684
rect 105596 83360 105648 83412
rect 108632 83360 108684 83412
rect 105504 82000 105556 82052
rect 108540 82000 108592 82052
rect 177724 82000 177776 82052
rect 180300 82000 180352 82052
rect 106516 81932 106568 81984
rect 107896 81932 107948 81984
rect 105228 80572 105280 80624
rect 108080 80572 108132 80624
rect 177356 80572 177408 80624
rect 180024 80572 180076 80624
rect 105136 79688 105188 79740
rect 107528 79688 107580 79740
rect 132552 79280 132604 79332
rect 54812 79255 54864 79264
rect 54812 79221 54821 79255
rect 54821 79221 54855 79255
rect 54855 79221 54864 79255
rect 54812 79212 54864 79221
rect 178184 79212 178236 79264
rect 179380 79212 179432 79264
rect 132552 79144 132604 79196
rect 30524 77784 30576 77836
rect 37424 77784 37476 77836
rect 57480 77580 57532 77632
rect 59596 77580 59648 77632
rect 54812 76467 54864 76476
rect 54812 76433 54821 76467
rect 54821 76433 54855 76467
rect 54855 76433 54864 76467
rect 54812 76424 54864 76433
rect 222988 75064 223040 75116
rect 223540 75064 223592 75116
rect 222804 73568 222856 73620
rect 223080 73568 223132 73620
rect 103204 72344 103256 72396
rect 108356 72344 108408 72396
rect 177356 72344 177408 72396
rect 180576 72344 180628 72396
rect 178368 70848 178420 70900
rect 181128 70848 181180 70900
rect 106516 70508 106568 70560
rect 109276 70508 109328 70560
rect 90140 69760 90192 69812
rect 54812 69692 54864 69744
rect 22244 69488 22296 69540
rect 28684 69488 28736 69540
rect 36044 69488 36096 69540
rect 40276 69488 40328 69540
rect 53800 69488 53852 69540
rect 59044 69556 59096 69608
rect 126296 69488 126348 69540
rect 131632 69556 131684 69608
rect 198884 69488 198936 69540
rect 203944 69556 203996 69608
rect 202196 69488 202248 69540
rect 16632 69420 16684 69472
rect 31904 69420 31956 69472
rect 35584 69420 35636 69472
rect 39816 69420 39868 69472
rect 54260 69420 54312 69472
rect 59412 69420 59464 69472
rect 198516 69420 198568 69472
rect 202932 69420 202984 69472
rect 210568 69420 210620 69472
rect 34112 69352 34164 69404
rect 39080 69352 39132 69404
rect 55364 69352 55416 69404
rect 60148 69352 60200 69404
rect 196124 69352 196176 69404
rect 199988 69352 200040 69404
rect 34664 69284 34716 69336
rect 39448 69284 39500 69336
rect 53432 69284 53484 69336
rect 58124 69284 58176 69336
rect 120316 69284 120368 69336
rect 123076 69284 123128 69336
rect 201000 69284 201052 69336
rect 215904 69284 215956 69336
rect 52236 69216 52288 69268
rect 56376 69216 56428 69268
rect 125100 69216 125152 69268
rect 129884 69216 129936 69268
rect 194100 69216 194152 69268
rect 197136 69216 197188 69268
rect 197320 69216 197372 69268
rect 201644 69216 201696 69268
rect 40000 69148 40052 69200
rect 42668 69148 42720 69200
rect 51408 69148 51460 69200
rect 54996 69148 55048 69200
rect 118292 69148 118344 69200
rect 120316 69148 120368 69200
rect 125836 69148 125888 69200
rect 131264 69148 131316 69200
rect 182232 69148 182284 69200
rect 183244 69148 183296 69200
rect 192536 69148 192588 69200
rect 194836 69148 194888 69200
rect 197412 69148 197464 69200
rect 201828 69148 201880 69200
rect 36596 69080 36648 69132
rect 40644 69080 40696 69132
rect 41288 69080 41340 69132
rect 43404 69080 43456 69132
rect 49476 69080 49528 69132
rect 51592 69080 51644 69132
rect 51868 69080 51920 69132
rect 55640 69080 55692 69132
rect 117464 69080 117516 69132
rect 119028 69080 119080 69132
rect 122708 69080 122760 69132
rect 126480 69080 126532 69132
rect 126664 69080 126716 69132
rect 132184 69080 132236 69132
rect 181680 69080 181732 69132
rect 182784 69080 182836 69132
rect 189684 69080 189736 69132
rect 190696 69080 190748 69132
rect 191800 69080 191852 69132
rect 194284 69080 194336 69132
rect 194560 69080 194612 69132
rect 197688 69080 197740 69132
rect 198148 69080 198200 69132
rect 202840 69080 202892 69132
rect 37240 69012 37292 69064
rect 41012 69012 41064 69064
rect 42668 69012 42720 69064
rect 44232 69012 44284 69064
rect 53064 69012 53116 69064
rect 57664 69012 57716 69064
rect 62724 69012 62776 69064
rect 68980 69012 69032 69064
rect 92348 69012 92400 69064
rect 97040 69012 97092 69064
rect 118660 69012 118712 69064
rect 120592 69012 120644 69064
rect 123720 69012 123772 69064
rect 127584 69012 127636 69064
rect 192904 69012 192956 69064
rect 195388 69012 195440 69064
rect 196952 69012 197004 69064
rect 201092 69012 201144 69064
rect 40644 68944 40696 68996
rect 43036 68944 43088 68996
rect 43404 68944 43456 68996
rect 44600 68944 44652 68996
rect 47820 68944 47872 68996
rect 48556 68944 48608 68996
rect 48648 68944 48700 68996
rect 49936 68944 49988 68996
rect 50672 68944 50724 68996
rect 53616 68944 53668 68996
rect 54628 68944 54680 68996
rect 55364 68944 55416 68996
rect 88944 68944 88996 68996
rect 96856 68944 96908 68996
rect 125468 68944 125520 68996
rect 130436 68944 130488 68996
rect 158772 68944 158824 68996
rect 165120 68944 165172 68996
rect 193364 68944 193416 68996
rect 195940 68944 195992 68996
rect 196492 68944 196544 68996
rect 200540 68944 200592 68996
rect 42024 68876 42076 68928
rect 43864 68876 43916 68928
rect 52604 68876 52656 68928
rect 56744 68876 56796 68928
rect 62908 68876 62960 68928
rect 67876 68876 67928 68928
rect 83424 68876 83476 68928
rect 87196 68876 87248 68928
rect 87840 68876 87892 68928
rect 94740 68876 94792 68928
rect 124272 68876 124324 68928
rect 128688 68876 128740 68928
rect 151044 68876 151096 68928
rect 152056 68876 152108 68928
rect 159876 68876 159928 68928
rect 167052 68876 167104 68928
rect 168800 68876 168852 68928
rect 173860 68876 173912 68928
rect 190604 68876 190656 68928
rect 192536 68876 192588 68928
rect 195756 68876 195808 68928
rect 199344 68876 199396 68928
rect 31904 68808 31956 68860
rect 39264 68808 39316 68860
rect 42208 68808 42260 68860
rect 51040 68808 51092 68860
rect 54260 68808 54312 68860
rect 62816 68808 62868 68860
rect 70084 68808 70136 68860
rect 82320 68808 82372 68860
rect 85356 68808 85408 68860
rect 93452 68808 93504 68860
rect 102836 68808 102888 68860
rect 122248 68808 122300 68860
rect 125836 68808 125888 68860
rect 140832 68808 140884 68860
rect 144328 68808 144380 68860
rect 160980 68808 161032 68860
rect 168892 68808 168944 68860
rect 169904 68808 169956 68860
rect 173952 68808 174004 68860
rect 193732 68808 193784 68860
rect 196492 68808 196544 68860
rect 205140 68808 205192 68860
rect 221240 68808 221292 68860
rect 27580 68740 27632 68792
rect 50212 68740 50264 68792
rect 52972 68740 53024 68792
rect 121880 68740 121932 68792
rect 125192 68740 125244 68792
rect 195296 68740 195348 68792
rect 198792 68740 198844 68792
rect 37884 68536 37936 68588
rect 41472 68536 41524 68588
rect 102284 68672 102336 68724
rect 174320 68672 174372 68724
rect 101180 68604 101232 68656
rect 173216 68604 173268 68656
rect 194652 68604 194704 68656
rect 198240 68604 198292 68656
rect 57480 68536 57532 68588
rect 120684 68536 120736 68588
rect 123444 68536 123496 68588
rect 125008 68536 125060 68588
rect 129332 68536 129384 68588
rect 191708 68536 191760 68588
rect 193640 68536 193692 68588
rect 38620 68468 38672 68520
rect 41840 68468 41892 68520
rect 110564 68468 110616 68520
rect 111484 68468 111536 68520
rect 116636 68468 116688 68520
rect 117648 68468 117700 68520
rect 119488 68468 119540 68520
rect 121696 68468 121748 68520
rect 123904 68468 123956 68520
rect 128136 68468 128188 68520
rect 49844 68400 49896 68452
rect 52236 68400 52288 68452
rect 74592 68400 74644 68452
rect 75604 68400 75656 68452
rect 94556 68400 94608 68452
rect 102744 68400 102796 68452
rect 110104 68400 110156 68452
rect 111116 68400 111168 68452
rect 116268 68400 116320 68452
rect 117096 68400 117148 68452
rect 182876 68400 182928 68452
rect 183612 68400 183664 68452
rect 86736 68332 86788 68384
rect 92808 68332 92860 68384
rect 97868 68332 97920 68384
rect 102560 68332 102612 68384
rect 119856 68332 119908 68384
rect 122340 68332 122392 68384
rect 123352 68332 123404 68384
rect 127308 68332 127360 68384
rect 155460 68332 155512 68384
rect 159508 68332 159560 68384
rect 63000 68264 63052 68316
rect 64564 68264 64616 68316
rect 62356 68196 62408 68248
rect 63460 68196 63512 68248
rect 63368 68128 63420 68180
rect 70820 68264 70872 68316
rect 71004 68264 71056 68316
rect 73396 68264 73448 68316
rect 81216 68264 81268 68316
rect 83516 68264 83568 68316
rect 85632 68264 85684 68316
rect 90968 68264 91020 68316
rect 95660 68264 95712 68316
rect 102652 68264 102704 68316
rect 121512 68264 121564 68316
rect 124640 68264 124692 68316
rect 132552 68264 132604 68316
rect 144512 68264 144564 68316
rect 146536 68264 146588 68316
rect 153252 68264 153304 68316
rect 155828 68264 155880 68316
rect 156564 68264 156616 68316
rect 161440 68264 161492 68316
rect 69164 68196 69216 68248
rect 72292 68196 72344 68248
rect 72844 68196 72896 68248
rect 74500 68196 74552 68248
rect 80112 68196 80164 68248
rect 81676 68196 81728 68248
rect 84528 68196 84580 68248
rect 89128 68196 89180 68248
rect 98972 68196 99024 68248
rect 100352 68196 100404 68248
rect 121052 68196 121104 68248
rect 124456 68196 124508 68248
rect 134484 68196 134536 68248
rect 136600 68196 136652 68248
rect 142672 68196 142724 68248
rect 145432 68196 145484 68248
rect 146444 68196 146496 68248
rect 147640 68196 147692 68248
rect 152148 68196 152200 68248
rect 153896 68196 153948 68248
rect 154356 68196 154408 68248
rect 157668 68196 157720 68248
rect 157944 68196 157996 68248
rect 163280 68264 163332 68316
rect 165488 68264 165540 68316
rect 167144 68264 167196 68316
rect 167696 68264 167748 68316
rect 169536 68264 169588 68316
rect 171008 68264 171060 68316
rect 174044 68264 174096 68316
rect 164384 68196 164436 68248
rect 169260 68196 169312 68248
rect 172112 68196 172164 68248
rect 135312 68128 135364 68180
rect 143224 68128 143276 68180
rect 174688 68128 174740 68180
rect 100076 68060 100128 68112
rect 102468 68060 102520 68112
rect 135036 68060 135088 68112
rect 142120 68060 142172 68112
rect 100352 67516 100404 67568
rect 102376 67516 102428 67568
rect 134668 66700 134720 66752
rect 139544 66700 139596 66752
rect 135312 66428 135364 66480
rect 141016 66428 141068 66480
rect 96764 65952 96816 66004
rect 102376 65952 102428 66004
rect 63276 65544 63328 65596
rect 66404 65544 66456 65596
rect 166592 65544 166644 65596
rect 167144 65544 167196 65596
rect 100904 65408 100956 65460
rect 102560 65408 102612 65460
rect 134668 65408 134720 65460
rect 136876 65408 136928 65460
rect 62816 65340 62868 65392
rect 66312 65340 66364 65392
rect 135036 65340 135088 65392
rect 137704 65340 137756 65392
rect 62724 65272 62776 65324
rect 65668 65272 65720 65324
rect 174228 65340 174280 65392
rect 174136 65272 174188 65324
rect 135312 65204 135364 65256
rect 138164 65204 138216 65256
rect 63552 64320 63604 64372
rect 66404 64320 66456 64372
rect 100628 64320 100680 64372
rect 102468 64320 102520 64372
rect 63460 64184 63512 64236
rect 66404 64184 66456 64236
rect 135404 64116 135456 64168
rect 136968 64116 137020 64168
rect 100904 64048 100956 64100
rect 102652 64048 102704 64100
rect 135036 64048 135088 64100
rect 136876 64048 136928 64100
rect 169260 63980 169312 64032
rect 174136 63980 174188 64032
rect 97040 63776 97092 63828
rect 102376 63776 102428 63828
rect 171836 63708 171888 63760
rect 174228 63708 174280 63760
rect 172020 63232 172072 63284
rect 173860 63232 173912 63284
rect 62816 62960 62868 63012
rect 66404 62960 66456 63012
rect 100444 62960 100496 63012
rect 102376 62960 102428 63012
rect 63184 62688 63236 62740
rect 66312 62688 66364 62740
rect 100904 62688 100956 62740
rect 102560 62688 102612 62740
rect 134484 62688 134536 62740
rect 136968 62688 137020 62740
rect 13320 62620 13372 62672
rect 29236 62620 29288 62672
rect 135312 62620 135364 62672
rect 136876 62620 136928 62672
rect 171652 62552 171704 62604
rect 174320 62552 174372 62604
rect 171744 62484 171796 62536
rect 174136 62484 174188 62536
rect 171652 62008 171704 62060
rect 174044 62008 174096 62060
rect 62724 61736 62776 61788
rect 66404 61736 66456 61788
rect 63736 61464 63788 61516
rect 66312 61464 66364 61516
rect 100904 61328 100956 61380
rect 102744 61328 102796 61380
rect 172664 61328 172716 61380
rect 173952 61328 174004 61380
rect 100260 61260 100312 61312
rect 102468 61260 102520 61312
rect 135220 61260 135272 61312
rect 136876 61260 136928 61312
rect 172756 61192 172808 61244
rect 174136 61192 174188 61244
rect 134852 60920 134904 60972
rect 136784 60920 136836 60972
rect 100628 60308 100680 60360
rect 102652 60308 102704 60360
rect 100904 60172 100956 60224
rect 102376 60172 102428 60224
rect 62632 60104 62684 60156
rect 66404 60104 66456 60156
rect 134484 60036 134536 60088
rect 136968 60036 137020 60088
rect 62816 59968 62868 60020
rect 66312 59968 66364 60020
rect 99708 59968 99760 60020
rect 102560 59968 102612 60020
rect 172664 59968 172716 60020
rect 173768 59968 173820 60020
rect 63736 59900 63788 59952
rect 66220 59900 66272 59952
rect 135404 59900 135456 59952
rect 136876 59900 136928 59952
rect 172204 59900 172256 59952
rect 174044 59900 174096 59952
rect 134392 59832 134444 59884
rect 136784 59832 136836 59884
rect 172664 58812 172716 58864
rect 174044 58812 174096 58864
rect 100628 58744 100680 58796
rect 102468 58744 102520 58796
rect 62908 58608 62960 58660
rect 66404 58608 66456 58660
rect 100628 58608 100680 58660
rect 102652 58608 102704 58660
rect 172664 58608 172716 58660
rect 173860 58608 173912 58660
rect 63552 58540 63604 58592
rect 66312 58540 66364 58592
rect 135220 58540 135272 58592
rect 136876 58540 136928 58592
rect 172756 58472 172808 58524
rect 174136 58472 174188 58524
rect 135036 58404 135088 58456
rect 136784 58404 136836 58456
rect 62816 57384 62868 57436
rect 66404 57384 66456 57436
rect 100628 57384 100680 57436
rect 102376 57384 102428 57436
rect 172664 57248 172716 57300
rect 173952 57248 174004 57300
rect 100628 57180 100680 57232
rect 102468 57180 102520 57232
rect 135404 57180 135456 57232
rect 136968 57180 137020 57232
rect 172572 57180 172624 57232
rect 173768 57180 173820 57232
rect 62724 57112 62776 57164
rect 66404 57112 66456 57164
rect 100536 57112 100588 57164
rect 102560 57112 102612 57164
rect 135312 57112 135364 57164
rect 136876 57112 136928 57164
rect 172112 57112 172164 57164
rect 174044 57112 174096 57164
rect 134576 57044 134628 57096
rect 136784 57044 136836 57096
rect 62632 56976 62684 57028
rect 65024 56976 65076 57028
rect 172664 56024 172716 56076
rect 174044 56024 174096 56076
rect 63276 55888 63328 55940
rect 66404 55888 66456 55940
rect 100628 55888 100680 55940
rect 102376 55888 102428 55940
rect 63552 55752 63604 55804
rect 66312 55752 66364 55804
rect 100904 55752 100956 55804
rect 102652 55752 102704 55804
rect 134300 55752 134352 55804
rect 136876 55752 136928 55804
rect 135036 55412 135088 55464
rect 136784 55412 136836 55464
rect 100628 54800 100680 54852
rect 102468 54800 102520 54852
rect 63368 54664 63420 54716
rect 66404 54664 66456 54716
rect 100812 54528 100864 54580
rect 102560 54528 102612 54580
rect 134208 54528 134260 54580
rect 137152 54528 137204 54580
rect 63460 54392 63512 54444
rect 66312 54392 66364 54444
rect 171744 54392 171796 54444
rect 174228 54324 174280 54376
rect 172940 54052 172992 54104
rect 174136 54052 174188 54104
rect 135128 53916 135180 53968
rect 136784 53916 136836 53968
rect 62816 53304 62868 53356
rect 66404 53304 66456 53356
rect 100628 53236 100680 53288
rect 102744 53236 102796 53288
rect 172572 53168 172624 53220
rect 174044 53168 174096 53220
rect 100628 53032 100680 53084
rect 102376 53032 102428 53084
rect 172664 53032 172716 53084
rect 173860 53032 173912 53084
rect 63736 52964 63788 53016
rect 66312 52964 66364 53016
rect 135404 52964 135456 53016
rect 136876 52964 136928 53016
rect 172848 52896 172900 52948
rect 174136 52896 174188 52948
rect 135036 52828 135088 52880
rect 136784 52828 136836 52880
rect 100628 52216 100680 52268
rect 102652 52216 102704 52268
rect 62908 52080 62960 52132
rect 66404 52080 66456 52132
rect 172664 51808 172716 51860
rect 173952 51808 174004 51860
rect 62724 51672 62776 51724
rect 66404 51672 66456 51724
rect 100628 51672 100680 51724
rect 102468 51672 102520 51724
rect 172664 51672 172716 51724
rect 173768 51672 173820 51724
rect 63736 51604 63788 51656
rect 65668 51604 65720 51656
rect 100536 51604 100588 51656
rect 102560 51604 102612 51656
rect 135312 51604 135364 51656
rect 136876 51604 136928 51656
rect 172020 51604 172072 51656
rect 174044 51604 174096 51656
rect 135036 51332 135088 51384
rect 136784 51332 136836 51384
rect 135404 51060 135456 51112
rect 136692 51060 136744 51112
rect 63828 50584 63880 50636
rect 66404 50584 66456 50636
rect 171652 50584 171704 50636
rect 174044 50584 174096 50636
rect 62816 50448 62868 50500
rect 66404 50448 66456 50500
rect 100628 50448 100680 50500
rect 102652 50448 102704 50500
rect 100628 50312 100680 50364
rect 102376 50312 102428 50364
rect 135404 50244 135456 50296
rect 136876 50244 136928 50296
rect 134852 50176 134904 50228
rect 136784 50176 136836 50228
rect 100628 49224 100680 49276
rect 102468 49224 102520 49276
rect 63736 48952 63788 49004
rect 65484 48952 65536 49004
rect 100628 48952 100680 49004
rect 102560 48952 102612 49004
rect 172664 48952 172716 49004
rect 173952 48952 174004 49004
rect 62908 48884 62960 48936
rect 66404 48884 66456 48936
rect 135312 48816 135364 48868
rect 136876 48884 136928 48936
rect 171836 48884 171888 48936
rect 174044 48884 174096 48936
rect 172756 48816 172808 48868
rect 174136 48816 174188 48868
rect 134760 48408 134812 48460
rect 136784 48408 136836 48460
rect 100628 47864 100680 47916
rect 102652 47864 102704 47916
rect 100628 47592 100680 47644
rect 102376 47592 102428 47644
rect 172112 47592 172164 47644
rect 174044 47592 174096 47644
rect 172572 47524 172624 47576
rect 173860 47524 173912 47576
rect 62816 47456 62868 47508
rect 66404 47456 66456 47508
rect 100628 47456 100680 47508
rect 102468 47456 102520 47508
rect 135404 47456 135456 47508
rect 136876 47456 136928 47508
rect 172664 47456 172716 47508
rect 174228 47388 174280 47440
rect 134852 47320 134904 47372
rect 136784 47320 136836 47372
rect 62724 47184 62776 47236
rect 65024 47184 65076 47236
rect 62908 47116 62960 47168
rect 64932 47116 64984 47168
rect 135312 47116 135364 47168
rect 136692 47116 136744 47168
rect 63736 46368 63788 46420
rect 66404 46368 66456 46420
rect 172664 46368 172716 46420
rect 174044 46368 174096 46420
rect 100628 46232 100680 46284
rect 102560 46232 102612 46284
rect 100904 46096 100956 46148
rect 102376 46096 102428 46148
rect 134668 46028 134720 46080
rect 136784 46028 136836 46080
rect 100536 45212 100588 45264
rect 102468 45212 102520 45264
rect 99984 44940 100036 44992
rect 102560 44940 102612 44992
rect 63736 44804 63788 44856
rect 66404 44804 66456 44856
rect 63644 44736 63696 44788
rect 65668 44736 65720 44788
rect 171836 44736 171888 44788
rect 62816 44668 62868 44720
rect 65300 44668 65352 44720
rect 135036 44668 135088 44720
rect 137520 44668 137572 44720
rect 172848 44668 172900 44720
rect 174136 44668 174188 44720
rect 174688 44600 174740 44652
rect 135404 44396 135456 44448
rect 136692 44396 136744 44448
rect 135036 44260 135088 44312
rect 136784 44260 136836 44312
rect 172756 44260 172808 44312
rect 174504 44260 174556 44312
rect 99892 44056 99944 44108
rect 102284 44056 102336 44108
rect 63920 43512 63972 43564
rect 66404 43512 66456 43564
rect 171836 43512 171888 43564
rect 174044 43512 174096 43564
rect 63736 43308 63788 43360
rect 65300 43308 65352 43360
rect 100628 43308 100680 43360
rect 102376 43240 102428 43292
rect 134944 43240 134996 43292
rect 136876 43308 136928 43360
rect 172664 43308 172716 43360
rect 174228 43240 174280 43292
rect 135404 43036 135456 43088
rect 136784 43036 136836 43088
rect 63828 42832 63880 42884
rect 66404 42832 66456 42884
rect 100628 42628 100680 42680
rect 102560 42628 102612 42680
rect 172388 42288 172440 42340
rect 173952 42288 174004 42340
rect 100628 42152 100680 42204
rect 102468 42152 102520 42204
rect 100628 42016 100680 42068
rect 102376 42016 102428 42068
rect 172664 42016 172716 42068
rect 174044 42016 174096 42068
rect 63736 41948 63788 42000
rect 66404 41948 66456 42000
rect 135404 41880 135456 41932
rect 136876 41948 136928 42000
rect 172572 41948 172624 42000
rect 174136 41880 174188 41932
rect 135312 41812 135364 41864
rect 136692 41812 136744 41864
rect 134852 41472 134904 41524
rect 136784 41472 136836 41524
rect 62816 40520 62868 40572
rect 65300 40520 65352 40572
rect 71924 39908 71976 39960
rect 82504 39908 82556 39960
rect 143592 39908 143644 39960
rect 154816 39908 154868 39960
rect 66312 39840 66364 39892
rect 86276 39840 86328 39892
rect 138072 39840 138124 39892
rect 158588 39840 158640 39892
rect 62816 39160 62868 39212
rect 72568 39160 72620 39212
rect 93176 39160 93228 39212
rect 102376 39160 102428 39212
rect 134484 39160 134536 39212
rect 144880 39160 144932 39212
rect 164844 39160 164896 39212
rect 174136 39160 174188 39212
rect 79376 37732 79428 37784
rect 127768 37732 127820 37784
rect 151044 37732 151096 37784
rect 200080 37732 200132 37784
rect 222528 37775 222580 37784
rect 222528 37741 222537 37775
rect 222537 37741 222571 37775
rect 222571 37741 222580 37775
rect 222528 37732 222580 37741
rect 190788 37664 190840 37716
rect 205140 37664 205192 37716
rect 30524 33584 30576 33636
rect 66220 33584 66272 33636
rect 118844 33584 118896 33636
rect 136876 33584 136928 33636
rect 222712 28144 222764 28196
rect 77996 12572 78048 12624
rect 79054 12572 79106 12624
rect 86920 11688 86972 11740
rect 132552 11688 132604 11740
rect 166040 11688 166092 11740
rect 214248 11688 214300 11740
rect 94004 11620 94056 11672
rect 187016 11620 187068 11672
rect 23532 10940 23584 10992
rect 71280 10940 71332 10992
rect 105228 10940 105280 10992
rect 151044 10940 151096 10992
rect 50764 10872 50816 10924
rect 143592 10872 143644 10924
rect 158588 10396 158640 10448
rect 159784 10396 159836 10448
<< metal2 >>
rect 23530 246344 23586 246824
rect 50762 246344 50818 246824
rect 77994 246344 78050 246824
rect 105226 246344 105282 246824
rect 132550 246344 132606 246824
rect 159782 246344 159838 246824
rect 187014 246344 187070 246824
rect 214246 246344 214302 246824
rect 23544 244918 23572 246344
rect 23532 244912 23584 244918
rect 23532 244854 23584 244860
rect 50776 244850 50804 246344
rect 70544 244912 70596 244918
rect 70544 244854 70596 244860
rect 50764 244844 50816 244850
rect 50764 244786 50816 244792
rect 70556 242812 70584 244854
rect 78008 242812 78036 246344
rect 105240 244918 105268 246344
rect 105228 244912 105280 244918
rect 105228 244854 105280 244860
rect 85632 242464 85684 242470
rect 85566 242412 85632 242418
rect 85566 242406 85684 242412
rect 85566 242390 85672 242406
rect 93018 242390 93400 242418
rect 93372 242130 93400 242390
rect 132564 242198 132592 246344
rect 149664 244912 149716 244918
rect 149664 244854 149716 244860
rect 142396 244844 142448 244850
rect 142396 244786 142448 244792
rect 142408 242826 142436 244786
rect 149676 242826 149704 244854
rect 159796 244850 159824 246344
rect 157484 244844 157536 244850
rect 157484 244786 157536 244792
rect 159784 244844 159836 244850
rect 159784 244786 159836 244792
rect 157496 242826 157524 244786
rect 142408 242798 142560 242826
rect 149676 242798 150012 242826
rect 157496 242798 157556 242826
rect 165008 242390 165344 242418
rect 165316 242198 165344 242390
rect 132552 242192 132604 242198
rect 132552 242134 132604 242140
rect 165304 242192 165356 242198
rect 165304 242134 165356 242140
rect 187028 242130 187056 246344
rect 214260 242198 214288 246344
rect 214248 242192 214300 242198
rect 214248 242134 214300 242140
rect 93360 242124 93412 242130
rect 93360 242066 93412 242072
rect 187016 242124 187068 242130
rect 187016 242066 187068 242072
rect 98234 238760 98290 238769
rect 98234 238695 98290 238704
rect 169994 238760 170050 238769
rect 169994 238695 170050 238704
rect 71280 217984 71332 217990
rect 71280 217926 71332 217932
rect 46532 217916 46584 217922
rect 46532 217858 46584 217864
rect 37240 217236 37292 217242
rect 37240 217178 37292 217184
rect 37252 215748 37280 217178
rect 46544 215748 46572 217858
rect 55822 217272 55878 217281
rect 71292 217242 71320 217926
rect 55822 217207 55878 217216
rect 71280 217236 71332 217242
rect 55836 215748 55864 217207
rect 71280 217178 71332 217184
rect 62540 215808 62592 215814
rect 62540 215750 62592 215756
rect 62552 215377 62580 215750
rect 62538 215368 62594 215377
rect 62538 215303 62594 215312
rect 62630 214688 62686 214697
rect 62630 214623 62686 214632
rect 62644 214522 62672 214623
rect 62632 214516 62684 214522
rect 62632 214458 62684 214464
rect 65024 214516 65076 214522
rect 65024 214458 65076 214464
rect 10466 214280 10522 214289
rect 10466 214215 10522 214224
rect 10480 213201 10508 214215
rect 63642 214008 63698 214017
rect 63698 213966 63776 213994
rect 63642 213943 63698 213952
rect 62538 213328 62594 213337
rect 62538 213263 62540 213272
rect 62592 213263 62594 213272
rect 62540 213234 62592 213240
rect 10466 213192 10522 213201
rect 10466 213127 10522 213136
rect 63748 213094 63776 213966
rect 65036 213609 65064 214458
rect 71292 213722 71320 217178
rect 71844 215814 71872 218876
rect 79376 217236 79428 217242
rect 79376 217178 79428 217184
rect 71832 215808 71884 215814
rect 71832 215750 71884 215756
rect 79388 213722 79416 217178
rect 81780 216630 81808 218876
rect 81768 216624 81820 216630
rect 81768 216566 81820 216572
rect 91808 216562 91836 218876
rect 98248 217922 98276 238695
rect 98326 230736 98382 230745
rect 98326 230671 98382 230680
rect 98236 217916 98288 217922
rect 98236 217858 98288 217864
rect 94004 216624 94056 216630
rect 94004 216566 94056 216572
rect 91796 216556 91848 216562
rect 91796 216498 91848 216504
rect 86920 216488 86972 216494
rect 86920 216430 86972 216436
rect 86932 213722 86960 216430
rect 71292 213694 71628 213722
rect 79080 213694 79416 213722
rect 86624 213694 86960 213722
rect 94016 213722 94044 216566
rect 98340 216494 98368 230671
rect 168522 230192 168578 230201
rect 168522 230127 168578 230136
rect 168536 229822 168564 230127
rect 167788 229816 167840 229822
rect 167708 229764 167788 229770
rect 167708 229758 167840 229764
rect 168524 229816 168576 229822
rect 168524 229758 168576 229764
rect 167708 229742 167828 229758
rect 98418 222848 98474 222857
rect 98418 222783 98474 222792
rect 98432 217922 98460 222783
rect 167708 218890 167736 229742
rect 143788 218862 143848 218890
rect 153784 218862 154120 218890
rect 163812 218862 164148 218890
rect 143684 217984 143736 217990
rect 143684 217926 143736 217932
rect 98420 217916 98472 217922
rect 98420 217858 98472 217864
rect 109276 217916 109328 217922
rect 109276 217858 109328 217864
rect 118844 217916 118896 217922
rect 118844 217858 118896 217864
rect 109288 217310 109316 217858
rect 109276 217304 109328 217310
rect 109276 217246 109328 217252
rect 102376 216556 102428 216562
rect 102376 216498 102428 216504
rect 98328 216488 98380 216494
rect 98328 216430 98380 216436
rect 102388 215377 102416 216498
rect 109288 215762 109316 217246
rect 118856 215762 118884 217858
rect 143696 217310 143724 217926
rect 143684 217304 143736 217310
rect 143684 217246 143736 217252
rect 127768 217236 127820 217242
rect 127768 217178 127820 217184
rect 109288 215734 109532 215762
rect 118824 215734 118884 215762
rect 127780 215762 127808 217178
rect 135404 215808 135456 215814
rect 127780 215734 128116 215762
rect 135404 215750 135456 215756
rect 135416 215649 135444 215750
rect 135402 215640 135458 215649
rect 135402 215575 135458 215584
rect 102374 215368 102430 215377
rect 102374 215303 102430 215312
rect 102374 214688 102430 214697
rect 100996 214652 101048 214658
rect 102374 214623 102376 214632
rect 100996 214594 101048 214600
rect 102428 214623 102430 214632
rect 135402 214688 135458 214697
rect 135402 214623 135458 214632
rect 102376 214594 102428 214600
rect 94016 213694 94076 213722
rect 65022 213600 65078 213609
rect 65022 213535 65078 213544
rect 101008 213473 101036 214594
rect 135416 214522 135444 214623
rect 135404 214516 135456 214522
rect 135404 214458 135456 214464
rect 136784 214516 136836 214522
rect 136784 214458 136836 214464
rect 102374 214008 102430 214017
rect 102374 213943 102430 213952
rect 135034 214008 135090 214017
rect 135034 213943 135090 213952
rect 100994 213464 101050 213473
rect 100994 213399 101050 213408
rect 102388 213366 102416 213943
rect 135048 213366 135076 213943
rect 136796 213473 136824 214458
rect 143696 213722 143724 217246
rect 143788 215814 143816 218862
rect 154092 216494 154120 218862
rect 158588 216624 158640 216630
rect 158588 216566 158640 216572
rect 154080 216488 154132 216494
rect 154080 216430 154132 216436
rect 151042 215912 151098 215921
rect 151042 215847 151098 215856
rect 143776 215808 143828 215814
rect 143776 215750 143828 215756
rect 143618 213694 143724 213722
rect 151056 213708 151084 215847
rect 158600 213708 158628 216566
rect 164120 216562 164148 218862
rect 167432 218862 167736 218890
rect 167432 218618 167460 218862
rect 167248 218590 167460 218618
rect 167248 216630 167276 218590
rect 170008 217922 170036 238695
rect 223078 234952 223134 234961
rect 223078 234887 223134 234896
rect 223092 223430 223120 234887
rect 207256 223424 207308 223430
rect 207256 223366 207308 223372
rect 223080 223424 223132 223430
rect 223080 223366 223132 223372
rect 170086 222848 170142 222857
rect 207268 222818 207296 223366
rect 170086 222783 170088 222792
rect 170140 222783 170142 222792
rect 207256 222812 207308 222818
rect 170088 222754 170140 222760
rect 207256 222754 207308 222760
rect 170100 217990 170128 222754
rect 170088 217984 170140 217990
rect 170088 217926 170140 217932
rect 169996 217916 170048 217922
rect 169996 217858 170048 217864
rect 167236 216624 167288 216630
rect 167236 216566 167288 216572
rect 164108 216556 164160 216562
rect 164108 216498 164160 216504
rect 174228 216556 174280 216562
rect 174228 216498 174280 216504
rect 166040 216488 166092 216494
rect 166040 216430 166092 216436
rect 166052 213708 166080 216430
rect 174240 215785 174268 216498
rect 174226 215776 174282 215785
rect 174226 215711 174282 215720
rect 174042 214688 174098 214697
rect 174042 214623 174098 214632
rect 174056 214046 174084 214623
rect 171836 214040 171888 214046
rect 171834 214008 171836 214017
rect 174044 214040 174096 214046
rect 171888 214008 171890 214017
rect 174044 213982 174096 213988
rect 174226 214008 174282 214017
rect 171834 213943 171890 213952
rect 174226 213943 174282 213952
rect 136782 213464 136838 213473
rect 136782 213399 136838 213408
rect 100996 213360 101048 213366
rect 100996 213302 101048 213308
rect 102376 213360 102428 213366
rect 135036 213360 135088 213366
rect 102376 213302 102428 213308
rect 102466 213328 102522 213337
rect 65024 213292 65076 213298
rect 65024 213234 65076 213240
rect 63736 213088 63788 213094
rect 63736 213030 63788 213036
rect 62354 212648 62410 212657
rect 62354 212583 62410 212592
rect 62368 211734 62396 212583
rect 65036 212249 65064 213234
rect 66220 213088 66272 213094
rect 66220 213030 66272 213036
rect 100536 213088 100588 213094
rect 100536 213030 100588 213036
rect 66232 212929 66260 213030
rect 66218 212920 66274 212929
rect 66218 212855 66274 212864
rect 100548 212249 100576 213030
rect 101008 212929 101036 213302
rect 136784 213360 136836 213366
rect 135036 213302 135088 213308
rect 135402 213328 135458 213337
rect 102466 213263 102522 213272
rect 136784 213302 136836 213308
rect 174042 213328 174098 213337
rect 135402 213263 135458 213272
rect 102480 213162 102508 213263
rect 135416 213162 135444 213263
rect 102468 213156 102520 213162
rect 102468 213098 102520 213104
rect 135404 213156 135456 213162
rect 135404 213098 135456 213104
rect 136796 212929 136824 213302
rect 174042 213263 174098 213272
rect 136876 213088 136928 213094
rect 172664 213088 172716 213094
rect 136876 213030 136928 213036
rect 172662 213056 172664 213065
rect 172716 213056 172718 213065
rect 100994 212920 101050 212929
rect 100994 212855 101050 212864
rect 136782 212920 136838 212929
rect 136782 212855 136838 212864
rect 102374 212648 102430 212657
rect 102374 212583 102430 212592
rect 134666 212648 134722 212657
rect 134666 212583 134722 212592
rect 102388 212278 102416 212583
rect 101088 212272 101140 212278
rect 65022 212240 65078 212249
rect 65022 212175 65078 212184
rect 100534 212240 100590 212249
rect 101088 212214 101140 212220
rect 102376 212272 102428 212278
rect 102376 212214 102428 212220
rect 100534 212175 100590 212184
rect 62630 211968 62686 211977
rect 62630 211903 62686 211912
rect 100996 211932 101048 211938
rect 62644 211802 62672 211903
rect 100996 211874 101048 211880
rect 62632 211796 62684 211802
rect 62632 211738 62684 211744
rect 65024 211796 65076 211802
rect 65024 211738 65076 211744
rect 62356 211728 62408 211734
rect 62356 211670 62408 211676
rect 64932 211728 64984 211734
rect 64932 211670 64984 211676
rect 62630 211288 62686 211297
rect 62630 211223 62686 211232
rect 62644 211122 62672 211223
rect 62632 211116 62684 211122
rect 62632 211058 62684 211064
rect 64944 210753 64972 211670
rect 65036 211161 65064 211738
rect 66402 211696 66458 211705
rect 66402 211631 66458 211640
rect 65022 211152 65078 211161
rect 65022 211087 65078 211096
rect 65484 211116 65536 211122
rect 65484 211058 65536 211064
rect 64930 210744 64986 210753
rect 64930 210679 64986 210688
rect 62630 210608 62686 210617
rect 62630 210543 62686 210552
rect 62644 210442 62672 210543
rect 65496 210481 65524 211058
rect 66416 210753 66444 211631
rect 101008 211161 101036 211874
rect 101100 211705 101128 212214
rect 134680 212142 134708 212583
rect 136888 212249 136916 213030
rect 171744 213020 171796 213026
rect 174056 213026 174084 213263
rect 174240 213162 174268 213943
rect 174228 213156 174280 213162
rect 174228 213098 174280 213104
rect 172662 212991 172718 213000
rect 174044 213020 174096 213026
rect 171744 212962 171796 212968
rect 174044 212962 174096 212968
rect 171756 212657 171784 212962
rect 171742 212648 171798 212657
rect 171742 212583 171798 212592
rect 174226 212648 174282 212657
rect 174226 212583 174282 212592
rect 136874 212240 136930 212249
rect 136874 212175 136930 212184
rect 134668 212136 134720 212142
rect 134668 212078 134720 212084
rect 136968 212136 137020 212142
rect 136968 212078 137020 212084
rect 102374 211968 102430 211977
rect 102374 211903 102376 211912
rect 102428 211903 102430 211912
rect 134298 211968 134354 211977
rect 134298 211903 134354 211912
rect 102376 211874 102428 211880
rect 134312 211802 134340 211903
rect 134300 211796 134352 211802
rect 134300 211738 134352 211744
rect 136876 211796 136928 211802
rect 136876 211738 136928 211744
rect 101086 211696 101142 211705
rect 101086 211631 101142 211640
rect 136888 211161 136916 211738
rect 136980 211705 137008 212078
rect 174042 211968 174098 211977
rect 174042 211903 174098 211912
rect 136966 211696 137022 211705
rect 136966 211631 137022 211640
rect 172664 211660 172716 211666
rect 172664 211602 172716 211608
rect 172676 211569 172704 211602
rect 172662 211560 172718 211569
rect 172662 211495 172718 211504
rect 174056 211462 174084 211903
rect 174240 211734 174268 212583
rect 174228 211728 174280 211734
rect 174228 211670 174280 211676
rect 172572 211456 172624 211462
rect 172570 211424 172572 211433
rect 174044 211456 174096 211462
rect 172624 211424 172626 211433
rect 174044 211398 174096 211404
rect 172570 211359 172626 211368
rect 174134 211288 174190 211297
rect 174134 211223 174190 211232
rect 100994 211152 101050 211161
rect 100994 211087 101050 211096
rect 136874 211152 136930 211161
rect 136874 211087 136930 211096
rect 174148 210782 174176 211223
rect 171836 210776 171888 210782
rect 66402 210744 66458 210753
rect 66402 210679 66458 210688
rect 171834 210744 171836 210753
rect 174136 210776 174188 210782
rect 171888 210744 171890 210753
rect 174136 210718 174188 210724
rect 171834 210679 171890 210688
rect 65482 210472 65538 210481
rect 62632 210436 62684 210442
rect 62632 210378 62684 210384
rect 65024 210436 65076 210442
rect 65482 210407 65538 210416
rect 65024 210378 65076 210384
rect 62630 209928 62686 209937
rect 62630 209863 62686 209872
rect 62644 209558 62672 209863
rect 62632 209552 62684 209558
rect 65036 209529 65064 210378
rect 174134 209928 174190 209937
rect 174134 209863 174190 209872
rect 174148 209694 174176 209863
rect 171928 209688 171980 209694
rect 171928 209630 171980 209636
rect 174136 209688 174188 209694
rect 174136 209630 174188 209636
rect 65484 209552 65536 209558
rect 62632 209494 62684 209500
rect 65022 209520 65078 209529
rect 65484 209494 65536 209500
rect 65022 209455 65078 209464
rect 65496 209257 65524 209494
rect 171940 209393 171968 209630
rect 171926 209384 171982 209393
rect 171926 209319 171982 209328
rect 62722 209248 62778 209257
rect 62722 209183 62778 209192
rect 65482 209248 65538 209257
rect 65482 209183 65538 209192
rect 135310 209248 135366 209257
rect 135310 209183 135366 209192
rect 174594 209248 174650 209257
rect 174594 209183 174650 209192
rect 62736 209082 62764 209183
rect 135324 209082 135352 209183
rect 62724 209076 62776 209082
rect 62724 209018 62776 209024
rect 65024 209076 65076 209082
rect 65024 209018 65076 209024
rect 135312 209076 135364 209082
rect 135312 209018 135364 209024
rect 137704 209076 137756 209082
rect 137704 209018 137756 209024
rect 65036 208713 65064 209018
rect 137716 208713 137744 209018
rect 174608 209014 174636 209183
rect 174596 209008 174648 209014
rect 174596 208950 174648 208956
rect 171468 208940 171520 208946
rect 171468 208882 171520 208888
rect 171480 208849 171508 208882
rect 171466 208840 171522 208849
rect 171466 208775 171522 208784
rect 65022 208704 65078 208713
rect 65022 208639 65078 208648
rect 137702 208704 137758 208713
rect 137702 208639 137758 208648
rect 62538 208568 62594 208577
rect 62538 208503 62594 208512
rect 62552 208130 62580 208503
rect 65666 208160 65722 208169
rect 62540 208124 62592 208130
rect 65666 208095 65668 208104
rect 62540 208066 62592 208072
rect 65720 208095 65722 208104
rect 65668 208066 65720 208072
rect 135402 207888 135458 207897
rect 135402 207823 135458 207832
rect 174042 207888 174098 207897
rect 174042 207823 174098 207832
rect 135416 207722 135444 207823
rect 135404 207716 135456 207722
rect 135404 207658 135456 207664
rect 136876 207716 136928 207722
rect 136876 207658 136928 207664
rect 136888 207489 136916 207658
rect 136874 207480 136930 207489
rect 136874 207415 136930 207424
rect 174056 207382 174084 207823
rect 172572 207376 172624 207382
rect 172570 207344 172572 207353
rect 174044 207376 174096 207382
rect 172624 207344 172626 207353
rect 174044 207318 174096 207324
rect 172570 207279 172626 207288
rect 62630 207208 62686 207217
rect 62630 207143 62686 207152
rect 62644 206906 62672 207143
rect 65666 206936 65722 206945
rect 62632 206900 62684 206906
rect 65666 206871 65668 206880
rect 62632 206842 62684 206848
rect 65720 206871 65722 206880
rect 65668 206842 65720 206848
rect 172662 202312 172718 202321
rect 172662 202247 172664 202256
rect 172716 202247 172718 202256
rect 174228 202276 174280 202282
rect 172664 202218 172716 202224
rect 174228 202218 174280 202224
rect 65022 202176 65078 202185
rect 65022 202111 65078 202120
rect 65036 201942 65064 202111
rect 174240 202049 174268 202218
rect 174226 202040 174282 202049
rect 174226 201975 174282 201984
rect 62632 201936 62684 201942
rect 62632 201878 62684 201884
rect 65024 201936 65076 201942
rect 65024 201878 65076 201884
rect 62644 201777 62672 201878
rect 62630 201768 62686 201777
rect 62630 201703 62686 201712
rect 65022 200952 65078 200961
rect 65022 200887 65078 200896
rect 65036 200446 65064 200887
rect 172662 200816 172718 200825
rect 172662 200751 172664 200760
rect 172716 200751 172718 200760
rect 174136 200780 174188 200786
rect 172664 200722 172716 200728
rect 174136 200722 174188 200728
rect 100904 200712 100956 200718
rect 100902 200680 100904 200689
rect 102376 200712 102428 200718
rect 100956 200680 100958 200689
rect 102376 200654 102428 200660
rect 136782 200680 136838 200689
rect 100902 200615 100958 200624
rect 62632 200440 62684 200446
rect 62630 200408 62632 200417
rect 65024 200440 65076 200446
rect 62684 200408 62686 200417
rect 102388 200417 102416 200654
rect 136782 200615 136838 200624
rect 136796 200514 136824 200615
rect 135404 200508 135456 200514
rect 135404 200450 135456 200456
rect 136784 200508 136836 200514
rect 136784 200450 136836 200456
rect 135416 200417 135444 200450
rect 174148 200417 174176 200722
rect 65024 200382 65076 200388
rect 102374 200408 102430 200417
rect 62630 200343 62686 200352
rect 102374 200343 102430 200352
rect 135402 200408 135458 200417
rect 135402 200343 135458 200352
rect 174134 200408 174190 200417
rect 174134 200343 174190 200352
rect 65022 199728 65078 199737
rect 65022 199663 65078 199672
rect 65036 199086 65064 199663
rect 171650 199592 171706 199601
rect 171650 199527 171706 199536
rect 136782 199456 136838 199465
rect 171664 199426 171692 199527
rect 136782 199391 136838 199400
rect 171652 199420 171704 199426
rect 100904 199352 100956 199358
rect 100902 199320 100904 199329
rect 102376 199352 102428 199358
rect 100956 199320 100958 199329
rect 102376 199294 102428 199300
rect 100902 199255 100958 199264
rect 62356 199080 62408 199086
rect 62354 199048 62356 199057
rect 65024 199080 65076 199086
rect 62408 199048 62410 199057
rect 102388 199057 102416 199294
rect 136796 199154 136824 199391
rect 171652 199362 171704 199368
rect 175240 199420 175292 199426
rect 175240 199362 175292 199368
rect 134760 199148 134812 199154
rect 134760 199090 134812 199096
rect 136784 199148 136836 199154
rect 136784 199090 136836 199096
rect 134772 199057 134800 199090
rect 175252 199057 175280 199362
rect 65024 199022 65076 199028
rect 102374 199048 102430 199057
rect 62354 198983 62410 198992
rect 102374 198983 102430 198992
rect 134758 199048 134814 199057
rect 134758 198983 134814 198992
rect 175238 199048 175294 199057
rect 175238 198983 175294 198992
rect 65022 198504 65078 198513
rect 65022 198439 65078 198448
rect 62540 197856 62592 197862
rect 62540 197798 62592 197804
rect 62552 197017 62580 197798
rect 65036 197794 65064 198439
rect 172662 198232 172718 198241
rect 172662 198167 172664 198176
rect 172716 198167 172718 198176
rect 174136 198196 174188 198202
rect 172664 198138 172716 198144
rect 174136 198138 174188 198144
rect 100810 198096 100866 198105
rect 136782 198096 136838 198105
rect 100810 198031 100812 198040
rect 100864 198031 100866 198040
rect 102376 198060 102428 198066
rect 100812 198002 100864 198008
rect 136782 198031 136838 198040
rect 172662 198096 172718 198105
rect 172662 198031 172664 198040
rect 102376 198002 102428 198008
rect 65666 197960 65722 197969
rect 65666 197895 65668 197904
rect 65720 197895 65722 197904
rect 100902 197960 100958 197969
rect 100902 197895 100904 197904
rect 65668 197866 65720 197872
rect 100956 197895 100958 197904
rect 100904 197866 100956 197872
rect 62632 197788 62684 197794
rect 62632 197730 62684 197736
rect 65024 197788 65076 197794
rect 65024 197730 65076 197736
rect 62644 197697 62672 197730
rect 102388 197697 102416 198002
rect 136690 197960 136746 197969
rect 102468 197924 102520 197930
rect 136690 197895 136746 197904
rect 102468 197866 102520 197872
rect 62630 197688 62686 197697
rect 62630 197623 62686 197632
rect 102374 197688 102430 197697
rect 102374 197623 102430 197632
rect 65022 197280 65078 197289
rect 65022 197215 65078 197224
rect 62538 197008 62594 197017
rect 62538 196943 62594 196952
rect 62632 196496 62684 196502
rect 62632 196438 62684 196444
rect 62540 196360 62592 196366
rect 62538 196328 62540 196337
rect 62592 196328 62594 196337
rect 62538 196263 62594 196272
rect 62644 195657 62672 196438
rect 65036 196366 65064 197215
rect 102480 197017 102508 197866
rect 135404 197788 135456 197794
rect 135404 197730 135456 197736
rect 135416 197697 135444 197730
rect 135402 197688 135458 197697
rect 135402 197623 135458 197632
rect 136704 197454 136732 197895
rect 136796 197794 136824 198031
rect 172716 198031 172718 198040
rect 172664 198002 172716 198008
rect 136784 197788 136836 197794
rect 136784 197730 136836 197736
rect 174148 197697 174176 198138
rect 174228 198060 174280 198066
rect 174228 198002 174280 198008
rect 174134 197688 174190 197697
rect 174134 197623 174190 197632
rect 174240 197561 174268 198002
rect 174226 197552 174282 197561
rect 174226 197487 174282 197496
rect 135404 197448 135456 197454
rect 135402 197416 135404 197425
rect 136692 197448 136744 197454
rect 135456 197416 135458 197425
rect 136692 197390 136744 197396
rect 135402 197351 135458 197360
rect 102466 197008 102522 197017
rect 102466 196943 102522 196952
rect 100718 196872 100774 196881
rect 100718 196807 100774 196816
rect 136782 196872 136838 196881
rect 136782 196807 136838 196816
rect 172570 196872 172626 196881
rect 172570 196807 172572 196816
rect 66218 196736 66274 196745
rect 100732 196706 100760 196807
rect 66218 196671 66274 196680
rect 100720 196700 100772 196706
rect 66232 196570 66260 196671
rect 100720 196642 100772 196648
rect 102376 196700 102428 196706
rect 102376 196642 102428 196648
rect 100902 196600 100958 196609
rect 66220 196564 66272 196570
rect 100902 196535 100904 196544
rect 66220 196506 66272 196512
rect 100956 196535 100958 196544
rect 100904 196506 100956 196512
rect 65024 196360 65076 196366
rect 102388 196337 102416 196642
rect 136690 196600 136746 196609
rect 102468 196564 102520 196570
rect 136690 196535 136746 196544
rect 102468 196506 102520 196512
rect 65024 196302 65076 196308
rect 102374 196328 102430 196337
rect 102374 196263 102430 196272
rect 65022 195784 65078 195793
rect 65022 195719 65078 195728
rect 62630 195648 62686 195657
rect 62630 195583 62686 195592
rect 62540 195136 62592 195142
rect 62540 195078 62592 195084
rect 62552 194297 62580 195078
rect 65036 195074 65064 195719
rect 102480 195657 102508 196506
rect 135404 196428 135456 196434
rect 135404 196370 135456 196376
rect 135416 196337 135444 196370
rect 135402 196328 135458 196337
rect 135402 196263 135458 196272
rect 136704 196230 136732 196535
rect 136796 196434 136824 196807
rect 172624 196807 172626 196816
rect 174136 196836 174188 196842
rect 172572 196778 172624 196784
rect 174136 196778 174188 196784
rect 172662 196600 172718 196609
rect 172662 196535 172664 196544
rect 172716 196535 172718 196544
rect 172664 196506 172716 196512
rect 136784 196428 136836 196434
rect 136784 196370 136836 196376
rect 174148 196337 174176 196778
rect 174228 196564 174280 196570
rect 174228 196506 174280 196512
rect 174134 196328 174190 196337
rect 174134 196263 174190 196272
rect 135404 196224 135456 196230
rect 135402 196192 135404 196201
rect 136692 196224 136744 196230
rect 135456 196192 135458 196201
rect 174240 196201 174268 196506
rect 136692 196166 136744 196172
rect 174226 196192 174282 196201
rect 135402 196127 135458 196136
rect 174226 196127 174282 196136
rect 172386 195784 172442 195793
rect 172386 195719 172442 195728
rect 100902 195648 100958 195657
rect 100902 195583 100958 195592
rect 102466 195648 102522 195657
rect 102466 195583 102522 195592
rect 136874 195648 136930 195657
rect 136874 195583 136930 195592
rect 66402 195512 66458 195521
rect 100916 195482 100944 195583
rect 66402 195447 66458 195456
rect 100904 195476 100956 195482
rect 66416 195210 66444 195447
rect 100904 195418 100956 195424
rect 102560 195476 102612 195482
rect 102560 195418 102612 195424
rect 100902 195240 100958 195249
rect 66404 195204 66456 195210
rect 100902 195175 100904 195184
rect 66404 195146 66456 195152
rect 100956 195175 100958 195184
rect 102376 195204 102428 195210
rect 100904 195146 100956 195152
rect 102376 195146 102428 195152
rect 62632 195068 62684 195074
rect 62632 195010 62684 195016
rect 65024 195068 65076 195074
rect 65024 195010 65076 195016
rect 62644 194977 62672 195010
rect 62630 194968 62686 194977
rect 62630 194903 62686 194912
rect 65022 194560 65078 194569
rect 65022 194495 65078 194504
rect 62538 194288 62594 194297
rect 62538 194223 62594 194232
rect 64930 193744 64986 193753
rect 62632 193708 62684 193714
rect 64930 193679 64986 193688
rect 62632 193650 62684 193656
rect 62540 193640 62592 193646
rect 62538 193608 62540 193617
rect 62592 193608 62594 193617
rect 62538 193543 62594 193552
rect 62644 192937 62672 193650
rect 62630 192928 62686 192937
rect 62630 192863 62686 192872
rect 11938 192656 11994 192665
rect 11938 192591 11994 192600
rect 11952 179745 11980 192591
rect 62632 192484 62684 192490
rect 62632 192426 62684 192432
rect 62540 192280 62592 192286
rect 62538 192248 62540 192257
rect 62592 192248 62594 192257
rect 62538 192183 62594 192192
rect 62356 191668 62408 191674
rect 62356 191610 62408 191616
rect 62368 191577 62396 191610
rect 62354 191568 62410 191577
rect 62354 191503 62410 191512
rect 62644 190897 62672 192426
rect 64944 192286 64972 193679
rect 65036 193646 65064 194495
rect 100626 194424 100682 194433
rect 100626 194359 100628 194368
rect 100680 194359 100682 194368
rect 100628 194330 100680 194336
rect 102388 194297 102416 195146
rect 102572 194977 102600 195418
rect 136782 195240 136838 195249
rect 136888 195210 136916 195583
rect 172400 195278 172428 195719
rect 172662 195376 172718 195385
rect 172662 195311 172664 195320
rect 172716 195311 172718 195320
rect 174136 195340 174188 195346
rect 172664 195282 172716 195288
rect 174136 195282 174188 195288
rect 172388 195272 172440 195278
rect 172388 195214 172440 195220
rect 136782 195175 136838 195184
rect 136876 195204 136928 195210
rect 135404 195136 135456 195142
rect 135404 195078 135456 195084
rect 135416 194977 135444 195078
rect 102558 194968 102614 194977
rect 102558 194903 102614 194912
rect 135402 194968 135458 194977
rect 135402 194903 135458 194912
rect 136796 194870 136824 195175
rect 136876 195146 136928 195152
rect 135404 194864 135456 194870
rect 135402 194832 135404 194841
rect 136784 194864 136836 194870
rect 135456 194832 135458 194841
rect 174148 194841 174176 195282
rect 174228 195272 174280 195278
rect 174228 195214 174280 195220
rect 174240 194977 174268 195214
rect 174226 194968 174282 194977
rect 174226 194903 174282 194912
rect 136784 194806 136836 194812
rect 174134 194832 174190 194841
rect 135402 194767 135458 194776
rect 174134 194767 174190 194776
rect 136782 194424 136838 194433
rect 102468 194388 102520 194394
rect 136782 194359 136838 194368
rect 171742 194424 171798 194433
rect 171742 194359 171798 194368
rect 102468 194330 102520 194336
rect 66402 194288 66458 194297
rect 66402 194223 66458 194232
rect 102374 194288 102430 194297
rect 102374 194223 102430 194232
rect 66416 193782 66444 194223
rect 100626 193880 100682 193889
rect 100626 193815 100628 193824
rect 100680 193815 100682 193824
rect 102376 193844 102428 193850
rect 100628 193786 100680 193792
rect 102376 193786 102428 193792
rect 66404 193776 66456 193782
rect 66404 193718 66456 193724
rect 65024 193640 65076 193646
rect 65024 193582 65076 193588
rect 99890 193336 99946 193345
rect 99890 193271 99946 193280
rect 99904 192966 99932 193271
rect 99892 192960 99944 192966
rect 102388 192937 102416 193786
rect 102480 193617 102508 194330
rect 136690 193880 136746 193889
rect 136690 193815 136746 193824
rect 135404 193708 135456 193714
rect 135404 193650 135456 193656
rect 135416 193617 135444 193650
rect 102466 193608 102522 193617
rect 102466 193543 102522 193552
rect 135402 193608 135458 193617
rect 135402 193543 135458 193552
rect 136704 193510 136732 193815
rect 136796 193714 136824 194359
rect 171756 193986 171784 194359
rect 172662 194016 172718 194025
rect 171744 193980 171796 193986
rect 172662 193951 172718 193960
rect 174136 193980 174188 193986
rect 171744 193922 171796 193928
rect 172676 193918 172704 193951
rect 174136 193922 174188 193928
rect 172664 193912 172716 193918
rect 172664 193854 172716 193860
rect 136784 193708 136836 193714
rect 136784 193650 136836 193656
rect 174148 193617 174176 193922
rect 174228 193912 174280 193918
rect 174228 193854 174280 193860
rect 174134 193608 174190 193617
rect 174134 193543 174190 193552
rect 135404 193504 135456 193510
rect 135402 193472 135404 193481
rect 136692 193504 136744 193510
rect 135456 193472 135458 193481
rect 174240 193481 174268 193854
rect 136692 193446 136744 193452
rect 174226 193472 174282 193481
rect 135402 193407 135458 193416
rect 174226 193407 174282 193416
rect 136782 193336 136838 193345
rect 136782 193271 136838 193280
rect 172018 193336 172074 193345
rect 172018 193271 172074 193280
rect 102468 192960 102520 192966
rect 99892 192902 99944 192908
rect 102374 192928 102430 192937
rect 102468 192902 102520 192908
rect 102374 192863 102430 192872
rect 65022 192792 65078 192801
rect 65022 192727 65078 192736
rect 64932 192280 64984 192286
rect 64932 192222 64984 192228
rect 65036 191674 65064 192727
rect 100626 192656 100682 192665
rect 100626 192591 100682 192600
rect 65666 192520 65722 192529
rect 65666 192455 65668 192464
rect 65720 192455 65722 192464
rect 100534 192520 100590 192529
rect 100640 192490 100668 192591
rect 100534 192455 100590 192464
rect 100628 192484 100680 192490
rect 65668 192426 65720 192432
rect 100548 192422 100576 192455
rect 100628 192426 100680 192432
rect 102376 192484 102428 192490
rect 102376 192426 102428 192432
rect 100536 192416 100588 192422
rect 100536 192358 100588 192364
rect 65024 191668 65076 191674
rect 65024 191610 65076 191616
rect 102388 191577 102416 192426
rect 102480 192257 102508 192902
rect 136690 192656 136746 192665
rect 136690 192591 136746 192600
rect 102652 192416 102704 192422
rect 102652 192358 102704 192364
rect 135312 192416 135364 192422
rect 135312 192358 135364 192364
rect 102466 192248 102522 192257
rect 102466 192183 102522 192192
rect 65022 191568 65078 191577
rect 65022 191503 65078 191512
rect 102374 191568 102430 191577
rect 102374 191503 102430 191512
rect 62630 190888 62686 190897
rect 62356 190852 62408 190858
rect 65036 190858 65064 191503
rect 100626 191432 100682 191441
rect 100626 191367 100682 191376
rect 65206 191296 65262 191305
rect 100640 191266 100668 191367
rect 65206 191231 65262 191240
rect 100628 191260 100680 191266
rect 62630 190823 62686 190832
rect 65024 190852 65076 190858
rect 62356 190794 62408 190800
rect 65024 190794 65076 190800
rect 62368 190217 62396 190794
rect 62354 190208 62410 190217
rect 62354 190143 62410 190152
rect 63644 189696 63696 189702
rect 63644 189638 63696 189644
rect 65022 189664 65078 189673
rect 62632 189560 62684 189566
rect 62630 189528 62632 189537
rect 62684 189528 62686 189537
rect 62630 189463 62686 189472
rect 62632 189084 62684 189090
rect 62632 189026 62684 189032
rect 62644 188857 62672 189026
rect 62630 188848 62686 188857
rect 62630 188783 62686 188792
rect 63656 188177 63684 189638
rect 65022 189599 65078 189608
rect 65036 189090 65064 189599
rect 65220 189566 65248 191231
rect 100628 191202 100680 191208
rect 102284 191260 102336 191266
rect 102284 191202 102336 191208
rect 100902 191160 100958 191169
rect 100902 191095 100958 191104
rect 100916 191062 100944 191095
rect 100904 191056 100956 191062
rect 100904 190998 100956 191004
rect 66310 190752 66366 190761
rect 66310 190687 66366 190696
rect 66324 189673 66352 190687
rect 100442 190344 100498 190353
rect 100442 190279 100498 190288
rect 66402 190208 66458 190217
rect 100456 190178 100484 190279
rect 102296 190217 102324 191202
rect 102560 191056 102612 191062
rect 102560 190998 102612 191004
rect 102282 190208 102338 190217
rect 66402 190143 66458 190152
rect 100444 190172 100496 190178
rect 66416 189702 66444 190143
rect 102282 190143 102338 190152
rect 102376 190172 102428 190178
rect 100444 190114 100496 190120
rect 102376 190114 102428 190120
rect 99982 189936 100038 189945
rect 99982 189871 99984 189880
rect 100036 189871 100038 189880
rect 99984 189842 100036 189848
rect 66404 189696 66456 189702
rect 66310 189664 66366 189673
rect 66404 189638 66456 189644
rect 66310 189599 66366 189608
rect 65208 189560 65260 189566
rect 65208 189502 65260 189508
rect 65024 189084 65076 189090
rect 65024 189026 65076 189032
rect 102388 188857 102416 190114
rect 102468 189900 102520 189906
rect 102468 189842 102520 189848
rect 102374 188848 102430 188857
rect 102374 188783 102430 188792
rect 102480 188177 102508 189842
rect 102572 189537 102600 190998
rect 102664 190897 102692 192358
rect 135220 192144 135272 192150
rect 135218 192112 135220 192121
rect 135272 192112 135274 192121
rect 135218 192047 135274 192056
rect 134208 191056 134260 191062
rect 134208 190998 134260 191004
rect 102650 190888 102706 190897
rect 102650 190823 102706 190832
rect 134220 189537 134248 190998
rect 135324 190897 135352 192358
rect 135404 192348 135456 192354
rect 135404 192290 135456 192296
rect 135416 192257 135444 192290
rect 135402 192248 135458 192257
rect 135402 192183 135458 192192
rect 136704 192150 136732 192591
rect 136796 192354 136824 193271
rect 172032 192694 172060 193271
rect 172662 192792 172718 192801
rect 172662 192727 172664 192736
rect 172716 192727 172718 192736
rect 174228 192756 174280 192762
rect 172664 192698 172716 192704
rect 174228 192698 174280 192704
rect 172020 192688 172072 192694
rect 171650 192656 171706 192665
rect 172020 192630 172072 192636
rect 174136 192688 174188 192694
rect 174136 192630 174188 192636
rect 171650 192591 171652 192600
rect 171704 192591 171706 192600
rect 171652 192562 171704 192568
rect 136874 192520 136930 192529
rect 136874 192455 136930 192464
rect 136888 192422 136916 192455
rect 136876 192416 136928 192422
rect 136876 192358 136928 192364
rect 136784 192348 136836 192354
rect 136784 192290 136836 192296
rect 174148 192257 174176 192630
rect 174134 192248 174190 192257
rect 174134 192183 174190 192192
rect 136692 192144 136744 192150
rect 174240 192121 174268 192698
rect 174320 192620 174372 192626
rect 174320 192562 174372 192568
rect 136692 192086 136744 192092
rect 174226 192112 174282 192121
rect 174226 192047 174282 192056
rect 136782 191432 136838 191441
rect 136782 191367 136838 191376
rect 172662 191432 172718 191441
rect 172662 191367 172718 191376
rect 135310 190888 135366 190897
rect 135310 190823 135366 190832
rect 136796 190790 136824 191367
rect 172676 191266 172704 191367
rect 172664 191260 172716 191266
rect 172664 191202 172716 191208
rect 174044 191260 174096 191266
rect 174044 191202 174096 191208
rect 137150 191160 137206 191169
rect 137150 191095 137206 191104
rect 171834 191160 171890 191169
rect 171834 191095 171836 191104
rect 137164 191062 137192 191095
rect 171888 191095 171890 191104
rect 171836 191066 171888 191072
rect 137152 191056 137204 191062
rect 137152 190998 137204 191004
rect 135404 190784 135456 190790
rect 135402 190752 135404 190761
rect 136784 190784 136836 190790
rect 135456 190752 135458 190761
rect 174056 190761 174084 191202
rect 174332 190897 174360 192562
rect 207268 192529 207296 222754
rect 223538 211152 223594 211161
rect 223538 211087 223594 211096
rect 223552 210374 223580 211087
rect 207900 210368 207952 210374
rect 207900 210310 207952 210316
rect 223540 210368 223592 210374
rect 223540 210310 223592 210316
rect 207912 201777 207940 210310
rect 207898 201768 207954 201777
rect 207898 201703 207954 201712
rect 207254 192520 207310 192529
rect 207254 192455 207310 192464
rect 207254 192384 207310 192393
rect 207254 192319 207310 192328
rect 175332 191124 175384 191130
rect 175332 191066 175384 191072
rect 174318 190888 174374 190897
rect 174318 190823 174374 190832
rect 136784 190726 136836 190732
rect 174042 190752 174098 190761
rect 135402 190687 135458 190696
rect 174042 190687 174098 190696
rect 136782 190344 136838 190353
rect 136782 190279 136838 190288
rect 171650 190344 171706 190353
rect 171650 190279 171706 190288
rect 102558 189528 102614 189537
rect 102558 189463 102614 189472
rect 134206 189528 134262 189537
rect 134206 189463 134262 189472
rect 136796 189294 136824 190279
rect 171664 189974 171692 190279
rect 171652 189968 171704 189974
rect 137242 189936 137298 189945
rect 174412 189968 174464 189974
rect 171652 189910 171704 189916
rect 171834 189936 171890 189945
rect 137242 189871 137298 189880
rect 174412 189910 174464 189916
rect 171834 189871 171890 189880
rect 134760 189288 134812 189294
rect 134758 189256 134760 189265
rect 136784 189288 136836 189294
rect 134812 189256 134814 189265
rect 136784 189230 136836 189236
rect 134758 189191 134814 189200
rect 137256 188206 137284 189871
rect 171848 189770 171876 189871
rect 171836 189764 171888 189770
rect 171836 189706 171888 189712
rect 174424 189265 174452 189910
rect 175344 189537 175372 191066
rect 175424 189764 175476 189770
rect 175424 189706 175476 189712
rect 175330 189528 175386 189537
rect 175330 189463 175386 189472
rect 174410 189256 174466 189265
rect 174410 189191 174466 189200
rect 134944 188200 134996 188206
rect 63642 188168 63698 188177
rect 63642 188103 63698 188112
rect 102466 188168 102522 188177
rect 102466 188103 102522 188112
rect 134942 188168 134944 188177
rect 137244 188200 137296 188206
rect 134996 188168 134998 188177
rect 175436 188177 175464 189706
rect 137244 188142 137296 188148
rect 175422 188168 175478 188177
rect 134942 188103 134998 188112
rect 175422 188103 175478 188112
rect 32008 187854 32942 187882
rect 11938 179736 11994 179745
rect 11938 179671 11994 179680
rect 32008 178249 32036 187854
rect 33572 184126 33600 187868
rect 34216 184330 34244 187868
rect 34952 185146 34980 187868
rect 34940 185140 34992 185146
rect 34940 185082 34992 185088
rect 35596 184466 35624 187868
rect 36332 185486 36360 187868
rect 36320 185480 36372 185486
rect 36320 185422 36372 185428
rect 36976 185214 37004 187868
rect 37620 185350 37648 187868
rect 37608 185344 37660 185350
rect 37608 185286 37660 185292
rect 36964 185208 37016 185214
rect 36964 185150 37016 185156
rect 38356 185010 38384 187868
rect 39000 185078 39028 187868
rect 39736 185282 39764 187868
rect 40380 185418 40408 187868
rect 41024 185486 41052 187868
rect 40644 185480 40696 185486
rect 40644 185422 40696 185428
rect 41012 185480 41064 185486
rect 41012 185422 41064 185428
rect 40368 185412 40420 185418
rect 40368 185354 40420 185360
rect 39724 185276 39776 185282
rect 39724 185218 39776 185224
rect 39540 185140 39592 185146
rect 39540 185082 39592 185088
rect 38988 185072 39040 185078
rect 38988 185014 39040 185020
rect 38344 185004 38396 185010
rect 38344 184946 38396 184952
rect 39552 184754 39580 185082
rect 39552 184726 39842 184754
rect 40656 184740 40684 185422
rect 41760 185350 41788 187868
rect 41472 185344 41524 185350
rect 41472 185286 41524 185292
rect 41748 185344 41800 185350
rect 41748 185286 41800 185292
rect 41012 185208 41064 185214
rect 41012 185150 41064 185156
rect 41024 184740 41052 185150
rect 41484 184740 41512 185286
rect 42404 185146 42432 187868
rect 43140 185418 43168 187868
rect 43784 185486 43812 187868
rect 44534 187854 45100 187882
rect 45178 187854 45652 187882
rect 45822 187854 46112 187882
rect 43404 185480 43456 185486
rect 43404 185422 43456 185428
rect 43772 185480 43824 185486
rect 43772 185422 43824 185428
rect 44692 185480 44744 185486
rect 44692 185422 44744 185428
rect 43036 185412 43088 185418
rect 43036 185354 43088 185360
rect 43128 185412 43180 185418
rect 43128 185354 43180 185360
rect 42668 185276 42720 185282
rect 42668 185218 42720 185224
rect 42392 185140 42444 185146
rect 42392 185082 42444 185088
rect 42208 185072 42260 185078
rect 42208 185014 42260 185020
rect 41840 185004 41892 185010
rect 41840 184946 41892 184952
rect 41852 184740 41880 184946
rect 42220 184740 42248 185014
rect 42680 184740 42708 185218
rect 43048 184740 43076 185354
rect 43416 184740 43444 185422
rect 44600 185412 44652 185418
rect 44600 185354 44652 185360
rect 43864 185344 43916 185350
rect 43864 185286 43916 185292
rect 43876 184740 43904 185286
rect 44232 185140 44284 185146
rect 44232 185082 44284 185088
rect 44244 184740 44272 185082
rect 44612 184740 44640 185354
rect 44704 184754 44732 185422
rect 45072 184890 45100 187854
rect 45072 184862 45192 184890
rect 45164 184754 45192 184862
rect 45624 184754 45652 187854
rect 46084 184754 46112 187854
rect 46544 184754 46572 187868
rect 47188 184754 47216 187868
rect 47648 187854 47938 187882
rect 48200 187854 48582 187882
rect 48660 187854 49226 187882
rect 47648 184754 47676 187854
rect 48200 184754 48228 187854
rect 48660 185162 48688 187854
rect 49016 185480 49068 185486
rect 49016 185422 49068 185428
rect 48568 185134 48688 185162
rect 48568 184754 48596 185134
rect 48648 185072 48700 185078
rect 48648 185014 48700 185020
rect 44704 184726 45086 184754
rect 45164 184726 45454 184754
rect 45624 184726 45822 184754
rect 46084 184726 46282 184754
rect 46544 184726 46650 184754
rect 47110 184726 47216 184754
rect 47478 184726 47676 184754
rect 47846 184726 48228 184754
rect 48306 184726 48596 184754
rect 48660 184740 48688 185014
rect 49028 184740 49056 185422
rect 49844 185412 49896 185418
rect 49844 185354 49896 185360
rect 49476 185276 49528 185282
rect 49476 185218 49528 185224
rect 49488 184740 49516 185218
rect 49856 184740 49884 185354
rect 49948 185078 49976 187868
rect 50592 185486 50620 187868
rect 50580 185480 50632 185486
rect 50580 185422 50632 185428
rect 50672 185480 50724 185486
rect 50672 185422 50724 185428
rect 50212 185208 50264 185214
rect 50212 185150 50264 185156
rect 49936 185072 49988 185078
rect 49936 185014 49988 185020
rect 50224 184740 50252 185150
rect 50684 184740 50712 185422
rect 51328 185282 51356 187868
rect 51972 185418 52000 187868
rect 51960 185412 52012 185418
rect 51960 185354 52012 185360
rect 52236 185344 52288 185350
rect 52236 185286 52288 185292
rect 51316 185276 51368 185282
rect 51316 185218 51368 185224
rect 51040 185072 51092 185078
rect 51040 185014 51092 185020
rect 51052 184740 51080 185014
rect 51408 185004 51460 185010
rect 51408 184946 51460 184952
rect 51420 184740 51448 184946
rect 51868 184936 51920 184942
rect 51868 184878 51920 184884
rect 51880 184740 51908 184878
rect 52248 184740 52276 185286
rect 52708 185214 52736 187868
rect 53352 185486 53380 187868
rect 53340 185480 53392 185486
rect 53340 185422 53392 185428
rect 53432 185480 53484 185486
rect 53432 185422 53484 185428
rect 53064 185276 53116 185282
rect 53064 185218 53116 185224
rect 52696 185208 52748 185214
rect 52696 185150 52748 185156
rect 52604 185140 52656 185146
rect 52604 185082 52656 185088
rect 52616 184740 52644 185082
rect 53076 184740 53104 185218
rect 53444 184740 53472 185422
rect 53996 185078 54024 187868
rect 53984 185072 54036 185078
rect 53984 185014 54036 185020
rect 54732 185010 54760 187868
rect 54720 185004 54772 185010
rect 54720 184946 54772 184952
rect 55376 184942 55404 187868
rect 56112 185350 56140 187868
rect 56100 185344 56152 185350
rect 56100 185286 56152 185292
rect 56756 185146 56784 187868
rect 57400 185282 57428 187868
rect 58136 185486 58164 187868
rect 58124 185480 58176 185486
rect 58124 185422 58176 185428
rect 57388 185276 57440 185282
rect 57388 185218 57440 185224
rect 56744 185140 56796 185146
rect 56744 185082 56796 185088
rect 55364 184936 55416 184942
rect 55364 184878 55416 184884
rect 38158 184496 38214 184505
rect 35584 184460 35636 184466
rect 40182 184496 40238 184505
rect 38158 184431 38160 184440
rect 35584 184402 35636 184408
rect 38212 184431 38214 184440
rect 38908 184454 39106 184482
rect 39276 184466 39474 184482
rect 39264 184460 39474 184466
rect 38160 184402 38212 184408
rect 34204 184324 34256 184330
rect 34204 184266 34256 184272
rect 38908 184126 38936 184454
rect 39316 184454 39474 184460
rect 40238 184454 40302 184482
rect 53826 184466 54024 184482
rect 54286 184466 54576 184482
rect 53826 184460 54036 184466
rect 53826 184454 53984 184460
rect 40182 184431 40238 184440
rect 39264 184402 39316 184408
rect 54286 184460 54588 184466
rect 54286 184454 54536 184460
rect 53984 184402 54036 184408
rect 54654 184454 54944 184482
rect 54536 184402 54588 184408
rect 54916 184233 54944 184454
rect 54902 184224 54958 184233
rect 54902 184159 54958 184168
rect 58780 184126 58808 187868
rect 59516 184262 59544 187868
rect 59504 184256 59556 184262
rect 60160 184233 60188 187868
rect 105194 187610 105222 187868
rect 105148 187582 105222 187610
rect 105332 187854 105760 187882
rect 105884 187854 106312 187882
rect 106620 187854 106956 187882
rect 107172 187854 107508 187882
rect 107908 187854 108060 187882
rect 108368 187854 108704 187882
rect 109256 187854 109316 187882
rect 109808 187854 110144 187882
rect 110452 187854 110788 187882
rect 111004 187854 111432 187882
rect 111556 187854 111984 187882
rect 112200 187854 112444 187882
rect 112752 187854 113088 187882
rect 113304 187854 113456 187882
rect 59504 184198 59556 184204
rect 60146 184224 60202 184233
rect 60146 184159 60202 184168
rect 33560 184120 33612 184126
rect 33560 184062 33612 184068
rect 38896 184120 38948 184126
rect 38896 184062 38948 184068
rect 58768 184120 58820 184126
rect 58768 184062 58820 184068
rect 31994 178240 32050 178249
rect 31994 178175 32050 178184
rect 37422 178240 37478 178249
rect 37422 178175 37478 178184
rect 59594 178240 59650 178249
rect 59594 178175 59650 178184
rect 37436 177258 37464 178175
rect 32640 177252 32692 177258
rect 32640 177194 32692 177200
rect 37424 177252 37476 177258
rect 37424 177194 37476 177200
rect 12030 171032 12086 171041
rect 12030 170967 12086 170976
rect 11938 149816 11994 149825
rect 11938 149751 11994 149760
rect 11952 62921 11980 149751
rect 12044 105761 12072 170967
rect 12122 169264 12178 169273
rect 12122 169199 12178 169208
rect 12136 149417 12164 169199
rect 32652 164921 32680 177194
rect 59608 175830 59636 178175
rect 105148 176753 105176 187582
rect 105332 183938 105360 187854
rect 105596 185276 105648 185282
rect 105596 185218 105648 185224
rect 105608 184777 105636 185218
rect 105594 184768 105650 184777
rect 105594 184703 105650 184712
rect 105240 183910 105360 183938
rect 105240 177977 105268 183910
rect 105596 182420 105648 182426
rect 105596 182362 105648 182368
rect 105608 182329 105636 182362
rect 105594 182320 105650 182329
rect 105594 182255 105650 182264
rect 105884 181218 105912 187854
rect 106056 184392 106108 184398
rect 106056 184334 106108 184340
rect 105964 184120 106016 184126
rect 105964 184062 106016 184068
rect 105332 181190 105912 181218
rect 105332 178521 105360 181190
rect 105412 180380 105464 180386
rect 105412 180322 105464 180328
rect 105318 178512 105374 178521
rect 105318 178447 105374 178456
rect 105226 177968 105282 177977
rect 105226 177903 105282 177912
rect 105134 176744 105190 176753
rect 105134 176679 105190 176688
rect 57388 175824 57440 175830
rect 57388 175766 57440 175772
rect 59596 175824 59648 175830
rect 59596 175766 59648 175772
rect 57400 174849 57428 175766
rect 57386 174840 57442 174849
rect 57386 174775 57442 174784
rect 105424 174441 105452 180322
rect 105976 179881 106004 184062
rect 106068 181241 106096 184334
rect 106620 184126 106648 187854
rect 107172 184398 107200 187854
rect 107160 184392 107212 184398
rect 107160 184334 107212 184340
rect 106608 184120 106660 184126
rect 106608 184062 106660 184068
rect 106148 184052 106200 184058
rect 106148 183994 106200 184000
rect 106160 183689 106188 183994
rect 106146 183680 106202 183689
rect 106146 183615 106202 183624
rect 107908 182426 107936 187854
rect 108368 184126 108396 187854
rect 109288 185282 109316 187854
rect 110116 185486 110144 187854
rect 110104 185480 110156 185486
rect 110104 185422 110156 185428
rect 110760 185418 110788 187854
rect 111404 185570 111432 187854
rect 111404 185542 111616 185570
rect 111116 185480 111168 185486
rect 111116 185422 111168 185428
rect 110748 185412 110800 185418
rect 110748 185354 110800 185360
rect 109276 185276 109328 185282
rect 109276 185218 109328 185224
rect 111128 184740 111156 185422
rect 111484 185412 111536 185418
rect 111484 185354 111536 185360
rect 111496 184740 111524 185354
rect 111588 184754 111616 185542
rect 111956 184754 111984 187854
rect 112416 184754 112444 187854
rect 111588 184726 111878 184754
rect 111956 184726 112338 184754
rect 112416 184726 112706 184754
rect 113060 184740 113088 187854
rect 113428 184754 113456 187854
rect 113934 187610 113962 187868
rect 113888 187582 113962 187610
rect 114256 187854 114500 187882
rect 114716 187854 115052 187882
rect 115360 187854 115696 187882
rect 115820 187854 116248 187882
rect 116372 187854 116800 187882
rect 113428 184726 113534 184754
rect 113888 184740 113916 187582
rect 114256 184740 114284 187854
rect 114716 184740 114744 187854
rect 115360 184754 115388 187854
rect 115820 184754 115848 187854
rect 116372 184890 116400 187854
rect 117430 187662 117458 187868
rect 117660 187854 117996 187882
rect 118212 187854 118548 187882
rect 118948 187854 119192 187882
rect 119592 187854 119744 187882
rect 120296 187854 120356 187882
rect 116452 187656 116504 187662
rect 116452 187598 116504 187604
rect 117418 187656 117470 187662
rect 117418 187598 117470 187604
rect 116188 184862 116400 184890
rect 116188 184754 116216 184862
rect 116464 184754 116492 187598
rect 117556 185480 117608 185486
rect 117094 185448 117150 185457
rect 117556 185422 117608 185428
rect 117094 185383 117150 185392
rect 116910 184768 116966 184777
rect 115098 184726 115388 184754
rect 115466 184726 115848 184754
rect 115926 184726 116216 184754
rect 116294 184726 116492 184754
rect 116662 184726 116910 184754
rect 117108 184740 117136 185383
rect 117568 184754 117596 185422
rect 117660 184777 117688 187854
rect 118212 185457 118240 187854
rect 118948 185486 118976 187854
rect 118936 185480 118988 185486
rect 118198 185448 118254 185457
rect 118936 185422 118988 185428
rect 119118 185448 119174 185457
rect 118198 185383 118254 185392
rect 118568 185412 118620 185418
rect 119118 185383 119174 185392
rect 118568 185354 118620 185360
rect 117490 184726 117596 184754
rect 117646 184768 117702 184777
rect 116910 184703 116966 184712
rect 118106 184768 118162 184777
rect 117858 184726 118106 184754
rect 117646 184703 117702 184712
rect 118580 184754 118608 185354
rect 118936 185276 118988 185282
rect 118936 185218 118988 185224
rect 118948 184754 118976 185218
rect 118318 184726 118608 184754
rect 118686 184726 118976 184754
rect 119132 184740 119160 185383
rect 119486 185312 119542 185321
rect 119486 185247 119542 185256
rect 119500 184740 119528 185247
rect 119592 184777 119620 187854
rect 120224 185480 120276 185486
rect 120224 185422 120276 185428
rect 119578 184768 119634 184777
rect 118106 184703 118162 184712
rect 120236 184754 120264 185422
rect 120328 185418 120356 187854
rect 120604 187854 120940 187882
rect 121156 187854 121492 187882
rect 121708 187854 122044 187882
rect 122352 187854 122688 187882
rect 123088 187854 123240 187882
rect 123456 187854 123792 187882
rect 124436 187854 124496 187882
rect 120316 185412 120368 185418
rect 120316 185354 120368 185360
rect 120604 185282 120632 187854
rect 121156 185457 121184 187854
rect 121142 185448 121198 185457
rect 121142 185383 121198 185392
rect 121602 185312 121658 185321
rect 120592 185276 120644 185282
rect 121708 185298 121736 187854
rect 122352 185486 122380 187854
rect 122340 185480 122392 185486
rect 122340 185422 122392 185428
rect 122432 185480 122484 185486
rect 122432 185422 122484 185428
rect 121658 185270 121736 185298
rect 121602 185247 121658 185256
rect 120592 185218 120644 185224
rect 122444 185185 122472 185422
rect 123088 185298 123116 187854
rect 123456 185486 123484 187854
rect 123444 185480 123496 185486
rect 123444 185422 123496 185428
rect 124180 185480 124232 185486
rect 124180 185422 124232 185428
rect 122904 185270 123116 185298
rect 123812 185344 123864 185350
rect 123812 185286 123864 185292
rect 123352 185276 123404 185282
rect 122616 185208 122668 185214
rect 120682 185176 120738 185185
rect 120682 185111 120738 185120
rect 122430 185176 122486 185185
rect 122616 185150 122668 185156
rect 122430 185111 122486 185120
rect 120314 185040 120370 185049
rect 120314 184975 120370 184984
rect 119882 184726 120264 184754
rect 120328 184740 120356 184975
rect 120696 184740 120724 185111
rect 121328 185072 121380 185078
rect 121328 185014 121380 185020
rect 121340 184754 121368 185014
rect 121788 185004 121840 185010
rect 121788 184946 121840 184952
rect 121800 184754 121828 184946
rect 122156 184936 122208 184942
rect 122156 184878 122208 184884
rect 122168 184754 122196 184878
rect 122628 184754 122656 185150
rect 122904 185049 122932 185270
rect 123352 185218 123404 185224
rect 122984 185140 123036 185146
rect 122984 185082 123036 185088
rect 122890 185040 122946 185049
rect 122890 184975 122946 184984
rect 122996 184754 123024 185082
rect 123364 184754 123392 185218
rect 123824 184754 123852 185286
rect 124192 184754 124220 185422
rect 124468 185078 124496 187854
rect 124652 187854 124988 187882
rect 125204 187854 125540 187882
rect 125848 187854 126184 187882
rect 126400 187854 126736 187882
rect 127288 187854 127348 187882
rect 124548 185412 124600 185418
rect 124548 185354 124600 185360
rect 124456 185072 124508 185078
rect 124456 185014 124508 185020
rect 124560 184754 124588 185354
rect 124652 185010 124680 187854
rect 125098 185312 125154 185321
rect 125098 185247 125154 185256
rect 124640 185004 124692 185010
rect 124640 184946 124692 184952
rect 124914 184904 124970 184913
rect 124914 184839 124970 184848
rect 124928 184754 124956 184839
rect 121078 184726 121368 184754
rect 121538 184726 121828 184754
rect 121906 184726 122196 184754
rect 122274 184726 122656 184754
rect 122734 184726 123024 184754
rect 123102 184726 123392 184754
rect 123470 184726 123852 184754
rect 123930 184726 124220 184754
rect 124298 184726 124588 184754
rect 124666 184726 124956 184754
rect 125112 184740 125140 185247
rect 125204 184942 125232 187854
rect 125848 185214 125876 187854
rect 125836 185208 125888 185214
rect 125466 185176 125522 185185
rect 125836 185150 125888 185156
rect 126400 185146 126428 187854
rect 126662 185448 126718 185457
rect 126662 185383 126718 185392
rect 125466 185111 125522 185120
rect 126388 185140 126440 185146
rect 125192 184936 125244 184942
rect 125192 184878 125244 184884
rect 125480 184740 125508 185111
rect 126388 185082 126440 185088
rect 125834 185040 125890 185049
rect 125834 184975 125890 184984
rect 125848 184740 125876 184975
rect 126478 184768 126534 184777
rect 126322 184726 126478 184754
rect 119578 184703 119634 184712
rect 126676 184740 126704 185383
rect 127320 185282 127348 187854
rect 127596 187854 127932 187882
rect 128148 187854 128484 187882
rect 128700 187854 129036 187882
rect 129344 187854 129680 187882
rect 129988 187854 130232 187882
rect 130448 187854 130784 187882
rect 131428 187854 131488 187882
rect 127596 185350 127624 187854
rect 128148 185486 128176 187854
rect 128136 185480 128188 185486
rect 128136 185422 128188 185428
rect 128700 185418 128728 187854
rect 128688 185412 128740 185418
rect 128688 185354 128740 185360
rect 127584 185344 127636 185350
rect 127584 185286 127636 185292
rect 127308 185276 127360 185282
rect 127308 185218 127360 185224
rect 129344 184913 129372 187854
rect 129988 185321 130016 187854
rect 129974 185312 130030 185321
rect 129974 185247 130030 185256
rect 130448 185185 130476 187854
rect 130434 185176 130490 185185
rect 130434 185111 130490 185120
rect 131460 185049 131488 187854
rect 131644 187854 131980 187882
rect 132196 187854 132532 187882
rect 177092 187854 177198 187882
rect 131446 185040 131502 185049
rect 131446 184975 131502 184984
rect 129330 184904 129386 184913
rect 129330 184839 129386 184848
rect 131644 184777 131672 187854
rect 132196 185457 132224 187854
rect 132182 185448 132238 185457
rect 132182 185383 132238 185392
rect 176896 185344 176948 185350
rect 176896 185286 176948 185292
rect 131630 184768 131686 184777
rect 126478 184703 126534 184712
rect 131630 184703 131686 184712
rect 108356 184120 108408 184126
rect 108356 184062 108408 184068
rect 108538 183544 108594 183553
rect 108538 183479 108594 183488
rect 107896 182420 107948 182426
rect 107896 182362 107948 182368
rect 106054 181232 106110 181241
rect 106054 181167 106110 181176
rect 108078 181232 108134 181241
rect 108078 181167 108134 181176
rect 108092 180386 108120 181167
rect 108080 180380 108132 180386
rect 108080 180322 108132 180328
rect 105962 179872 106018 179881
rect 105962 179807 106018 179816
rect 107894 178920 107950 178929
rect 107894 178855 107950 178864
rect 107908 178618 107936 178855
rect 106332 178612 106384 178618
rect 106332 178554 106384 178560
rect 107896 178612 107948 178618
rect 107896 178554 107948 178560
rect 106148 175416 106200 175422
rect 106146 175384 106148 175393
rect 106200 175384 106202 175393
rect 106146 175319 106202 175328
rect 105410 174432 105466 174441
rect 105410 174367 105466 174376
rect 105964 173104 106016 173110
rect 105964 173046 106016 173052
rect 105688 171744 105740 171750
rect 105688 171686 105740 171692
rect 105700 169953 105728 171686
rect 105976 171041 106004 173046
rect 106344 172945 106372 178554
rect 107894 176472 107950 176481
rect 107894 176407 107950 176416
rect 107908 175898 107936 176407
rect 106424 175892 106476 175898
rect 106424 175834 106476 175840
rect 107896 175892 107948 175898
rect 107896 175834 107948 175840
rect 106330 172936 106386 172945
rect 106330 172871 106386 172880
rect 106436 172265 106464 175834
rect 108552 175422 108580 183479
rect 176908 177433 176936 185286
rect 176988 184392 177040 184398
rect 176988 184334 177040 184340
rect 177000 180833 177028 184334
rect 176986 180824 177042 180833
rect 176986 180759 177042 180768
rect 176894 177424 176950 177433
rect 176894 177359 176950 177368
rect 177092 176209 177120 187854
rect 177736 185350 177764 187868
rect 177724 185344 177776 185350
rect 177724 185286 177776 185292
rect 177724 185208 177776 185214
rect 177724 185150 177776 185156
rect 177736 184233 177764 185150
rect 177722 184224 177778 184233
rect 177632 184188 177684 184194
rect 178288 184194 178316 187868
rect 177722 184159 177778 184168
rect 178276 184188 178328 184194
rect 177632 184130 177684 184136
rect 178276 184130 178328 184136
rect 177356 184052 177408 184058
rect 177356 183994 177408 184000
rect 177368 183145 177396 183994
rect 177354 183136 177410 183145
rect 177354 183071 177410 183080
rect 177172 182216 177224 182222
rect 177172 182158 177224 182164
rect 177184 181921 177212 182158
rect 177170 181912 177226 181921
rect 177170 181847 177226 181856
rect 177644 178521 177672 184130
rect 178840 184126 178868 187868
rect 179392 184398 179420 187868
rect 179380 184392 179432 184398
rect 179380 184334 179432 184340
rect 177816 184120 177868 184126
rect 177816 184062 177868 184068
rect 178828 184120 178880 184126
rect 178828 184062 178880 184068
rect 177828 179745 177856 184062
rect 180036 182222 180064 187868
rect 180588 184126 180616 187868
rect 181140 185214 181168 187868
rect 181128 185208 181180 185214
rect 181128 185150 181180 185156
rect 181692 185010 181720 187868
rect 182244 185486 182272 187868
rect 182232 185480 182284 185486
rect 182232 185422 182284 185428
rect 181680 185004 181732 185010
rect 181680 184946 181732 184952
rect 182888 184942 182916 187868
rect 183244 185480 183296 185486
rect 183244 185422 183296 185428
rect 183106 185004 183158 185010
rect 183106 184946 183158 184952
rect 182876 184936 182928 184942
rect 182876 184878 182928 184884
rect 183118 184740 183146 184946
rect 183256 184754 183284 185422
rect 183440 185010 183468 187868
rect 183992 186914 184020 187868
rect 183980 186908 184032 186914
rect 183980 186850 184032 186856
rect 184440 186908 184492 186914
rect 184440 186850 184492 186856
rect 183428 185004 183480 185010
rect 183428 184946 183480 184952
rect 184302 185004 184354 185010
rect 184302 184946 184354 184952
rect 183842 184936 183894 184942
rect 183842 184878 183894 184884
rect 183256 184726 183500 184754
rect 183854 184740 183882 184878
rect 184314 184740 184342 184946
rect 184452 184754 184480 186850
rect 184544 184890 184572 187868
rect 185096 184890 185124 187868
rect 184544 184862 184848 184890
rect 185096 184862 185216 184890
rect 184820 184754 184848 184862
rect 185188 184754 185216 184862
rect 185740 184754 185768 187868
rect 186292 185026 186320 187868
rect 186246 184998 186320 185026
rect 184452 184726 184696 184754
rect 184820 184726 185064 184754
rect 185188 184726 185524 184754
rect 185740 184726 185892 184754
rect 186246 184740 186274 184998
rect 186844 184754 186872 187868
rect 187396 184890 187424 187868
rect 187948 184890 187976 187868
rect 188488 186908 188540 186914
rect 188488 186850 188540 186856
rect 188120 185480 188172 185486
rect 188120 185422 188172 185428
rect 187304 184862 187424 184890
rect 187764 184862 187976 184890
rect 187304 184754 187332 184862
rect 187764 184754 187792 184862
rect 188132 184754 188160 185422
rect 188500 184754 188528 186850
rect 188592 185486 188620 187868
rect 189144 186914 189172 187868
rect 189132 186908 189184 186914
rect 189132 186850 189184 186856
rect 188580 185480 188632 185486
rect 188580 185422 188632 185428
rect 189696 185010 189724 187868
rect 188626 185004 188678 185010
rect 188626 184946 188678 184952
rect 189684 185004 189736 185010
rect 189684 184946 189736 184952
rect 189822 185004 189874 185010
rect 189822 184946 189874 184952
rect 186720 184726 186872 184754
rect 187088 184726 187332 184754
rect 187456 184726 187792 184754
rect 187916 184726 188160 184754
rect 188284 184726 188528 184754
rect 188638 184740 188666 184946
rect 189086 184936 189138 184942
rect 189086 184878 189138 184884
rect 189098 184740 189126 184878
rect 189684 184868 189736 184874
rect 189684 184810 189736 184816
rect 189696 184754 189724 184810
rect 189480 184726 189724 184754
rect 189834 184740 189862 184946
rect 190248 184942 190276 187868
rect 190604 185480 190656 185486
rect 190604 185422 190656 185428
rect 190420 185140 190472 185146
rect 190420 185082 190472 185088
rect 190236 184936 190288 184942
rect 190236 184878 190288 184884
rect 190432 184754 190460 185082
rect 190308 184726 190460 184754
rect 190616 184754 190644 185422
rect 190800 184874 190828 187868
rect 191444 185010 191472 187868
rect 191708 185412 191760 185418
rect 191708 185354 191760 185360
rect 191432 185004 191484 185010
rect 191432 184946 191484 184952
rect 191110 184936 191162 184942
rect 191110 184878 191162 184884
rect 190788 184868 190840 184874
rect 190788 184810 190840 184816
rect 190616 184726 190676 184754
rect 191122 184740 191150 184878
rect 191720 184754 191748 185354
rect 191996 185146 192024 187868
rect 192548 185486 192576 187868
rect 192536 185480 192588 185486
rect 192536 185422 192588 185428
rect 192904 185480 192956 185486
rect 192904 185422 192956 185428
rect 192536 185344 192588 185350
rect 192536 185286 192588 185292
rect 191984 185140 192036 185146
rect 191984 185082 192036 185088
rect 191846 185004 191898 185010
rect 191846 184946 191898 184952
rect 191504 184726 191748 184754
rect 191858 184740 191886 184946
rect 192548 184754 192576 185286
rect 192916 184754 192944 185422
rect 193100 184942 193128 187868
rect 193652 185418 193680 187868
rect 193640 185412 193692 185418
rect 193640 185354 193692 185360
rect 194100 185412 194152 185418
rect 194100 185354 194152 185360
rect 193364 185276 193416 185282
rect 193364 185218 193416 185224
rect 193088 184936 193140 184942
rect 193088 184878 193140 184884
rect 193376 184754 193404 185218
rect 193732 185140 193784 185146
rect 193732 185082 193784 185088
rect 193744 184754 193772 185082
rect 194112 184754 194140 185354
rect 194296 185010 194324 187868
rect 194848 185350 194876 187868
rect 195400 185486 195428 187868
rect 195388 185480 195440 185486
rect 195388 185422 195440 185428
rect 194836 185344 194888 185350
rect 194836 185286 194888 185292
rect 195756 185344 195808 185350
rect 195756 185286 195808 185292
rect 194560 185208 194612 185214
rect 194560 185150 194612 185156
rect 194284 185004 194336 185010
rect 194284 184946 194336 184952
rect 194572 184754 194600 185150
rect 194652 185072 194704 185078
rect 194652 185014 194704 185020
rect 192332 184726 192576 184754
rect 192700 184726 192944 184754
rect 193068 184726 193404 184754
rect 193528 184726 193772 184754
rect 193896 184726 194140 184754
rect 194264 184726 194600 184754
rect 194664 184618 194692 185014
rect 195296 184800 195348 184806
rect 195092 184748 195296 184754
rect 195768 184754 195796 185286
rect 195952 185282 195980 187868
rect 195940 185276 195992 185282
rect 195940 185218 195992 185224
rect 196124 185276 196176 185282
rect 196124 185218 196176 185224
rect 196136 184754 196164 185218
rect 196504 185146 196532 187868
rect 197148 185418 197176 187868
rect 197320 185480 197372 185486
rect 197320 185422 197372 185428
rect 197136 185412 197188 185418
rect 197136 185354 197188 185360
rect 196492 185140 196544 185146
rect 196492 185082 196544 185088
rect 196630 184936 196682 184942
rect 196630 184878 196682 184884
rect 196492 184868 196544 184874
rect 196492 184810 196544 184816
rect 196504 184754 196532 184810
rect 195092 184742 195348 184748
rect 195092 184726 195336 184742
rect 195460 184726 195796 184754
rect 195920 184726 196164 184754
rect 196288 184726 196532 184754
rect 196642 184740 196670 184878
rect 197332 184754 197360 185422
rect 197700 185214 197728 187868
rect 197688 185208 197740 185214
rect 197688 185150 197740 185156
rect 198252 185078 198280 187868
rect 198240 185072 198292 185078
rect 197456 185040 197512 185049
rect 198240 185014 198292 185020
rect 197456 184975 197512 184984
rect 197826 185004 197878 185010
rect 197116 184726 197360 184754
rect 197470 184740 197498 184975
rect 197826 184946 197878 184952
rect 197838 184740 197866 184946
rect 198804 184806 198832 187868
rect 199356 185350 199384 187868
rect 199344 185344 199396 185350
rect 199344 185286 199396 185292
rect 200000 185282 200028 187868
rect 199988 185276 200040 185282
rect 199988 185218 200040 185224
rect 200552 184874 200580 187868
rect 201104 184942 201132 187868
rect 201656 185486 201684 187868
rect 201644 185480 201696 185486
rect 201644 185422 201696 185428
rect 202208 185049 202236 187868
rect 202194 185040 202250 185049
rect 202852 185010 202880 187868
rect 202194 184975 202250 184984
rect 202840 185004 202892 185010
rect 202840 184946 202892 184952
rect 201092 184936 201144 184942
rect 201092 184878 201144 184884
rect 200540 184868 200592 184874
rect 200540 184810 200592 184816
rect 198792 184800 198844 184806
rect 198792 184742 198844 184748
rect 194664 184590 194724 184618
rect 203404 184505 203432 187868
rect 198514 184496 198570 184505
rect 198312 184454 198514 184482
rect 203390 184496 203446 184505
rect 198680 184454 198924 184482
rect 198514 184431 198570 184440
rect 198896 184233 198924 184454
rect 203390 184431 203446 184440
rect 203956 184233 203984 187868
rect 198882 184224 198938 184233
rect 198882 184159 198938 184168
rect 203942 184224 203998 184233
rect 203942 184159 203998 184168
rect 180576 184120 180628 184126
rect 180576 184062 180628 184068
rect 180298 183544 180354 183553
rect 180298 183479 180354 183488
rect 180024 182216 180076 182222
rect 180024 182158 180076 182164
rect 179654 181232 179710 181241
rect 179654 181167 179710 181176
rect 179668 180386 179696 181167
rect 178092 180380 178144 180386
rect 178092 180322 178144 180328
rect 179656 180380 179708 180386
rect 179656 180322 179708 180328
rect 177814 179736 177870 179745
rect 177814 179671 177870 179680
rect 177816 178612 177868 178618
rect 177816 178554 177868 178560
rect 177630 178512 177686 178521
rect 177630 178447 177686 178456
rect 177078 176200 177134 176209
rect 177078 176135 177134 176144
rect 177724 175892 177776 175898
rect 177724 175834 177776 175840
rect 177172 175620 177224 175626
rect 177172 175562 177224 175568
rect 108540 175416 108592 175422
rect 108540 175358 108592 175364
rect 177184 175121 177212 175562
rect 177170 175112 177226 175121
rect 177170 175047 177226 175056
rect 107894 174160 107950 174169
rect 107894 174095 107950 174104
rect 107908 173110 107936 174095
rect 107896 173104 107948 173110
rect 107896 173046 107948 173052
rect 177540 173104 177592 173110
rect 177540 173046 177592 173052
rect 106422 172256 106478 172265
rect 106422 172191 106478 172200
rect 108078 171848 108134 171857
rect 108078 171783 108134 171792
rect 108092 171750 108120 171783
rect 108080 171744 108132 171750
rect 108080 171686 108132 171692
rect 105962 171032 106018 171041
rect 105962 170967 106018 170976
rect 177552 170497 177580 173046
rect 177736 171721 177764 175834
rect 177828 172809 177856 178554
rect 178104 174033 178132 180322
rect 179654 178920 179710 178929
rect 179654 178855 179710 178864
rect 179668 178618 179696 178855
rect 179656 178612 179708 178618
rect 179656 178554 179708 178560
rect 179654 176472 179710 176481
rect 179654 176407 179710 176416
rect 179668 175898 179696 176407
rect 179656 175892 179708 175898
rect 179656 175834 179708 175840
rect 180312 175626 180340 183479
rect 204508 178249 204536 187868
rect 207268 183009 207296 192319
rect 225194 187352 225250 187361
rect 225194 187287 225250 187296
rect 207254 183000 207310 183009
rect 207254 182935 207310 182944
rect 225208 179745 225236 187287
rect 225194 179736 225250 179745
rect 225194 179671 225250 179680
rect 204494 178240 204550 178249
rect 204494 178175 204550 178184
rect 201090 177696 201146 177705
rect 201090 177631 201146 177640
rect 180300 175620 180352 175626
rect 180300 175562 180352 175568
rect 179654 174160 179710 174169
rect 179654 174095 179710 174104
rect 178090 174024 178146 174033
rect 178090 173959 178146 173968
rect 179668 173110 179696 174095
rect 179656 173104 179708 173110
rect 179656 173046 179708 173052
rect 177814 172800 177870 172809
rect 177814 172735 177870 172744
rect 179654 171848 179710 171857
rect 179654 171783 179710 171792
rect 179668 171750 179696 171783
rect 178184 171744 178236 171750
rect 177722 171712 177778 171721
rect 178184 171686 178236 171692
rect 179656 171744 179708 171750
rect 179656 171686 179708 171692
rect 177722 171647 177778 171656
rect 177538 170488 177594 170497
rect 177538 170423 177594 170432
rect 105686 169944 105742 169953
rect 105686 169879 105742 169888
rect 178196 169409 178224 171686
rect 178182 169400 178238 169409
rect 178182 169335 178238 169344
rect 106606 167360 106662 167369
rect 106606 167295 106662 167304
rect 106514 166952 106570 166961
rect 106514 166887 106570 166896
rect 106528 166802 106556 166887
rect 106620 166802 106648 167295
rect 106528 166774 106648 166802
rect 201104 166174 201132 177631
rect 223538 169264 223594 169273
rect 223538 169199 223594 169208
rect 223552 169166 223580 169199
rect 222804 169160 222856 169166
rect 222724 169120 222804 169148
rect 201092 166168 201144 166174
rect 201092 166110 201144 166116
rect 204496 166168 204548 166174
rect 222724 166122 222752 169120
rect 222804 169102 222856 169108
rect 223540 169160 223592 169166
rect 223540 169102 223592 169108
rect 204496 166110 204548 166116
rect 177170 166000 177226 166009
rect 177170 165935 177226 165944
rect 105226 165456 105282 165465
rect 105226 165391 105282 165400
rect 105240 165290 105268 165391
rect 177184 165358 177212 165935
rect 177172 165352 177224 165358
rect 177172 165294 177224 165300
rect 179564 165352 179616 165358
rect 179564 165294 179616 165300
rect 105228 165284 105280 165290
rect 105228 165226 105280 165232
rect 107804 165284 107856 165290
rect 107804 165226 107856 165232
rect 32638 164912 32694 164921
rect 32638 164847 32694 164856
rect 37422 164912 37478 164921
rect 37422 164847 37478 164856
rect 59594 164912 59650 164921
rect 59594 164847 59650 164856
rect 37436 164814 37464 164847
rect 59608 164814 59636 164847
rect 28868 164808 28920 164814
rect 28868 164750 28920 164756
rect 37424 164808 37476 164814
rect 37424 164750 37476 164756
rect 54812 164808 54864 164814
rect 54812 164750 54864 164756
rect 59596 164808 59648 164814
rect 107816 164785 107844 165226
rect 179576 164785 179604 165294
rect 204508 164921 204536 166110
rect 222632 166094 222752 166122
rect 200998 164912 201054 164921
rect 200998 164847 201054 164856
rect 204494 164912 204550 164921
rect 204494 164847 204550 164856
rect 59596 164750 59648 164756
rect 107802 164776 107858 164785
rect 12214 159336 12270 159345
rect 12214 159271 12270 159280
rect 12122 149408 12178 149417
rect 12122 149343 12178 149352
rect 12122 127784 12178 127793
rect 12122 127719 12178 127728
rect 12030 105752 12086 105761
rect 12030 105687 12086 105696
rect 12136 95833 12164 127719
rect 12228 106169 12256 159271
rect 28880 153746 28908 164750
rect 28696 153718 28908 153746
rect 28696 145230 28724 153718
rect 31994 151584 32050 151593
rect 31994 151519 32050 151528
rect 22244 145224 22296 145230
rect 21948 145172 22244 145178
rect 21948 145166 22296 145172
rect 28684 145224 28736 145230
rect 28684 145166 28736 145172
rect 21948 145150 22284 145166
rect 16612 144878 16764 144906
rect 27284 144878 27620 144906
rect 16736 142646 16764 144878
rect 16724 142640 16776 142646
rect 16724 142582 16776 142588
rect 27592 142510 27620 144878
rect 31904 142640 31956 142646
rect 31904 142582 31956 142588
rect 27580 142504 27632 142510
rect 27580 142446 27632 142452
rect 31916 142306 31944 142582
rect 32008 142322 32036 151519
rect 54824 151026 54852 164750
rect 107802 164711 107858 164720
rect 177538 164776 177594 164785
rect 177538 164711 177594 164720
rect 179562 164776 179618 164785
rect 179562 164711 179618 164720
rect 105778 164232 105834 164241
rect 105778 164167 105834 164176
rect 105594 163552 105650 163561
rect 105594 163487 105596 163496
rect 105648 163487 105650 163496
rect 105596 163458 105648 163464
rect 105792 163454 105820 164167
rect 176986 163688 177042 163697
rect 177552 163658 177580 164711
rect 176986 163623 177042 163632
rect 177540 163652 177592 163658
rect 107436 163516 107488 163522
rect 107436 163458 107488 163464
rect 105780 163448 105832 163454
rect 105780 163390 105832 163396
rect 105686 162328 105742 162337
rect 105686 162263 105742 162272
rect 105700 162094 105728 162263
rect 105688 162088 105740 162094
rect 105688 162030 105740 162036
rect 105226 161104 105282 161113
rect 105226 161039 105228 161048
rect 105280 161039 105282 161048
rect 105228 161010 105280 161016
rect 107448 160025 107476 163458
rect 177000 163454 177028 163623
rect 177540 163594 177592 163600
rect 179564 163652 179616 163658
rect 179564 163594 179616 163600
rect 107804 163448 107856 163454
rect 107804 163390 107856 163396
rect 176988 163448 177040 163454
rect 176988 163390 177040 163396
rect 179196 163448 179248 163454
rect 179196 163390 179248 163396
rect 107816 162473 107844 163390
rect 176986 162600 177042 162609
rect 176986 162535 177042 162544
rect 107802 162464 107858 162473
rect 107802 162399 107858 162408
rect 177000 162094 177028 162535
rect 107804 162088 107856 162094
rect 107804 162030 107856 162036
rect 176988 162088 177040 162094
rect 176988 162030 177040 162036
rect 107712 161068 107764 161074
rect 107712 161010 107764 161016
rect 107434 160016 107490 160025
rect 107434 159951 107490 159960
rect 105594 159744 105650 159753
rect 105594 159679 105650 159688
rect 105608 159578 105636 159679
rect 105596 159572 105648 159578
rect 105596 159514 105648 159520
rect 107620 159572 107672 159578
rect 107620 159514 107672 159520
rect 105778 158520 105834 158529
rect 105778 158455 105834 158464
rect 105792 158354 105820 158455
rect 105780 158348 105832 158354
rect 105780 158290 105832 158296
rect 106146 157976 106202 157985
rect 106146 157911 106148 157920
rect 106200 157911 106202 157920
rect 106148 157882 106200 157888
rect 106146 156752 106202 156761
rect 106146 156687 106148 156696
rect 106200 156687 106202 156696
rect 106148 156658 106200 156664
rect 105778 155392 105834 155401
rect 105778 155327 105780 155336
rect 105832 155327 105834 155336
rect 105780 155298 105832 155304
rect 57478 154848 57534 154857
rect 57478 154783 57534 154792
rect 57492 151554 57520 154783
rect 106422 154168 106478 154177
rect 106478 154126 106556 154154
rect 106422 154103 106478 154112
rect 105226 151720 105282 151729
rect 105226 151655 105282 151664
rect 59594 151584 59650 151593
rect 57480 151548 57532 151554
rect 59594 151519 59596 151528
rect 57480 151490 57532 151496
rect 59648 151519 59650 151528
rect 59596 151490 59648 151496
rect 54824 150998 54944 151026
rect 39092 142714 39120 144892
rect 34112 142708 34164 142714
rect 34112 142650 34164 142656
rect 39080 142708 39132 142714
rect 39080 142650 39132 142656
rect 39264 142708 39316 142714
rect 39264 142650 39316 142656
rect 31904 142300 31956 142306
rect 32008 142294 32956 142322
rect 31904 142242 31956 142248
rect 31916 141393 31944 142242
rect 32928 141778 32956 142294
rect 34124 141778 34152 142650
rect 34664 142640 34716 142646
rect 34664 142582 34716 142588
rect 34676 141778 34704 142582
rect 37240 142572 37292 142578
rect 37240 142514 37292 142520
rect 36596 142436 36648 142442
rect 36596 142378 36648 142384
rect 32928 141750 33218 141778
rect 33862 141750 34152 141778
rect 34506 141750 34704 141778
rect 35242 141762 35624 141778
rect 36608 141764 36636 142378
rect 37252 141764 37280 142514
rect 38620 142232 38672 142238
rect 38620 142174 38672 142180
rect 37884 142164 37936 142170
rect 37884 142106 37936 142112
rect 37896 141764 37924 142106
rect 38632 141764 38660 142174
rect 39276 141764 39304 142650
rect 39460 142646 39488 144892
rect 39448 142640 39500 142646
rect 39448 142582 39500 142588
rect 39828 141762 39856 144892
rect 40000 142300 40052 142306
rect 40000 142242 40052 142248
rect 40012 141764 40040 142242
rect 35242 141756 35636 141762
rect 35242 141750 35584 141756
rect 35584 141698 35636 141704
rect 39816 141756 39868 141762
rect 39816 141698 39868 141704
rect 35952 141688 36004 141694
rect 35886 141636 35952 141642
rect 35886 141630 36004 141636
rect 40184 141688 40236 141694
rect 40288 141676 40316 144892
rect 40380 144878 40670 144906
rect 40380 142442 40408 144878
rect 40644 144204 40696 144210
rect 40644 144146 40696 144152
rect 40368 142436 40420 142442
rect 40368 142378 40420 142384
rect 40656 141764 40684 144146
rect 41024 142578 41052 144892
rect 41288 144136 41340 144142
rect 41288 144078 41340 144084
rect 41012 142572 41064 142578
rect 41012 142514 41064 142520
rect 41300 141764 41328 144078
rect 41484 142170 41512 144892
rect 41852 142238 41880 144892
rect 42220 142714 42248 144892
rect 42312 144878 42694 144906
rect 42208 142708 42260 142714
rect 42208 142650 42260 142656
rect 42312 142306 42340 144878
rect 43048 144210 43076 144892
rect 43036 144204 43088 144210
rect 43036 144146 43088 144152
rect 43416 144142 43444 144892
rect 43404 144136 43456 144142
rect 43404 144078 43456 144084
rect 43404 142708 43456 142714
rect 43404 142650 43456 142656
rect 42668 142640 42720 142646
rect 42668 142582 42720 142588
rect 42300 142300 42352 142306
rect 42300 142242 42352 142248
rect 41840 142232 41892 142238
rect 41840 142174 41892 142180
rect 41472 142164 41524 142170
rect 41472 142106 41524 142112
rect 42024 142164 42076 142170
rect 42024 142106 42076 142112
rect 42036 141764 42064 142106
rect 42680 141764 42708 142582
rect 43416 141764 43444 142650
rect 43876 142170 43904 144892
rect 44244 142646 44272 144892
rect 44612 142714 44640 144892
rect 44704 144878 45086 144906
rect 45164 144878 45454 144906
rect 45624 144878 45822 144906
rect 44600 142708 44652 142714
rect 44600 142650 44652 142656
rect 44232 142640 44284 142646
rect 44232 142582 44284 142588
rect 43864 142164 43916 142170
rect 43864 142106 43916 142112
rect 44704 141914 44732 144878
rect 44520 141886 44732 141914
rect 44520 141778 44548 141886
rect 45164 141778 45192 144878
rect 45624 141778 45652 144878
rect 46268 141778 46296 144892
rect 44074 141750 44548 141778
rect 44810 141750 45192 141778
rect 45454 141750 45652 141778
rect 46098 141750 46296 141778
rect 46636 141778 46664 144892
rect 47096 141778 47124 144892
rect 47478 144878 47768 144906
rect 47740 141778 47768 144878
rect 47832 142646 47860 144892
rect 48292 142714 48320 144892
rect 48280 142708 48332 142714
rect 48280 142650 48332 142656
rect 47820 142640 47872 142646
rect 47820 142582 47872 142588
rect 48660 142442 48688 144892
rect 48832 142640 48884 142646
rect 48832 142582 48884 142588
rect 48648 142436 48700 142442
rect 48648 142378 48700 142384
rect 46636 141750 46834 141778
rect 47096 141750 47478 141778
rect 47740 141750 48214 141778
rect 48844 141764 48872 142582
rect 49028 142238 49056 144892
rect 49502 144878 49792 144906
rect 49476 142708 49528 142714
rect 49476 142650 49528 142656
rect 49016 142232 49068 142238
rect 49016 142174 49068 142180
rect 49488 141764 49516 142650
rect 49764 142646 49792 144878
rect 49752 142640 49804 142646
rect 49752 142582 49804 142588
rect 49856 142102 49884 144892
rect 50224 142578 50252 144892
rect 50212 142572 50264 142578
rect 50212 142514 50264 142520
rect 50684 142510 50712 144892
rect 51052 142714 51080 144892
rect 51040 142708 51092 142714
rect 51040 142650 51092 142656
rect 50672 142504 50724 142510
rect 50672 142446 50724 142452
rect 50212 142436 50264 142442
rect 50212 142378 50264 142384
rect 49844 142096 49896 142102
rect 49844 142038 49896 142044
rect 50224 141764 50252 142378
rect 51420 142306 51448 144892
rect 51592 142640 51644 142646
rect 51592 142582 51644 142588
rect 51408 142300 51460 142306
rect 51408 142242 51460 142248
rect 50856 142232 50908 142238
rect 50856 142174 50908 142180
rect 50868 141764 50896 142174
rect 51604 141764 51632 142582
rect 51880 142374 51908 144892
rect 52248 142442 52276 144892
rect 52236 142436 52288 142442
rect 52236 142378 52288 142384
rect 51868 142368 51920 142374
rect 51868 142310 51920 142316
rect 52236 142232 52288 142238
rect 52236 142174 52288 142180
rect 52248 141764 52276 142174
rect 52616 142034 52644 144892
rect 53076 142646 53104 144892
rect 53064 142640 53116 142646
rect 53064 142582 53116 142588
rect 53444 142578 53472 144892
rect 53812 142714 53840 144892
rect 54272 144210 54300 144892
rect 54260 144204 54312 144210
rect 54260 144146 54312 144152
rect 54640 144142 54668 144892
rect 54628 144136 54680 144142
rect 54628 144078 54680 144084
rect 53800 142708 53852 142714
rect 53800 142650 53852 142656
rect 52972 142572 53024 142578
rect 52972 142514 53024 142520
rect 53432 142572 53484 142578
rect 53432 142514 53484 142520
rect 52604 142028 52656 142034
rect 52604 141970 52656 141976
rect 52984 141764 53012 142514
rect 53616 142504 53668 142510
rect 53616 142446 53668 142452
rect 54260 142504 54312 142510
rect 54260 142446 54312 142452
rect 53628 141764 53656 142446
rect 54272 141764 54300 142446
rect 54916 142170 54944 150998
rect 56100 142436 56152 142442
rect 56100 142378 56152 142384
rect 55364 142368 55416 142374
rect 55364 142310 55416 142316
rect 54996 142300 55048 142306
rect 54996 142242 55048 142248
rect 54904 142164 54956 142170
rect 54904 142106 54956 142112
rect 55008 141764 55036 142242
rect 55376 141778 55404 142310
rect 56112 141778 56140 142378
rect 57492 142102 57520 151490
rect 105134 149680 105190 149689
rect 105134 149615 105190 149624
rect 59780 144204 59832 144210
rect 59780 144146 59832 144152
rect 58676 142708 58728 142714
rect 58676 142650 58728 142656
rect 57664 142640 57716 142646
rect 57664 142582 57716 142588
rect 57480 142096 57532 142102
rect 57480 142038 57532 142044
rect 57020 142028 57072 142034
rect 57020 141970 57072 141976
rect 55376 141750 55666 141778
rect 56112 141750 56402 141778
rect 57032 141764 57060 141970
rect 57676 141764 57704 142582
rect 58124 142572 58176 142578
rect 58124 142514 58176 142520
rect 58136 141778 58164 142514
rect 58688 141778 58716 142650
rect 58136 141750 58426 141778
rect 58688 141750 59070 141778
rect 59792 141764 59820 144146
rect 60424 144136 60476 144142
rect 60424 144078 60476 144084
rect 60436 141764 60464 144078
rect 62816 142708 62868 142714
rect 62816 142650 62868 142656
rect 62356 142300 62408 142306
rect 62356 142242 62408 142248
rect 40236 141648 40316 141676
rect 40184 141630 40236 141636
rect 35886 141614 35992 141630
rect 31902 141384 31958 141393
rect 31902 141319 31958 141328
rect 62368 137721 62396 142242
rect 62828 142073 62856 142650
rect 63472 142306 63500 144892
rect 63460 142300 63512 142306
rect 63460 142242 63512 142248
rect 64576 142170 64604 144892
rect 65128 144878 65694 144906
rect 66600 144878 66798 144906
rect 63460 142164 63512 142170
rect 63460 142106 63512 142112
rect 64564 142164 64616 142170
rect 64564 142106 64616 142112
rect 62814 142064 62870 142073
rect 62814 141999 62870 142008
rect 62816 141280 62868 141286
rect 62816 141222 62868 141228
rect 62724 141212 62776 141218
rect 62724 141154 62776 141160
rect 62736 140713 62764 141154
rect 62828 140985 62856 141222
rect 62814 140976 62870 140985
rect 62814 140911 62870 140920
rect 62722 140704 62778 140713
rect 62722 140639 62778 140648
rect 62816 139920 62868 139926
rect 62816 139862 62868 139868
rect 62724 139784 62776 139790
rect 62828 139761 62856 139862
rect 62724 139726 62776 139732
rect 62814 139752 62870 139761
rect 62736 138945 62764 139726
rect 62814 139687 62870 139696
rect 62816 139648 62868 139654
rect 62816 139590 62868 139596
rect 62828 139489 62856 139590
rect 62814 139480 62870 139489
rect 62814 139415 62870 139424
rect 62722 138936 62778 138945
rect 62722 138871 62778 138880
rect 62908 138696 62960 138702
rect 62908 138638 62960 138644
rect 62816 138628 62868 138634
rect 62816 138570 62868 138576
rect 62354 137712 62410 137721
rect 62354 137647 62410 137656
rect 62724 137268 62776 137274
rect 62724 137210 62776 137216
rect 62632 137200 62684 137206
rect 30522 137168 30578 137177
rect 62632 137142 62684 137148
rect 30522 137103 30578 137112
rect 30430 127784 30486 127793
rect 30430 127719 30486 127728
rect 30444 114358 30472 127719
rect 30432 114352 30484 114358
rect 30432 114294 30484 114300
rect 12214 106160 12270 106169
rect 12214 106095 12270 106104
rect 12122 95824 12178 95833
rect 12122 95759 12178 95768
rect 28512 90342 28908 90370
rect 28512 88874 28540 90342
rect 28880 90286 28908 90342
rect 28868 90280 28920 90286
rect 28868 90222 28920 90228
rect 28512 88846 28632 88874
rect 28604 79218 28632 88846
rect 28604 79190 28724 79218
rect 12030 75152 12086 75161
rect 12030 75087 12086 75096
rect 11938 62912 11994 62921
rect 11938 62847 11994 62856
rect 12044 41297 12072 75087
rect 16598 70650 16626 70908
rect 21948 70894 22284 70922
rect 27284 70894 27620 70922
rect 16598 70622 16672 70650
rect 16644 69478 16672 70622
rect 22256 69546 22284 70894
rect 22244 69540 22296 69546
rect 22244 69482 22296 69488
rect 16632 69472 16684 69478
rect 16632 69414 16684 69420
rect 27592 68798 27620 70894
rect 28696 69546 28724 79190
rect 30536 77842 30564 137103
rect 62644 135409 62672 137142
rect 62736 135681 62764 137210
rect 62828 137177 62856 138570
rect 62814 137168 62870 137177
rect 62814 137103 62870 137112
rect 62920 136633 62948 138638
rect 63472 138401 63500 142106
rect 65128 139790 65156 144878
rect 66496 142708 66548 142714
rect 66496 142650 66548 142656
rect 66508 139926 66536 142650
rect 66496 139920 66548 139926
rect 66496 139862 66548 139868
rect 65116 139784 65168 139790
rect 65116 139726 65168 139732
rect 66600 139654 66628 144878
rect 67888 142714 67916 144892
rect 68072 144878 69006 144906
rect 69268 144878 70110 144906
rect 67876 142708 67928 142714
rect 67876 142650 67928 142656
rect 68072 141218 68100 144878
rect 69164 142436 69216 142442
rect 69164 142378 69216 142384
rect 68060 141212 68112 141218
rect 68060 141154 68112 141160
rect 69176 139738 69204 142378
rect 69268 141286 69296 144878
rect 71200 142578 71228 144892
rect 71188 142572 71240 142578
rect 71188 142514 71240 142520
rect 72304 142442 72332 144892
rect 72844 142708 72896 142714
rect 72844 142650 72896 142656
rect 72292 142436 72344 142442
rect 72292 142378 72344 142384
rect 71004 141892 71056 141898
rect 71004 141834 71056 141840
rect 69256 141280 69308 141286
rect 69256 141222 69308 141228
rect 71016 139738 71044 141834
rect 72856 139738 72884 142650
rect 73408 141898 73436 144892
rect 74512 142714 74540 144892
rect 75616 142714 75644 144892
rect 76260 144878 76826 144906
rect 77930 144878 78128 144906
rect 79034 144878 80060 144906
rect 74500 142708 74552 142714
rect 74500 142650 74552 142656
rect 74776 142708 74828 142714
rect 74776 142650 74828 142656
rect 75604 142708 75656 142714
rect 75604 142650 75656 142656
rect 73396 141892 73448 141898
rect 73396 141834 73448 141840
rect 74788 141370 74816 142650
rect 74696 141342 74816 141370
rect 74696 139738 74724 141342
rect 68868 139710 69204 139738
rect 70708 139710 71044 139738
rect 72548 139710 72884 139738
rect 74480 139710 74724 139738
rect 76260 139738 76288 144878
rect 78100 139738 78128 144878
rect 80032 139738 80060 144878
rect 80124 142714 80152 144892
rect 80112 142708 80164 142714
rect 80112 142650 80164 142656
rect 81228 142646 81256 144892
rect 81676 142708 81728 142714
rect 81676 142650 81728 142656
rect 81216 142640 81268 142646
rect 81216 142582 81268 142588
rect 81688 139738 81716 142650
rect 82332 141558 82360 144892
rect 83436 142034 83464 144892
rect 84540 142714 84568 144892
rect 84528 142708 84580 142714
rect 84528 142650 84580 142656
rect 83516 142640 83568 142646
rect 83516 142582 83568 142588
rect 83424 142028 83476 142034
rect 83424 141970 83476 141976
rect 82320 141552 82372 141558
rect 82320 141494 82372 141500
rect 83528 139738 83556 142582
rect 85644 142442 85672 144892
rect 86748 142646 86776 144892
rect 86736 142640 86788 142646
rect 86736 142582 86788 142588
rect 85632 142436 85684 142442
rect 85632 142378 85684 142384
rect 87852 142170 87880 144892
rect 87840 142164 87892 142170
rect 87840 142106 87892 142112
rect 88956 142034 88984 144892
rect 89128 142708 89180 142714
rect 89128 142650 89180 142656
rect 87288 142028 87340 142034
rect 87288 141970 87340 141976
rect 88944 142028 88996 142034
rect 88944 141970 88996 141976
rect 85356 141552 85408 141558
rect 85356 141494 85408 141500
rect 85368 139738 85396 141494
rect 87300 139738 87328 141970
rect 89140 139738 89168 142650
rect 90152 141354 90180 144892
rect 90968 142436 91020 142442
rect 90968 142378 91020 142384
rect 90140 141348 90192 141354
rect 90140 141290 90192 141296
rect 90980 139738 91008 142378
rect 91256 141937 91284 144892
rect 91242 141928 91298 141937
rect 91242 141863 91298 141872
rect 92360 141354 92388 144892
rect 92808 142640 92860 142646
rect 92808 142582 92860 142588
rect 92348 141348 92400 141354
rect 92348 141290 92400 141296
rect 92820 139738 92848 142582
rect 93464 141354 93492 144892
rect 94108 144878 94582 144906
rect 95580 144878 95686 144906
rect 93452 141348 93504 141354
rect 93452 141290 93504 141296
rect 94108 139790 94136 144878
rect 95476 142708 95528 142714
rect 95476 142650 95528 142656
rect 94740 142164 94792 142170
rect 94740 142106 94792 142112
rect 94096 139784 94148 139790
rect 76260 139710 76320 139738
rect 78100 139710 78160 139738
rect 80032 139710 80092 139738
rect 81688 139710 81932 139738
rect 83528 139710 83864 139738
rect 85368 139710 85704 139738
rect 87300 139710 87544 139738
rect 89140 139710 89476 139738
rect 90980 139710 91316 139738
rect 92820 139710 93156 139738
rect 94096 139726 94148 139732
rect 94752 139738 94780 142106
rect 95488 139926 95516 142650
rect 95476 139920 95528 139926
rect 95476 139862 95528 139868
rect 95580 139858 95608 144878
rect 96776 142714 96804 144892
rect 96764 142708 96816 142714
rect 96764 142650 96816 142656
rect 96856 142028 96908 142034
rect 96856 141970 96908 141976
rect 95568 139852 95620 139858
rect 95568 139794 95620 139800
rect 96868 139738 96896 141970
rect 97880 141354 97908 144892
rect 98984 142374 99012 144892
rect 98972 142368 99024 142374
rect 98972 142310 99024 142316
rect 100088 142034 100116 144892
rect 101192 142481 101220 144892
rect 102296 142617 102324 144892
rect 102282 142608 102338 142617
rect 102282 142543 102338 142552
rect 102296 142510 102324 142543
rect 102284 142504 102336 142510
rect 101178 142472 101234 142481
rect 102284 142446 102336 142452
rect 101178 142407 101234 142416
rect 100076 142028 100128 142034
rect 100076 141970 100128 141976
rect 101192 141966 101220 142407
rect 102284 142368 102336 142374
rect 102284 142310 102336 142316
rect 101180 141960 101232 141966
rect 101180 141902 101232 141908
rect 97868 141348 97920 141354
rect 97868 141290 97920 141296
rect 94752 139710 95088 139738
rect 96868 139710 96928 139738
rect 66588 139648 66640 139654
rect 66588 139590 66640 139596
rect 66218 139480 66274 139489
rect 66218 139415 66274 139424
rect 66232 138634 66260 139415
rect 100626 139072 100682 139081
rect 100626 139007 100682 139016
rect 66402 138936 66458 138945
rect 66402 138871 66458 138880
rect 66416 138702 66444 138871
rect 66404 138696 66456 138702
rect 66404 138638 66456 138644
rect 100534 138664 100590 138673
rect 66220 138628 66272 138634
rect 100534 138599 100590 138608
rect 66220 138570 66272 138576
rect 63458 138392 63514 138401
rect 63458 138327 63514 138336
rect 66218 138256 66274 138265
rect 66218 138191 66274 138200
rect 66232 137274 66260 138191
rect 66402 137712 66458 137721
rect 66402 137647 66458 137656
rect 66220 137268 66272 137274
rect 66220 137210 66272 137216
rect 66416 137206 66444 137647
rect 100350 137304 100406 137313
rect 100350 137239 100406 137248
rect 66404 137200 66456 137206
rect 66404 137142 66456 137148
rect 62906 136624 62962 136633
rect 62906 136559 62962 136568
rect 66034 136488 66090 136497
rect 66034 136423 66090 136432
rect 65022 136216 65078 136225
rect 65022 136151 65078 136160
rect 62908 135908 62960 135914
rect 62908 135850 62960 135856
rect 62722 135672 62778 135681
rect 62722 135607 62778 135616
rect 62630 135400 62686 135409
rect 62630 135335 62686 135344
rect 62724 135024 62776 135030
rect 62724 134966 62776 134972
rect 62736 134865 62764 134966
rect 62722 134856 62778 134865
rect 62722 134791 62778 134800
rect 62816 134684 62868 134690
rect 62816 134626 62868 134632
rect 62724 134480 62776 134486
rect 62724 134422 62776 134428
rect 62736 132553 62764 134422
rect 62828 132825 62856 134626
rect 62920 134321 62948 135850
rect 63000 135840 63052 135846
rect 63000 135782 63052 135788
rect 62906 134312 62962 134321
rect 62906 134247 62962 134256
rect 63012 133641 63040 135782
rect 65036 135030 65064 136151
rect 66048 135914 66076 136423
rect 66402 135944 66458 135953
rect 66036 135908 66088 135914
rect 66402 135879 66458 135888
rect 66036 135850 66088 135856
rect 66416 135846 66444 135879
rect 66404 135840 66456 135846
rect 66404 135782 66456 135788
rect 100364 135642 100392 137239
rect 100548 136730 100576 138599
rect 100640 137070 100668 139007
rect 100996 138424 101048 138430
rect 100994 138392 100996 138401
rect 101048 138392 101050 138401
rect 100994 138327 101050 138336
rect 100718 137848 100774 137857
rect 100718 137783 100774 137792
rect 100628 137064 100680 137070
rect 100628 137006 100680 137012
rect 100536 136724 100588 136730
rect 100536 136666 100588 136672
rect 100626 136080 100682 136089
rect 100626 136015 100628 136024
rect 100680 136015 100682 136024
rect 100628 135986 100680 135992
rect 100732 135778 100760 137783
rect 100902 136624 100958 136633
rect 100958 136582 101036 136610
rect 100902 136559 100958 136568
rect 100902 135944 100958 135953
rect 100902 135879 100904 135888
rect 100956 135879 100958 135888
rect 100904 135850 100956 135856
rect 100720 135772 100772 135778
rect 100720 135714 100772 135720
rect 101008 135710 101036 136582
rect 100996 135704 101048 135710
rect 100996 135646 101048 135652
rect 100352 135636 100404 135642
rect 100352 135578 100404 135584
rect 66310 135264 66366 135273
rect 66310 135199 66366 135208
rect 65024 135024 65076 135030
rect 65024 134966 65076 134972
rect 66324 134690 66352 135199
rect 100074 134856 100130 134865
rect 100074 134791 100130 134800
rect 66402 134720 66458 134729
rect 66312 134684 66364 134690
rect 100088 134690 100116 134791
rect 100902 134720 100958 134729
rect 66402 134655 66458 134664
rect 100076 134684 100128 134690
rect 66312 134626 66364 134632
rect 66416 134486 66444 134655
rect 100958 134678 101036 134706
rect 100902 134655 100958 134664
rect 100076 134626 100128 134632
rect 66404 134480 66456 134486
rect 66404 134422 66456 134428
rect 65850 134176 65906 134185
rect 65850 134111 65906 134120
rect 62998 133632 63054 133641
rect 62998 133567 63054 133576
rect 63552 133120 63604 133126
rect 63552 133062 63604 133068
rect 62814 132816 62870 132825
rect 62814 132751 62870 132760
rect 62722 132544 62778 132553
rect 62722 132479 62778 132488
rect 63276 131760 63328 131766
rect 63276 131702 63328 131708
rect 62816 130808 62868 130814
rect 62814 130776 62816 130785
rect 62868 130776 62870 130785
rect 62814 130711 62870 130720
rect 62632 130400 62684 130406
rect 62632 130342 62684 130348
rect 62644 128473 62672 130342
rect 62724 130332 62776 130338
rect 62724 130274 62776 130280
rect 62736 128745 62764 130274
rect 63288 129561 63316 131702
rect 63460 131692 63512 131698
rect 63460 131634 63512 131640
rect 63472 130241 63500 131634
rect 63564 131329 63592 133062
rect 65864 133058 65892 134111
rect 100074 133632 100130 133641
rect 100074 133567 100130 133576
rect 66402 133496 66458 133505
rect 66402 133431 66458 133440
rect 66416 133126 66444 133431
rect 66404 133120 66456 133126
rect 66404 133062 66456 133068
rect 100088 133058 100116 133567
rect 100902 133224 100958 133233
rect 100902 133159 100904 133168
rect 100956 133159 100958 133168
rect 100904 133130 100956 133136
rect 63644 133052 63696 133058
rect 63644 132994 63696 133000
rect 65852 133052 65904 133058
rect 65852 132994 65904 133000
rect 100076 133052 100128 133058
rect 100076 132994 100128 133000
rect 63656 131601 63684 132994
rect 101008 132990 101036 134678
rect 101192 134593 101220 141902
rect 102296 140985 102324 142310
rect 105148 142050 105176 149615
rect 105240 144142 105268 151655
rect 105410 151040 105466 151049
rect 105410 150975 105466 150984
rect 105228 144136 105280 144142
rect 105228 144078 105280 144084
rect 103112 142028 103164 142034
rect 105148 142022 105222 142050
rect 103112 141970 103164 141976
rect 103124 141529 103152 141970
rect 105194 141764 105222 142022
rect 105424 141778 105452 150975
rect 105962 147232 106018 147241
rect 105962 147167 106018 147176
rect 105976 147066 106004 147167
rect 105964 147060 106016 147066
rect 105964 147002 106016 147008
rect 106528 144142 106556 154126
rect 107632 152953 107660 159514
rect 107724 155401 107752 161010
rect 107816 157713 107844 162030
rect 177538 161376 177594 161385
rect 177538 161311 177594 161320
rect 177552 160938 177580 161311
rect 177540 160932 177592 160938
rect 177540 160874 177592 160880
rect 177354 160288 177410 160297
rect 177354 160223 177410 160232
rect 177368 159306 177396 160223
rect 179208 160025 179236 163390
rect 179576 162473 179604 163594
rect 179562 162464 179618 162473
rect 179562 162399 179618 162408
rect 179564 162088 179616 162094
rect 179564 162030 179616 162036
rect 179472 160932 179524 160938
rect 179472 160874 179524 160880
rect 179194 160016 179250 160025
rect 179194 159951 179250 159960
rect 177356 159300 177408 159306
rect 177356 159242 177408 159248
rect 179380 159300 179432 159306
rect 179380 159242 179432 159248
rect 177630 159064 177686 159073
rect 177630 158999 177686 159008
rect 108724 158348 108776 158354
rect 108724 158290 108776 158296
rect 108632 157940 108684 157946
rect 108632 157882 108684 157888
rect 107802 157704 107858 157713
rect 107802 157639 107858 157648
rect 108540 156716 108592 156722
rect 108540 156658 108592 156664
rect 107710 155392 107766 155401
rect 107710 155327 107766 155336
rect 107896 155356 107948 155362
rect 107896 155298 107948 155304
rect 106606 152944 106662 152953
rect 106606 152879 106662 152888
rect 107618 152944 107674 152953
rect 107618 152879 107674 152888
rect 105964 144136 106016 144142
rect 105964 144078 106016 144084
rect 106516 144136 106568 144142
rect 106516 144078 106568 144084
rect 105976 141778 106004 144078
rect 106620 141778 106648 152879
rect 106698 148320 106754 148329
rect 106698 148255 106754 148264
rect 106712 144890 106740 148255
rect 106700 144884 106752 144890
rect 106700 144826 106752 144832
rect 107160 144136 107212 144142
rect 107160 144078 107212 144084
rect 107172 141778 107200 144078
rect 107908 141778 107936 155298
rect 108356 147060 108408 147066
rect 108356 147002 108408 147008
rect 108368 141778 108396 147002
rect 108552 146017 108580 156658
rect 108644 148329 108672 157882
rect 108736 150641 108764 158290
rect 177644 158014 177672 158999
rect 177632 158008 177684 158014
rect 177632 157950 177684 157956
rect 178182 157976 178238 157985
rect 178182 157911 178184 157920
rect 178236 157911 178238 157920
rect 178184 157882 178236 157888
rect 177354 156888 177410 156897
rect 177354 156823 177410 156832
rect 177368 156518 177396 156823
rect 177356 156512 177408 156518
rect 177356 156454 177408 156460
rect 178090 155664 178146 155673
rect 178090 155599 178146 155608
rect 178104 155158 178132 155599
rect 178092 155152 178144 155158
rect 178092 155094 178144 155100
rect 178274 154576 178330 154585
rect 178274 154511 178330 154520
rect 132366 151584 132422 151593
rect 132366 151519 132422 151528
rect 108722 150632 108778 150641
rect 108722 150567 108778 150576
rect 108630 148320 108686 148329
rect 108630 148255 108686 148264
rect 108538 146008 108594 146017
rect 108538 145943 108594 145952
rect 109276 144884 109328 144890
rect 109276 144826 109328 144832
rect 109288 141778 109316 144826
rect 111128 142714 111156 144892
rect 110104 142708 110156 142714
rect 110104 142650 110156 142656
rect 111116 142708 111168 142714
rect 111116 142650 111168 142656
rect 110116 141778 110144 142650
rect 111496 142034 111524 144892
rect 111588 144878 111878 144906
rect 111956 144878 112338 144906
rect 112416 144878 112706 144906
rect 110426 142028 110478 142034
rect 110426 141970 110478 141976
rect 111484 142028 111536 142034
rect 111484 141970 111536 141976
rect 105424 141750 105760 141778
rect 105976 141750 106312 141778
rect 106620 141750 106956 141778
rect 107172 141750 107508 141778
rect 107908 141750 108060 141778
rect 108368 141750 108704 141778
rect 109256 141750 109316 141778
rect 109808 141750 110144 141778
rect 110438 141764 110466 141970
rect 111588 141880 111616 144878
rect 111404 141852 111616 141880
rect 111404 141778 111432 141852
rect 111956 141778 111984 144878
rect 112416 141778 112444 144878
rect 113060 141778 113088 144892
rect 113520 142034 113548 144892
rect 113902 144878 114008 144906
rect 113278 142028 113330 142034
rect 113278 141970 113330 141976
rect 113508 142028 113560 142034
rect 113508 141970 113560 141976
rect 111004 141750 111432 141778
rect 111556 141750 111984 141778
rect 112200 141750 112444 141778
rect 112752 141750 113088 141778
rect 113290 141764 113318 141970
rect 113980 141642 114008 144878
rect 114256 141778 114284 144892
rect 114716 141778 114744 144892
rect 115098 144878 115388 144906
rect 115466 144878 115848 144906
rect 115926 144878 116216 144906
rect 115360 141778 115388 144878
rect 115820 141778 115848 144878
rect 116188 141914 116216 144878
rect 116280 142034 116308 144892
rect 116648 142306 116676 144892
rect 116636 142300 116688 142306
rect 116636 142242 116688 142248
rect 117108 142170 117136 144892
rect 117476 142442 117504 144892
rect 117464 142436 117516 142442
rect 117464 142378 117516 142384
rect 117648 142300 117700 142306
rect 117648 142242 117700 142248
rect 117096 142164 117148 142170
rect 117096 142106 117148 142112
rect 116268 142028 116320 142034
rect 116268 141970 116320 141976
rect 117418 142028 117470 142034
rect 117418 141970 117470 141976
rect 116188 141886 116400 141914
rect 116372 141778 116400 141886
rect 114256 141750 114500 141778
rect 114716 141750 115052 141778
rect 115360 141750 115696 141778
rect 115820 141750 116248 141778
rect 116372 141750 116800 141778
rect 117430 141764 117458 141970
rect 117660 141778 117688 142242
rect 117844 142034 117872 144892
rect 118304 142170 118332 144892
rect 118686 144878 118976 144906
rect 118948 144142 118976 144878
rect 118936 144136 118988 144142
rect 118936 144078 118988 144084
rect 119132 142646 119160 144892
rect 119120 142640 119172 142646
rect 119120 142582 119172 142588
rect 119500 142442 119528 144892
rect 119882 144878 120264 144906
rect 120236 144210 120264 144878
rect 120224 144204 120276 144210
rect 120224 144146 120276 144152
rect 118844 142436 118896 142442
rect 118844 142378 118896 142384
rect 119488 142436 119540 142442
rect 119488 142378 119540 142384
rect 118200 142164 118252 142170
rect 118200 142106 118252 142112
rect 118292 142164 118344 142170
rect 118292 142106 118344 142112
rect 117832 142028 117884 142034
rect 117832 141970 117884 141976
rect 118212 141778 118240 142106
rect 118856 141778 118884 142378
rect 120328 142306 120356 144892
rect 120592 144136 120644 144142
rect 120592 144078 120644 144084
rect 120316 142300 120368 142306
rect 120316 142242 120368 142248
rect 119948 142164 120000 142170
rect 119948 142106 120000 142112
rect 119718 142028 119770 142034
rect 119718 141970 119770 141976
rect 117660 141750 117996 141778
rect 118212 141750 118548 141778
rect 118856 141750 119192 141778
rect 119730 141764 119758 141970
rect 119960 141778 119988 142106
rect 120604 141778 120632 144078
rect 120696 142714 120724 144892
rect 120684 142708 120736 142714
rect 120684 142650 120736 142656
rect 121064 142578 121092 144892
rect 121144 142640 121196 142646
rect 121144 142582 121196 142588
rect 121052 142572 121104 142578
rect 121052 142514 121104 142520
rect 121156 141778 121184 142582
rect 121524 142238 121552 144892
rect 121696 142436 121748 142442
rect 121696 142378 121748 142384
rect 121512 142232 121564 142238
rect 121512 142174 121564 142180
rect 121708 141778 121736 142378
rect 121892 142034 121920 144892
rect 121880 142028 121932 142034
rect 121880 141970 121932 141976
rect 119960 141750 120296 141778
rect 120604 141750 120940 141778
rect 121156 141750 121492 141778
rect 121708 141750 122044 141778
rect 122260 141762 122288 144892
rect 122734 144878 122932 144906
rect 123102 144878 123392 144906
rect 123470 144878 123760 144906
rect 122340 144204 122392 144210
rect 122340 144146 122392 144152
rect 122352 141778 122380 144146
rect 122904 141830 122932 144878
rect 123076 142300 123128 142306
rect 123076 142242 123128 142248
rect 122892 141824 122944 141830
rect 122248 141756 122300 141762
rect 122352 141750 122688 141778
rect 122892 141766 122944 141772
rect 123088 141778 123116 142242
rect 123364 142170 123392 144878
rect 123444 142708 123496 142714
rect 123444 142650 123496 142656
rect 123352 142164 123404 142170
rect 123352 142106 123404 142112
rect 123456 141778 123484 142650
rect 123732 142374 123760 144878
rect 123916 142646 123944 144892
rect 123904 142640 123956 142646
rect 123904 142582 123956 142588
rect 124284 142442 124312 144892
rect 124652 142578 124680 144892
rect 124456 142572 124508 142578
rect 124456 142514 124508 142520
rect 124640 142572 124692 142578
rect 124640 142514 124692 142520
rect 124272 142436 124324 142442
rect 124272 142378 124324 142384
rect 123720 142368 123772 142374
rect 123720 142310 123772 142316
rect 124468 141778 124496 142514
rect 125112 142306 125140 144892
rect 125480 142714 125508 144892
rect 125848 144278 125876 144892
rect 125836 144272 125888 144278
rect 125836 144214 125888 144220
rect 126308 144142 126336 144892
rect 126676 144210 126704 144892
rect 131448 144272 131500 144278
rect 131448 144214 131500 144220
rect 126664 144204 126716 144210
rect 126664 144146 126716 144152
rect 126296 144136 126348 144142
rect 126296 144078 126348 144084
rect 125468 142708 125520 142714
rect 125468 142650 125520 142656
rect 130436 142708 130488 142714
rect 130436 142650 130488 142656
rect 128136 142640 128188 142646
rect 128136 142582 128188 142588
rect 127584 142368 127636 142374
rect 127584 142310 127636 142316
rect 125100 142300 125152 142306
rect 125100 142242 125152 142248
rect 124640 142232 124692 142238
rect 124640 142174 124692 142180
rect 123088 141750 123240 141778
rect 123456 141750 123792 141778
rect 124436 141750 124496 141778
rect 124652 141778 124680 142174
rect 126940 142164 126992 142170
rect 126940 142106 126992 142112
rect 125514 142028 125566 142034
rect 125514 141970 125566 141976
rect 124652 141750 124988 141778
rect 125526 141764 125554 141970
rect 126388 141824 126440 141830
rect 125848 141762 126184 141778
rect 126952 141778 126980 142106
rect 127596 141778 127624 142310
rect 128148 141778 128176 142582
rect 129332 142572 129384 142578
rect 129332 142514 129384 142520
rect 128688 142436 128740 142442
rect 128688 142378 128740 142384
rect 128700 141778 128728 142378
rect 129344 141778 129372 142514
rect 129884 142300 129936 142306
rect 129884 142242 129936 142248
rect 129896 141778 129924 142242
rect 130448 141778 130476 142650
rect 126440 141772 126736 141778
rect 126388 141766 126736 141772
rect 125836 141756 126184 141762
rect 122248 141698 122300 141704
rect 125888 141750 126184 141756
rect 126400 141750 126736 141766
rect 126952 141750 127288 141778
rect 127596 141750 127932 141778
rect 128148 141750 128484 141778
rect 128700 141750 129036 141778
rect 129344 141750 129680 141778
rect 129896 141750 130232 141778
rect 130448 141750 130784 141778
rect 125836 141698 125888 141704
rect 131460 141642 131488 144214
rect 132184 144204 132236 144210
rect 132184 144146 132236 144152
rect 131632 144136 131684 144142
rect 131632 144078 131684 144084
rect 131644 141778 131672 144078
rect 132196 141778 132224 144146
rect 132380 141898 132408 151519
rect 176894 151176 176950 151185
rect 176894 151111 176950 151120
rect 176908 150074 176936 151111
rect 176908 150046 177488 150074
rect 177170 149952 177226 149961
rect 177170 149887 177226 149896
rect 174134 144920 174190 144929
rect 135522 144878 135628 144906
rect 135496 144476 135548 144482
rect 135496 144418 135548 144424
rect 132644 144136 132696 144142
rect 132644 144078 132696 144084
rect 132656 143462 132684 144078
rect 132644 143456 132696 143462
rect 132644 143398 132696 143404
rect 134116 142572 134168 142578
rect 134116 142514 134168 142520
rect 134128 142073 134156 142514
rect 135508 142238 135536 144418
rect 134484 142232 134536 142238
rect 134484 142174 134536 142180
rect 135496 142232 135548 142238
rect 135496 142174 135548 142180
rect 134114 142064 134170 142073
rect 134114 141999 134170 142008
rect 134300 142028 134352 142034
rect 134300 141970 134352 141976
rect 132368 141892 132420 141898
rect 132368 141834 132420 141840
rect 131644 141750 131980 141778
rect 132196 141750 132532 141778
rect 113948 141614 114008 141642
rect 131428 141614 131488 141642
rect 103110 141520 103166 141529
rect 103110 141455 103166 141464
rect 132644 141348 132696 141354
rect 132644 141290 132696 141296
rect 102376 141212 102428 141218
rect 102376 141154 102428 141160
rect 102282 140976 102338 140985
rect 102282 140911 102338 140920
rect 102388 140441 102416 141154
rect 102374 140432 102430 140441
rect 102374 140367 102430 140376
rect 102376 139920 102428 139926
rect 102376 139862 102428 139868
rect 102388 139761 102416 139862
rect 102468 139852 102520 139858
rect 102468 139794 102520 139800
rect 102374 139752 102430 139761
rect 102374 139687 102430 139696
rect 102480 139217 102508 139794
rect 102560 139784 102612 139790
rect 102560 139726 102612 139732
rect 102466 139208 102522 139217
rect 102466 139143 102522 139152
rect 102572 138673 102600 139726
rect 102558 138664 102614 138673
rect 102558 138599 102614 138608
rect 102376 138560 102428 138566
rect 102376 138502 102428 138508
rect 102388 137993 102416 138502
rect 102468 138492 102520 138498
rect 102468 138434 102520 138440
rect 102374 137984 102430 137993
rect 102374 137919 102430 137928
rect 102480 137449 102508 138434
rect 102466 137440 102522 137449
rect 102466 137375 102522 137384
rect 102836 137064 102888 137070
rect 102836 137006 102888 137012
rect 102848 136905 102876 137006
rect 102834 136896 102890 136905
rect 102834 136831 102890 136840
rect 102468 136724 102520 136730
rect 102468 136666 102520 136672
rect 102480 136361 102508 136666
rect 102466 136352 102522 136361
rect 102466 136287 102522 136296
rect 102192 136044 102244 136050
rect 102192 135986 102244 135992
rect 102100 135908 102152 135914
rect 102100 135850 102152 135856
rect 101178 134584 101234 134593
rect 101178 134519 101234 134528
rect 102112 133369 102140 135850
rect 102204 133913 102232 135986
rect 102376 135772 102428 135778
rect 102376 135714 102428 135720
rect 102388 135681 102416 135714
rect 102468 135704 102520 135710
rect 102374 135672 102430 135681
rect 102468 135646 102520 135652
rect 102374 135607 102430 135616
rect 102284 134684 102336 134690
rect 102284 134626 102336 134632
rect 102190 133904 102246 133913
rect 102190 133839 102246 133848
rect 102098 133360 102154 133369
rect 102098 133295 102154 133304
rect 102192 133188 102244 133194
rect 102192 133130 102244 133136
rect 102100 133052 102152 133058
rect 102100 132994 102152 133000
rect 100996 132984 101048 132990
rect 100996 132926 101048 132932
rect 65022 132544 65078 132553
rect 65022 132479 65078 132488
rect 63642 131592 63698 131601
rect 63642 131527 63698 131536
rect 63550 131320 63606 131329
rect 63550 131255 63606 131264
rect 65036 130814 65064 132479
rect 100442 132408 100498 132417
rect 100442 132343 100498 132352
rect 66402 132272 66458 132281
rect 66402 132207 66458 132216
rect 65668 131760 65720 131766
rect 65666 131728 65668 131737
rect 65720 131728 65722 131737
rect 66416 131698 66444 132207
rect 100456 131698 100484 132343
rect 100902 132000 100958 132009
rect 100958 131958 101036 131986
rect 100902 131935 100958 131944
rect 100904 131760 100956 131766
rect 100902 131728 100904 131737
rect 100956 131728 100958 131737
rect 65666 131663 65722 131672
rect 66404 131692 66456 131698
rect 66404 131634 66456 131640
rect 100444 131692 100496 131698
rect 100902 131663 100958 131672
rect 100444 131634 100496 131640
rect 66310 131184 66366 131193
rect 66310 131119 66366 131128
rect 65024 130808 65076 130814
rect 65024 130750 65076 130756
rect 66324 130338 66352 131119
rect 100442 130640 100498 130649
rect 100442 130575 100444 130584
rect 100496 130575 100498 130584
rect 100444 130546 100496 130552
rect 66402 130504 66458 130513
rect 66402 130439 66458 130448
rect 100902 130504 100958 130513
rect 100902 130439 100958 130448
rect 66416 130406 66444 130439
rect 100916 130406 100944 130439
rect 66404 130400 66456 130406
rect 66404 130342 66456 130348
rect 100904 130400 100956 130406
rect 100904 130342 100956 130348
rect 66312 130332 66364 130338
rect 66312 130274 66364 130280
rect 101008 130270 101036 131958
rect 102008 131760 102060 131766
rect 102008 131702 102060 131708
rect 100996 130264 101048 130270
rect 63458 130232 63514 130241
rect 100996 130206 101048 130212
rect 63458 130167 63514 130176
rect 65482 129960 65538 129969
rect 65482 129895 65538 129904
rect 63274 129552 63330 129561
rect 63274 129487 63330 129496
rect 62908 129040 62960 129046
rect 62908 128982 62960 128988
rect 62816 128972 62868 128978
rect 62816 128914 62868 128920
rect 62722 128736 62778 128745
rect 62722 128671 62778 128680
rect 62630 128464 62686 128473
rect 62630 128399 62686 128408
rect 62632 127544 62684 127550
rect 62828 127521 62856 128914
rect 62632 127486 62684 127492
rect 62814 127512 62870 127521
rect 62644 126025 62672 127486
rect 62814 127447 62870 127456
rect 62920 127249 62948 128982
rect 65496 128978 65524 129895
rect 100074 129416 100130 129425
rect 100074 129351 100130 129360
rect 66402 129280 66458 129289
rect 66402 129215 66458 129224
rect 66416 129046 66444 129215
rect 66404 129040 66456 129046
rect 66404 128982 66456 128988
rect 100088 128978 100116 129351
rect 102020 129289 102048 131702
rect 102112 131601 102140 132994
rect 102098 131592 102154 131601
rect 102098 131527 102154 131536
rect 102204 131057 102232 133130
rect 102296 132825 102324 134626
rect 102480 134593 102508 135646
rect 102652 135636 102704 135642
rect 102652 135578 102704 135584
rect 102664 135137 102692 135578
rect 102650 135128 102706 135137
rect 102650 135063 102706 135072
rect 102466 134584 102522 134593
rect 102466 134519 102522 134528
rect 102376 132984 102428 132990
rect 102376 132926 102428 132932
rect 102282 132816 102338 132825
rect 102282 132751 102338 132760
rect 102388 132281 102416 132926
rect 102374 132272 102430 132281
rect 102374 132207 102430 132216
rect 102376 131624 102428 131630
rect 102376 131566 102428 131572
rect 102190 131048 102246 131057
rect 102190 130983 102246 130992
rect 102284 130604 102336 130610
rect 102284 130546 102336 130552
rect 102192 130400 102244 130406
rect 102192 130342 102244 130348
rect 102006 129280 102062 129289
rect 102006 129215 102062 129224
rect 100904 129040 100956 129046
rect 100902 129008 100904 129017
rect 102008 129040 102060 129046
rect 100956 129008 100958 129017
rect 65484 128972 65536 128978
rect 65484 128914 65536 128920
rect 100076 128972 100128 128978
rect 102008 128982 102060 128988
rect 100902 128943 100958 128952
rect 101916 128972 101968 128978
rect 100076 128914 100128 128920
rect 101916 128914 101968 128920
rect 100350 128328 100406 128337
rect 100350 128263 100406 128272
rect 66402 128192 66458 128201
rect 66402 128127 66458 128136
rect 65022 127920 65078 127929
rect 65022 127855 65078 127864
rect 62906 127240 62962 127249
rect 62906 127175 62962 127184
rect 65036 126938 65064 127855
rect 66416 127550 66444 128127
rect 100364 127890 100392 128263
rect 101928 127906 101956 128914
rect 102020 128042 102048 128982
rect 102204 128201 102232 130342
rect 102296 128745 102324 130546
rect 102388 130513 102416 131566
rect 102374 130504 102430 130513
rect 102374 130439 102430 130448
rect 102376 130264 102428 130270
rect 102376 130206 102428 130212
rect 102388 129833 102416 130206
rect 102374 129824 102430 129833
rect 102374 129759 102430 129768
rect 102282 128736 102338 128745
rect 102282 128671 102338 128680
rect 102190 128192 102246 128201
rect 102190 128127 102246 128136
rect 102020 128014 102232 128042
rect 100352 127884 100404 127890
rect 101928 127878 102140 127906
rect 100352 127826 100404 127832
rect 100534 127648 100590 127657
rect 100534 127583 100536 127592
rect 100588 127583 100590 127592
rect 102008 127612 102060 127618
rect 100536 127554 100588 127560
rect 102008 127554 102060 127560
rect 66404 127544 66456 127550
rect 66404 127486 66456 127492
rect 100442 127104 100498 127113
rect 100442 127039 100498 127048
rect 66310 126968 66366 126977
rect 62816 126932 62868 126938
rect 62816 126874 62868 126880
rect 65024 126932 65076 126938
rect 66310 126903 66366 126912
rect 65024 126874 65076 126880
rect 62828 126705 62856 126874
rect 62814 126696 62870 126705
rect 62814 126631 62870 126640
rect 65022 126560 65078 126569
rect 65022 126495 65078 126504
rect 62724 126252 62776 126258
rect 62724 126194 62776 126200
rect 62630 126016 62686 126025
rect 62630 125951 62686 125960
rect 62632 124824 62684 124830
rect 62632 124766 62684 124772
rect 62644 123169 62672 124766
rect 62736 124665 62764 126194
rect 62908 126184 62960 126190
rect 62908 126126 62960 126132
rect 62816 125572 62868 125578
rect 62816 125514 62868 125520
rect 62828 125481 62856 125514
rect 62814 125472 62870 125481
rect 62814 125407 62870 125416
rect 62722 124656 62778 124665
rect 62722 124591 62778 124600
rect 62920 124393 62948 126126
rect 65036 125578 65064 126495
rect 66324 126258 66352 126903
rect 66402 126288 66458 126297
rect 66312 126252 66364 126258
rect 66402 126223 66458 126232
rect 66312 126194 66364 126200
rect 66416 126190 66444 126223
rect 100456 126190 100484 127039
rect 100902 126424 100958 126433
rect 100902 126359 100958 126368
rect 100812 126320 100864 126326
rect 100810 126288 100812 126297
rect 100864 126288 100866 126297
rect 100916 126258 100944 126359
rect 100810 126223 100866 126232
rect 100904 126252 100956 126258
rect 100904 126194 100956 126200
rect 66404 126184 66456 126190
rect 66404 126126 66456 126132
rect 100444 126184 100496 126190
rect 100444 126126 100496 126132
rect 102020 125753 102048 127554
rect 102112 127521 102140 127878
rect 102098 127512 102154 127521
rect 102098 127447 102154 127456
rect 102204 126977 102232 128014
rect 102284 127884 102336 127890
rect 102284 127826 102336 127832
rect 102190 126968 102246 126977
rect 102190 126903 102246 126912
rect 102296 126433 102324 127826
rect 102282 126424 102338 126433
rect 102282 126359 102338 126368
rect 102100 126320 102152 126326
rect 102100 126262 102152 126268
rect 66310 125744 66366 125753
rect 66310 125679 66366 125688
rect 102006 125744 102062 125753
rect 102006 125679 102062 125688
rect 65024 125572 65076 125578
rect 65024 125514 65076 125520
rect 66324 124801 66352 125679
rect 100902 125336 100958 125345
rect 100902 125271 100958 125280
rect 66402 125200 66458 125209
rect 66402 125135 66458 125144
rect 66416 124830 66444 125135
rect 100810 124928 100866 124937
rect 100810 124863 100812 124872
rect 100864 124863 100866 124872
rect 100812 124834 100864 124840
rect 100916 124830 100944 125271
rect 66404 124824 66456 124830
rect 65022 124792 65078 124801
rect 65022 124727 65078 124736
rect 66310 124792 66366 124801
rect 66404 124766 66456 124772
rect 100904 124824 100956 124830
rect 100904 124766 100956 124772
rect 66310 124727 66366 124736
rect 62906 124384 62962 124393
rect 62906 124319 62962 124328
rect 65036 123810 65064 124727
rect 100258 124112 100314 124121
rect 100258 124047 100314 124056
rect 66402 123976 66458 123985
rect 66402 123911 66458 123920
rect 62816 123804 62868 123810
rect 62816 123746 62868 123752
rect 65024 123804 65076 123810
rect 65024 123746 65076 123752
rect 62828 123713 62856 123746
rect 62814 123704 62870 123713
rect 62814 123639 62870 123648
rect 65022 123704 65078 123713
rect 65022 123639 65078 123648
rect 63552 123396 63604 123402
rect 63552 123338 63604 123344
rect 62630 123160 62686 123169
rect 62630 123095 62686 123104
rect 62816 122716 62868 122722
rect 62816 122658 62868 122664
rect 62828 122625 62856 122658
rect 62814 122616 62870 122625
rect 62814 122551 62870 122560
rect 63460 122104 63512 122110
rect 63460 122046 63512 122052
rect 62816 121492 62868 121498
rect 62816 121434 62868 121440
rect 62828 121401 62856 121434
rect 62814 121392 62870 121401
rect 62814 121327 62870 121336
rect 63472 120585 63500 122046
rect 63564 121673 63592 123338
rect 65036 122722 65064 123639
rect 66416 123402 66444 123911
rect 100272 123402 100300 124047
rect 102112 123985 102140 126262
rect 102284 126252 102336 126258
rect 102284 126194 102336 126200
rect 102192 124892 102244 124898
rect 102192 124834 102244 124840
rect 102098 123976 102154 123985
rect 102098 123911 102154 123920
rect 100902 123432 100958 123441
rect 66404 123396 66456 123402
rect 66404 123338 66456 123344
rect 100260 123396 100312 123402
rect 100958 123390 101036 123418
rect 100902 123367 100958 123376
rect 100260 123338 100312 123344
rect 100166 122888 100222 122897
rect 100166 122823 100222 122832
rect 66310 122752 66366 122761
rect 65024 122716 65076 122722
rect 66310 122687 66366 122696
rect 65024 122658 65076 122664
rect 65022 122480 65078 122489
rect 65022 122415 65078 122424
rect 63644 122036 63696 122042
rect 63644 121978 63696 121984
rect 63550 121664 63606 121673
rect 63550 121599 63606 121608
rect 63458 120576 63514 120585
rect 63458 120511 63514 120520
rect 63656 120313 63684 121978
rect 65036 121498 65064 122415
rect 66324 122110 66352 122687
rect 100180 122246 100208 122823
rect 100626 122480 100682 122489
rect 100626 122415 100682 122424
rect 100168 122240 100220 122246
rect 66402 122208 66458 122217
rect 100168 122182 100220 122188
rect 66402 122143 66458 122152
rect 66312 122104 66364 122110
rect 66312 122046 66364 122052
rect 66416 122042 66444 122143
rect 100640 122042 100668 122415
rect 100902 122208 100958 122217
rect 100902 122143 100904 122152
rect 100956 122143 100958 122152
rect 100904 122114 100956 122120
rect 66404 122036 66456 122042
rect 66404 121978 66456 121984
rect 100628 122036 100680 122042
rect 100628 121978 100680 121984
rect 101008 121974 101036 123390
rect 101822 123024 101878 123033
rect 101822 122959 101878 122968
rect 100996 121968 101048 121974
rect 100996 121910 101048 121916
rect 65024 121492 65076 121498
rect 65024 121434 65076 121440
rect 100074 121120 100130 121129
rect 100074 121055 100130 121064
rect 66218 120984 66274 120993
rect 66218 120919 66274 120928
rect 65022 120712 65078 120721
rect 65022 120647 65078 120656
rect 63642 120304 63698 120313
rect 63642 120239 63698 120248
rect 65036 120002 65064 120647
rect 62816 119996 62868 120002
rect 62816 119938 62868 119944
rect 65024 119996 65076 120002
rect 65024 119938 65076 119944
rect 62828 119633 62856 119938
rect 65482 119760 65538 119769
rect 65482 119695 65538 119704
rect 62814 119624 62870 119633
rect 62814 119559 62870 119568
rect 65022 119488 65078 119497
rect 65022 119423 65078 119432
rect 62908 119316 62960 119322
rect 62908 119258 62960 119264
rect 62724 119180 62776 119186
rect 62724 119122 62776 119128
rect 62736 118817 62764 119122
rect 62722 118808 62778 118817
rect 62722 118743 62778 118752
rect 62816 118772 62868 118778
rect 62816 118714 62868 118720
rect 62828 118545 62856 118714
rect 62814 118536 62870 118545
rect 62814 118471 62870 118480
rect 62724 117888 62776 117894
rect 62920 117865 62948 119258
rect 65036 118778 65064 119423
rect 65496 119322 65524 119695
rect 65484 119316 65536 119322
rect 65484 119258 65536 119264
rect 66232 119186 66260 120919
rect 100088 120682 100116 121055
rect 100902 120984 100958 120993
rect 100902 120919 100904 120928
rect 100956 120919 100958 120928
rect 100904 120890 100956 120896
rect 100076 120676 100128 120682
rect 100076 120618 100128 120624
rect 100442 119896 100498 119905
rect 100442 119831 100498 119840
rect 100456 119322 100484 119831
rect 100902 119352 100958 119361
rect 100444 119316 100496 119322
rect 100958 119310 101036 119338
rect 100902 119287 100958 119296
rect 100444 119258 100496 119264
rect 66402 119216 66458 119225
rect 66220 119180 66272 119186
rect 66402 119151 66458 119160
rect 66220 119122 66272 119128
rect 65024 118772 65076 118778
rect 65024 118714 65076 118720
rect 64930 118536 64986 118545
rect 64930 118471 64986 118480
rect 62724 117830 62776 117836
rect 62906 117856 62962 117865
rect 62736 116233 62764 117830
rect 62906 117791 62962 117800
rect 62816 117344 62868 117350
rect 62814 117312 62816 117321
rect 62868 117312 62870 117321
rect 62814 117247 62870 117256
rect 64944 117214 64972 118471
rect 66416 118273 66444 119151
rect 100626 118672 100682 118681
rect 100626 118607 100682 118616
rect 65022 118264 65078 118273
rect 65022 118199 65078 118208
rect 66402 118264 66458 118273
rect 66402 118199 66458 118208
rect 65036 117350 65064 118199
rect 100640 118166 100668 118607
rect 100628 118160 100680 118166
rect 100258 118128 100314 118137
rect 100628 118102 100680 118108
rect 100258 118063 100314 118072
rect 66402 117992 66458 118001
rect 66402 117927 66458 117936
rect 66416 117894 66444 117927
rect 100272 117894 100300 118063
rect 100534 117992 100590 118001
rect 100534 117927 100590 117936
rect 66404 117888 66456 117894
rect 66404 117830 66456 117836
rect 100260 117888 100312 117894
rect 100260 117830 100312 117836
rect 65024 117344 65076 117350
rect 65024 117286 65076 117292
rect 62816 117208 62868 117214
rect 62816 117150 62868 117156
rect 64932 117208 64984 117214
rect 64932 117150 64984 117156
rect 62828 116777 62856 117150
rect 62814 116768 62870 116777
rect 62814 116703 62870 116712
rect 66402 116768 66458 116777
rect 66402 116703 66458 116712
rect 100258 116768 100314 116777
rect 100258 116703 100260 116712
rect 65022 116496 65078 116505
rect 65022 116431 65078 116440
rect 62722 116224 62778 116233
rect 62722 116159 62778 116168
rect 65036 115786 65064 116431
rect 62816 115780 62868 115786
rect 62816 115722 62868 115728
rect 65024 115780 65076 115786
rect 65024 115722 65076 115728
rect 62828 115553 62856 115722
rect 62814 115544 62870 115553
rect 62814 115479 62870 115488
rect 65022 115136 65078 115145
rect 65022 115071 65078 115080
rect 62816 114896 62868 114902
rect 62816 114838 62868 114844
rect 62828 114737 62856 114838
rect 62814 114728 62870 114737
rect 62814 114663 62870 114672
rect 65036 114630 65064 115071
rect 66416 114902 66444 116703
rect 100312 116703 100314 116712
rect 100260 116674 100312 116680
rect 100548 116398 100576 117927
rect 101008 117758 101036 119310
rect 100996 117752 101048 117758
rect 100996 117694 101048 117700
rect 100902 116904 100958 116913
rect 100902 116839 100958 116848
rect 100916 116534 100944 116839
rect 100904 116528 100956 116534
rect 100904 116470 100956 116476
rect 100536 116392 100588 116398
rect 100536 116334 100588 116340
rect 72856 115910 72916 115938
rect 82516 115910 82852 115938
rect 92728 115910 92880 115938
rect 66404 114896 66456 114902
rect 66404 114838 66456 114844
rect 62816 114624 62868 114630
rect 62816 114566 62868 114572
rect 65024 114624 65076 114630
rect 65024 114566 65076 114572
rect 62828 114465 62856 114566
rect 62814 114456 62870 114465
rect 62814 114391 62870 114400
rect 32008 113870 33218 113898
rect 32008 104265 32036 113870
rect 33848 111638 33876 113884
rect 34492 111774 34520 113884
rect 35228 111910 35256 113884
rect 35216 111904 35268 111910
rect 35216 111846 35268 111852
rect 34480 111768 34532 111774
rect 34480 111710 34532 111716
rect 35872 111706 35900 113884
rect 35860 111700 35912 111706
rect 35860 111642 35912 111648
rect 33836 111632 33888 111638
rect 33836 111574 33888 111580
rect 36608 111230 36636 113884
rect 37252 111298 37280 113884
rect 37896 111570 37924 113884
rect 37884 111564 37936 111570
rect 37884 111506 37936 111512
rect 37240 111292 37292 111298
rect 37240 111234 37292 111240
rect 36596 111224 36648 111230
rect 36596 111166 36648 111172
rect 38632 111094 38660 113884
rect 39080 111632 39132 111638
rect 39080 111574 39132 111580
rect 38620 111088 38672 111094
rect 38620 111030 38672 111036
rect 39092 110756 39120 111574
rect 39276 111502 39304 113884
rect 39816 111904 39868 111910
rect 39816 111846 39868 111852
rect 39448 111768 39500 111774
rect 39448 111710 39500 111716
rect 39264 111496 39316 111502
rect 39264 111438 39316 111444
rect 39460 110756 39488 111710
rect 39828 110756 39856 111846
rect 40012 111434 40040 113884
rect 40276 111700 40328 111706
rect 40276 111642 40328 111648
rect 40000 111428 40052 111434
rect 40000 111370 40052 111376
rect 40288 110756 40316 111642
rect 40656 111366 40684 113884
rect 40644 111360 40696 111366
rect 40644 111302 40696 111308
rect 41012 111292 41064 111298
rect 41012 111234 41064 111240
rect 40644 111224 40696 111230
rect 40644 111166 40696 111172
rect 40656 110756 40684 111166
rect 41024 110756 41052 111234
rect 41300 111230 41328 113884
rect 41472 111564 41524 111570
rect 41472 111506 41524 111512
rect 41288 111224 41340 111230
rect 41288 111166 41340 111172
rect 41484 110756 41512 111506
rect 42036 111162 42064 113884
rect 42208 111496 42260 111502
rect 42208 111438 42260 111444
rect 42024 111156 42076 111162
rect 42024 111098 42076 111104
rect 41840 111088 41892 111094
rect 41840 111030 41892 111036
rect 41852 110756 41880 111030
rect 42220 110756 42248 111438
rect 42300 111428 42352 111434
rect 42300 111370 42352 111376
rect 42312 110770 42340 111370
rect 42680 111026 42708 113884
rect 43416 111366 43444 113884
rect 44074 113870 44364 113898
rect 44810 113870 45192 113898
rect 45454 113870 45744 113898
rect 43036 111360 43088 111366
rect 43036 111302 43088 111308
rect 43404 111360 43456 111366
rect 43404 111302 43456 111308
rect 42668 111020 42720 111026
rect 42668 110962 42720 110968
rect 42312 110742 42694 110770
rect 43048 110756 43076 111302
rect 44336 111230 44364 113870
rect 44600 111360 44652 111366
rect 44600 111302 44652 111308
rect 43404 111224 43456 111230
rect 43404 111166 43456 111172
rect 44324 111224 44376 111230
rect 44324 111166 44376 111172
rect 43416 110756 43444 111166
rect 43864 111156 43916 111162
rect 43864 111098 43916 111104
rect 43876 110756 43904 111098
rect 44232 111020 44284 111026
rect 44232 110962 44284 110968
rect 44244 110756 44272 110962
rect 44612 110756 44640 111302
rect 45060 111224 45112 111230
rect 45060 111166 45112 111172
rect 45072 110756 45100 111166
rect 45164 110770 45192 113870
rect 45716 112130 45744 113870
rect 45716 112102 45836 112130
rect 45164 110742 45454 110770
rect 45808 110756 45836 112102
rect 46084 110770 46112 113884
rect 46820 110770 46848 113884
rect 46084 110742 46282 110770
rect 46650 110742 46848 110770
rect 47188 113870 47478 113898
rect 47740 113870 48214 113898
rect 47188 110634 47216 113870
rect 47740 110770 47768 113870
rect 48280 111428 48332 111434
rect 48280 111370 48332 111376
rect 47820 111360 47872 111366
rect 47820 111302 47872 111308
rect 47478 110742 47768 110770
rect 47832 110756 47860 111302
rect 48292 110756 48320 111370
rect 48844 111366 48872 113884
rect 49488 111434 49516 113884
rect 49476 111428 49528 111434
rect 49476 111370 49528 111376
rect 48832 111360 48884 111366
rect 48832 111302 48884 111308
rect 49844 111360 49896 111366
rect 49844 111302 49896 111308
rect 48648 111292 48700 111298
rect 48648 111234 48700 111240
rect 48660 110756 48688 111234
rect 49476 111224 49528 111230
rect 49476 111166 49528 111172
rect 49016 111088 49068 111094
rect 49016 111030 49068 111036
rect 49028 110756 49056 111030
rect 49488 110756 49516 111166
rect 49856 110756 49884 111302
rect 50224 111298 50252 113884
rect 50672 111428 50724 111434
rect 50672 111370 50724 111376
rect 50212 111292 50264 111298
rect 50212 111234 50264 111240
rect 50212 111156 50264 111162
rect 50212 111098 50264 111104
rect 50224 110756 50252 111098
rect 50684 110756 50712 111370
rect 50868 111094 50896 113884
rect 51040 112108 51092 112114
rect 51040 112050 51092 112056
rect 50856 111088 50908 111094
rect 50856 111030 50908 111036
rect 51052 110756 51080 112050
rect 51408 111292 51460 111298
rect 51408 111234 51460 111240
rect 51420 110756 51448 111234
rect 51604 111230 51632 113884
rect 51868 111972 51920 111978
rect 51868 111914 51920 111920
rect 51592 111224 51644 111230
rect 51592 111166 51644 111172
rect 51880 110756 51908 111914
rect 52248 111366 52276 113884
rect 52604 112176 52656 112182
rect 52604 112118 52656 112124
rect 52512 111904 52564 111910
rect 52512 111846 52564 111852
rect 52236 111360 52288 111366
rect 52236 111302 52288 111308
rect 52524 110770 52552 111846
rect 52262 110742 52552 110770
rect 52616 110756 52644 112118
rect 52984 111162 53012 113884
rect 53064 112040 53116 112046
rect 53064 111982 53116 111988
rect 52972 111156 53024 111162
rect 52972 111098 53024 111104
rect 53076 110756 53104 111982
rect 53432 111700 53484 111706
rect 53432 111642 53484 111648
rect 53444 110756 53472 111642
rect 53628 111434 53656 113884
rect 54272 112114 54300 113884
rect 54260 112108 54312 112114
rect 54260 112050 54312 112056
rect 53800 111836 53852 111842
rect 53800 111778 53852 111784
rect 53616 111428 53668 111434
rect 53616 111370 53668 111376
rect 53812 110756 53840 111778
rect 54260 111768 54312 111774
rect 54260 111710 54312 111716
rect 54272 110756 54300 111710
rect 54628 111632 54680 111638
rect 54628 111574 54680 111580
rect 54640 110756 54668 111574
rect 55008 111298 55036 113884
rect 55652 111978 55680 113884
rect 55640 111972 55692 111978
rect 55640 111914 55692 111920
rect 56388 111910 56416 113884
rect 56926 113232 56982 113241
rect 56926 113167 56982 113176
rect 56376 111904 56428 111910
rect 56376 111846 56428 111852
rect 54996 111292 55048 111298
rect 54996 111234 55048 111240
rect 47110 110606 47216 110634
rect 31994 104256 32050 104265
rect 31994 104191 32050 104200
rect 37422 104256 37478 104265
rect 37422 104191 37478 104200
rect 37436 104090 37464 104191
rect 32640 104084 32692 104090
rect 32640 104026 32692 104032
rect 37424 104084 37476 104090
rect 37424 104026 37476 104032
rect 56836 104084 56888 104090
rect 56836 104026 56888 104032
rect 32652 90937 32680 104026
rect 56848 100865 56876 104026
rect 56834 100856 56890 100865
rect 56834 100791 56890 100800
rect 32638 90928 32694 90937
rect 32638 90863 32694 90872
rect 36410 90928 36466 90937
rect 36410 90863 36466 90872
rect 36424 90286 36452 90863
rect 36412 90280 36464 90286
rect 36412 90222 36464 90228
rect 54812 86132 54864 86138
rect 54812 86074 54864 86080
rect 54824 79270 54852 86074
rect 56940 81961 56968 113167
rect 57032 112182 57060 113884
rect 57020 112176 57072 112182
rect 57020 112118 57072 112124
rect 57676 112046 57704 113884
rect 57664 112040 57716 112046
rect 57664 111982 57716 111988
rect 58412 111706 58440 113884
rect 59056 111842 59084 113884
rect 59044 111836 59096 111842
rect 59044 111778 59096 111784
rect 59792 111774 59820 113884
rect 59780 111768 59832 111774
rect 59780 111710 59832 111716
rect 58400 111700 58452 111706
rect 58400 111642 58452 111648
rect 60436 111638 60464 113884
rect 72014 113232 72070 113241
rect 72014 113167 72070 113176
rect 72028 112998 72056 113167
rect 72856 112998 72884 115910
rect 72016 112992 72068 112998
rect 72016 112934 72068 112940
rect 72844 112992 72896 112998
rect 72844 112934 72896 112940
rect 82516 112794 82544 115910
rect 92728 114358 92756 115910
rect 100902 115544 100958 115553
rect 100902 115479 100904 115488
rect 100956 115479 100958 115488
rect 100904 115450 100956 115456
rect 92716 114352 92768 114358
rect 92716 114294 92768 114300
rect 101836 113785 101864 122959
rect 102204 122897 102232 124834
rect 102296 124665 102324 126194
rect 102376 126116 102428 126122
rect 102376 126058 102428 126064
rect 102388 125209 102416 126058
rect 102374 125200 102430 125209
rect 102374 125135 102430 125144
rect 102376 124756 102428 124762
rect 102376 124698 102428 124704
rect 102282 124656 102338 124665
rect 102282 124591 102338 124600
rect 102388 123441 102416 124698
rect 102374 123432 102430 123441
rect 102284 123396 102336 123402
rect 102374 123367 102430 123376
rect 102284 123338 102336 123344
rect 102190 122888 102246 122897
rect 102190 122823 102246 122832
rect 102296 122353 102324 123338
rect 102282 122344 102338 122353
rect 102282 122279 102338 122288
rect 102284 122240 102336 122246
rect 102284 122182 102336 122188
rect 102008 122172 102060 122178
rect 102008 122114 102060 122120
rect 102020 119905 102048 122114
rect 102100 122036 102152 122042
rect 102100 121978 102152 121984
rect 102112 120585 102140 121978
rect 102296 121129 102324 122182
rect 102376 121968 102428 121974
rect 102376 121910 102428 121916
rect 102388 121673 102416 121910
rect 102374 121664 102430 121673
rect 102374 121599 102430 121608
rect 102282 121120 102338 121129
rect 102282 121055 102338 121064
rect 102192 120948 102244 120954
rect 102192 120890 102244 120896
rect 102098 120576 102154 120585
rect 102098 120511 102154 120520
rect 102006 119896 102062 119905
rect 102006 119831 102062 119840
rect 102204 118817 102232 120890
rect 102376 120608 102428 120614
rect 102376 120550 102428 120556
rect 102388 119361 102416 120550
rect 102374 119352 102430 119361
rect 102284 119316 102336 119322
rect 102374 119287 102430 119296
rect 102284 119258 102336 119264
rect 102190 118808 102246 118817
rect 102190 118743 102246 118752
rect 102296 118273 102324 119258
rect 102282 118264 102338 118273
rect 102282 118199 102338 118208
rect 102284 118160 102336 118166
rect 102284 118102 102336 118108
rect 102296 117049 102324 118102
rect 132656 117826 132684 141290
rect 134312 138945 134340 141970
rect 134298 138936 134354 138945
rect 134298 138871 134354 138880
rect 134496 138401 134524 142174
rect 135600 142102 135628 144878
rect 136336 144878 136626 144906
rect 136888 144878 137730 144906
rect 138268 144878 138834 144906
rect 139648 144878 139938 144906
rect 136336 144482 136364 144878
rect 136324 144476 136376 144482
rect 136324 144418 136376 144424
rect 134576 142096 134628 142102
rect 134576 142038 134628 142044
rect 135588 142096 135640 142102
rect 135588 142038 135640 142044
rect 134482 138392 134538 138401
rect 134482 138327 134538 138336
rect 134588 137721 134616 142038
rect 136888 142034 136916 144878
rect 136876 142028 136928 142034
rect 136876 141970 136928 141976
rect 135404 141144 135456 141150
rect 135404 141086 135456 141092
rect 135416 140985 135444 141086
rect 135402 140976 135458 140985
rect 135402 140911 135458 140920
rect 135404 140736 135456 140742
rect 135402 140704 135404 140713
rect 135456 140704 135458 140713
rect 135402 140639 135458 140648
rect 135404 139852 135456 139858
rect 135404 139794 135456 139800
rect 135416 139761 135444 139794
rect 135402 139752 135458 139761
rect 135402 139687 135458 139696
rect 138268 139518 138296 144878
rect 139648 141370 139676 144878
rect 139556 141342 139676 141370
rect 140832 141348 140884 141354
rect 139556 139858 139584 141342
rect 140832 141290 140884 141296
rect 139544 139852 139596 139858
rect 139544 139794 139596 139800
rect 140844 139724 140872 141290
rect 141028 140742 141056 144892
rect 141120 144878 142146 144906
rect 141120 141150 141148 144878
rect 143236 142578 143264 144892
rect 143224 142572 143276 142578
rect 143224 142514 143276 142520
rect 142672 142232 142724 142238
rect 142672 142174 142724 142180
rect 141108 141144 141160 141150
rect 141108 141086 141160 141092
rect 141016 140736 141068 140742
rect 141016 140678 141068 140684
rect 142684 139724 142712 142174
rect 144340 141354 144368 144892
rect 145444 142238 145472 144892
rect 145432 142232 145484 142238
rect 145432 142174 145484 142180
rect 146548 141694 146576 144892
rect 144512 141688 144564 141694
rect 144512 141630 144564 141636
rect 146536 141688 146588 141694
rect 146536 141630 146588 141636
rect 144328 141348 144380 141354
rect 144328 141290 144380 141296
rect 144524 139724 144552 141630
rect 147652 141558 147680 144892
rect 148296 144878 148862 144906
rect 149966 144878 150164 144906
rect 146444 141552 146496 141558
rect 146444 141494 146496 141500
rect 147640 141552 147692 141558
rect 147640 141494 147692 141500
rect 146456 139724 146484 141494
rect 148296 139724 148324 144878
rect 150136 139724 150164 144878
rect 151056 141558 151084 144892
rect 152160 141830 152188 144892
rect 153264 142714 153292 144892
rect 153252 142708 153304 142714
rect 153252 142650 153304 142656
rect 154368 142646 154396 144892
rect 154356 142640 154408 142646
rect 154356 142582 154408 142588
rect 155472 142578 155500 144892
rect 156576 142714 156604 144892
rect 157694 144878 157984 144906
rect 155828 142708 155880 142714
rect 155828 142650 155880 142656
rect 156564 142708 156616 142714
rect 156564 142650 156616 142656
rect 155460 142572 155512 142578
rect 155460 142514 155512 142520
rect 152148 141824 152200 141830
rect 152148 141766 152200 141772
rect 153896 141824 153948 141830
rect 153896 141766 153948 141772
rect 151044 141552 151096 141558
rect 151044 141494 151096 141500
rect 152056 141552 152108 141558
rect 152056 141494 152108 141500
rect 152068 139724 152096 141494
rect 153908 139724 153936 141766
rect 155840 139724 155868 142650
rect 157668 142640 157720 142646
rect 157668 142582 157720 142588
rect 157680 139724 157708 142582
rect 157956 141626 157984 144878
rect 158784 142170 158812 144892
rect 159508 142572 159560 142578
rect 159508 142514 159560 142520
rect 158772 142164 158824 142170
rect 158772 142106 158824 142112
rect 157944 141620 157996 141626
rect 157944 141562 157996 141568
rect 159520 139724 159548 142514
rect 159888 142442 159916 144892
rect 159876 142436 159928 142442
rect 159876 142378 159928 142384
rect 160992 142374 161020 144892
rect 161440 142708 161492 142714
rect 161440 142650 161492 142656
rect 160980 142368 161032 142374
rect 160980 142310 161032 142316
rect 161452 139724 161480 142650
rect 162188 141937 162216 144892
rect 163292 142646 163320 144892
rect 163280 142640 163332 142646
rect 163280 142582 163332 142588
rect 162174 141928 162230 141937
rect 162174 141863 162230 141872
rect 163280 141620 163332 141626
rect 163280 141562 163332 141568
rect 163292 139724 163320 141562
rect 164396 141354 164424 144892
rect 165120 142164 165172 142170
rect 165120 142106 165172 142112
rect 164384 141348 164436 141354
rect 164384 141290 164436 141296
rect 165132 139724 165160 142106
rect 165500 142102 165528 144892
rect 166604 142170 166632 144892
rect 167052 142436 167104 142442
rect 167052 142378 167104 142384
rect 166592 142164 166644 142170
rect 166592 142106 166644 142112
rect 165488 142096 165540 142102
rect 165488 142038 165540 142044
rect 167064 139724 167092 142378
rect 167708 142306 167736 144892
rect 167696 142300 167748 142306
rect 167696 142242 167748 142248
rect 168812 142034 168840 144892
rect 168892 142368 168944 142374
rect 168892 142310 168944 142316
rect 168800 142028 168852 142034
rect 168800 141970 168852 141976
rect 168904 139724 168932 142310
rect 169916 141422 169944 144892
rect 169904 141416 169956 141422
rect 169904 141358 169956 141364
rect 171020 141354 171048 144892
rect 172124 142238 172152 144892
rect 172112 142232 172164 142238
rect 172112 142174 172164 142180
rect 172848 142028 172900 142034
rect 172848 141970 172900 141976
rect 171008 141348 171060 141354
rect 171008 141290 171060 141296
rect 172860 139926 172888 141970
rect 173228 141966 173256 144892
rect 174134 144855 174190 144864
rect 174148 144142 174176 144855
rect 174136 144136 174188 144142
rect 174136 144078 174188 144084
rect 174332 142510 174360 144892
rect 174412 142640 174464 142646
rect 174412 142582 174464 142588
rect 174320 142504 174372 142510
rect 174320 142446 174372 142452
rect 174320 142300 174372 142306
rect 174320 142242 174372 142248
rect 173216 141960 173268 141966
rect 173216 141902 173268 141908
rect 174228 141280 174280 141286
rect 174228 141222 174280 141228
rect 174240 140713 174268 141222
rect 174226 140704 174282 140713
rect 174226 140639 174282 140648
rect 172848 139920 172900 139926
rect 172848 139862 172900 139868
rect 135404 139512 135456 139518
rect 135402 139480 135404 139489
rect 138256 139512 138308 139518
rect 135456 139480 135458 139489
rect 174332 139489 174360 142242
rect 138256 139454 138308 139460
rect 174318 139480 174374 139489
rect 135402 139415 135458 139424
rect 174318 139415 174374 139424
rect 136874 139072 136930 139081
rect 136874 139007 136930 139016
rect 172478 139072 172534 139081
rect 172478 139007 172534 139016
rect 135128 138696 135180 138702
rect 135128 138638 135180 138644
rect 134574 137712 134630 137721
rect 134574 137647 134630 137656
rect 135140 136633 135168 138638
rect 136888 138634 136916 139007
rect 136966 138936 137022 138945
rect 136966 138871 137022 138880
rect 136980 138702 137008 138871
rect 172492 138770 172520 139007
rect 172662 138800 172718 138809
rect 172480 138764 172532 138770
rect 172662 138735 172718 138744
rect 174228 138764 174280 138770
rect 172480 138706 172532 138712
rect 172676 138702 172704 138735
rect 174228 138706 174280 138712
rect 136968 138696 137020 138702
rect 136968 138638 137020 138644
rect 172664 138696 172716 138702
rect 172664 138638 172716 138644
rect 135404 138628 135456 138634
rect 135404 138570 135456 138576
rect 136876 138628 136928 138634
rect 136876 138570 136928 138576
rect 135220 137268 135272 137274
rect 135220 137210 135272 137216
rect 135126 136624 135182 136633
rect 135126 136559 135182 136568
rect 134944 135908 134996 135914
rect 134944 135850 134996 135856
rect 132920 134480 132972 134486
rect 132920 134422 132972 134428
rect 132932 117894 132960 134422
rect 134956 133641 134984 135850
rect 135128 135840 135180 135846
rect 135128 135782 135180 135788
rect 135036 134956 135088 134962
rect 135036 134898 135088 134904
rect 135048 134865 135076 134898
rect 135034 134856 135090 134865
rect 135034 134791 135090 134800
rect 135140 134321 135168 135782
rect 135232 135409 135260 137210
rect 135312 137200 135364 137206
rect 135312 137142 135364 137148
rect 135324 135681 135352 137142
rect 135416 136905 135444 138570
rect 174136 138492 174188 138498
rect 174136 138434 174188 138440
rect 136874 137848 136930 137857
rect 136874 137783 136930 137792
rect 172202 137848 172258 137857
rect 172202 137783 172258 137792
rect 136888 137206 136916 137783
rect 136966 137304 137022 137313
rect 136966 137239 136968 137248
rect 137020 137239 137022 137248
rect 136968 137210 137020 137216
rect 172216 137206 172244 137783
rect 174148 137721 174176 138434
rect 174134 137712 174190 137721
rect 174134 137647 174190 137656
rect 172662 137304 172718 137313
rect 172662 137239 172664 137248
rect 172716 137239 172718 137248
rect 174044 137268 174096 137274
rect 172664 137210 172716 137216
rect 174044 137210 174096 137216
rect 136876 137200 136928 137206
rect 136876 137142 136928 137148
rect 172204 137200 172256 137206
rect 172204 137142 172256 137148
rect 173952 137200 174004 137206
rect 173952 137142 174004 137148
rect 135402 136896 135458 136905
rect 135402 136831 135458 136840
rect 136782 136624 136838 136633
rect 136782 136559 136838 136568
rect 172018 136624 172074 136633
rect 172018 136559 172074 136568
rect 135310 135672 135366 135681
rect 135310 135607 135366 135616
rect 135218 135400 135274 135409
rect 135218 135335 135274 135344
rect 136796 134962 136824 136559
rect 136874 136080 136930 136089
rect 136874 136015 136930 136024
rect 136888 135846 136916 136015
rect 136966 135944 137022 135953
rect 136966 135879 136968 135888
rect 137020 135879 137022 135888
rect 136968 135850 137020 135856
rect 172032 135846 172060 136559
rect 172570 136216 172626 136225
rect 172570 136151 172572 136160
rect 172624 136151 172626 136160
rect 172572 136122 172624 136128
rect 172662 136080 172718 136089
rect 172662 136015 172664 136024
rect 172716 136015 172718 136024
rect 172664 135986 172716 135992
rect 136876 135840 136928 135846
rect 136876 135782 136928 135788
rect 172020 135840 172072 135846
rect 172020 135782 172072 135788
rect 173964 135681 173992 137142
rect 173950 135672 174006 135681
rect 173950 135607 174006 135616
rect 174056 135409 174084 137210
rect 174240 137177 174268 138706
rect 174320 138696 174372 138702
rect 174320 138638 174372 138644
rect 174226 137168 174282 137177
rect 174226 137103 174282 137112
rect 174332 136633 174360 138638
rect 174318 136624 174374 136633
rect 174318 136559 174374 136568
rect 174136 136180 174188 136186
rect 174136 136122 174188 136128
rect 174042 135400 174098 135409
rect 174042 135335 174098 135344
rect 136784 134956 136836 134962
rect 136784 134898 136836 134904
rect 136874 134856 136930 134865
rect 136874 134791 136930 134800
rect 171834 134856 171890 134865
rect 171834 134791 171890 134800
rect 135220 134548 135272 134554
rect 135220 134490 135272 134496
rect 135126 134312 135182 134321
rect 135126 134247 135182 134256
rect 134942 133632 134998 133641
rect 134942 133567 134998 133576
rect 135128 133120 135180 133126
rect 135128 133062 135180 133068
rect 134944 131760 134996 131766
rect 134944 131702 134996 131708
rect 134956 129561 134984 131702
rect 135140 131601 135168 133062
rect 135232 132553 135260 134490
rect 136888 134486 136916 134791
rect 136966 134720 137022 134729
rect 171848 134690 171876 134791
rect 136966 134655 137022 134664
rect 171836 134684 171888 134690
rect 136980 134554 137008 134655
rect 171836 134626 171888 134632
rect 172662 134584 172718 134593
rect 136968 134548 137020 134554
rect 172662 134519 172664 134528
rect 136968 134490 137020 134496
rect 172716 134519 172718 134528
rect 172664 134490 172716 134496
rect 135404 134480 135456 134486
rect 135404 134422 135456 134428
rect 136876 134480 136928 134486
rect 136876 134422 136928 134428
rect 135312 133052 135364 133058
rect 135312 132994 135364 133000
rect 135218 132544 135274 132553
rect 135218 132479 135274 132488
rect 135220 131692 135272 131698
rect 135220 131634 135272 131640
rect 135126 131592 135182 131601
rect 135126 131527 135182 131536
rect 135036 130400 135088 130406
rect 135036 130342 135088 130348
rect 134942 129552 134998 129561
rect 134942 129487 134998 129496
rect 135048 128473 135076 130342
rect 135232 130241 135260 131634
rect 135324 131329 135352 132994
rect 135416 132825 135444 134422
rect 174148 134321 174176 136122
rect 174320 135840 174372 135846
rect 174320 135782 174372 135788
rect 174332 134865 174360 135782
rect 174318 134856 174374 134865
rect 174318 134791 174374 134800
rect 174228 134684 174280 134690
rect 174228 134626 174280 134632
rect 174134 134312 174190 134321
rect 174134 134247 174190 134256
rect 136966 133632 137022 133641
rect 136966 133567 137022 133576
rect 172202 133632 172258 133641
rect 172202 133567 172204 133576
rect 136980 133126 137008 133567
rect 172256 133567 172258 133576
rect 172204 133538 172256 133544
rect 172662 133224 172718 133233
rect 172662 133159 172718 133168
rect 172676 133126 172704 133159
rect 136968 133120 137020 133126
rect 136874 133088 136930 133097
rect 136968 133062 137020 133068
rect 172664 133120 172716 133126
rect 172664 133062 172716 133068
rect 136874 133023 136876 133032
rect 136928 133023 136930 133032
rect 136876 132994 136928 133000
rect 174240 132825 174268 134626
rect 174320 134548 174372 134554
rect 174320 134490 174372 134496
rect 135402 132816 135458 132825
rect 135402 132751 135458 132760
rect 174226 132816 174282 132825
rect 174226 132751 174282 132760
rect 174332 132553 174360 134490
rect 174318 132544 174374 132553
rect 174318 132479 174374 132488
rect 136782 132408 136838 132417
rect 136782 132343 136838 132352
rect 172386 132408 172442 132417
rect 172386 132343 172442 132352
rect 135310 131320 135366 131329
rect 135310 131255 135366 131264
rect 136796 131086 136824 132343
rect 136874 132000 136930 132009
rect 136874 131935 136930 131944
rect 172018 132000 172074 132009
rect 172400 131970 172428 132343
rect 172018 131935 172074 131944
rect 172388 131964 172440 131970
rect 136888 131698 136916 131935
rect 172032 131766 172060 131935
rect 172388 131906 172440 131912
rect 172662 131864 172718 131873
rect 172662 131799 172664 131808
rect 172716 131799 172718 131808
rect 172664 131770 172716 131776
rect 136968 131760 137020 131766
rect 136966 131728 136968 131737
rect 172020 131760 172072 131766
rect 137020 131728 137022 131737
rect 136876 131692 136928 131698
rect 172020 131702 172072 131708
rect 136966 131663 137022 131672
rect 136876 131634 136928 131640
rect 135312 131080 135364 131086
rect 135312 131022 135364 131028
rect 136784 131080 136836 131086
rect 136784 131022 136836 131028
rect 135324 130785 135352 131022
rect 135310 130776 135366 130785
rect 135310 130711 135366 130720
rect 172662 130776 172718 130785
rect 172662 130711 172718 130720
rect 136874 130640 136930 130649
rect 172676 130610 172704 130711
rect 136874 130575 136930 130584
rect 172664 130604 172716 130610
rect 136888 130338 136916 130575
rect 172664 130546 172716 130552
rect 174228 130604 174280 130610
rect 174228 130546 174280 130552
rect 136966 130504 137022 130513
rect 136966 130439 137022 130448
rect 136980 130406 137008 130439
rect 136968 130400 137020 130406
rect 136968 130342 137020 130348
rect 172662 130368 172718 130377
rect 135404 130332 135456 130338
rect 135404 130274 135456 130280
rect 136876 130332 136928 130338
rect 172662 130303 172664 130312
rect 136876 130274 136928 130280
rect 172716 130303 172718 130312
rect 172664 130274 172716 130280
rect 135218 130232 135274 130241
rect 135218 130167 135274 130176
rect 135128 129040 135180 129046
rect 135128 128982 135180 128988
rect 135034 128464 135090 128473
rect 135034 128399 135090 128408
rect 135140 127521 135168 128982
rect 135312 128972 135364 128978
rect 135312 128914 135364 128920
rect 135220 127612 135272 127618
rect 135220 127554 135272 127560
rect 135126 127512 135182 127521
rect 135126 127447 135182 127456
rect 134668 127204 134720 127210
rect 134668 127146 134720 127152
rect 134680 126705 134708 127146
rect 134666 126696 134722 126705
rect 134666 126631 134722 126640
rect 135036 126252 135088 126258
rect 135036 126194 135088 126200
rect 135048 124393 135076 126194
rect 135232 126025 135260 127554
rect 135324 127249 135352 128914
rect 135416 128745 135444 130274
rect 171834 129552 171890 129561
rect 171834 129487 171890 129496
rect 136966 129416 137022 129425
rect 171848 129386 171876 129487
rect 136966 129351 137022 129360
rect 171836 129380 171888 129386
rect 136980 129046 137008 129351
rect 171836 129322 171888 129328
rect 174136 129380 174188 129386
rect 174136 129322 174188 129328
rect 171834 129144 171890 129153
rect 171834 129079 171836 129088
rect 171888 129079 171890 129088
rect 171836 129050 171888 129056
rect 136968 129040 137020 129046
rect 136874 129008 136930 129017
rect 136968 128982 137020 128988
rect 136874 128943 136876 128952
rect 136928 128943 136930 128952
rect 136876 128914 136928 128920
rect 135402 128736 135458 128745
rect 135402 128671 135458 128680
rect 136782 128328 136838 128337
rect 136782 128263 136838 128272
rect 172570 128328 172626 128337
rect 172570 128263 172626 128272
rect 135310 127240 135366 127249
rect 136796 127210 136824 128263
rect 171558 127920 171614 127929
rect 172584 127890 172612 128263
rect 171558 127855 171614 127864
rect 172572 127884 172624 127890
rect 136874 127648 136930 127657
rect 171572 127618 171600 127855
rect 172572 127826 172624 127832
rect 136874 127583 136876 127592
rect 136928 127583 136930 127592
rect 171560 127612 171612 127618
rect 136876 127554 136928 127560
rect 171560 127554 171612 127560
rect 174148 127521 174176 129322
rect 174240 128745 174268 130546
rect 174320 130332 174372 130338
rect 174320 130274 174372 130280
rect 174226 128736 174282 128745
rect 174226 128671 174282 128680
rect 174332 128473 174360 130274
rect 174318 128464 174374 128473
rect 174318 128399 174374 128408
rect 174228 127884 174280 127890
rect 174228 127826 174280 127832
rect 174134 127512 174190 127521
rect 174134 127447 174190 127456
rect 135310 127175 135366 127184
rect 136784 127204 136836 127210
rect 136784 127146 136836 127152
rect 136782 127104 136838 127113
rect 136782 127039 136838 127048
rect 172018 127104 172074 127113
rect 172018 127039 172074 127048
rect 135312 126184 135364 126190
rect 135312 126126 135364 126132
rect 135218 126016 135274 126025
rect 135218 125951 135274 125960
rect 135128 124824 135180 124830
rect 135128 124766 135180 124772
rect 135034 124384 135090 124393
rect 135034 124319 135090 124328
rect 135140 123169 135168 124766
rect 135324 124665 135352 126126
rect 136796 125714 136824 127039
rect 136874 126424 136930 126433
rect 136874 126359 136930 126368
rect 136888 126190 136916 126359
rect 136966 126288 137022 126297
rect 136966 126223 136968 126232
rect 137020 126223 137022 126232
rect 136968 126194 137020 126200
rect 172032 126190 172060 127039
rect 174240 126705 174268 127826
rect 172202 126696 172258 126705
rect 172202 126631 172258 126640
rect 174226 126696 174282 126705
rect 174226 126631 174282 126640
rect 172216 126530 172244 126631
rect 172204 126524 172256 126530
rect 172204 126466 172256 126472
rect 174320 126524 174372 126530
rect 174320 126466 174372 126472
rect 172664 126252 172716 126258
rect 172664 126194 172716 126200
rect 136876 126184 136928 126190
rect 136876 126126 136928 126132
rect 172020 126184 172072 126190
rect 172676 126161 172704 126194
rect 174136 126184 174188 126190
rect 172020 126126 172072 126132
rect 172662 126152 172718 126161
rect 174136 126126 174188 126132
rect 172662 126087 172718 126096
rect 135404 125708 135456 125714
rect 135404 125650 135456 125656
rect 136784 125708 136836 125714
rect 136784 125650 136836 125656
rect 135416 125481 135444 125650
rect 174148 125481 174176 126126
rect 135402 125472 135458 125481
rect 135402 125407 135458 125416
rect 174134 125472 174190 125481
rect 174134 125407 174190 125416
rect 136782 125336 136838 125345
rect 136782 125271 136838 125280
rect 171834 125336 171890 125345
rect 171834 125271 171836 125280
rect 135310 124656 135366 124665
rect 135310 124591 135366 124600
rect 136796 124286 136824 125271
rect 171888 125271 171890 125280
rect 174228 125300 174280 125306
rect 171836 125242 171888 125248
rect 174228 125242 174280 125248
rect 172202 125064 172258 125073
rect 172202 124999 172258 125008
rect 136874 124928 136930 124937
rect 172216 124898 172244 124999
rect 136874 124863 136930 124872
rect 172204 124892 172256 124898
rect 136888 124830 136916 124863
rect 172204 124834 172256 124840
rect 136876 124824 136928 124830
rect 136876 124766 136928 124772
rect 135220 124280 135272 124286
rect 135220 124222 135272 124228
rect 136784 124280 136836 124286
rect 136784 124222 136836 124228
rect 135232 123713 135260 124222
rect 136782 124112 136838 124121
rect 136782 124047 136838 124056
rect 171834 124112 171890 124121
rect 171834 124047 171890 124056
rect 135218 123704 135274 123713
rect 135218 123639 135274 123648
rect 135404 123396 135456 123402
rect 135404 123338 135456 123344
rect 135126 123160 135182 123169
rect 135126 123095 135182 123104
rect 135312 122920 135364 122926
rect 135312 122862 135364 122868
rect 135324 122625 135352 122862
rect 135310 122616 135366 122625
rect 135310 122551 135366 122560
rect 135128 122172 135180 122178
rect 135128 122114 135180 122120
rect 135140 120313 135168 122114
rect 135220 122104 135272 122110
rect 135220 122046 135272 122052
rect 135232 120585 135260 122046
rect 135312 121968 135364 121974
rect 135416 121945 135444 123338
rect 136796 122926 136824 124047
rect 136874 123432 136930 123441
rect 171848 123402 171876 124047
rect 174240 123713 174268 125242
rect 174332 124665 174360 126466
rect 174318 124656 174374 124665
rect 174318 124591 174374 124600
rect 172570 123704 172626 123713
rect 172570 123639 172626 123648
rect 174226 123704 174282 123713
rect 174226 123639 174282 123648
rect 172584 123538 172612 123639
rect 172572 123532 172624 123538
rect 172572 123474 172624 123480
rect 136874 123367 136876 123376
rect 136928 123367 136930 123376
rect 171836 123396 171888 123402
rect 136876 123338 136928 123344
rect 171836 123338 171888 123344
rect 174136 123396 174188 123402
rect 174136 123338 174188 123344
rect 136784 122920 136836 122926
rect 136784 122862 136836 122868
rect 136874 122888 136930 122897
rect 136874 122823 136930 122832
rect 171834 122888 171890 122897
rect 171834 122823 171890 122832
rect 136888 122042 136916 122823
rect 136966 122480 137022 122489
rect 171848 122450 171876 122823
rect 174148 122625 174176 123338
rect 174134 122616 174190 122625
rect 174134 122551 174190 122560
rect 172018 122480 172074 122489
rect 136966 122415 137022 122424
rect 171836 122444 171888 122450
rect 136980 122110 137008 122415
rect 172018 122415 172074 122424
rect 171836 122386 171888 122392
rect 137058 122208 137114 122217
rect 172032 122178 172060 122415
rect 137058 122143 137060 122152
rect 137112 122143 137114 122152
rect 172020 122172 172072 122178
rect 137060 122114 137112 122120
rect 172020 122114 172072 122120
rect 136968 122104 137020 122110
rect 136968 122046 137020 122052
rect 172662 122072 172718 122081
rect 136876 122036 136928 122042
rect 172662 122007 172664 122016
rect 136876 121978 136928 121984
rect 172716 122007 172718 122016
rect 172664 121978 172716 121984
rect 135312 121910 135364 121916
rect 135402 121936 135458 121945
rect 135324 121401 135352 121910
rect 135402 121871 135458 121880
rect 135310 121392 135366 121401
rect 135310 121327 135366 121336
rect 136782 121120 136838 121129
rect 136782 121055 136838 121064
rect 172110 121120 172166 121129
rect 172110 121055 172166 121064
rect 135218 120576 135274 120585
rect 135218 120511 135274 120520
rect 135126 120304 135182 120313
rect 134852 120268 134904 120274
rect 136796 120274 136824 121055
rect 172124 120954 172152 121055
rect 172112 120948 172164 120954
rect 172112 120890 172164 120896
rect 174320 120948 174372 120954
rect 174320 120890 174372 120896
rect 172662 120848 172718 120857
rect 172662 120783 172664 120792
rect 172716 120783 172718 120792
rect 174228 120812 174280 120818
rect 172664 120754 172716 120760
rect 174228 120754 174280 120760
rect 136966 120712 137022 120721
rect 136966 120647 137022 120656
rect 135126 120239 135182 120248
rect 136784 120268 136836 120274
rect 134852 120210 134904 120216
rect 136784 120210 136836 120216
rect 134864 119633 134892 120210
rect 136782 119896 136838 119905
rect 136782 119831 136838 119840
rect 134850 119624 134906 119633
rect 134850 119559 134906 119568
rect 135220 119316 135272 119322
rect 135220 119258 135272 119264
rect 135128 117956 135180 117962
rect 135128 117898 135180 117904
rect 132920 117888 132972 117894
rect 132920 117830 132972 117836
rect 102468 117820 102520 117826
rect 102468 117762 102520 117768
rect 132644 117820 132696 117826
rect 132644 117762 132696 117768
rect 134116 117820 134168 117826
rect 134116 117762 134168 117768
rect 102376 117752 102428 117758
rect 102376 117694 102428 117700
rect 102388 117593 102416 117694
rect 102374 117584 102430 117593
rect 102374 117519 102430 117528
rect 102282 117040 102338 117049
rect 102282 116975 102338 116984
rect 102192 116732 102244 116738
rect 102192 116674 102244 116680
rect 102204 114737 102232 116674
rect 102480 116505 102508 117762
rect 132644 117684 132696 117690
rect 132644 117626 132696 117632
rect 102466 116496 102522 116505
rect 102376 116460 102428 116466
rect 102466 116431 102522 116440
rect 102376 116402 102428 116408
rect 102284 115508 102336 115514
rect 102284 115450 102336 115456
rect 102190 114728 102246 114737
rect 102190 114663 102246 114672
rect 102296 114193 102324 115450
rect 102388 115281 102416 116402
rect 102652 116392 102704 116398
rect 102652 116334 102704 116340
rect 102664 115825 102692 116334
rect 102650 115816 102706 115825
rect 102650 115751 102706 115760
rect 102374 115272 102430 115281
rect 102374 115207 102430 115216
rect 102282 114184 102338 114193
rect 102282 114119 102338 114128
rect 101822 113776 101878 113785
rect 101822 113711 101878 113720
rect 105102 113626 105130 113884
rect 105562 113626 105590 113884
rect 106114 113626 106142 113884
rect 106666 113626 106694 113884
rect 107218 113626 107246 113884
rect 107770 113626 107798 113884
rect 108322 113626 108350 113884
rect 108874 113626 108902 113884
rect 105102 113598 105176 113626
rect 105562 113598 105636 113626
rect 103664 112992 103716 112998
rect 103664 112934 103716 112940
rect 81676 112788 81728 112794
rect 81676 112730 81728 112736
rect 82504 112788 82556 112794
rect 82504 112730 82556 112736
rect 81688 112182 81716 112730
rect 103676 112318 103704 112934
rect 103664 112312 103716 112318
rect 103664 112254 103716 112260
rect 81676 112176 81728 112182
rect 81676 112118 81728 112124
rect 60424 111632 60476 111638
rect 60424 111574 60476 111580
rect 59870 104256 59926 104265
rect 59870 104191 59926 104200
rect 59884 104090 59912 104191
rect 59872 104084 59924 104090
rect 59872 104026 59924 104032
rect 105148 102225 105176 113598
rect 105412 111156 105464 111162
rect 105412 111098 105464 111104
rect 105228 111020 105280 111026
rect 105228 110962 105280 110968
rect 105240 105761 105268 110962
rect 105320 109184 105372 109190
rect 105318 109152 105320 109161
rect 105372 109152 105374 109161
rect 105318 109087 105374 109096
rect 105424 106849 105452 111098
rect 105410 106840 105466 106849
rect 105410 106775 105466 106784
rect 105226 105752 105282 105761
rect 105226 105687 105282 105696
rect 105608 103449 105636 113598
rect 106068 113598 106142 113626
rect 106620 113598 106694 113626
rect 107172 113598 107246 113626
rect 107724 113598 107798 113626
rect 108276 113598 108350 113626
rect 108828 113598 108902 113626
rect 109426 113626 109454 113884
rect 109978 113626 110006 113884
rect 110530 113626 110558 113884
rect 109426 113598 109500 113626
rect 109978 113598 110052 113626
rect 105688 111088 105740 111094
rect 105688 111030 105740 111036
rect 105700 107937 105728 111030
rect 105780 110952 105832 110958
rect 105780 110894 105832 110900
rect 105792 110249 105820 110894
rect 105778 110240 105834 110249
rect 105778 110175 105834 110184
rect 105686 107928 105742 107937
rect 105686 107863 105742 107872
rect 106068 104537 106096 113598
rect 106620 111026 106648 113598
rect 107172 111162 107200 113598
rect 107160 111156 107212 111162
rect 107160 111098 107212 111104
rect 107724 111094 107752 113598
rect 107712 111088 107764 111094
rect 107712 111030 107764 111036
rect 106608 111020 106660 111026
rect 106608 110962 106660 110968
rect 108276 109190 108304 113598
rect 108828 111026 108856 113598
rect 109472 112318 109500 113598
rect 109460 112312 109512 112318
rect 109460 112254 109512 112260
rect 110024 112250 110052 113598
rect 110484 113598 110558 113626
rect 111082 113626 111110 113884
rect 111634 113626 111662 113884
rect 112186 113626 112214 113884
rect 112738 113626 112766 113884
rect 113290 113626 113318 113884
rect 111082 113598 111156 113626
rect 110012 112244 110064 112250
rect 110012 112186 110064 112192
rect 110484 112182 110512 113598
rect 110472 112176 110524 112182
rect 110472 112118 110524 112124
rect 108816 111020 108868 111026
rect 108816 110962 108868 110968
rect 111128 110756 111156 113598
rect 111588 113598 111662 113626
rect 112140 113598 112214 113626
rect 112600 113598 112766 113626
rect 112968 113598 113318 113626
rect 113508 113672 113560 113678
rect 113842 113626 113870 113884
rect 114394 113678 114422 113884
rect 113508 113614 113560 113620
rect 111588 110770 111616 113598
rect 112140 110770 112168 113598
rect 112600 110770 112628 113598
rect 112968 110770 112996 113598
rect 113048 111836 113100 111842
rect 113048 111778 113100 111784
rect 111510 110742 111616 110770
rect 111878 110742 112168 110770
rect 112338 110742 112628 110770
rect 112706 110742 112996 110770
rect 113060 110756 113088 111778
rect 113520 110756 113548 113614
rect 113796 113598 113870 113626
rect 114382 113672 114434 113678
rect 114946 113626 114974 113884
rect 115498 113626 115526 113884
rect 116050 113626 116078 113884
rect 116602 113626 116630 113884
rect 117154 113626 117182 113884
rect 117706 113626 117734 113884
rect 118258 113626 118286 113884
rect 118810 113626 118838 113884
rect 119270 113626 119298 113884
rect 119822 113626 119850 113884
rect 120374 113626 120402 113884
rect 120926 113626 120954 113884
rect 121478 113626 121506 113884
rect 122030 113626 122058 113884
rect 122582 113626 122610 113884
rect 123134 113626 123162 113884
rect 123686 113626 123714 113884
rect 124238 113626 124266 113884
rect 124790 113626 124818 113884
rect 125342 113626 125370 113884
rect 125894 113626 125922 113884
rect 126446 113626 126474 113884
rect 126998 113626 127026 113884
rect 127550 113626 127578 113884
rect 128102 113626 128130 113884
rect 128654 113626 128682 113884
rect 129206 113626 129234 113884
rect 129758 113626 129786 113884
rect 130310 113626 130338 113884
rect 130862 113626 130890 113884
rect 131414 113626 131442 113884
rect 131966 113626 131994 113884
rect 114382 113614 114434 113620
rect 114900 113598 114974 113626
rect 115452 113598 115526 113626
rect 116004 113598 116078 113626
rect 116556 113598 116630 113626
rect 117108 113598 117182 113626
rect 117660 113598 117734 113626
rect 118212 113598 118286 113626
rect 118764 113598 118838 113626
rect 119224 113598 119298 113626
rect 119776 113598 119850 113626
rect 120328 113598 120402 113626
rect 120880 113598 120954 113626
rect 121432 113598 121506 113626
rect 121984 113598 122058 113626
rect 122536 113598 122610 113626
rect 123088 113598 123162 113626
rect 123640 113598 123714 113626
rect 124192 113598 124266 113626
rect 124744 113598 124818 113626
rect 125296 113598 125370 113626
rect 125848 113598 125922 113626
rect 126400 113598 126474 113626
rect 126952 113598 127026 113626
rect 127504 113598 127578 113626
rect 128056 113598 128130 113626
rect 128608 113598 128682 113626
rect 129160 113598 129234 113626
rect 129712 113598 129786 113626
rect 130264 113598 130338 113626
rect 130816 113598 130890 113626
rect 131368 113598 131442 113626
rect 131920 113598 131994 113626
rect 132092 113672 132144 113678
rect 132518 113626 132546 113884
rect 132092 113614 132144 113620
rect 113796 111842 113824 113598
rect 113784 111836 113836 111842
rect 113784 111778 113836 111784
rect 114244 111428 114296 111434
rect 114244 111370 114296 111376
rect 113876 111360 113928 111366
rect 113876 111302 113928 111308
rect 113888 110756 113916 111302
rect 114256 110756 114284 111370
rect 114900 111366 114928 113598
rect 115452 111434 115480 113598
rect 115440 111428 115492 111434
rect 115440 111370 115492 111376
rect 114888 111360 114940 111366
rect 114888 111302 114940 111308
rect 116004 111298 116032 113598
rect 116268 111360 116320 111366
rect 116268 111302 116320 111308
rect 114704 111292 114756 111298
rect 114704 111234 114756 111240
rect 115992 111292 116044 111298
rect 115992 111234 116044 111240
rect 114716 110756 114744 111234
rect 115440 111224 115492 111230
rect 115440 111166 115492 111172
rect 115072 111020 115124 111026
rect 115072 110962 115124 110968
rect 115084 110756 115112 110962
rect 115452 110756 115480 111166
rect 115900 111088 115952 111094
rect 115900 111030 115952 111036
rect 115912 110756 115940 111030
rect 116280 110756 116308 111302
rect 116556 111026 116584 113598
rect 116636 111428 116688 111434
rect 116636 111370 116688 111376
rect 116544 111020 116596 111026
rect 116544 110962 116596 110968
rect 116648 110756 116676 111370
rect 117108 111230 117136 113598
rect 117464 111292 117516 111298
rect 117464 111234 117516 111240
rect 117096 111224 117148 111230
rect 117096 111166 117148 111172
rect 117096 111020 117148 111026
rect 117096 110962 117148 110968
rect 117108 110756 117136 110962
rect 117476 110756 117504 111234
rect 117660 111094 117688 113598
rect 117832 111904 117884 111910
rect 117832 111846 117884 111852
rect 117648 111088 117700 111094
rect 117648 111030 117700 111036
rect 117844 110756 117872 111846
rect 118212 111366 118240 113598
rect 118660 111496 118712 111502
rect 118660 111438 118712 111444
rect 118200 111360 118252 111366
rect 118200 111302 118252 111308
rect 118292 111360 118344 111366
rect 118292 111302 118344 111308
rect 118304 110756 118332 111302
rect 118672 110756 118700 111438
rect 118764 111434 118792 113598
rect 118752 111428 118804 111434
rect 118752 111370 118804 111376
rect 119120 111156 119172 111162
rect 119120 111098 119172 111104
rect 119132 110756 119160 111098
rect 119224 111026 119252 113598
rect 119776 111298 119804 113598
rect 120328 111910 120356 113598
rect 120316 111904 120368 111910
rect 120316 111846 120368 111852
rect 119856 111836 119908 111842
rect 119856 111778 119908 111784
rect 119764 111292 119816 111298
rect 119764 111234 119816 111240
rect 119488 111224 119540 111230
rect 119488 111166 119540 111172
rect 119212 111020 119264 111026
rect 119212 110962 119264 110968
rect 119500 110756 119528 111166
rect 119868 110756 119896 111778
rect 120316 111768 120368 111774
rect 120316 111710 120368 111716
rect 120328 110756 120356 111710
rect 120880 111366 120908 113598
rect 121052 112176 121104 112182
rect 121052 112118 121104 112124
rect 120868 111360 120920 111366
rect 120868 111302 120920 111308
rect 120684 111292 120736 111298
rect 120684 111234 120736 111240
rect 120696 110756 120724 111234
rect 121064 110756 121092 112118
rect 121432 111502 121460 113598
rect 121420 111496 121472 111502
rect 121420 111438 121472 111444
rect 121512 111428 121564 111434
rect 121512 111370 121564 111376
rect 121524 110756 121552 111370
rect 121880 111360 121932 111366
rect 121880 111302 121932 111308
rect 121892 110756 121920 111302
rect 121984 111162 122012 113598
rect 122248 111972 122300 111978
rect 122248 111914 122300 111920
rect 121972 111156 122024 111162
rect 121972 111098 122024 111104
rect 122260 110756 122288 111914
rect 122536 111230 122564 113598
rect 123088 111910 123116 113598
rect 123076 111904 123128 111910
rect 123076 111846 123128 111852
rect 122708 111836 122760 111842
rect 122708 111778 122760 111784
rect 122524 111224 122576 111230
rect 122524 111166 122576 111172
rect 122720 110756 122748 111778
rect 123640 111774 123668 113598
rect 123628 111768 123680 111774
rect 123628 111710 123680 111716
rect 123076 111632 123128 111638
rect 123076 111574 123128 111580
rect 123088 110756 123116 111574
rect 123444 111564 123496 111570
rect 123444 111506 123496 111512
rect 123456 110756 123484 111506
rect 124192 111298 124220 113598
rect 124744 112182 124772 113598
rect 124732 112176 124784 112182
rect 124732 112118 124784 112124
rect 124272 111496 124324 111502
rect 124272 111438 124324 111444
rect 124180 111292 124232 111298
rect 124180 111234 124232 111240
rect 123904 111156 123956 111162
rect 123904 111098 123956 111104
rect 123916 110756 123944 111098
rect 124284 110756 124312 111438
rect 125296 111434 125324 113598
rect 125848 111434 125876 113598
rect 126400 111978 126428 113598
rect 126388 111972 126440 111978
rect 126388 111914 126440 111920
rect 126952 111842 126980 113598
rect 126940 111836 126992 111842
rect 126940 111778 126992 111784
rect 127504 111638 127532 113598
rect 127492 111632 127544 111638
rect 127492 111574 127544 111580
rect 128056 111570 128084 113598
rect 128044 111564 128096 111570
rect 128044 111506 128096 111512
rect 125284 111428 125336 111434
rect 125284 111370 125336 111376
rect 125836 111428 125888 111434
rect 125836 111370 125888 111376
rect 126296 111428 126348 111434
rect 126296 111370 126348 111376
rect 125468 111360 125520 111366
rect 125468 111302 125520 111308
rect 125100 111292 125152 111298
rect 125100 111234 125152 111240
rect 124640 111224 124692 111230
rect 124640 111166 124692 111172
rect 124652 110756 124680 111166
rect 125112 110756 125140 111234
rect 125480 110756 125508 111302
rect 125836 111020 125888 111026
rect 125836 110962 125888 110968
rect 125848 110756 125876 110962
rect 126308 110756 126336 111370
rect 128608 111162 128636 113598
rect 129160 111502 129188 113598
rect 129148 111496 129200 111502
rect 129148 111438 129200 111444
rect 129712 111230 129740 113598
rect 130264 111298 130292 113598
rect 130816 111366 130844 113598
rect 130804 111360 130856 111366
rect 130804 111302 130856 111308
rect 130252 111292 130304 111298
rect 130252 111234 130304 111240
rect 129700 111224 129752 111230
rect 129700 111166 129752 111172
rect 128596 111156 128648 111162
rect 128596 111098 128648 111104
rect 126664 111088 126716 111094
rect 126664 111030 126716 111036
rect 126676 110756 126704 111030
rect 131368 111026 131396 113598
rect 131920 111434 131948 113598
rect 132104 112318 132132 113614
rect 132196 113598 132546 113626
rect 132092 112312 132144 112318
rect 132092 112254 132144 112260
rect 131908 111428 131960 111434
rect 131908 111370 131960 111376
rect 132196 111094 132224 113598
rect 132656 113082 132684 117626
rect 134128 117321 134156 117762
rect 134114 117312 134170 117321
rect 134114 117247 134170 117256
rect 134668 117208 134720 117214
rect 134668 117150 134720 117156
rect 134680 116777 134708 117150
rect 134666 116768 134722 116777
rect 134666 116703 134722 116712
rect 135140 116233 135168 117898
rect 135232 117593 135260 119258
rect 135312 119180 135364 119186
rect 135312 119122 135364 119128
rect 135324 119089 135352 119122
rect 135310 119080 135366 119089
rect 135310 119015 135366 119024
rect 136796 118574 136824 119831
rect 136874 119352 136930 119361
rect 136874 119287 136876 119296
rect 136928 119287 136930 119296
rect 136876 119258 136928 119264
rect 136980 119186 137008 120647
rect 171834 119896 171890 119905
rect 171834 119831 171890 119840
rect 171848 119730 171876 119831
rect 171836 119724 171888 119730
rect 171836 119666 171888 119672
rect 174136 119724 174188 119730
rect 174136 119666 174188 119672
rect 171834 119624 171890 119633
rect 171834 119559 171890 119568
rect 171848 119458 171876 119559
rect 171836 119452 171888 119458
rect 171836 119394 171888 119400
rect 136968 119180 137020 119186
rect 136968 119122 137020 119128
rect 136966 118672 137022 118681
rect 136966 118607 137022 118616
rect 171834 118672 171890 118681
rect 171834 118607 171890 118616
rect 135312 118568 135364 118574
rect 135310 118536 135312 118545
rect 136784 118568 136836 118574
rect 135364 118536 135366 118545
rect 136784 118510 136836 118516
rect 135310 118471 135366 118480
rect 136782 118128 136838 118137
rect 136782 118063 136838 118072
rect 135218 117584 135274 117593
rect 135218 117519 135274 117528
rect 136796 117214 136824 118063
rect 136874 117992 136930 118001
rect 136874 117927 136876 117936
rect 136928 117927 136930 117936
rect 136876 117898 136928 117904
rect 136980 117894 137008 118607
rect 171650 118264 171706 118273
rect 171650 118199 171652 118208
rect 171704 118199 171706 118208
rect 171652 118170 171704 118176
rect 171848 117894 171876 118607
rect 174148 118545 174176 119666
rect 174240 119089 174268 120754
rect 174332 119633 174360 120890
rect 174318 119624 174374 119633
rect 174318 119559 174374 119568
rect 174226 119080 174282 119089
rect 174226 119015 174282 119024
rect 174134 118536 174190 118545
rect 174134 118471 174190 118480
rect 173952 118228 174004 118234
rect 173952 118170 174004 118176
rect 172662 118128 172718 118137
rect 172662 118063 172664 118072
rect 172716 118063 172718 118072
rect 172664 118034 172716 118040
rect 136968 117888 137020 117894
rect 136968 117830 137020 117836
rect 171836 117888 171888 117894
rect 171836 117830 171888 117836
rect 136784 117208 136836 117214
rect 136784 117150 136836 117156
rect 136782 116904 136838 116913
rect 136782 116839 136838 116848
rect 172662 116904 172718 116913
rect 172662 116839 172718 116848
rect 135312 116528 135364 116534
rect 135312 116470 135364 116476
rect 135126 116224 135182 116233
rect 135126 116159 135182 116168
rect 134852 115644 134904 115650
rect 134852 115586 134904 115592
rect 134864 115553 134892 115586
rect 134850 115544 134906 115553
rect 134850 115479 134906 115488
rect 135324 115009 135352 116470
rect 136796 115650 136824 116839
rect 136874 116768 136930 116777
rect 136874 116703 136930 116712
rect 136888 116534 136916 116703
rect 172570 116632 172626 116641
rect 172676 116602 172704 116839
rect 173964 116777 173992 118170
rect 174320 118092 174372 118098
rect 174320 118034 174372 118040
rect 174044 117888 174096 117894
rect 174044 117830 174096 117836
rect 174056 117321 174084 117830
rect 174042 117312 174098 117321
rect 174042 117247 174098 117256
rect 173950 116768 174006 116777
rect 173950 116703 174006 116712
rect 172570 116567 172626 116576
rect 172664 116596 172716 116602
rect 172584 116534 172612 116567
rect 172664 116538 172716 116544
rect 174136 116596 174188 116602
rect 174136 116538 174188 116544
rect 136876 116528 136928 116534
rect 136876 116470 136928 116476
rect 172572 116528 172624 116534
rect 172572 116470 172624 116476
rect 136784 115644 136836 115650
rect 136784 115586 136836 115592
rect 136782 115544 136838 115553
rect 136782 115479 136838 115488
rect 135310 115000 135366 115009
rect 135310 114935 135366 114944
rect 136796 114494 136824 115479
rect 134852 114488 134904 114494
rect 134850 114456 134852 114465
rect 136784 114488 136836 114494
rect 134904 114456 134906 114465
rect 136784 114430 136836 114436
rect 134850 114391 134906 114400
rect 144892 113678 144920 115924
rect 144880 113672 144932 113678
rect 144880 113614 144932 113620
rect 154828 113610 154856 115924
rect 154816 113604 154868 113610
rect 154816 113546 154868 113552
rect 132564 113054 132684 113082
rect 132184 111088 132236 111094
rect 132184 111030 132236 111036
rect 131356 111020 131408 111026
rect 131356 110962 131408 110968
rect 108538 109560 108594 109569
rect 108538 109495 108594 109504
rect 108264 109184 108316 109190
rect 108264 109126 108316 109132
rect 107894 107248 107950 107257
rect 106424 107212 106476 107218
rect 107894 107183 107896 107192
rect 106424 107154 106476 107160
rect 107948 107183 107950 107192
rect 107896 107154 107948 107160
rect 106054 104528 106110 104537
rect 106054 104463 106110 104472
rect 105780 104084 105832 104090
rect 105780 104026 105832 104032
rect 105594 103440 105650 103449
rect 105594 103375 105650 103384
rect 105134 102216 105190 102225
rect 105134 102151 105190 102160
rect 105792 98825 105820 104026
rect 106332 101364 106384 101370
rect 106332 101306 106384 101312
rect 105964 101296 106016 101302
rect 105964 101238 106016 101244
rect 105976 101137 106004 101238
rect 105962 101128 106018 101137
rect 105962 101063 106018 101072
rect 105778 98816 105834 98825
rect 105778 98751 105834 98760
rect 106344 97737 106372 101306
rect 106436 100049 106464 107154
rect 108446 104936 108502 104945
rect 108446 104871 108502 104880
rect 108460 104090 108488 104871
rect 108448 104084 108500 104090
rect 108448 104026 108500 104032
rect 107894 102488 107950 102497
rect 107894 102423 107950 102432
rect 107908 101370 107936 102423
rect 107896 101364 107948 101370
rect 107896 101306 107948 101312
rect 108552 101302 108580 109495
rect 132564 105489 132592 113054
rect 164856 112998 164884 115924
rect 171834 115680 171890 115689
rect 171834 115615 171836 115624
rect 171888 115615 171890 115624
rect 174044 115644 174096 115650
rect 171836 115586 171888 115592
rect 174044 115586 174096 115592
rect 174056 114465 174084 115586
rect 174148 115553 174176 116538
rect 174228 116528 174280 116534
rect 174228 116470 174280 116476
rect 174134 115544 174190 115553
rect 174134 115479 174190 115488
rect 174240 115009 174268 116470
rect 174332 116233 174360 118034
rect 174318 116224 174374 116233
rect 174318 116159 174374 116168
rect 174226 115000 174282 115009
rect 174226 114935 174282 114944
rect 174042 114456 174098 114465
rect 174042 114391 174098 114400
rect 132644 112992 132696 112998
rect 132644 112934 132696 112940
rect 164844 112992 164896 112998
rect 164844 112934 164896 112940
rect 132656 112250 132684 112934
rect 132644 112244 132696 112250
rect 132644 112186 132696 112192
rect 132274 105480 132330 105489
rect 132274 105415 132330 105424
rect 132550 105480 132606 105489
rect 132550 105415 132606 105424
rect 108540 101296 108592 101302
rect 108540 101238 108592 101244
rect 107894 100176 107950 100185
rect 107894 100111 107950 100120
rect 106422 100040 106478 100049
rect 106422 99975 106478 99984
rect 107908 99942 107936 100111
rect 106424 99936 106476 99942
rect 106424 99878 106476 99884
rect 107896 99936 107948 99942
rect 107896 99878 107948 99884
rect 106330 97728 106386 97737
rect 106240 97692 106292 97698
rect 106330 97663 106386 97672
rect 106240 97634 106292 97640
rect 106252 95425 106280 97634
rect 106436 96513 106464 99878
rect 132288 98530 132316 105415
rect 132288 98502 132408 98530
rect 107894 97864 107950 97873
rect 107894 97799 107950 97808
rect 107908 97698 107936 97799
rect 107896 97692 107948 97698
rect 107896 97634 107948 97640
rect 106422 96504 106478 96513
rect 106422 96439 106478 96448
rect 132380 95794 132408 98502
rect 132368 95788 132420 95794
rect 132368 95730 132420 95736
rect 106238 95416 106294 95425
rect 106238 95351 106294 95360
rect 108446 95416 108502 95425
rect 108446 95351 108502 95360
rect 108460 94842 108488 95351
rect 106516 94836 106568 94842
rect 106516 94778 106568 94784
rect 108448 94836 108500 94842
rect 108448 94778 108500 94784
rect 106528 94337 106556 94778
rect 106514 94328 106570 94337
rect 106514 94263 106570 94272
rect 105870 91744 105926 91753
rect 105870 91679 105872 91688
rect 105924 91679 105926 91688
rect 107804 91708 107856 91714
rect 105872 91650 105924 91656
rect 107804 91650 107856 91656
rect 59594 90928 59650 90937
rect 59594 90863 59650 90872
rect 59608 90286 59636 90863
rect 107816 90801 107844 91650
rect 107802 90792 107858 90801
rect 107802 90727 107858 90736
rect 105226 90384 105282 90393
rect 105226 90319 105282 90328
rect 105240 90286 105268 90319
rect 59596 90280 59648 90286
rect 59596 90222 59648 90228
rect 105228 90280 105280 90286
rect 105228 90222 105280 90228
rect 107896 90280 107948 90286
rect 107896 90222 107948 90228
rect 105134 89296 105190 89305
rect 105134 89231 105136 89240
rect 105188 89231 105190 89240
rect 107804 89260 107856 89266
rect 105136 89202 105188 89208
rect 107804 89202 107856 89208
rect 105870 87936 105926 87945
rect 105870 87871 105926 87880
rect 105884 87770 105912 87871
rect 105872 87764 105924 87770
rect 105872 87706 105924 87712
rect 107712 87764 107764 87770
rect 107712 87706 107764 87712
rect 106422 86712 106478 86721
rect 106478 86670 106556 86698
rect 106422 86647 106478 86656
rect 105594 86304 105650 86313
rect 105594 86239 105650 86248
rect 105608 86138 105636 86239
rect 105596 86132 105648 86138
rect 105596 86074 105648 86080
rect 106330 84808 106386 84817
rect 106330 84743 106332 84752
rect 106384 84743 106386 84752
rect 106332 84714 106384 84720
rect 105594 83448 105650 83457
rect 105594 83383 105596 83392
rect 105648 83383 105650 83392
rect 105596 83354 105648 83360
rect 105502 82224 105558 82233
rect 105502 82159 105558 82168
rect 105516 82058 105544 82159
rect 105504 82052 105556 82058
rect 105504 81994 105556 82000
rect 106528 81990 106556 86670
rect 107724 83729 107752 87706
rect 107816 86041 107844 89202
rect 107908 88489 107936 90222
rect 132552 88784 132604 88790
rect 132552 88726 132604 88732
rect 107894 88480 107950 88489
rect 107894 88415 107950 88424
rect 108724 86132 108776 86138
rect 108724 86074 108776 86080
rect 107802 86032 107858 86041
rect 107802 85967 107858 85976
rect 107710 83720 107766 83729
rect 107710 83655 107766 83664
rect 108632 83412 108684 83418
rect 108632 83354 108684 83360
rect 108540 82052 108592 82058
rect 108540 81994 108592 82000
rect 106516 81984 106568 81990
rect 56926 81952 56982 81961
rect 56926 81887 56982 81896
rect 57478 81952 57534 81961
rect 106516 81926 106568 81932
rect 107896 81984 107948 81990
rect 107896 81926 107948 81932
rect 57478 81887 57534 81896
rect 57492 80873 57520 81887
rect 107908 81417 107936 81926
rect 107894 81408 107950 81417
rect 107894 81343 107950 81352
rect 105226 81000 105282 81009
rect 105226 80935 105282 80944
rect 57478 80864 57534 80873
rect 57478 80799 57534 80808
rect 54812 79264 54864 79270
rect 54812 79206 54864 79212
rect 30524 77836 30576 77842
rect 30524 77778 30576 77784
rect 37424 77836 37476 77842
rect 37424 77778 37476 77784
rect 37436 77609 37464 77778
rect 57492 77638 57520 80799
rect 105240 80630 105268 80935
rect 105228 80624 105280 80630
rect 105228 80566 105280 80572
rect 108080 80624 108132 80630
rect 108080 80566 108132 80572
rect 105134 79912 105190 79921
rect 105134 79847 105190 79856
rect 105148 79746 105176 79847
rect 105136 79740 105188 79746
rect 105136 79682 105188 79688
rect 107528 79740 107580 79746
rect 107528 79682 107580 79688
rect 106974 79368 107030 79377
rect 106974 79303 107030 79312
rect 106330 77872 106386 77881
rect 106330 77807 106386 77816
rect 57480 77632 57532 77638
rect 31994 77600 32050 77609
rect 31994 77535 32050 77544
rect 37422 77600 37478 77609
rect 59596 77632 59648 77638
rect 57480 77574 57532 77580
rect 59594 77600 59596 77609
rect 59648 77600 59650 77609
rect 37422 77535 37478 77544
rect 28684 69540 28736 69546
rect 28684 69482 28736 69488
rect 31904 69472 31956 69478
rect 31904 69414 31956 69420
rect 31916 68866 31944 69414
rect 31904 68860 31956 68866
rect 31904 68802 31956 68808
rect 27580 68792 27632 68798
rect 31916 68769 31944 68802
rect 27580 68734 27632 68740
rect 31902 68760 31958 68769
rect 31902 68695 31958 68704
rect 32008 67658 32036 77535
rect 54812 76476 54864 76482
rect 54812 76418 54864 76424
rect 36044 69540 36096 69546
rect 36044 69482 36096 69488
rect 35584 69472 35636 69478
rect 35584 69414 35636 69420
rect 34112 69404 34164 69410
rect 34112 69346 34164 69352
rect 32008 67630 32956 67658
rect 32928 67522 32956 67630
rect 34124 67522 34152 69346
rect 34664 69336 34716 69342
rect 34664 69278 34716 69284
rect 34676 67522 34704 69278
rect 35596 67522 35624 69414
rect 36056 67522 36084 69482
rect 39092 69410 39120 70908
rect 39080 69404 39132 69410
rect 39080 69346 39132 69352
rect 39460 69342 39488 70908
rect 39828 69478 39856 70908
rect 40288 69546 40316 70908
rect 40276 69540 40328 69546
rect 40276 69482 40328 69488
rect 39816 69472 39868 69478
rect 39816 69414 39868 69420
rect 39448 69336 39500 69342
rect 39448 69278 39500 69284
rect 40000 69200 40052 69206
rect 40000 69142 40052 69148
rect 36596 69132 36648 69138
rect 36596 69074 36648 69080
rect 32928 67494 33218 67522
rect 33862 67494 34152 67522
rect 34506 67494 34704 67522
rect 35242 67494 35624 67522
rect 35886 67494 36084 67522
rect 36608 67508 36636 69074
rect 37240 69064 37292 69070
rect 37240 69006 37292 69012
rect 37252 67508 37280 69006
rect 39264 68860 39316 68866
rect 39264 68802 39316 68808
rect 37884 68588 37936 68594
rect 37884 68530 37936 68536
rect 37896 67508 37924 68530
rect 38620 68520 38672 68526
rect 38620 68462 38672 68468
rect 38632 67508 38660 68462
rect 39276 67508 39304 68802
rect 40012 67508 40040 69142
rect 40656 69138 40684 70908
rect 40644 69132 40696 69138
rect 40644 69074 40696 69080
rect 41024 69070 41052 70908
rect 41288 69132 41340 69138
rect 41288 69074 41340 69080
rect 41012 69064 41064 69070
rect 41012 69006 41064 69012
rect 40644 68996 40696 69002
rect 40644 68938 40696 68944
rect 40656 67508 40684 68938
rect 41300 67508 41328 69074
rect 41484 68594 41512 70908
rect 41472 68588 41524 68594
rect 41472 68530 41524 68536
rect 41852 68526 41880 70908
rect 42024 68928 42076 68934
rect 42024 68870 42076 68876
rect 41840 68520 41892 68526
rect 41840 68462 41892 68468
rect 42036 67508 42064 68870
rect 42220 68866 42248 70908
rect 42680 69206 42708 70908
rect 42668 69200 42720 69206
rect 42668 69142 42720 69148
rect 42668 69064 42720 69070
rect 42668 69006 42720 69012
rect 42208 68860 42260 68866
rect 42208 68802 42260 68808
rect 42680 67508 42708 69006
rect 43048 69002 43076 70908
rect 43416 69138 43444 70908
rect 43404 69132 43456 69138
rect 43404 69074 43456 69080
rect 43036 68996 43088 69002
rect 43036 68938 43088 68944
rect 43404 68996 43456 69002
rect 43404 68938 43456 68944
rect 43416 67508 43444 68938
rect 43876 68934 43904 70908
rect 44244 69070 44272 70908
rect 44232 69064 44284 69070
rect 44232 69006 44284 69012
rect 44612 69002 44640 70908
rect 44704 70894 45086 70922
rect 45164 70894 45454 70922
rect 45716 70894 45822 70922
rect 44600 68996 44652 69002
rect 44600 68938 44652 68944
rect 43864 68928 43916 68934
rect 43864 68870 43916 68876
rect 44704 68338 44732 70894
rect 44336 68310 44732 68338
rect 44336 67522 44364 68310
rect 45164 67522 45192 70894
rect 45716 67522 45744 70894
rect 46268 67522 46296 70908
rect 44074 67494 44364 67522
rect 44810 67494 45192 67522
rect 45454 67494 45744 67522
rect 46098 67494 46296 67522
rect 46636 67522 46664 70908
rect 47110 70894 47308 70922
rect 47478 70894 47768 70922
rect 47280 67522 47308 70894
rect 47740 67522 47768 70894
rect 47832 69002 47860 70908
rect 48292 69041 48320 70908
rect 48278 69032 48334 69041
rect 47820 68996 47872 69002
rect 48660 69002 48688 70908
rect 48278 68967 48334 68976
rect 48556 68996 48608 69002
rect 47820 68938 47872 68944
rect 48556 68938 48608 68944
rect 48648 68996 48700 69002
rect 48648 68938 48700 68944
rect 48568 67522 48596 68938
rect 49028 68905 49056 70908
rect 49488 69138 49516 70908
rect 49476 69132 49528 69138
rect 49476 69074 49528 69080
rect 49474 69032 49530 69041
rect 49474 68967 49530 68976
rect 49014 68896 49070 68905
rect 49014 68831 49070 68840
rect 46636 67494 46834 67522
rect 47280 67494 47478 67522
rect 47740 67494 48214 67522
rect 48568 67494 48858 67522
rect 49488 67508 49516 68967
rect 49856 68458 49884 70908
rect 49936 68996 49988 69002
rect 49936 68938 49988 68944
rect 49844 68452 49896 68458
rect 49844 68394 49896 68400
rect 49948 67522 49976 68938
rect 50224 68798 50252 70908
rect 50684 69002 50712 70908
rect 50672 68996 50724 69002
rect 50672 68938 50724 68944
rect 50854 68896 50910 68905
rect 51052 68866 51080 70908
rect 51420 69206 51448 70908
rect 51408 69200 51460 69206
rect 51408 69142 51460 69148
rect 51880 69138 51908 70908
rect 52248 69274 52276 70908
rect 52236 69268 52288 69274
rect 52236 69210 52288 69216
rect 51592 69132 51644 69138
rect 51592 69074 51644 69080
rect 51868 69132 51920 69138
rect 51868 69074 51920 69080
rect 50854 68831 50910 68840
rect 51040 68860 51092 68866
rect 50212 68792 50264 68798
rect 50212 68734 50264 68740
rect 49948 67494 50238 67522
rect 50868 67508 50896 68831
rect 51040 68802 51092 68808
rect 51604 67508 51632 69074
rect 52616 68934 52644 70908
rect 53076 69070 53104 70908
rect 53444 69342 53472 70908
rect 53812 69546 53840 70908
rect 53800 69540 53852 69546
rect 53800 69482 53852 69488
rect 54272 69478 54300 70908
rect 54260 69472 54312 69478
rect 54260 69414 54312 69420
rect 53432 69336 53484 69342
rect 53432 69278 53484 69284
rect 53064 69064 53116 69070
rect 53064 69006 53116 69012
rect 54640 69002 54668 70908
rect 54824 69750 54852 76418
rect 54812 69744 54864 69750
rect 54812 69686 54864 69692
rect 55364 69404 55416 69410
rect 55364 69346 55416 69352
rect 54996 69200 55048 69206
rect 54996 69142 55048 69148
rect 53616 68996 53668 69002
rect 53616 68938 53668 68944
rect 54628 68996 54680 69002
rect 54628 68938 54680 68944
rect 52604 68928 52656 68934
rect 52604 68870 52656 68876
rect 52972 68792 53024 68798
rect 52972 68734 53024 68740
rect 52236 68452 52288 68458
rect 52236 68394 52288 68400
rect 52248 67508 52276 68394
rect 52984 67508 53012 68734
rect 53628 67508 53656 68938
rect 54260 68860 54312 68866
rect 54260 68802 54312 68808
rect 54272 67508 54300 68802
rect 55008 67508 55036 69142
rect 55376 69002 55404 69346
rect 56376 69268 56428 69274
rect 56376 69210 56428 69216
rect 55640 69132 55692 69138
rect 55640 69074 55692 69080
rect 55364 68996 55416 69002
rect 55364 68938 55416 68944
rect 55652 67508 55680 69074
rect 56388 67508 56416 69210
rect 56744 68928 56796 68934
rect 56796 68876 56876 68882
rect 56744 68870 56876 68876
rect 56756 68854 56876 68870
rect 56848 67522 56876 68854
rect 57492 68594 57520 77574
rect 59594 77535 59650 77544
rect 105410 76512 105466 76521
rect 105410 76447 105466 76456
rect 105226 75288 105282 75297
rect 105226 75223 105282 75232
rect 103202 73588 103258 73597
rect 103202 73523 103258 73532
rect 102558 73384 102614 73393
rect 102558 73319 102614 73328
rect 102572 72033 102600 73319
rect 103216 72402 103244 73523
rect 103204 72396 103256 72402
rect 103204 72338 103256 72344
rect 102558 72024 102614 72033
rect 102558 71959 102614 71968
rect 102650 71888 102706 71897
rect 102650 71823 102706 71832
rect 101362 71208 101418 71217
rect 101206 71180 101362 71194
rect 101192 71166 101362 71180
rect 59044 69608 59096 69614
rect 59044 69550 59096 69556
rect 58124 69336 58176 69342
rect 58176 69284 58256 69290
rect 58124 69278 58256 69284
rect 58136 69262 58256 69278
rect 57664 69064 57716 69070
rect 57664 69006 57716 69012
rect 57480 68588 57532 68594
rect 57480 68530 57532 68536
rect 56848 67494 57046 67522
rect 57676 67508 57704 69006
rect 58228 67522 58256 69262
rect 58228 67494 58426 67522
rect 59056 67508 59084 69550
rect 59412 69472 59464 69478
rect 59412 69414 59464 69420
rect 59424 69290 59452 69414
rect 60148 69404 60200 69410
rect 60148 69346 60200 69352
rect 59424 69262 59636 69290
rect 59608 67522 59636 69262
rect 60160 67522 60188 69346
rect 62724 69064 62776 69070
rect 62724 69006 62776 69012
rect 62356 68248 62408 68254
rect 62356 68190 62408 68196
rect 59608 67494 59806 67522
rect 60160 67494 60450 67522
rect 62368 63329 62396 68190
rect 62736 66185 62764 69006
rect 62908 68928 62960 68934
rect 62908 68870 62960 68876
rect 62816 68860 62868 68866
rect 62816 68802 62868 68808
rect 62828 66729 62856 68802
rect 62814 66720 62870 66729
rect 62814 66655 62870 66664
rect 62722 66176 62778 66185
rect 62722 66111 62778 66120
rect 62920 65641 62948 68870
rect 63000 68316 63052 68322
rect 63000 68258 63052 68264
rect 62906 65632 62962 65641
rect 62906 65567 62962 65576
rect 62816 65392 62868 65398
rect 62816 65334 62868 65340
rect 62724 65324 62776 65330
rect 62724 65266 62776 65272
rect 62736 64417 62764 65266
rect 62828 64961 62856 65334
rect 62814 64952 62870 64961
rect 62814 64887 62870 64896
rect 62722 64408 62778 64417
rect 62722 64343 62778 64352
rect 63012 63873 63040 68258
rect 63472 68254 63500 70908
rect 64576 68322 64604 70908
rect 64564 68316 64616 68322
rect 64564 68258 64616 68264
rect 63460 68248 63512 68254
rect 63460 68190 63512 68196
rect 63368 68180 63420 68186
rect 63368 68122 63420 68128
rect 63380 67273 63408 68122
rect 63366 67264 63422 67273
rect 63366 67199 63422 67208
rect 63276 65596 63328 65602
rect 63276 65538 63328 65544
rect 62998 63864 63054 63873
rect 62998 63799 63054 63808
rect 62354 63320 62410 63329
rect 62354 63255 62410 63264
rect 62816 63012 62868 63018
rect 62816 62954 62868 62960
rect 29234 62912 29290 62921
rect 29234 62847 29290 62856
rect 29248 62678 29276 62847
rect 13320 62672 13372 62678
rect 13320 62614 13372 62620
rect 29236 62672 29288 62678
rect 29236 62614 29288 62620
rect 12030 41288 12086 41297
rect 12030 41223 12086 41232
rect 13332 19673 13360 62614
rect 62724 61788 62776 61794
rect 62724 61730 62776 61736
rect 62632 60156 62684 60162
rect 62632 60098 62684 60104
rect 62644 57617 62672 60098
rect 62736 59249 62764 61730
rect 62828 60473 62856 62954
rect 63288 62785 63316 65538
rect 65680 65330 65708 70908
rect 66508 70894 66798 70922
rect 66508 68202 66536 70894
rect 67888 68934 67916 70908
rect 68992 69070 69020 70908
rect 68980 69064 69032 69070
rect 68980 69006 69032 69012
rect 67876 68928 67928 68934
rect 67876 68870 67928 68876
rect 70096 68866 70124 70908
rect 70832 70894 71214 70922
rect 70084 68860 70136 68866
rect 70084 68802 70136 68808
rect 70832 68322 70860 70894
rect 70820 68316 70872 68322
rect 70820 68258 70872 68264
rect 71004 68316 71056 68322
rect 71004 68258 71056 68264
rect 66324 68174 66536 68202
rect 69164 68248 69216 68254
rect 69164 68190 69216 68196
rect 66324 65398 66352 68174
rect 69176 65754 69204 68190
rect 71016 65754 71044 68258
rect 72304 68254 72332 70908
rect 73408 68322 73436 70908
rect 73396 68316 73448 68322
rect 73396 68258 73448 68264
rect 74512 68254 74540 70908
rect 75616 68458 75644 70908
rect 76536 70894 76826 70922
rect 74592 68452 74644 68458
rect 74592 68394 74644 68400
rect 75604 68452 75656 68458
rect 75604 68394 75656 68400
rect 72292 68248 72344 68254
rect 72292 68190 72344 68196
rect 72844 68248 72896 68254
rect 72844 68190 72896 68196
rect 74500 68248 74552 68254
rect 74500 68190 74552 68196
rect 72856 65754 72884 68190
rect 74604 65754 74632 68394
rect 76536 65754 76564 70894
rect 68868 65726 69204 65754
rect 70708 65726 71044 65754
rect 72548 65726 72884 65754
rect 74480 65726 74632 65754
rect 76320 65726 76564 65754
rect 77916 65754 77944 70908
rect 79034 70894 79692 70922
rect 79664 65754 79692 70894
rect 80124 68254 80152 70908
rect 81228 68322 81256 70908
rect 82332 68866 82360 70908
rect 83436 68934 83464 70908
rect 83424 68928 83476 68934
rect 83424 68870 83476 68876
rect 82320 68860 82372 68866
rect 82320 68802 82372 68808
rect 81216 68316 81268 68322
rect 81216 68258 81268 68264
rect 83516 68316 83568 68322
rect 83516 68258 83568 68264
rect 80112 68248 80164 68254
rect 80112 68190 80164 68196
rect 81676 68248 81728 68254
rect 81676 68190 81728 68196
rect 81688 65754 81716 68190
rect 83528 65754 83556 68258
rect 84540 68254 84568 70908
rect 85356 68860 85408 68866
rect 85356 68802 85408 68808
rect 84528 68248 84580 68254
rect 84528 68190 84580 68196
rect 85368 65754 85396 68802
rect 85644 68322 85672 70908
rect 86748 68390 86776 70908
rect 87852 68934 87880 70908
rect 88956 69002 88984 70908
rect 90152 69818 90180 70908
rect 90140 69812 90192 69818
rect 90140 69754 90192 69760
rect 91256 69313 91284 70908
rect 91242 69304 91298 69313
rect 91242 69239 91298 69248
rect 92360 69070 92388 70908
rect 92348 69064 92400 69070
rect 92348 69006 92400 69012
rect 88944 68996 88996 69002
rect 88944 68938 88996 68944
rect 87196 68928 87248 68934
rect 87196 68870 87248 68876
rect 87840 68928 87892 68934
rect 87840 68870 87892 68876
rect 86736 68384 86788 68390
rect 86736 68326 86788 68332
rect 85632 68316 85684 68322
rect 85632 68258 85684 68264
rect 87208 65754 87236 68870
rect 93464 68866 93492 70908
rect 93452 68860 93504 68866
rect 93452 68802 93504 68808
rect 94568 68458 94596 70908
rect 94740 68928 94792 68934
rect 94740 68870 94792 68876
rect 94556 68452 94608 68458
rect 94556 68394 94608 68400
rect 92808 68384 92860 68390
rect 92808 68326 92860 68332
rect 90968 68316 91020 68322
rect 90968 68258 91020 68264
rect 89128 68248 89180 68254
rect 89128 68190 89180 68196
rect 89140 65754 89168 68190
rect 90980 65754 91008 68258
rect 92820 65754 92848 68326
rect 94752 65754 94780 68870
rect 95672 68322 95700 70908
rect 95660 68316 95712 68322
rect 95660 68258 95712 68264
rect 96776 66010 96804 70908
rect 97040 69064 97092 69070
rect 97040 69006 97092 69012
rect 96856 68996 96908 69002
rect 96856 68938 96908 68944
rect 96764 66004 96816 66010
rect 96764 65946 96816 65952
rect 96868 65754 96896 68938
rect 77916 65726 78160 65754
rect 79664 65726 80092 65754
rect 81688 65726 81932 65754
rect 83528 65726 83864 65754
rect 85368 65726 85704 65754
rect 87208 65726 87544 65754
rect 89140 65726 89476 65754
rect 90980 65726 91316 65754
rect 92820 65726 93156 65754
rect 94752 65726 95088 65754
rect 96868 65726 96928 65754
rect 66404 65596 66456 65602
rect 66404 65538 66456 65544
rect 66416 65505 66444 65538
rect 66402 65496 66458 65505
rect 66402 65431 66458 65440
rect 66312 65392 66364 65398
rect 66312 65334 66364 65340
rect 65668 65324 65720 65330
rect 65668 65266 65720 65272
rect 66402 64952 66458 64961
rect 66402 64887 66458 64896
rect 66416 64378 66444 64887
rect 63552 64372 63604 64378
rect 63552 64314 63604 64320
rect 66404 64372 66456 64378
rect 66404 64314 66456 64320
rect 63460 64236 63512 64242
rect 63460 64178 63512 64184
rect 63274 62776 63330 62785
rect 63184 62740 63236 62746
rect 63274 62711 63330 62720
rect 63184 62682 63236 62688
rect 63196 61017 63224 62682
rect 63472 61561 63500 64178
rect 63564 62105 63592 64314
rect 66402 64272 66458 64281
rect 66402 64207 66404 64216
rect 66456 64207 66458 64216
rect 66404 64178 66456 64184
rect 97052 63834 97080 69006
rect 97880 68390 97908 70908
rect 97868 68384 97920 68390
rect 97868 68326 97920 68332
rect 98984 68254 99012 70908
rect 98972 68248 99024 68254
rect 98972 68190 99024 68196
rect 100088 68118 100116 70908
rect 101192 68662 101220 71166
rect 101362 71143 101418 71152
rect 101914 71072 101970 71081
rect 101970 71044 102310 71058
rect 101970 71030 102324 71044
rect 101914 71007 101970 71016
rect 102296 68730 102324 71030
rect 102664 70945 102692 71823
rect 102650 70936 102706 70945
rect 102650 70871 102706 70880
rect 102836 68860 102888 68866
rect 102836 68802 102888 68808
rect 102284 68724 102336 68730
rect 102284 68666 102336 68672
rect 101180 68656 101232 68662
rect 101180 68598 101232 68604
rect 102744 68452 102796 68458
rect 102744 68394 102796 68400
rect 102560 68384 102612 68390
rect 102560 68326 102612 68332
rect 100352 68248 100404 68254
rect 100352 68190 100404 68196
rect 100076 68112 100128 68118
rect 100076 68054 100128 68060
rect 100364 67574 100392 68190
rect 102468 68112 102520 68118
rect 102468 68054 102520 68060
rect 100352 67568 100404 67574
rect 100352 67510 100404 67516
rect 102376 67568 102428 67574
rect 102480 67545 102508 68054
rect 102376 67510 102428 67516
rect 102466 67536 102522 67545
rect 102388 67001 102416 67510
rect 102466 67471 102522 67480
rect 102374 66992 102430 67001
rect 102374 66927 102430 66936
rect 102572 66457 102600 68326
rect 102652 68316 102704 68322
rect 102652 68258 102704 68264
rect 102558 66448 102614 66457
rect 102558 66383 102614 66392
rect 102376 66004 102428 66010
rect 102376 65946 102428 65952
rect 102388 65913 102416 65946
rect 102374 65904 102430 65913
rect 102374 65839 102430 65848
rect 100902 65496 100958 65505
rect 100902 65431 100904 65440
rect 100956 65431 100958 65440
rect 102560 65460 102612 65466
rect 100904 65402 100956 65408
rect 102560 65402 102612 65408
rect 100626 64544 100682 64553
rect 100626 64479 100682 64488
rect 100640 64378 100668 64479
rect 100628 64372 100680 64378
rect 100628 64314 100680 64320
rect 102468 64372 102520 64378
rect 102468 64314 102520 64320
rect 100902 64136 100958 64145
rect 100902 64071 100904 64080
rect 100956 64071 100958 64080
rect 100904 64042 100956 64048
rect 97040 63828 97092 63834
rect 97040 63770 97092 63776
rect 102376 63828 102428 63834
rect 102376 63770 102428 63776
rect 66310 63728 66366 63737
rect 66310 63663 66366 63672
rect 66324 62746 66352 63663
rect 102388 63601 102416 63770
rect 102374 63592 102430 63601
rect 102374 63527 102430 63536
rect 100442 63320 100498 63329
rect 100442 63255 100498 63264
rect 66402 63184 66458 63193
rect 66402 63119 66458 63128
rect 66416 63018 66444 63119
rect 100456 63018 100484 63255
rect 66404 63012 66456 63018
rect 66404 62954 66456 62960
rect 100444 63012 100496 63018
rect 100444 62954 100496 62960
rect 102376 63012 102428 63018
rect 102376 62954 102428 62960
rect 100902 62776 100958 62785
rect 66312 62740 66364 62746
rect 100902 62711 100904 62720
rect 66312 62682 66364 62688
rect 100956 62711 100958 62720
rect 100904 62682 100956 62688
rect 66310 62504 66366 62513
rect 66310 62439 66366 62448
rect 63550 62096 63606 62105
rect 63550 62031 63606 62040
rect 63458 61552 63514 61561
rect 66324 61522 66352 62439
rect 100258 62096 100314 62105
rect 100258 62031 100314 62040
rect 66402 61960 66458 61969
rect 66402 61895 66458 61904
rect 66416 61794 66444 61895
rect 66404 61788 66456 61794
rect 66404 61730 66456 61736
rect 63458 61487 63514 61496
rect 63736 61516 63788 61522
rect 63736 61458 63788 61464
rect 66312 61516 66364 61522
rect 66312 61458 66364 61464
rect 63182 61008 63238 61017
rect 63182 60943 63238 60952
rect 62814 60464 62870 60473
rect 62814 60399 62870 60408
rect 63748 60201 63776 61458
rect 100272 61318 100300 62031
rect 100902 61416 100958 61425
rect 100902 61351 100904 61360
rect 100956 61351 100958 61360
rect 100904 61322 100956 61328
rect 100260 61312 100312 61318
rect 66218 61280 66274 61289
rect 102388 61289 102416 62954
rect 102480 62377 102508 64314
rect 102572 63057 102600 65402
rect 102664 65233 102692 68258
rect 102650 65224 102706 65233
rect 102650 65159 102706 65168
rect 102756 64689 102784 68394
rect 102742 64680 102798 64689
rect 102742 64615 102798 64624
rect 102848 64145 102876 68802
rect 105240 67794 105268 75223
rect 105208 67766 105268 67794
rect 105424 67794 105452 76447
rect 106344 67794 106372 77807
rect 106422 74200 106478 74209
rect 106478 74158 106556 74186
rect 106422 74135 106478 74144
rect 106528 70566 106556 74158
rect 106516 70560 106568 70566
rect 106516 70502 106568 70508
rect 106988 67794 107016 79303
rect 107540 67794 107568 79682
rect 108092 67794 108120 80566
rect 108356 72396 108408 72402
rect 108356 72338 108408 72344
rect 105424 67766 105760 67794
rect 106312 67766 106372 67794
rect 106956 67766 107016 67794
rect 107508 67766 107568 67794
rect 108060 67766 108120 67794
rect 108368 67794 108396 72338
rect 108552 72033 108580 81994
rect 108644 74345 108672 83354
rect 108736 78969 108764 86074
rect 108816 84772 108868 84778
rect 108816 84714 108868 84720
rect 108722 78960 108778 78969
rect 108722 78895 108778 78904
rect 108828 76657 108856 84714
rect 132564 79338 132592 88726
rect 132552 79332 132604 79338
rect 132552 79274 132604 79280
rect 132552 79196 132604 79202
rect 132552 79138 132604 79144
rect 108814 76648 108870 76657
rect 108814 76583 108870 76592
rect 108630 74336 108686 74345
rect 108630 74271 108686 74280
rect 108538 72024 108594 72033
rect 108538 71959 108594 71968
rect 109276 70560 109328 70566
rect 109276 70502 109328 70508
rect 109288 67794 109316 70502
rect 110564 68520 110616 68526
rect 110564 68462 110616 68468
rect 110104 68452 110156 68458
rect 110104 68394 110156 68400
rect 110116 67794 110144 68394
rect 110576 67794 110604 68462
rect 111128 68458 111156 70908
rect 111496 68526 111524 70908
rect 111588 70894 111878 70922
rect 111956 70894 112338 70922
rect 112416 70894 112706 70922
rect 111484 68520 111536 68526
rect 111484 68462 111536 68468
rect 111116 68452 111168 68458
rect 111116 68394 111168 68400
rect 111588 67930 111616 70894
rect 111404 67902 111616 67930
rect 111404 67794 111432 67902
rect 111956 67794 111984 70894
rect 112416 67794 112444 70894
rect 113060 67794 113088 70908
rect 113336 70894 113534 70922
rect 113902 70894 114008 70922
rect 113336 67794 113364 70894
rect 113980 67794 114008 70894
rect 108368 67766 108704 67794
rect 109256 67766 109316 67794
rect 109808 67766 110144 67794
rect 110452 67766 110604 67794
rect 111004 67766 111432 67794
rect 111556 67766 111984 67794
rect 112200 67766 112444 67794
rect 112752 67766 113088 67794
rect 113304 67766 113364 67794
rect 113948 67766 114008 67794
rect 114256 67794 114284 70908
rect 114730 70894 114928 70922
rect 115098 70894 115388 70922
rect 115466 70894 115848 70922
rect 115926 70894 116216 70922
rect 114900 67794 114928 70894
rect 115360 67794 115388 70894
rect 115820 68338 115848 70894
rect 116188 68338 116216 70894
rect 116280 68458 116308 70908
rect 116648 68526 116676 70908
rect 117108 68633 117136 70908
rect 117476 69138 117504 70908
rect 117844 69177 117872 70908
rect 118304 69206 118332 70908
rect 118292 69200 118344 69206
rect 117830 69168 117886 69177
rect 117464 69132 117516 69138
rect 118292 69142 118344 69148
rect 117830 69103 117886 69112
rect 117464 69074 117516 69080
rect 118672 69070 118700 70908
rect 119028 69132 119080 69138
rect 119028 69074 119080 69080
rect 118660 69064 118712 69070
rect 118660 69006 118712 69012
rect 117094 68624 117150 68633
rect 117094 68559 117150 68568
rect 118198 68624 118254 68633
rect 118198 68559 118254 68568
rect 116636 68520 116688 68526
rect 116636 68462 116688 68468
rect 117648 68520 117700 68526
rect 117648 68462 117700 68468
rect 116268 68452 116320 68458
rect 116268 68394 116320 68400
rect 117096 68452 117148 68458
rect 117096 68394 117148 68400
rect 115820 68310 115940 68338
rect 116188 68310 116400 68338
rect 115912 67794 115940 68310
rect 116372 67794 116400 68310
rect 117108 67794 117136 68394
rect 117660 67794 117688 68462
rect 118212 67794 118240 68559
rect 119040 67794 119068 69074
rect 119132 68497 119160 70908
rect 119394 69168 119450 69177
rect 119394 69103 119450 69112
rect 119118 68488 119174 68497
rect 119118 68423 119174 68432
rect 119408 67794 119436 69103
rect 119500 68526 119528 70908
rect 119488 68520 119540 68526
rect 119488 68462 119540 68468
rect 119868 68390 119896 70908
rect 120328 69342 120356 70908
rect 120316 69336 120368 69342
rect 120316 69278 120368 69284
rect 120316 69200 120368 69206
rect 120316 69142 120368 69148
rect 119856 68384 119908 68390
rect 119856 68326 119908 68332
rect 120328 67794 120356 69142
rect 120592 69064 120644 69070
rect 120592 69006 120644 69012
rect 114256 67766 114500 67794
rect 114900 67766 115052 67794
rect 115360 67766 115696 67794
rect 115912 67766 116032 67794
rect 116372 67766 116800 67794
rect 117108 67766 117444 67794
rect 117660 67766 117996 67794
rect 118212 67766 118548 67794
rect 119040 67766 119192 67794
rect 119408 67766 119744 67794
rect 120296 67766 120356 67794
rect 120604 67794 120632 69006
rect 120696 68594 120724 70908
rect 120684 68588 120736 68594
rect 120684 68530 120736 68536
rect 121064 68254 121092 70908
rect 121142 68488 121198 68497
rect 121142 68423 121198 68432
rect 121052 68248 121104 68254
rect 121052 68190 121104 68196
rect 121156 67794 121184 68423
rect 121524 68322 121552 70908
rect 121892 68798 121920 70908
rect 122260 68866 122288 70908
rect 122720 69138 122748 70908
rect 123102 70894 123392 70922
rect 123470 70894 123760 70922
rect 123076 69336 123128 69342
rect 123076 69278 123128 69284
rect 122708 69132 122760 69138
rect 122708 69074 122760 69080
rect 122248 68860 122300 68866
rect 122248 68802 122300 68808
rect 121880 68792 121932 68798
rect 121880 68734 121932 68740
rect 121696 68520 121748 68526
rect 121696 68462 121748 68468
rect 121512 68316 121564 68322
rect 121512 68258 121564 68264
rect 121708 67794 121736 68462
rect 122340 68384 122392 68390
rect 122340 68326 122392 68332
rect 122352 67794 122380 68326
rect 123088 67794 123116 69278
rect 123364 68390 123392 70894
rect 123732 69070 123760 70894
rect 123720 69064 123772 69070
rect 123720 69006 123772 69012
rect 123444 68588 123496 68594
rect 123444 68530 123496 68536
rect 123352 68384 123404 68390
rect 123352 68326 123404 68332
rect 123456 67794 123484 68530
rect 123916 68526 123944 70908
rect 124284 68934 124312 70908
rect 124666 70894 125048 70922
rect 124272 68928 124324 68934
rect 124272 68870 124324 68876
rect 125020 68594 125048 70894
rect 125112 69274 125140 70908
rect 125100 69268 125152 69274
rect 125100 69210 125152 69216
rect 125480 69002 125508 70908
rect 125848 69206 125876 70908
rect 126308 69546 126336 70908
rect 126296 69540 126348 69546
rect 126296 69482 126348 69488
rect 125836 69200 125888 69206
rect 125836 69142 125888 69148
rect 126676 69138 126704 70908
rect 131632 69608 131684 69614
rect 131632 69550 131684 69556
rect 129884 69268 129936 69274
rect 129884 69210 129936 69216
rect 129896 69154 129924 69210
rect 131264 69200 131316 69206
rect 126480 69132 126532 69138
rect 126480 69074 126532 69080
rect 126664 69132 126716 69138
rect 129896 69126 130016 69154
rect 131316 69148 131396 69154
rect 131264 69142 131396 69148
rect 131276 69126 131396 69142
rect 126664 69074 126716 69080
rect 125468 68996 125520 69002
rect 125468 68938 125520 68944
rect 125836 68860 125888 68866
rect 125836 68802 125888 68808
rect 125192 68792 125244 68798
rect 125192 68734 125244 68740
rect 125008 68588 125060 68594
rect 125008 68530 125060 68536
rect 123904 68520 123956 68526
rect 123904 68462 123956 68468
rect 124640 68316 124692 68322
rect 124640 68258 124692 68264
rect 124456 68248 124508 68254
rect 124456 68190 124508 68196
rect 124468 67794 124496 68190
rect 120604 67766 120940 67794
rect 121156 67766 121492 67794
rect 121708 67766 122044 67794
rect 122352 67766 122688 67794
rect 123088 67766 123240 67794
rect 123456 67766 123792 67794
rect 124436 67766 124496 67794
rect 124652 67794 124680 68258
rect 125204 67794 125232 68734
rect 125848 67794 125876 68802
rect 126492 67794 126520 69074
rect 127584 69064 127636 69070
rect 127584 69006 127636 69012
rect 127308 68384 127360 68390
rect 127308 68326 127360 68332
rect 124652 67766 124988 67794
rect 125204 67766 125540 67794
rect 125848 67766 126184 67794
rect 126492 67766 126736 67794
rect 116004 67658 116032 67766
rect 127320 67658 127348 68326
rect 127596 67794 127624 69006
rect 128688 68928 128740 68934
rect 128688 68870 128740 68876
rect 128136 68520 128188 68526
rect 128136 68462 128188 68468
rect 128148 67794 128176 68462
rect 128700 67794 128728 68870
rect 129332 68588 129384 68594
rect 129332 68530 129384 68536
rect 129344 67794 129372 68530
rect 129988 67794 130016 69126
rect 130436 68996 130488 69002
rect 130436 68938 130488 68944
rect 130448 67794 130476 68938
rect 131368 68066 131396 69126
rect 131368 68038 131442 68066
rect 127596 67766 127932 67794
rect 128148 67766 128484 67794
rect 128700 67766 129036 67794
rect 129344 67766 129680 67794
rect 129988 67766 130232 67794
rect 130448 67766 130784 67794
rect 131414 67780 131442 68038
rect 116004 67630 116248 67658
rect 127288 67630 127348 67658
rect 131644 67658 131672 69550
rect 132184 69132 132236 69138
rect 132184 69074 132236 69080
rect 132196 67794 132224 69074
rect 132564 68322 132592 79138
rect 174424 72962 174452 142582
rect 175240 142232 175292 142238
rect 175238 142200 175240 142209
rect 175292 142200 175294 142209
rect 175238 142135 175294 142144
rect 175424 142164 175476 142170
rect 175424 142106 175476 142112
rect 175148 142096 175200 142102
rect 175148 142038 175200 142044
rect 174780 141212 174832 141218
rect 174780 141154 174832 141160
rect 174792 140985 174820 141154
rect 174778 140976 174834 140985
rect 174778 140911 174834 140920
rect 174964 139920 175016 139926
rect 174964 139862 175016 139868
rect 174976 139761 175004 139862
rect 174962 139752 175018 139761
rect 174962 139687 175018 139696
rect 175160 138401 175188 142038
rect 175436 138945 175464 142106
rect 177184 141764 177212 149887
rect 177354 147640 177410 147649
rect 177354 147575 177410 147584
rect 177368 146930 177396 147575
rect 177356 146924 177408 146930
rect 177356 146866 177408 146872
rect 177460 141778 177488 150046
rect 178288 146182 178316 154511
rect 178550 153352 178606 153361
rect 178550 153287 178606 153296
rect 178458 152264 178514 152273
rect 178458 152199 178514 152208
rect 178366 148864 178422 148873
rect 178366 148799 178422 148808
rect 178276 146176 178328 146182
rect 178276 146118 178328 146124
rect 178380 145162 178408 148799
rect 178368 145156 178420 145162
rect 178368 145098 178420 145104
rect 178472 141778 178500 152199
rect 177460 141750 177750 141778
rect 178302 141750 178500 141778
rect 178564 141778 178592 153287
rect 179392 152953 179420 159242
rect 179484 155401 179512 160874
rect 179576 157713 179604 162030
rect 180484 158008 180536 158014
rect 180484 157950 180536 157956
rect 180392 157940 180444 157946
rect 180392 157882 180444 157888
rect 179562 157704 179618 157713
rect 179562 157639 179618 157648
rect 180300 156512 180352 156518
rect 180300 156454 180352 156460
rect 179470 155392 179526 155401
rect 179470 155327 179526 155336
rect 179656 155152 179708 155158
rect 179656 155094 179708 155100
rect 179378 152944 179434 152953
rect 179378 152879 179434 152888
rect 179012 146176 179064 146182
rect 179012 146118 179064 146124
rect 179024 141778 179052 146118
rect 179668 141778 179696 155094
rect 180312 146017 180340 156454
rect 180404 148329 180432 157882
rect 180496 150641 180524 157950
rect 200538 151584 200594 151593
rect 200538 151519 200540 151528
rect 200592 151519 200594 151528
rect 200540 151490 200592 151496
rect 180482 150632 180538 150641
rect 180482 150567 180538 150576
rect 180390 148320 180446 148329
rect 180390 148255 180446 148264
rect 180576 146924 180628 146930
rect 180576 146866 180628 146872
rect 180298 146008 180354 146017
rect 180298 145943 180354 145952
rect 178564 141750 178854 141778
rect 179024 141750 179406 141778
rect 179668 141750 180050 141778
rect 180588 141764 180616 146866
rect 181128 145156 181180 145162
rect 181128 145098 181180 145104
rect 181140 141764 181168 145098
rect 182796 144878 183132 144906
rect 183256 144878 183500 144906
rect 183624 144878 183868 144906
rect 183992 144878 184328 144906
rect 184452 144878 184696 144906
rect 184820 144878 185064 144906
rect 185280 144878 185524 144906
rect 185740 144878 185892 144906
rect 182232 142708 182284 142714
rect 182232 142650 182284 142656
rect 181680 142572 181732 142578
rect 181680 142514 181732 142520
rect 181692 141764 181720 142514
rect 182244 141764 182272 142650
rect 182796 142578 182824 144878
rect 183256 142714 183284 144878
rect 183244 142708 183296 142714
rect 183244 142650 183296 142656
rect 182784 142572 182836 142578
rect 182784 142514 182836 142520
rect 183624 142306 183652 144878
rect 182876 142300 182928 142306
rect 182876 142242 182928 142248
rect 183612 142300 183664 142306
rect 183612 142242 183664 142248
rect 182888 141764 182916 142242
rect 183992 142186 184020 144878
rect 183808 142158 184020 142186
rect 183808 141778 183836 142158
rect 184452 141778 184480 144878
rect 184820 141778 184848 144878
rect 185280 141778 185308 144878
rect 183454 141750 183836 141778
rect 184006 141750 184480 141778
rect 184558 141750 184848 141778
rect 185110 141750 185308 141778
rect 185740 141764 185768 144878
rect 186246 144634 186274 144892
rect 186720 144878 186872 144906
rect 187088 144878 187240 144906
rect 187456 144878 187700 144906
rect 187916 144878 188160 144906
rect 188284 144878 188528 144906
rect 188652 144878 188988 144906
rect 189112 144878 189356 144906
rect 189480 144878 189724 144906
rect 189848 144878 190184 144906
rect 190308 144878 190552 144906
rect 186246 144606 186320 144634
rect 186292 141764 186320 144606
rect 186844 141764 186872 144878
rect 187212 141778 187240 144878
rect 187672 141778 187700 144878
rect 188132 141778 188160 144878
rect 188500 141914 188528 144878
rect 188960 141914 188988 144878
rect 189328 142646 189356 144878
rect 189696 142714 189724 144878
rect 189684 142708 189736 142714
rect 189684 142650 189736 142656
rect 189316 142640 189368 142646
rect 189316 142582 189368 142588
rect 190156 142034 190184 144878
rect 190524 142646 190552 144878
rect 190616 144878 190676 144906
rect 191136 144878 191380 144906
rect 190616 144278 190644 144878
rect 190604 144272 190656 144278
rect 190604 144214 190656 144220
rect 191352 142714 191380 144878
rect 191490 144686 191518 144892
rect 191858 144754 191886 144892
rect 192332 144878 192484 144906
rect 192700 144878 192944 144906
rect 193068 144878 193404 144906
rect 193528 144878 193772 144906
rect 193896 144878 194140 144906
rect 194264 144878 194600 144906
rect 191846 144748 191898 144754
rect 191846 144690 191898 144696
rect 191478 144680 191530 144686
rect 191478 144622 191530 144628
rect 190788 142708 190840 142714
rect 190788 142650 190840 142656
rect 191340 142708 191392 142714
rect 191340 142650 191392 142656
rect 190236 142640 190288 142646
rect 190236 142582 190288 142588
rect 190512 142640 190564 142646
rect 190512 142582 190564 142588
rect 190144 142028 190196 142034
rect 190144 141970 190196 141976
rect 188500 141886 188804 141914
rect 188960 141886 189264 141914
rect 188776 141778 188804 141886
rect 189236 141778 189264 141886
rect 187212 141750 187410 141778
rect 187672 141750 187962 141778
rect 188132 141750 188606 141778
rect 188776 141750 189158 141778
rect 189236 141750 189710 141778
rect 190248 141764 190276 142582
rect 190800 141764 190828 142650
rect 191984 142640 192036 142646
rect 191984 142582 192036 142588
rect 191432 142028 191484 142034
rect 191432 141970 191484 141976
rect 191444 141764 191472 141970
rect 191996 141764 192024 142582
rect 192456 142374 192484 144878
rect 192536 144272 192588 144278
rect 192536 144214 192588 144220
rect 192444 142368 192496 142374
rect 192444 142310 192496 142316
rect 192548 141764 192576 144214
rect 192916 142442 192944 144878
rect 193088 142708 193140 142714
rect 193088 142650 193140 142656
rect 192904 142436 192956 142442
rect 192904 142378 192956 142384
rect 193100 141764 193128 142650
rect 193376 142306 193404 144878
rect 193640 144680 193692 144686
rect 193640 144622 193692 144628
rect 193364 142300 193416 142306
rect 193364 142242 193416 142248
rect 193652 141764 193680 144622
rect 193744 142578 193772 144878
rect 194112 142646 194140 144878
rect 194284 144748 194336 144754
rect 194284 144690 194336 144696
rect 194100 142640 194152 142646
rect 194100 142582 194152 142588
rect 193732 142572 193784 142578
rect 193732 142514 193784 142520
rect 194296 141764 194324 144690
rect 194572 142510 194600 144878
rect 194664 144878 194724 144906
rect 195092 144878 195336 144906
rect 195460 144878 195796 144906
rect 195920 144878 196164 144906
rect 196288 144878 196532 144906
rect 196656 144878 196992 144906
rect 197116 144878 197360 144906
rect 194560 142504 194612 142510
rect 194560 142446 194612 142452
rect 194664 142170 194692 144878
rect 194836 142368 194888 142374
rect 194836 142310 194888 142316
rect 194652 142164 194704 142170
rect 194652 142106 194704 142112
rect 194848 141764 194876 142310
rect 195308 142102 195336 144878
rect 195768 142442 195796 144878
rect 195388 142436 195440 142442
rect 195388 142378 195440 142384
rect 195756 142436 195808 142442
rect 195756 142378 195808 142384
rect 195296 142096 195348 142102
rect 195296 142038 195348 142044
rect 195400 141764 195428 142378
rect 195940 142300 195992 142306
rect 195940 142242 195992 142248
rect 195952 141764 195980 142242
rect 196136 142238 196164 144878
rect 196504 142714 196532 144878
rect 196492 142708 196544 142714
rect 196492 142650 196544 142656
rect 196492 142572 196544 142578
rect 196492 142514 196544 142520
rect 196124 142232 196176 142238
rect 196124 142174 196176 142180
rect 196504 141764 196532 142514
rect 196964 142374 196992 144878
rect 197136 142640 197188 142646
rect 197136 142582 197188 142588
rect 196952 142368 197004 142374
rect 196952 142310 197004 142316
rect 197148 141764 197176 142582
rect 197332 142306 197360 144878
rect 197470 144634 197498 144892
rect 197838 144686 197866 144892
rect 198312 144878 198556 144906
rect 198680 144878 198924 144906
rect 197826 144680 197878 144686
rect 197470 144606 197544 144634
rect 197826 144622 197878 144628
rect 197516 144142 197544 144606
rect 198528 144210 198556 144878
rect 198896 144278 198924 144878
rect 198884 144272 198936 144278
rect 198884 144214 198936 144220
rect 198516 144204 198568 144210
rect 198516 144146 198568 144152
rect 197504 144136 197556 144142
rect 197504 144078 197556 144084
rect 201012 142714 201040 164847
rect 222632 163402 222660 166094
rect 224458 163552 224514 163561
rect 224458 163487 224514 163496
rect 222632 163374 222752 163402
rect 207438 163280 207494 163289
rect 207438 163215 207494 163224
rect 207452 153769 207480 163215
rect 222724 159594 222752 163374
rect 222632 159566 222752 159594
rect 222632 158098 222660 159566
rect 223538 159200 223594 159209
rect 223538 159135 223594 159144
rect 222632 158070 222936 158098
rect 222804 156920 222856 156926
rect 222540 156868 222804 156874
rect 222540 156862 222856 156868
rect 222540 156846 222844 156862
rect 207438 153760 207494 153769
rect 207438 153695 207494 153704
rect 207346 153352 207402 153361
rect 207346 153287 207402 153296
rect 204494 151584 204550 151593
rect 207360 151554 207388 153287
rect 204494 151519 204550 151528
rect 207348 151548 207400 151554
rect 202840 144680 202892 144686
rect 202840 144622 202892 144628
rect 202196 144136 202248 144142
rect 202196 144078 202248 144084
rect 200540 142708 200592 142714
rect 200540 142650 200592 142656
rect 201000 142708 201052 142714
rect 201000 142650 201052 142656
rect 197688 142504 197740 142510
rect 197688 142446 197740 142452
rect 197320 142300 197372 142306
rect 197320 142242 197372 142248
rect 197700 141764 197728 142446
rect 199068 142436 199120 142442
rect 199068 142378 199120 142384
rect 198240 142164 198292 142170
rect 198240 142106 198292 142112
rect 198252 141764 198280 142106
rect 198792 142096 198844 142102
rect 198792 142038 198844 142044
rect 198804 141764 198832 142038
rect 199080 141778 199108 142378
rect 199620 142232 199672 142238
rect 199620 142174 199672 142180
rect 199632 141778 199660 142174
rect 199080 141750 199370 141778
rect 199632 141750 200014 141778
rect 200552 141764 200580 142650
rect 201092 142368 201144 142374
rect 201092 142310 201144 142316
rect 201104 141764 201132 142310
rect 201644 142300 201696 142306
rect 201644 142242 201696 142248
rect 201656 141764 201684 142242
rect 202208 141764 202236 144078
rect 202852 141764 202880 144622
rect 203944 144272 203996 144278
rect 203944 144214 203996 144220
rect 203392 144204 203444 144210
rect 203392 144146 203444 144152
rect 203404 141764 203432 144146
rect 203956 141764 203984 144214
rect 204508 141764 204536 151519
rect 207348 151490 207400 151496
rect 207360 145230 207388 151490
rect 207348 145224 207400 145230
rect 207348 145166 207400 145172
rect 210016 145224 210068 145230
rect 210016 145166 210068 145172
rect 210292 145224 210344 145230
rect 210344 145172 210594 145178
rect 210292 145166 210594 145172
rect 207992 142028 208044 142034
rect 207992 141970 208044 141976
rect 207900 141960 207952 141966
rect 207900 141902 207952 141908
rect 175422 138936 175478 138945
rect 175422 138871 175478 138880
rect 175146 138392 175202 138401
rect 175146 138327 175202 138336
rect 207254 137168 207310 137177
rect 207254 137103 207310 137112
rect 174504 136044 174556 136050
rect 174504 135986 174556 135992
rect 174516 133641 174544 135986
rect 174502 133632 174558 133641
rect 174502 133567 174558 133576
rect 175332 133596 175384 133602
rect 175332 133538 175384 133544
rect 174872 133120 174924 133126
rect 174872 133062 174924 133068
rect 174884 131329 174912 133062
rect 175148 131828 175200 131834
rect 175148 131770 175200 131776
rect 174870 131320 174926 131329
rect 174870 131255 174926 131264
rect 175160 129561 175188 131770
rect 175240 131760 175292 131766
rect 175240 131702 175292 131708
rect 175252 130241 175280 131702
rect 175344 131601 175372 133538
rect 175424 131964 175476 131970
rect 175424 131906 175476 131912
rect 175330 131592 175386 131601
rect 175330 131527 175386 131536
rect 175436 130785 175464 131906
rect 175422 130776 175478 130785
rect 175422 130711 175478 130720
rect 175238 130232 175294 130241
rect 175238 130167 175294 130176
rect 175146 129552 175202 129561
rect 175146 129487 175202 129496
rect 174504 129108 174556 129114
rect 174504 129050 174556 129056
rect 174516 127249 174544 129050
rect 174596 127612 174648 127618
rect 174596 127554 174648 127560
rect 174502 127240 174558 127249
rect 174502 127175 174558 127184
rect 174504 126252 174556 126258
rect 174504 126194 174556 126200
rect 174516 124393 174544 126194
rect 174608 126025 174636 127554
rect 174594 126016 174650 126025
rect 174594 125951 174650 125960
rect 174596 124892 174648 124898
rect 174596 124834 174648 124840
rect 174502 124384 174558 124393
rect 174502 124319 174558 124328
rect 174608 123169 174636 124834
rect 175332 123532 175384 123538
rect 175332 123474 175384 123480
rect 174594 123160 174650 123169
rect 174594 123095 174650 123104
rect 175056 122444 175108 122450
rect 175056 122386 175108 122392
rect 175068 121401 175096 122386
rect 175148 122036 175200 122042
rect 175148 121978 175200 121984
rect 175054 121392 175110 121401
rect 175054 121327 175110 121336
rect 175160 120313 175188 121978
rect 175344 121673 175372 123474
rect 175424 122172 175476 122178
rect 175424 122114 175476 122120
rect 175330 121664 175386 121673
rect 175330 121599 175386 121608
rect 175436 120585 175464 122114
rect 175422 120576 175478 120585
rect 175422 120511 175478 120520
rect 175146 120304 175202 120313
rect 175146 120239 175202 120248
rect 174504 119452 174556 119458
rect 174504 119394 174556 119400
rect 174516 117865 174544 119394
rect 204678 117992 204734 118001
rect 204678 117927 204734 117936
rect 174502 117856 174558 117865
rect 174502 117791 174558 117800
rect 176908 113870 177198 113898
rect 177368 113870 177750 113898
rect 176908 102225 176936 113870
rect 177080 111156 177132 111162
rect 177080 111098 177132 111104
rect 176988 111088 177040 111094
rect 176988 111030 177040 111036
rect 177000 106849 177028 111030
rect 176986 106840 177042 106849
rect 176986 106775 177042 106784
rect 177092 105761 177120 111098
rect 177264 111020 177316 111026
rect 177264 110962 177316 110968
rect 177172 109524 177224 109530
rect 177172 109466 177224 109472
rect 177184 109161 177212 109466
rect 177170 109152 177226 109161
rect 177170 109087 177226 109096
rect 177276 107937 177304 110962
rect 177262 107928 177318 107937
rect 177262 107863 177318 107872
rect 177078 105752 177134 105761
rect 177078 105687 177134 105696
rect 177368 103449 177396 113870
rect 178288 111230 178316 113884
rect 177448 111224 177500 111230
rect 177448 111166 177500 111172
rect 178276 111224 178328 111230
rect 178276 111166 178328 111172
rect 177460 104537 177488 111166
rect 178840 111162 178868 113884
rect 178828 111156 178880 111162
rect 178828 111098 178880 111104
rect 179392 111094 179420 113884
rect 179380 111088 179432 111094
rect 179380 111030 179432 111036
rect 180036 111026 180064 113884
rect 180024 111020 180076 111026
rect 180024 110962 180076 110968
rect 177724 110952 177776 110958
rect 177724 110894 177776 110900
rect 177736 110249 177764 110894
rect 177722 110240 177778 110249
rect 177722 110175 177778 110184
rect 180298 109560 180354 109569
rect 180588 109530 180616 113884
rect 181140 110958 181168 113884
rect 181692 111026 181720 113884
rect 182244 111434 182272 113884
rect 182232 111428 182284 111434
rect 182232 111370 182284 111376
rect 182888 111366 182916 113884
rect 183244 111428 183296 111434
rect 183244 111370 183296 111376
rect 182876 111360 182928 111366
rect 182876 111302 182928 111308
rect 181680 111020 181732 111026
rect 181680 110962 181732 110968
rect 183106 111020 183158 111026
rect 183106 110962 183158 110968
rect 181128 110952 181180 110958
rect 181128 110894 181180 110900
rect 183118 110756 183146 110962
rect 183256 110770 183284 111370
rect 183440 111026 183468 113884
rect 184006 113870 184480 113898
rect 184558 113870 184848 113898
rect 183796 111360 183848 111366
rect 183796 111302 183848 111308
rect 183428 111020 183480 111026
rect 183428 110962 183480 110968
rect 183808 110770 183836 111302
rect 184302 111020 184354 111026
rect 184302 110962 184354 110968
rect 183256 110742 183500 110770
rect 183808 110742 183868 110770
rect 184314 110756 184342 110962
rect 184452 110770 184480 113870
rect 184820 110770 184848 113870
rect 185096 111042 185124 113884
rect 185096 111014 185216 111042
rect 185188 110770 185216 111014
rect 185740 110770 185768 113884
rect 186292 111042 186320 113884
rect 186246 111014 186320 111042
rect 184452 110742 184696 110770
rect 184820 110742 185064 110770
rect 185188 110742 185524 110770
rect 185740 110742 185892 110770
rect 186246 110756 186274 111014
rect 186844 110770 186872 113884
rect 187212 113870 187410 113898
rect 187764 113870 187962 113898
rect 188132 113870 188606 113898
rect 188684 113870 189158 113898
rect 189328 113870 189710 113898
rect 187212 110770 187240 113870
rect 187764 110770 187792 113870
rect 188132 110770 188160 113870
rect 188684 110906 188712 113870
rect 189328 111314 189356 113870
rect 190248 113134 190276 113884
rect 189408 113128 189460 113134
rect 189408 113070 189460 113076
rect 190236 113128 190288 113134
rect 190236 113070 190288 113076
rect 188408 110878 188712 110906
rect 188868 111286 189356 111314
rect 188408 110770 188436 110878
rect 188868 110770 188896 111286
rect 189420 111042 189448 113070
rect 190512 112584 190564 112590
rect 190512 112526 190564 112532
rect 190144 112516 190196 112522
rect 190144 112458 190196 112464
rect 189684 112448 189736 112454
rect 189684 112390 189736 112396
rect 189236 111014 189448 111042
rect 189236 110770 189264 111014
rect 189696 110770 189724 112390
rect 190156 110770 190184 112458
rect 190524 110770 190552 112526
rect 190800 112454 190828 113884
rect 191340 113128 191392 113134
rect 191340 113070 191392 113076
rect 190788 112448 190840 112454
rect 190788 112390 190840 112396
rect 190604 112108 190656 112114
rect 190604 112050 190656 112056
rect 186720 110742 186872 110770
rect 187088 110742 187240 110770
rect 187456 110742 187792 110770
rect 187916 110742 188160 110770
rect 188284 110742 188436 110770
rect 188652 110742 188896 110770
rect 189112 110742 189264 110770
rect 189480 110742 189724 110770
rect 189848 110742 190184 110770
rect 190308 110742 190552 110770
rect 190616 110770 190644 112050
rect 191352 110770 191380 113070
rect 191444 112522 191472 113884
rect 191996 112590 192024 113884
rect 192272 113870 192562 113898
rect 191984 112584 192036 112590
rect 191984 112526 192036 112532
rect 191432 112516 191484 112522
rect 191432 112458 191484 112464
rect 192272 112114 192300 113870
rect 193100 113134 193128 113884
rect 193088 113128 193140 113134
rect 193088 113070 193140 113076
rect 192536 112584 192588 112590
rect 192536 112526 192588 112532
rect 192260 112108 192312 112114
rect 192260 112050 192312 112056
rect 191984 111428 192036 111434
rect 191984 111370 192036 111376
rect 191708 111360 191760 111366
rect 191708 111302 191760 111308
rect 191720 110770 191748 111302
rect 191996 110770 192024 111370
rect 192548 110770 192576 112526
rect 192904 112448 192956 112454
rect 192904 112390 192956 112396
rect 192916 110770 192944 112390
rect 193180 112380 193232 112386
rect 193180 112322 193232 112328
rect 193192 110770 193220 112322
rect 193652 111366 193680 113884
rect 193732 113128 193784 113134
rect 193732 113070 193784 113076
rect 193640 111360 193692 111366
rect 193640 111302 193692 111308
rect 193744 110770 193772 113070
rect 194192 112380 194244 112386
rect 194192 112322 194244 112328
rect 194204 112250 194232 112322
rect 194192 112244 194244 112250
rect 194192 112186 194244 112192
rect 194296 111434 194324 113884
rect 194652 113196 194704 113202
rect 194652 113138 194704 113144
rect 194560 112788 194612 112794
rect 194560 112730 194612 112736
rect 194284 111428 194336 111434
rect 194284 111370 194336 111376
rect 194100 111360 194152 111366
rect 194100 111302 194152 111308
rect 194112 110770 194140 111302
rect 194572 110770 194600 112730
rect 190616 110742 190676 110770
rect 191136 110742 191380 110770
rect 191504 110742 191748 110770
rect 191872 110742 192024 110770
rect 192332 110742 192576 110770
rect 192700 110742 192944 110770
rect 193068 110742 193220 110770
rect 193528 110742 193772 110770
rect 193896 110742 194140 110770
rect 194264 110742 194600 110770
rect 194664 110770 194692 113138
rect 194744 112584 194796 112590
rect 194848 112572 194876 113884
rect 194796 112544 194876 112572
rect 194744 112526 194796 112532
rect 195400 112318 195428 113884
rect 195756 113060 195808 113066
rect 195756 113002 195808 113008
rect 195388 112312 195440 112318
rect 195388 112254 195440 112260
rect 195296 111428 195348 111434
rect 195296 111370 195348 111376
rect 195308 110770 195336 111370
rect 195768 110770 195796 113002
rect 195952 112250 195980 113884
rect 196228 113870 196518 113898
rect 196124 113128 196176 113134
rect 196228 113116 196256 113870
rect 196176 113088 196256 113116
rect 196124 113070 196176 113076
rect 196124 112924 196176 112930
rect 196124 112866 196176 112872
rect 195940 112244 195992 112250
rect 195940 112186 195992 112192
rect 196136 110770 196164 112866
rect 196492 112584 196544 112590
rect 196492 112526 196544 112532
rect 196504 110770 196532 112526
rect 196952 112516 197004 112522
rect 196952 112458 197004 112464
rect 196964 110770 196992 112458
rect 197148 111366 197176 113884
rect 197700 112794 197728 113884
rect 198252 113202 198280 113884
rect 198240 113196 198292 113202
rect 198240 113138 198292 113144
rect 198516 113128 198568 113134
rect 198516 113070 198568 113076
rect 197688 112788 197740 112794
rect 197688 112730 197740 112736
rect 197320 112652 197372 112658
rect 197320 112594 197372 112600
rect 197136 111360 197188 111366
rect 197136 111302 197188 111308
rect 197332 110770 197360 112594
rect 197504 112448 197556 112454
rect 197504 112390 197556 112396
rect 197516 111042 197544 112390
rect 198148 112380 198200 112386
rect 198148 112322 198200 112328
rect 194664 110742 194724 110770
rect 195092 110742 195336 110770
rect 195460 110742 195796 110770
rect 195920 110742 196164 110770
rect 196288 110742 196532 110770
rect 196656 110742 196992 110770
rect 197116 110742 197360 110770
rect 197470 111014 197544 111042
rect 197470 110756 197498 111014
rect 198160 110770 198188 112322
rect 198528 110770 198556 113070
rect 198804 111434 198832 113884
rect 199356 113066 199384 113884
rect 199344 113060 199396 113066
rect 199344 113002 199396 113008
rect 198884 112992 198936 112998
rect 198884 112934 198936 112940
rect 198792 111428 198844 111434
rect 198792 111370 198844 111376
rect 198896 110770 198924 112934
rect 200000 112930 200028 113884
rect 199988 112924 200040 112930
rect 199988 112866 200040 112872
rect 200552 112590 200580 113884
rect 200540 112584 200592 112590
rect 200540 112526 200592 112532
rect 201104 112522 201132 113884
rect 201656 112658 201684 113884
rect 201748 113870 202222 113898
rect 201644 112652 201696 112658
rect 201644 112594 201696 112600
rect 201748 112538 201776 113870
rect 201092 112516 201144 112522
rect 201092 112458 201144 112464
rect 201656 112510 201776 112538
rect 201656 112454 201684 112510
rect 201644 112448 201696 112454
rect 201644 112390 201696 112396
rect 202852 112386 202880 113884
rect 203404 113134 203432 113884
rect 203392 113128 203444 113134
rect 203392 113070 203444 113076
rect 203956 112998 203984 113884
rect 204522 113870 204628 113898
rect 203944 112992 203996 112998
rect 203944 112934 203996 112940
rect 202840 112380 202892 112386
rect 202840 112322 202892 112328
rect 197852 110742 198188 110770
rect 198312 110742 198556 110770
rect 198680 110742 198924 110770
rect 180298 109495 180354 109504
rect 180576 109524 180628 109530
rect 179654 107248 179710 107257
rect 179654 107183 179710 107192
rect 179668 106878 179696 107183
rect 177540 106872 177592 106878
rect 177540 106814 177592 106820
rect 179656 106872 179708 106878
rect 179656 106814 179708 106820
rect 177446 104528 177502 104537
rect 177446 104463 177502 104472
rect 177354 103440 177410 103449
rect 177354 103375 177410 103384
rect 176894 102216 176950 102225
rect 176894 102151 176950 102160
rect 176988 101296 177040 101302
rect 176988 101238 177040 101244
rect 177000 101137 177028 101238
rect 176986 101128 177042 101137
rect 176986 101063 177042 101072
rect 177552 100049 177580 106814
rect 179654 104936 179710 104945
rect 179654 104871 179710 104880
rect 179668 104090 179696 104871
rect 177816 104084 177868 104090
rect 177816 104026 177868 104032
rect 179656 104084 179708 104090
rect 179656 104026 179708 104032
rect 177632 101364 177684 101370
rect 177632 101306 177684 101312
rect 177538 100040 177594 100049
rect 177538 99975 177594 99984
rect 177644 97737 177672 101306
rect 177724 99936 177776 99942
rect 177724 99878 177776 99884
rect 177630 97728 177686 97737
rect 177630 97663 177686 97672
rect 177540 97216 177592 97222
rect 177540 97158 177592 97164
rect 177552 95425 177580 97158
rect 177736 96513 177764 99878
rect 177828 98825 177856 104026
rect 179654 102488 179710 102497
rect 179654 102423 179710 102432
rect 179668 101370 179696 102423
rect 179656 101364 179708 101370
rect 179656 101306 179708 101312
rect 180312 101302 180340 109495
rect 180576 109466 180628 109472
rect 204600 104265 204628 113870
rect 204692 113678 204720 117927
rect 204680 113672 204732 113678
rect 204680 113614 204732 113620
rect 207268 113610 207296 137103
rect 207912 118545 207940 141902
rect 208004 127793 208032 141970
rect 210028 141966 210056 145166
rect 210304 145150 210594 145166
rect 215916 142714 215944 144892
rect 215904 142708 215956 142714
rect 215904 142650 215956 142656
rect 221252 142034 221280 144892
rect 222540 142102 222568 156846
rect 222908 156602 222936 158070
rect 223552 156926 223580 159135
rect 223540 156920 223592 156926
rect 223540 156862 223592 156868
rect 222724 156574 222936 156602
rect 222724 146946 222752 156574
rect 223538 149544 223594 149553
rect 223538 149479 223594 149488
rect 222632 146918 222752 146946
rect 222632 146810 222660 146918
rect 222632 146782 222936 146810
rect 222528 142096 222580 142102
rect 222528 142038 222580 142044
rect 222804 142096 222856 142102
rect 222804 142038 222856 142044
rect 221240 142028 221292 142034
rect 221240 141970 221292 141976
rect 210016 141960 210068 141966
rect 210016 141902 210068 141908
rect 222528 141960 222580 141966
rect 222528 141902 222580 141908
rect 207990 127784 208046 127793
rect 207990 127719 208046 127728
rect 207898 118536 207954 118545
rect 207898 118471 207954 118480
rect 207256 113604 207308 113610
rect 207256 113546 207308 113552
rect 201090 104256 201146 104265
rect 201090 104191 201146 104200
rect 204586 104256 204642 104265
rect 204586 104191 204642 104200
rect 180300 101296 180352 101302
rect 180300 101238 180352 101244
rect 179654 100176 179710 100185
rect 179654 100111 179710 100120
rect 179668 99942 179696 100111
rect 179656 99936 179708 99942
rect 179656 99878 179708 99884
rect 177814 98816 177870 98825
rect 177814 98751 177870 98760
rect 179654 97864 179710 97873
rect 179654 97799 179710 97808
rect 179668 97222 179696 97799
rect 179656 97216 179708 97222
rect 179656 97158 179708 97164
rect 177722 96504 177778 96513
rect 177722 96439 177778 96448
rect 177538 95416 177594 95425
rect 177538 95351 177594 95360
rect 179562 95416 179618 95425
rect 179562 95351 179618 95360
rect 179576 94366 179604 95351
rect 177448 94360 177500 94366
rect 177446 94328 177448 94337
rect 179564 94360 179616 94366
rect 177500 94328 177502 94337
rect 179564 94302 179616 94308
rect 177446 94263 177502 94272
rect 177538 92016 177594 92025
rect 177538 91951 177594 91960
rect 177552 91714 177580 91951
rect 177540 91708 177592 91714
rect 177540 91650 177592 91656
rect 179564 91708 179616 91714
rect 179564 91650 179616 91656
rect 179576 90801 179604 91650
rect 201104 91646 201132 104191
rect 201092 91640 201144 91646
rect 201092 91582 201144 91588
rect 204496 91640 204548 91646
rect 204496 91582 204548 91588
rect 204508 90937 204536 91582
rect 204494 90928 204550 90937
rect 204494 90863 204550 90872
rect 177354 90792 177410 90801
rect 177354 90727 177410 90736
rect 179562 90792 179618 90801
rect 179562 90727 179618 90736
rect 177368 90286 177396 90727
rect 200998 90384 201054 90393
rect 200998 90319 201054 90328
rect 177356 90280 177408 90286
rect 177356 90222 177408 90228
rect 179656 90280 179708 90286
rect 179656 90222 179708 90228
rect 177354 89704 177410 89713
rect 177354 89639 177410 89648
rect 177368 89198 177396 89639
rect 177356 89192 177408 89198
rect 177356 89134 177408 89140
rect 179564 89192 179616 89198
rect 179564 89134 179616 89140
rect 177354 88616 177410 88625
rect 177354 88551 177410 88560
rect 177368 88246 177396 88551
rect 177356 88240 177408 88246
rect 177356 88182 177408 88188
rect 179472 88240 179524 88246
rect 179472 88182 179524 88188
rect 178918 87392 178974 87401
rect 178918 87327 178974 87336
rect 178090 86304 178146 86313
rect 178090 86239 178146 86248
rect 178104 86138 178132 86239
rect 178092 86132 178144 86138
rect 178092 86074 178144 86080
rect 177538 85080 177594 85089
rect 177538 85015 177594 85024
rect 177552 84778 177580 85015
rect 177540 84772 177592 84778
rect 177540 84714 177592 84720
rect 178182 83992 178238 84001
rect 178182 83927 178238 83936
rect 178196 83690 178224 83927
rect 178184 83684 178236 83690
rect 178184 83626 178236 83632
rect 177722 82904 177778 82913
rect 177722 82839 177778 82848
rect 177736 82058 177764 82839
rect 177724 82052 177776 82058
rect 177724 81994 177776 82000
rect 177354 81680 177410 81689
rect 177354 81615 177410 81624
rect 177368 80630 177396 81615
rect 178932 81417 178960 87327
rect 179484 83729 179512 88182
rect 179576 86041 179604 89134
rect 179668 88489 179696 90222
rect 179654 88480 179710 88489
rect 179654 88415 179710 88424
rect 180484 86132 180536 86138
rect 180484 86074 180536 86080
rect 179562 86032 179618 86041
rect 179562 85967 179618 85976
rect 179656 84772 179708 84778
rect 179656 84714 179708 84720
rect 179470 83720 179526 83729
rect 179470 83655 179526 83664
rect 178918 81408 178974 81417
rect 178918 81343 178974 81352
rect 177356 80624 177408 80630
rect 177356 80566 177408 80572
rect 178182 80592 178238 80601
rect 178182 80527 178238 80536
rect 178196 79270 178224 80527
rect 178826 79368 178882 79377
rect 178826 79303 178882 79312
rect 178184 79264 178236 79270
rect 178184 79206 178236 79212
rect 178274 78280 178330 78289
rect 178274 78215 178330 78224
rect 177722 77192 177778 77201
rect 177722 77127 177778 77136
rect 177170 75968 177226 75977
rect 177170 75903 177226 75912
rect 174502 72976 174558 72985
rect 174424 72934 174502 72962
rect 174502 72911 174558 72920
rect 135522 70894 135628 70922
rect 132552 68316 132604 68322
rect 132552 68258 132604 68264
rect 134484 68248 134536 68254
rect 134484 68190 134536 68196
rect 132196 67766 132532 67794
rect 131644 67630 131980 67658
rect 134496 64145 134524 68190
rect 135312 68180 135364 68186
rect 135312 68122 135364 68128
rect 135036 68112 135088 68118
rect 135036 68054 135088 68060
rect 135048 67001 135076 68054
rect 135324 67545 135352 68122
rect 135310 67536 135366 67545
rect 135310 67471 135366 67480
rect 135034 66992 135090 67001
rect 135034 66927 135090 66936
rect 134668 66752 134720 66758
rect 134668 66694 134720 66700
rect 134680 65913 134708 66694
rect 135312 66480 135364 66486
rect 135310 66448 135312 66457
rect 135364 66448 135366 66457
rect 135310 66383 135366 66392
rect 134666 65904 134722 65913
rect 134666 65839 134722 65848
rect 134668 65460 134720 65466
rect 134668 65402 134720 65408
rect 102834 64136 102890 64145
rect 102652 64100 102704 64106
rect 102834 64071 102890 64080
rect 134482 64136 134538 64145
rect 134482 64071 134538 64080
rect 102652 64042 102704 64048
rect 102558 63048 102614 63057
rect 102558 62983 102614 62992
rect 102560 62740 102612 62746
rect 102560 62682 102612 62688
rect 102466 62368 102522 62377
rect 102466 62303 102522 62312
rect 102468 61312 102520 61318
rect 100260 61254 100312 61260
rect 102374 61280 102430 61289
rect 66218 61215 66274 61224
rect 102468 61254 102520 61260
rect 102374 61215 102430 61224
rect 63734 60192 63790 60201
rect 63734 60127 63790 60136
rect 62816 60020 62868 60026
rect 62816 59962 62868 59968
rect 62722 59240 62778 59249
rect 62722 59175 62778 59184
rect 62828 58161 62856 59962
rect 66232 59958 66260 61215
rect 100626 60872 100682 60881
rect 100626 60807 100682 60816
rect 66310 60736 66366 60745
rect 66310 60671 66366 60680
rect 66324 60026 66352 60671
rect 100640 60366 100668 60807
rect 100628 60360 100680 60366
rect 100628 60302 100680 60308
rect 100902 60328 100958 60337
rect 100902 60263 100958 60272
rect 100916 60230 100944 60263
rect 100904 60224 100956 60230
rect 66402 60192 66458 60201
rect 100904 60166 100956 60172
rect 102376 60224 102428 60230
rect 102480 60201 102508 61254
rect 102572 60745 102600 62682
rect 102664 61833 102692 64042
rect 134680 63057 134708 65402
rect 135036 65392 135088 65398
rect 135036 65334 135088 65340
rect 135048 64689 135076 65334
rect 135312 65256 135364 65262
rect 135310 65224 135312 65233
rect 135364 65224 135366 65233
rect 135310 65159 135366 65168
rect 135034 64680 135090 64689
rect 135034 64615 135090 64624
rect 135404 64168 135456 64174
rect 135404 64110 135456 64116
rect 135036 64100 135088 64106
rect 135036 64042 135088 64048
rect 134666 63048 134722 63057
rect 134666 62983 134722 62992
rect 134484 62740 134536 62746
rect 134484 62682 134536 62688
rect 102650 61824 102706 61833
rect 102650 61759 102706 61768
rect 102744 61380 102796 61386
rect 102744 61322 102796 61328
rect 102558 60736 102614 60745
rect 102558 60671 102614 60680
rect 102652 60360 102704 60366
rect 102652 60302 102704 60308
rect 102376 60166 102428 60172
rect 102466 60192 102522 60201
rect 66402 60127 66404 60136
rect 66456 60127 66458 60136
rect 66404 60098 66456 60104
rect 99706 60056 99762 60065
rect 66312 60020 66364 60026
rect 99706 59991 99708 60000
rect 66312 59962 66364 59968
rect 99760 59991 99762 60000
rect 99708 59962 99760 59968
rect 63736 59952 63788 59958
rect 63736 59894 63788 59900
rect 66220 59952 66272 59958
rect 66220 59894 66272 59900
rect 63748 58705 63776 59894
rect 66310 59512 66366 59521
rect 66310 59447 66366 59456
rect 63734 58696 63790 58705
rect 62908 58660 62960 58666
rect 63734 58631 63790 58640
rect 62908 58602 62960 58608
rect 62814 58152 62870 58161
rect 62814 58087 62870 58096
rect 62630 57608 62686 57617
rect 62630 57543 62686 57552
rect 62816 57436 62868 57442
rect 62816 57378 62868 57384
rect 62724 57164 62776 57170
rect 62724 57106 62776 57112
rect 62632 57028 62684 57034
rect 62632 56970 62684 56976
rect 62644 55849 62672 56970
rect 62630 55840 62686 55849
rect 62630 55775 62686 55784
rect 62736 54761 62764 57106
rect 62828 55305 62856 57378
rect 62920 56393 62948 58602
rect 66324 58598 66352 59447
rect 100626 59104 100682 59113
rect 100626 59039 100682 59048
rect 66402 58968 66458 58977
rect 66402 58903 66458 58912
rect 66416 58666 66444 58903
rect 100640 58802 100668 59039
rect 100628 58796 100680 58802
rect 100628 58738 100680 58744
rect 100626 58696 100682 58705
rect 66404 58660 66456 58666
rect 100626 58631 100628 58640
rect 66404 58602 66456 58608
rect 100680 58631 100682 58640
rect 100628 58602 100680 58608
rect 63552 58592 63604 58598
rect 63552 58534 63604 58540
rect 66312 58592 66364 58598
rect 66312 58534 66364 58540
rect 63564 57073 63592 58534
rect 102388 58433 102416 60166
rect 102466 60127 102522 60136
rect 102560 60020 102612 60026
rect 102560 59962 102612 59968
rect 102468 58796 102520 58802
rect 102468 58738 102520 58744
rect 102374 58424 102430 58433
rect 102374 58359 102430 58368
rect 65022 58288 65078 58297
rect 65022 58223 65078 58232
rect 63550 57064 63606 57073
rect 65036 57034 65064 58223
rect 100626 57880 100682 57889
rect 100626 57815 100682 57824
rect 66402 57744 66458 57753
rect 66402 57679 66458 57688
rect 66416 57442 66444 57679
rect 100640 57442 100668 57815
rect 66404 57436 66456 57442
rect 66404 57378 66456 57384
rect 100628 57436 100680 57442
rect 100628 57378 100680 57384
rect 102376 57436 102428 57442
rect 102376 57378 102428 57384
rect 100626 57336 100682 57345
rect 100626 57271 100682 57280
rect 100640 57238 100668 57271
rect 100628 57232 100680 57238
rect 66402 57200 66458 57209
rect 66402 57135 66404 57144
rect 66456 57135 66458 57144
rect 100534 57200 100590 57209
rect 100628 57174 100680 57180
rect 100534 57135 100536 57144
rect 66404 57106 66456 57112
rect 100588 57135 100590 57144
rect 100536 57106 100588 57112
rect 63550 56999 63606 57008
rect 65024 57028 65076 57034
rect 65024 56970 65076 56976
rect 66310 56520 66366 56529
rect 66310 56455 66366 56464
rect 62906 56384 62962 56393
rect 62906 56319 62962 56328
rect 63276 55940 63328 55946
rect 63276 55882 63328 55888
rect 62814 55296 62870 55305
rect 62814 55231 62870 55240
rect 62722 54752 62778 54761
rect 62722 54687 62778 54696
rect 63288 53537 63316 55882
rect 66324 55810 66352 56455
rect 102388 56121 102416 57378
rect 102480 57345 102508 58738
rect 102572 57889 102600 59962
rect 102664 58977 102692 60302
rect 102756 59521 102784 61322
rect 134496 60745 134524 62682
rect 135048 62377 135076 64042
rect 135312 62672 135364 62678
rect 135312 62614 135364 62620
rect 135034 62368 135090 62377
rect 135034 62303 135090 62312
rect 135220 61312 135272 61318
rect 135324 61289 135352 62614
rect 135416 61833 135444 64110
rect 135600 63601 135628 70894
rect 136612 68254 136640 70908
rect 136600 68248 136652 68254
rect 136600 68190 136652 68196
rect 136874 65496 136930 65505
rect 136874 65431 136876 65440
rect 136928 65431 136930 65440
rect 136876 65402 136928 65408
rect 137716 65398 137744 70908
rect 138268 70894 138834 70922
rect 139648 70894 139938 70922
rect 138268 68202 138296 70894
rect 139648 68338 139676 70894
rect 140832 68860 140884 68866
rect 140832 68802 140884 68808
rect 138176 68174 138296 68202
rect 139556 68310 139676 68338
rect 137704 65392 137756 65398
rect 137704 65334 137756 65340
rect 138176 65262 138204 68174
rect 139556 66758 139584 68310
rect 139544 66752 139596 66758
rect 139544 66694 139596 66700
rect 140844 65740 140872 68802
rect 141028 66486 141056 70908
rect 142132 68118 142160 70908
rect 142672 68248 142724 68254
rect 142672 68190 142724 68196
rect 142120 68112 142172 68118
rect 142120 68054 142172 68060
rect 141016 66480 141068 66486
rect 141016 66422 141068 66428
rect 142684 65740 142712 68190
rect 143236 68186 143264 70908
rect 144340 68866 144368 70908
rect 144328 68860 144380 68866
rect 144328 68802 144380 68808
rect 144512 68316 144564 68322
rect 144512 68258 144564 68264
rect 143224 68180 143276 68186
rect 143224 68122 143276 68128
rect 144524 65740 144552 68258
rect 145444 68254 145472 70908
rect 146548 68322 146576 70908
rect 146536 68316 146588 68322
rect 146536 68258 146588 68264
rect 147652 68254 147680 70908
rect 148572 70894 148862 70922
rect 145432 68248 145484 68254
rect 145432 68190 145484 68196
rect 146444 68248 146496 68254
rect 146444 68190 146496 68196
rect 147640 68248 147692 68254
rect 147640 68190 147692 68196
rect 146456 65740 146484 68190
rect 148572 65754 148600 70894
rect 148310 65726 148600 65754
rect 149952 65754 149980 70908
rect 151056 68934 151084 70908
rect 151044 68928 151096 68934
rect 151044 68870 151096 68876
rect 152056 68928 152108 68934
rect 152056 68870 152108 68876
rect 149952 65726 150150 65754
rect 152068 65740 152096 68870
rect 152160 68254 152188 70908
rect 153264 68322 153292 70908
rect 153252 68316 153304 68322
rect 153252 68258 153304 68264
rect 154368 68254 154396 70908
rect 155472 68390 155500 70908
rect 155460 68384 155512 68390
rect 155460 68326 155512 68332
rect 156576 68322 156604 70908
rect 157694 70894 157984 70922
rect 155828 68316 155880 68322
rect 155828 68258 155880 68264
rect 156564 68316 156616 68322
rect 156564 68258 156616 68264
rect 152148 68248 152200 68254
rect 152148 68190 152200 68196
rect 153896 68248 153948 68254
rect 153896 68190 153948 68196
rect 154356 68248 154408 68254
rect 154356 68190 154408 68196
rect 153908 65740 153936 68190
rect 155840 65740 155868 68258
rect 157956 68254 157984 70894
rect 158784 69002 158812 70908
rect 158772 68996 158824 69002
rect 158772 68938 158824 68944
rect 159888 68934 159916 70908
rect 159876 68928 159928 68934
rect 159876 68870 159928 68876
rect 160992 68866 161020 70908
rect 160980 68860 161032 68866
rect 160980 68802 161032 68808
rect 159508 68384 159560 68390
rect 159508 68326 159560 68332
rect 157668 68248 157720 68254
rect 157668 68190 157720 68196
rect 157944 68248 157996 68254
rect 157944 68190 157996 68196
rect 157680 65740 157708 68190
rect 159520 65740 159548 68326
rect 161440 68316 161492 68322
rect 161440 68258 161492 68264
rect 163280 68316 163332 68322
rect 163280 68258 163332 68264
rect 161452 65740 161480 68258
rect 163292 65740 163320 68258
rect 164396 68254 164424 70908
rect 165120 68996 165172 69002
rect 165120 68938 165172 68944
rect 164384 68248 164436 68254
rect 164384 68190 164436 68196
rect 165132 65740 165160 68938
rect 165500 68322 165528 70908
rect 165488 68316 165540 68322
rect 165488 68258 165540 68264
rect 166604 65602 166632 70908
rect 167052 68928 167104 68934
rect 167052 68870 167104 68876
rect 167064 65740 167092 68870
rect 167708 68322 167736 70908
rect 168812 68934 168840 70908
rect 168800 68928 168852 68934
rect 168800 68870 168852 68876
rect 169916 68866 169944 70908
rect 168892 68860 168944 68866
rect 168892 68802 168944 68808
rect 169904 68860 169956 68866
rect 169904 68802 169956 68808
rect 167144 68316 167196 68322
rect 167144 68258 167196 68264
rect 167696 68316 167748 68322
rect 167696 68258 167748 68264
rect 167156 65602 167184 68258
rect 168904 65740 168932 68802
rect 171020 68322 171048 70908
rect 169536 68316 169588 68322
rect 169536 68258 169588 68264
rect 171008 68316 171060 68322
rect 171008 68258 171060 68264
rect 169260 68248 169312 68254
rect 169260 68190 169312 68196
rect 166592 65596 166644 65602
rect 166592 65538 166644 65544
rect 167144 65596 167196 65602
rect 167144 65538 167196 65544
rect 138164 65256 138216 65262
rect 138164 65198 138216 65204
rect 136874 64544 136930 64553
rect 136874 64479 136930 64488
rect 136888 64106 136916 64479
rect 136968 64168 137020 64174
rect 136966 64136 136968 64145
rect 137020 64136 137022 64145
rect 136876 64100 136928 64106
rect 136966 64071 137022 64080
rect 136876 64042 136928 64048
rect 169272 64038 169300 68190
rect 169548 65233 169576 68258
rect 172124 68254 172152 70908
rect 173228 68662 173256 70908
rect 173860 68928 173912 68934
rect 173860 68870 173912 68876
rect 173216 68656 173268 68662
rect 173216 68598 173268 68604
rect 172112 68248 172164 68254
rect 172112 68190 172164 68196
rect 173872 65913 173900 68870
rect 173952 68860 174004 68866
rect 173952 68802 174004 68808
rect 173964 66457 173992 68802
rect 174332 68730 174360 70908
rect 174320 68724 174372 68730
rect 174320 68666 174372 68672
rect 174044 68316 174096 68322
rect 174044 68258 174096 68264
rect 174056 67001 174084 68258
rect 174688 68180 174740 68186
rect 174688 68122 174740 68128
rect 174700 67545 174728 68122
rect 177184 67780 177212 75903
rect 177354 73656 177410 73665
rect 177354 73591 177410 73600
rect 177368 72402 177396 73591
rect 177356 72396 177408 72402
rect 177356 72338 177408 72344
rect 177736 67780 177764 77127
rect 178288 67780 178316 78215
rect 178366 74880 178422 74889
rect 178366 74815 178422 74824
rect 178380 70906 178408 74815
rect 178368 70900 178420 70906
rect 178368 70842 178420 70848
rect 178840 67780 178868 79303
rect 179380 79264 179432 79270
rect 179380 79206 179432 79212
rect 179392 67780 179420 79206
rect 179668 76657 179696 84714
rect 180392 83684 180444 83690
rect 180392 83626 180444 83632
rect 180300 82052 180352 82058
rect 180300 81994 180352 82000
rect 180024 80624 180076 80630
rect 180024 80566 180076 80572
rect 179654 76648 179710 76657
rect 179654 76583 179710 76592
rect 180036 67780 180064 80566
rect 180312 72033 180340 81994
rect 180404 74345 180432 83626
rect 180496 78969 180524 86074
rect 180482 78960 180538 78969
rect 180482 78895 180538 78904
rect 180390 74336 180446 74345
rect 180390 74271 180446 74280
rect 180576 72396 180628 72402
rect 180576 72338 180628 72344
rect 180298 72024 180354 72033
rect 180298 71959 180354 71968
rect 180588 67780 180616 72338
rect 181128 70900 181180 70906
rect 181128 70842 181180 70848
rect 182796 70894 183132 70922
rect 183256 70894 183500 70922
rect 183624 70894 183868 70922
rect 183992 70894 184328 70922
rect 184452 70894 184696 70922
rect 184820 70894 185064 70922
rect 185188 70894 185524 70922
rect 185740 70894 185892 70922
rect 181140 67780 181168 70842
rect 182232 69200 182284 69206
rect 182232 69142 182284 69148
rect 181680 69132 181732 69138
rect 181680 69074 181732 69080
rect 181692 67780 181720 69074
rect 182244 67780 182272 69142
rect 182796 69138 182824 70894
rect 183256 69206 183284 70894
rect 183244 69200 183296 69206
rect 183244 69142 183296 69148
rect 182784 69132 182836 69138
rect 182784 69074 182836 69080
rect 183624 68458 183652 70894
rect 182876 68452 182928 68458
rect 182876 68394 182928 68400
rect 183612 68452 183664 68458
rect 183612 68394 183664 68400
rect 182888 67780 182916 68394
rect 183992 68338 184020 70894
rect 183716 68310 184020 68338
rect 183716 67794 183744 68310
rect 184452 67794 184480 70894
rect 184820 67794 184848 70894
rect 185188 69154 185216 70894
rect 183454 67766 183744 67794
rect 184006 67766 184480 67794
rect 184558 67766 184848 67794
rect 185096 69126 185216 69154
rect 185096 67780 185124 69126
rect 185740 67780 185768 70894
rect 186246 70650 186274 70908
rect 186720 70894 186872 70922
rect 187088 70894 187240 70922
rect 187456 70894 187792 70922
rect 187916 70894 188160 70922
rect 188284 70894 188528 70922
rect 188652 70894 188988 70922
rect 189112 70894 189356 70922
rect 189480 70894 189724 70922
rect 189848 70894 190184 70922
rect 190308 70894 190460 70922
rect 186246 70622 186320 70650
rect 186292 67780 186320 70622
rect 186844 67780 186872 70894
rect 187212 67794 187240 70894
rect 187764 69154 187792 70894
rect 187764 69126 187976 69154
rect 187212 67766 187410 67794
rect 187948 67780 187976 69126
rect 188132 67794 188160 70894
rect 188500 67930 188528 70894
rect 188960 68338 188988 70894
rect 189328 69177 189356 70894
rect 189314 69168 189370 69177
rect 189696 69138 189724 70894
rect 189314 69103 189370 69112
rect 189684 69132 189736 69138
rect 189684 69074 189736 69080
rect 190156 69041 190184 70894
rect 190432 69177 190460 70894
rect 190616 70894 190676 70922
rect 191136 70894 191380 70922
rect 191504 70894 191748 70922
rect 190234 69168 190290 69177
rect 190234 69103 190290 69112
rect 190418 69168 190474 69177
rect 190418 69103 190474 69112
rect 190142 69032 190198 69041
rect 190142 68967 190198 68976
rect 188960 68310 189356 68338
rect 188500 67902 188804 67930
rect 188776 67794 188804 67902
rect 189328 67794 189356 68310
rect 188132 67766 188606 67794
rect 188776 67766 189158 67794
rect 189328 67766 189710 67794
rect 190248 67780 190276 69103
rect 190616 68934 190644 70894
rect 191352 69313 191380 70894
rect 191338 69304 191394 69313
rect 191338 69239 191394 69248
rect 190696 69132 190748 69138
rect 190696 69074 190748 69080
rect 190604 68928 190656 68934
rect 190604 68870 190656 68876
rect 190708 67794 190736 69074
rect 191430 69032 191486 69041
rect 191430 68967 191486 68976
rect 190708 67766 190814 67794
rect 191444 67780 191472 68967
rect 191720 68594 191748 70894
rect 191812 70894 191872 70922
rect 192332 70894 192576 70922
rect 192700 70894 192944 70922
rect 193068 70894 193404 70922
rect 193528 70894 193772 70922
rect 193896 70894 194140 70922
rect 194264 70894 194600 70922
rect 191812 69138 191840 70894
rect 192548 69206 192576 70894
rect 192536 69200 192588 69206
rect 191982 69168 192038 69177
rect 191800 69132 191852 69138
rect 192536 69142 192588 69148
rect 191982 69103 192038 69112
rect 191800 69074 191852 69080
rect 191708 68588 191760 68594
rect 191708 68530 191760 68536
rect 191996 67780 192024 69103
rect 192916 69070 192944 70894
rect 193086 69304 193142 69313
rect 193086 69239 193142 69248
rect 192904 69064 192956 69070
rect 192904 69006 192956 69012
rect 192536 68928 192588 68934
rect 192536 68870 192588 68876
rect 192548 67780 192576 68870
rect 193100 67780 193128 69239
rect 193376 69002 193404 70894
rect 193364 68996 193416 69002
rect 193364 68938 193416 68944
rect 193744 68866 193772 70894
rect 194112 69274 194140 70894
rect 194100 69268 194152 69274
rect 194100 69210 194152 69216
rect 194572 69138 194600 70894
rect 194664 70894 194724 70922
rect 195092 70894 195336 70922
rect 195460 70894 195796 70922
rect 195920 70894 196164 70922
rect 196288 70894 196532 70922
rect 196656 70894 196992 70922
rect 197116 70894 197360 70922
rect 194284 69132 194336 69138
rect 194284 69074 194336 69080
rect 194560 69132 194612 69138
rect 194560 69074 194612 69080
rect 193732 68860 193784 68866
rect 193732 68802 193784 68808
rect 193640 68588 193692 68594
rect 193640 68530 193692 68536
rect 193652 67780 193680 68530
rect 194296 67780 194324 69074
rect 194664 68662 194692 70894
rect 194836 69200 194888 69206
rect 194836 69142 194888 69148
rect 194652 68656 194704 68662
rect 194652 68598 194704 68604
rect 194848 67780 194876 69142
rect 195308 68798 195336 70894
rect 195388 69064 195440 69070
rect 195388 69006 195440 69012
rect 195296 68792 195348 68798
rect 195296 68734 195348 68740
rect 195400 67780 195428 69006
rect 195768 68934 195796 70894
rect 196136 69410 196164 70894
rect 196124 69404 196176 69410
rect 196124 69346 196176 69352
rect 196504 69002 196532 70894
rect 196964 69070 196992 70894
rect 197332 69274 197360 70894
rect 197424 70894 197484 70922
rect 197852 70894 198188 70922
rect 198312 70894 198556 70922
rect 198680 70894 198924 70922
rect 197136 69268 197188 69274
rect 197136 69210 197188 69216
rect 197320 69268 197372 69274
rect 197320 69210 197372 69216
rect 196952 69064 197004 69070
rect 196952 69006 197004 69012
rect 195940 68996 195992 69002
rect 195940 68938 195992 68944
rect 196492 68996 196544 69002
rect 196492 68938 196544 68944
rect 195756 68928 195808 68934
rect 195756 68870 195808 68876
rect 195952 67780 195980 68938
rect 196492 68860 196544 68866
rect 196492 68802 196544 68808
rect 196504 67780 196532 68802
rect 197148 67780 197176 69210
rect 197424 69206 197452 70894
rect 197412 69200 197464 69206
rect 197412 69142 197464 69148
rect 198160 69138 198188 70894
rect 198528 69478 198556 70894
rect 198896 69546 198924 70894
rect 198884 69540 198936 69546
rect 198884 69482 198936 69488
rect 198516 69472 198568 69478
rect 198516 69414 198568 69420
rect 199988 69404 200040 69410
rect 199988 69346 200040 69352
rect 197688 69132 197740 69138
rect 197688 69074 197740 69080
rect 198148 69132 198200 69138
rect 198148 69074 198200 69080
rect 197700 67780 197728 69074
rect 199344 68928 199396 68934
rect 199344 68870 199396 68876
rect 198792 68792 198844 68798
rect 198792 68734 198844 68740
rect 198240 68656 198292 68662
rect 198240 68598 198292 68604
rect 198252 67780 198280 68598
rect 198804 67780 198832 68734
rect 199356 67780 199384 68870
rect 200000 67780 200028 69346
rect 201012 69342 201040 90319
rect 204494 77600 204550 77609
rect 204494 77535 204550 77544
rect 201090 77056 201146 77065
rect 201090 76991 201146 77000
rect 201104 69449 201132 76991
rect 203944 69608 203996 69614
rect 203944 69550 203996 69556
rect 202196 69540 202248 69546
rect 202196 69482 202248 69488
rect 202208 69449 202236 69482
rect 202932 69472 202984 69478
rect 201090 69440 201146 69449
rect 201090 69375 201146 69384
rect 202194 69440 202250 69449
rect 202932 69414 202984 69420
rect 202194 69375 202250 69384
rect 201000 69336 201052 69342
rect 201000 69278 201052 69284
rect 202944 69290 202972 69414
rect 201644 69268 201696 69274
rect 202944 69262 203156 69290
rect 201644 69210 201696 69216
rect 201092 69064 201144 69070
rect 201092 69006 201144 69012
rect 200540 68996 200592 69002
rect 200540 68938 200592 68944
rect 200552 67780 200580 68938
rect 201104 67780 201132 69006
rect 201656 67780 201684 69210
rect 201828 69200 201880 69206
rect 201828 69142 201880 69148
rect 201840 67794 201868 69142
rect 202840 69132 202892 69138
rect 202840 69074 202892 69080
rect 201840 67766 202222 67794
rect 202852 67780 202880 69074
rect 203128 67794 203156 69262
rect 203128 67766 203418 67794
rect 203956 67780 203984 69550
rect 204508 67780 204536 77535
rect 210580 69478 210608 70908
rect 210568 69472 210620 69478
rect 210568 69414 210620 69420
rect 215916 69342 215944 70908
rect 215904 69336 215956 69342
rect 215904 69278 215956 69284
rect 221252 68866 221280 70908
rect 205140 68860 205192 68866
rect 205140 68802 205192 68808
rect 221240 68860 221292 68866
rect 221240 68802 221292 68808
rect 174686 67536 174742 67545
rect 174686 67471 174742 67480
rect 174042 66992 174098 67001
rect 174042 66927 174098 66936
rect 173950 66448 174006 66457
rect 173950 66383 174006 66392
rect 173858 65904 173914 65913
rect 173858 65839 173914 65848
rect 171834 65632 171890 65641
rect 171834 65567 171890 65576
rect 169534 65224 169590 65233
rect 169534 65159 169590 65168
rect 171650 64408 171706 64417
rect 171650 64343 171706 64352
rect 169260 64032 169312 64038
rect 169260 63974 169312 63980
rect 135586 63592 135642 63601
rect 135586 63527 135642 63536
rect 136874 63320 136930 63329
rect 136874 63255 136930 63264
rect 136888 62678 136916 63255
rect 136966 62776 137022 62785
rect 136966 62711 136968 62720
rect 137020 62711 137022 62720
rect 136968 62682 137020 62688
rect 136876 62672 136928 62678
rect 136876 62614 136928 62620
rect 171664 62610 171692 64343
rect 171742 64136 171798 64145
rect 171742 64071 171798 64080
rect 171652 62604 171704 62610
rect 171652 62546 171704 62552
rect 171756 62542 171784 64071
rect 171848 63766 171876 65567
rect 174228 65392 174280 65398
rect 174228 65334 174280 65340
rect 174136 65324 174188 65330
rect 174136 65266 174188 65272
rect 174148 64689 174176 65266
rect 174134 64680 174190 64689
rect 174134 64615 174190 64624
rect 174240 64145 174268 65334
rect 174226 64136 174282 64145
rect 174226 64071 174282 64080
rect 174136 64032 174188 64038
rect 174136 63974 174188 63980
rect 171836 63760 171888 63766
rect 171836 63702 171888 63708
rect 174148 63601 174176 63974
rect 174228 63760 174280 63766
rect 174228 63702 174280 63708
rect 174134 63592 174190 63601
rect 174134 63527 174190 63536
rect 172018 63456 172074 63465
rect 172018 63391 172074 63400
rect 172032 63290 172060 63391
rect 172020 63284 172072 63290
rect 172020 63226 172072 63232
rect 173860 63284 173912 63290
rect 173860 63226 173912 63232
rect 172662 62776 172718 62785
rect 172718 62734 172796 62762
rect 172662 62711 172718 62720
rect 171744 62536 171796 62542
rect 171744 62478 171796 62484
rect 136782 62096 136838 62105
rect 136782 62031 136838 62040
rect 171650 62096 171706 62105
rect 171650 62031 171652 62040
rect 135402 61824 135458 61833
rect 135402 61759 135458 61768
rect 135220 61254 135272 61260
rect 135310 61280 135366 61289
rect 134852 60972 134904 60978
rect 134852 60914 134904 60920
rect 134482 60736 134538 60745
rect 134482 60671 134538 60680
rect 134864 60201 134892 60914
rect 134850 60192 134906 60201
rect 134850 60127 134906 60136
rect 134484 60088 134536 60094
rect 134484 60030 134536 60036
rect 134392 59884 134444 59890
rect 134392 59826 134444 59832
rect 102742 59512 102798 59521
rect 102742 59447 102798 59456
rect 134404 58977 134432 59826
rect 102650 58968 102706 58977
rect 102650 58903 102706 58912
rect 134390 58968 134446 58977
rect 134390 58903 134446 58912
rect 102652 58660 102704 58666
rect 102652 58602 102704 58608
rect 102558 57880 102614 57889
rect 102558 57815 102614 57824
rect 102466 57336 102522 57345
rect 102466 57271 102522 57280
rect 102468 57232 102520 57238
rect 102468 57174 102520 57180
rect 100626 56112 100682 56121
rect 100626 56047 100682 56056
rect 102374 56112 102430 56121
rect 102374 56047 102430 56056
rect 66402 55976 66458 55985
rect 100640 55946 100668 56047
rect 66402 55911 66404 55920
rect 66456 55911 66458 55920
rect 100628 55940 100680 55946
rect 66404 55882 66456 55888
rect 100628 55882 100680 55888
rect 102376 55940 102428 55946
rect 102376 55882 102428 55888
rect 100902 55840 100958 55849
rect 63552 55804 63604 55810
rect 63552 55746 63604 55752
rect 66312 55804 66364 55810
rect 100902 55775 100904 55784
rect 66312 55746 66364 55752
rect 100956 55775 100958 55784
rect 100904 55746 100956 55752
rect 63368 54716 63420 54722
rect 63368 54658 63420 54664
rect 30522 53528 30578 53537
rect 30522 53463 30578 53472
rect 63274 53528 63330 53537
rect 63274 53463 63330 53472
rect 30536 33642 30564 53463
rect 62816 53356 62868 53362
rect 62816 53298 62868 53304
rect 62724 51724 62776 51730
rect 62724 51666 62776 51672
rect 62736 49593 62764 51666
rect 62828 51361 62856 53298
rect 63380 52449 63408 54658
rect 63460 54444 63512 54450
rect 63460 54386 63512 54392
rect 63472 52993 63500 54386
rect 63564 54217 63592 55746
rect 66310 55296 66366 55305
rect 66310 55231 66366 55240
rect 66324 54450 66352 55231
rect 100626 54888 100682 54897
rect 100626 54823 100628 54832
rect 100680 54823 100682 54832
rect 100628 54794 100680 54800
rect 66402 54752 66458 54761
rect 66402 54687 66404 54696
rect 66456 54687 66458 54696
rect 66404 54658 66456 54664
rect 100810 54616 100866 54625
rect 100810 54551 100812 54560
rect 100864 54551 100866 54560
rect 100812 54522 100864 54528
rect 102388 54489 102416 55882
rect 102480 55577 102508 57174
rect 102560 57164 102612 57170
rect 102560 57106 102612 57112
rect 102466 55568 102522 55577
rect 102466 55503 102522 55512
rect 102572 55033 102600 57106
rect 102664 56665 102692 58602
rect 134496 58433 134524 60030
rect 135232 59521 135260 61254
rect 135310 61215 135366 61224
rect 136796 60978 136824 62031
rect 171704 62031 171706 62040
rect 171652 62002 171704 62008
rect 136874 61416 136930 61425
rect 136874 61351 136930 61360
rect 172662 61416 172718 61425
rect 172662 61351 172664 61360
rect 136888 61318 136916 61351
rect 172716 61351 172718 61360
rect 172664 61322 172716 61328
rect 136876 61312 136928 61318
rect 136876 61254 136928 61260
rect 172768 61250 172796 62734
rect 173872 61289 173900 63226
rect 174240 63057 174268 63702
rect 174226 63048 174282 63057
rect 174226 62983 174282 62992
rect 174320 62604 174372 62610
rect 174320 62546 174372 62552
rect 174136 62536 174188 62542
rect 174136 62478 174188 62484
rect 174044 62060 174096 62066
rect 174044 62002 174096 62008
rect 173952 61380 174004 61386
rect 173952 61322 174004 61328
rect 173858 61280 173914 61289
rect 172756 61244 172808 61250
rect 173858 61215 173914 61224
rect 172756 61186 172808 61192
rect 136784 60972 136836 60978
rect 136784 60914 136836 60920
rect 136782 60872 136838 60881
rect 136782 60807 136838 60816
rect 172202 60872 172258 60881
rect 172202 60807 172258 60816
rect 135404 59952 135456 59958
rect 135404 59894 135456 59900
rect 135218 59512 135274 59521
rect 135218 59447 135274 59456
rect 135220 58592 135272 58598
rect 135220 58534 135272 58540
rect 135036 58456 135088 58462
rect 134482 58424 134538 58433
rect 135036 58398 135088 58404
rect 134482 58359 134538 58368
rect 135048 57345 135076 58398
rect 135034 57336 135090 57345
rect 135034 57271 135090 57280
rect 134576 57096 134628 57102
rect 134576 57038 134628 57044
rect 102650 56656 102706 56665
rect 102650 56591 102706 56600
rect 134588 56121 134616 57038
rect 135232 56665 135260 58534
rect 135416 57889 135444 59894
rect 136796 59890 136824 60807
rect 136966 60328 137022 60337
rect 136966 60263 137022 60272
rect 136980 60094 137008 60263
rect 136968 60088 137020 60094
rect 136874 60056 136930 60065
rect 136968 60030 137020 60036
rect 136874 59991 136930 60000
rect 136888 59958 136916 59991
rect 172216 59958 172244 60807
rect 172662 60328 172718 60337
rect 172718 60286 172796 60314
rect 172662 60263 172718 60272
rect 172664 60020 172716 60026
rect 172664 59962 172716 59968
rect 136876 59952 136928 59958
rect 136876 59894 136928 59900
rect 172204 59952 172256 59958
rect 172676 59929 172704 59962
rect 172204 59894 172256 59900
rect 172662 59920 172718 59929
rect 136784 59884 136836 59890
rect 172662 59855 172718 59864
rect 136784 59826 136836 59832
rect 136782 59104 136838 59113
rect 136782 59039 136838 59048
rect 172662 59104 172718 59113
rect 172662 59039 172718 59048
rect 136796 58462 136824 59039
rect 172676 58870 172704 59039
rect 172664 58864 172716 58870
rect 172664 58806 172716 58812
rect 136874 58696 136930 58705
rect 136874 58631 136930 58640
rect 172662 58696 172718 58705
rect 172662 58631 172664 58640
rect 136888 58598 136916 58631
rect 172716 58631 172718 58640
rect 172664 58602 172716 58608
rect 136876 58592 136928 58598
rect 136876 58534 136928 58540
rect 172768 58530 172796 60286
rect 173768 60020 173820 60026
rect 173768 59962 173820 59968
rect 172756 58524 172808 58530
rect 172756 58466 172808 58472
rect 136784 58456 136836 58462
rect 136784 58398 136836 58404
rect 173780 57889 173808 59962
rect 173964 59521 173992 61322
rect 174056 60201 174084 62002
rect 174148 61833 174176 62478
rect 174332 62377 174360 62546
rect 174318 62368 174374 62377
rect 174318 62303 174374 62312
rect 174134 61824 174190 61833
rect 174134 61759 174190 61768
rect 174136 61244 174188 61250
rect 174136 61186 174188 61192
rect 174148 60745 174176 61186
rect 174134 60736 174190 60745
rect 174134 60671 174190 60680
rect 174042 60192 174098 60201
rect 174042 60127 174098 60136
rect 174044 59952 174096 59958
rect 174044 59894 174096 59900
rect 173950 59512 174006 59521
rect 173950 59447 174006 59456
rect 174056 58977 174084 59894
rect 174042 58968 174098 58977
rect 174042 58903 174098 58912
rect 174044 58864 174096 58870
rect 174044 58806 174096 58812
rect 173860 58660 173912 58666
rect 173860 58602 173912 58608
rect 135402 57880 135458 57889
rect 135402 57815 135458 57824
rect 136782 57880 136838 57889
rect 136782 57815 136838 57824
rect 172110 57880 172166 57889
rect 172110 57815 172166 57824
rect 173766 57880 173822 57889
rect 173766 57815 173822 57824
rect 135404 57232 135456 57238
rect 135404 57174 135456 57180
rect 135312 57164 135364 57170
rect 135312 57106 135364 57112
rect 135218 56656 135274 56665
rect 135218 56591 135274 56600
rect 134574 56112 134630 56121
rect 134574 56047 134630 56056
rect 102652 55804 102704 55810
rect 102652 55746 102704 55752
rect 134300 55804 134352 55810
rect 134300 55746 134352 55752
rect 102558 55024 102614 55033
rect 102558 54959 102614 54968
rect 102468 54852 102520 54858
rect 102468 54794 102520 54800
rect 102374 54480 102430 54489
rect 66312 54444 66364 54450
rect 102374 54415 102430 54424
rect 66312 54386 66364 54392
rect 63550 54208 63606 54217
rect 63550 54143 63606 54152
rect 66310 54208 66366 54217
rect 66310 54143 66366 54152
rect 66324 53022 66352 54143
rect 100626 53664 100682 53673
rect 100626 53599 100682 53608
rect 66402 53528 66458 53537
rect 66402 53463 66458 53472
rect 66416 53362 66444 53463
rect 66404 53356 66456 53362
rect 66404 53298 66456 53304
rect 100640 53294 100668 53599
rect 100628 53288 100680 53294
rect 102480 53265 102508 54794
rect 102560 54580 102612 54586
rect 102560 54522 102612 54528
rect 100628 53230 100680 53236
rect 102466 53256 102522 53265
rect 102466 53191 102522 53200
rect 100626 53120 100682 53129
rect 100626 53055 100628 53064
rect 100680 53055 100682 53064
rect 102376 53084 102428 53090
rect 100628 53026 100680 53032
rect 102376 53026 102428 53032
rect 63736 53016 63788 53022
rect 63458 52984 63514 52993
rect 66312 53016 66364 53022
rect 63736 52958 63788 52964
rect 65666 52984 65722 52993
rect 63458 52919 63514 52928
rect 63366 52440 63422 52449
rect 63366 52375 63422 52384
rect 62908 52132 62960 52138
rect 62908 52074 62960 52080
rect 62814 51352 62870 51361
rect 62814 51287 62870 51296
rect 62816 50500 62868 50506
rect 62816 50442 62868 50448
rect 62722 49584 62778 49593
rect 62722 49519 62778 49528
rect 62828 48505 62856 50442
rect 62920 50137 62948 52074
rect 63748 51905 63776 52958
rect 66312 52958 66364 52964
rect 65666 52919 65722 52928
rect 63734 51896 63790 51905
rect 63734 51831 63790 51840
rect 65680 51662 65708 52919
rect 100626 52440 100682 52449
rect 100626 52375 100682 52384
rect 66402 52304 66458 52313
rect 100640 52274 100668 52375
rect 66402 52239 66458 52248
rect 100628 52268 100680 52274
rect 66416 52138 66444 52239
rect 100628 52210 100680 52216
rect 66404 52132 66456 52138
rect 66404 52074 66456 52080
rect 100626 51896 100682 51905
rect 100626 51831 100682 51840
rect 66402 51760 66458 51769
rect 66402 51695 66404 51704
rect 66456 51695 66458 51704
rect 100534 51760 100590 51769
rect 100640 51730 100668 51831
rect 100534 51695 100590 51704
rect 100628 51724 100680 51730
rect 66404 51666 66456 51672
rect 100548 51662 100576 51695
rect 100628 51666 100680 51672
rect 63736 51656 63788 51662
rect 63736 51598 63788 51604
rect 65668 51656 65720 51662
rect 65668 51598 65720 51604
rect 100536 51656 100588 51662
rect 102388 51633 102416 53026
rect 102572 52721 102600 54522
rect 102664 53809 102692 55746
rect 134208 54580 134260 54586
rect 134208 54522 134260 54528
rect 102650 53800 102706 53809
rect 102650 53735 102706 53744
rect 102744 53288 102796 53294
rect 102744 53230 102796 53236
rect 102558 52712 102614 52721
rect 102558 52647 102614 52656
rect 102652 52268 102704 52274
rect 102652 52210 102704 52216
rect 102468 51724 102520 51730
rect 102468 51666 102520 51672
rect 100536 51598 100588 51604
rect 102374 51624 102430 51633
rect 63748 50681 63776 51598
rect 102374 51559 102430 51568
rect 66402 51216 66458 51225
rect 66402 51151 66458 51160
rect 63734 50672 63790 50681
rect 66416 50642 66444 51151
rect 100626 50672 100682 50681
rect 63734 50607 63790 50616
rect 63828 50636 63880 50642
rect 63828 50578 63880 50584
rect 66404 50636 66456 50642
rect 100626 50607 100682 50616
rect 66404 50578 66456 50584
rect 62906 50128 62962 50137
rect 62906 50063 62962 50072
rect 63840 49049 63868 50578
rect 66402 50536 66458 50545
rect 100640 50506 100668 50607
rect 66402 50471 66404 50480
rect 66456 50471 66458 50480
rect 100628 50500 100680 50506
rect 66404 50442 66456 50448
rect 100628 50442 100680 50448
rect 102480 50409 102508 51666
rect 102560 51656 102612 51662
rect 102560 51598 102612 51604
rect 100626 50400 100682 50409
rect 102466 50400 102522 50409
rect 100626 50335 100628 50344
rect 100680 50335 100682 50344
rect 102376 50364 102428 50370
rect 100628 50306 100680 50312
rect 102466 50335 102522 50344
rect 102376 50306 102428 50312
rect 65482 49992 65538 50001
rect 65482 49927 65538 49936
rect 63826 49040 63882 49049
rect 63736 49004 63788 49010
rect 65496 49010 65524 49927
rect 100626 49448 100682 49457
rect 100626 49383 100682 49392
rect 66402 49312 66458 49321
rect 100640 49282 100668 49383
rect 66402 49247 66458 49256
rect 100628 49276 100680 49282
rect 63826 48975 63882 48984
rect 65484 49004 65536 49010
rect 63736 48946 63788 48952
rect 65484 48946 65536 48952
rect 62908 48936 62960 48942
rect 62908 48878 62960 48884
rect 62814 48496 62870 48505
rect 62814 48431 62870 48440
rect 62816 47508 62868 47514
rect 62816 47450 62868 47456
rect 62724 47236 62776 47242
rect 62724 47178 62776 47184
rect 62736 46737 62764 47178
rect 62722 46728 62778 46737
rect 62722 46663 62778 46672
rect 62828 45649 62856 47450
rect 62920 47281 62948 48878
rect 63748 47825 63776 48946
rect 66416 48942 66444 49247
rect 100628 49218 100680 49224
rect 100626 49040 100682 49049
rect 100626 48975 100628 48984
rect 100680 48975 100682 48984
rect 100628 48946 100680 48952
rect 66404 48936 66456 48942
rect 66404 48878 66456 48884
rect 102388 48777 102416 50306
rect 102572 49865 102600 51598
rect 102664 50953 102692 52210
rect 102756 52177 102784 53230
rect 134220 52721 134248 54522
rect 134312 53809 134340 55746
rect 135324 55577 135352 57106
rect 135310 55568 135366 55577
rect 135310 55503 135366 55512
rect 135036 55464 135088 55470
rect 135036 55406 135088 55412
rect 135048 54489 135076 55406
rect 135416 55033 135444 57174
rect 136796 57102 136824 57815
rect 136874 57336 136930 57345
rect 136874 57271 136930 57280
rect 136888 57170 136916 57271
rect 136968 57232 137020 57238
rect 136966 57200 136968 57209
rect 137020 57200 137022 57209
rect 136876 57164 136928 57170
rect 172124 57170 172152 57815
rect 172662 57472 172718 57481
rect 172662 57407 172718 57416
rect 172570 57336 172626 57345
rect 172676 57306 172704 57407
rect 172570 57271 172626 57280
rect 172664 57300 172716 57306
rect 172584 57238 172612 57271
rect 172664 57242 172716 57248
rect 172572 57232 172624 57238
rect 172572 57174 172624 57180
rect 173768 57232 173820 57238
rect 173768 57174 173820 57180
rect 136966 57135 137022 57144
rect 172112 57164 172164 57170
rect 136876 57106 136928 57112
rect 172112 57106 172164 57112
rect 136784 57096 136836 57102
rect 136784 57038 136836 57044
rect 136782 56112 136838 56121
rect 136782 56047 136838 56056
rect 172662 56112 172718 56121
rect 172662 56047 172664 56056
rect 136796 55470 136824 56047
rect 172716 56047 172718 56056
rect 172664 56018 172716 56024
rect 136874 55840 136930 55849
rect 136874 55775 136876 55784
rect 136928 55775 136930 55784
rect 172662 55840 172718 55849
rect 172718 55798 172980 55826
rect 172662 55775 172718 55784
rect 136876 55746 136928 55752
rect 136784 55464 136836 55470
rect 136784 55406 136836 55412
rect 135402 55024 135458 55033
rect 135402 54959 135458 54968
rect 136782 54888 136838 54897
rect 136782 54823 136838 54832
rect 171742 54888 171798 54897
rect 171742 54823 171798 54832
rect 135034 54480 135090 54489
rect 135034 54415 135090 54424
rect 136796 53974 136824 54823
rect 137150 54616 137206 54625
rect 137150 54551 137152 54560
rect 137204 54551 137206 54560
rect 137152 54522 137204 54528
rect 171756 54450 171784 54823
rect 172846 54480 172902 54489
rect 171744 54444 171796 54450
rect 172846 54415 172902 54424
rect 171744 54386 171796 54392
rect 135128 53968 135180 53974
rect 135128 53910 135180 53916
rect 136784 53968 136836 53974
rect 136784 53910 136836 53916
rect 134298 53800 134354 53809
rect 134298 53735 134354 53744
rect 135140 53265 135168 53910
rect 136782 53664 136838 53673
rect 136782 53599 136838 53608
rect 172570 53664 172626 53673
rect 172570 53599 172626 53608
rect 135126 53256 135182 53265
rect 135126 53191 135182 53200
rect 135404 53016 135456 53022
rect 135404 52958 135456 52964
rect 135036 52880 135088 52886
rect 135036 52822 135088 52828
rect 134206 52712 134262 52721
rect 134206 52647 134262 52656
rect 135048 52177 135076 52822
rect 102742 52168 102798 52177
rect 102742 52103 102798 52112
rect 135034 52168 135090 52177
rect 135034 52103 135090 52112
rect 135312 51656 135364 51662
rect 135416 51633 135444 52958
rect 136796 52886 136824 53599
rect 172584 53226 172612 53599
rect 172572 53220 172624 53226
rect 172572 53162 172624 53168
rect 136874 53120 136930 53129
rect 136874 53055 136930 53064
rect 172662 53120 172718 53129
rect 172662 53055 172664 53064
rect 136888 53022 136916 53055
rect 172716 53055 172718 53064
rect 172664 53026 172716 53032
rect 136876 53016 136928 53022
rect 136876 52958 136928 52964
rect 172860 52954 172888 54415
rect 172952 54110 172980 55798
rect 173780 55033 173808 57174
rect 173872 56665 173900 58602
rect 174056 57345 174084 58806
rect 174136 58524 174188 58530
rect 174136 58466 174188 58472
rect 174148 58433 174176 58466
rect 174134 58424 174190 58433
rect 174134 58359 174190 58368
rect 174042 57336 174098 57345
rect 173952 57300 174004 57306
rect 174042 57271 174098 57280
rect 173952 57242 174004 57248
rect 173858 56656 173914 56665
rect 173858 56591 173914 56600
rect 173964 55577 173992 57242
rect 174044 57164 174096 57170
rect 174044 57106 174096 57112
rect 174056 56393 174084 57106
rect 174042 56384 174098 56393
rect 174042 56319 174098 56328
rect 174044 56076 174096 56082
rect 174044 56018 174096 56024
rect 173950 55568 174006 55577
rect 173950 55503 174006 55512
rect 173766 55024 173822 55033
rect 173766 54959 173822 54968
rect 174056 54489 174084 56018
rect 174042 54480 174098 54489
rect 174042 54415 174098 54424
rect 174228 54376 174280 54382
rect 174228 54318 174280 54324
rect 172940 54104 172992 54110
rect 172940 54046 172992 54052
rect 174136 54104 174188 54110
rect 174136 54046 174188 54052
rect 174148 53809 174176 54046
rect 174134 53800 174190 53809
rect 174134 53735 174190 53744
rect 174240 53265 174268 54318
rect 174226 53256 174282 53265
rect 174044 53220 174096 53226
rect 174226 53191 174282 53200
rect 174044 53162 174096 53168
rect 173860 53084 173912 53090
rect 173860 53026 173912 53032
rect 172848 52948 172900 52954
rect 172848 52890 172900 52896
rect 136784 52880 136836 52886
rect 136784 52822 136836 52828
rect 136690 52440 136746 52449
rect 136690 52375 136746 52384
rect 172018 52440 172074 52449
rect 172018 52375 172074 52384
rect 135312 51598 135364 51604
rect 135402 51624 135458 51633
rect 135036 51384 135088 51390
rect 135036 51326 135088 51332
rect 102650 50944 102706 50953
rect 102650 50879 102706 50888
rect 102652 50500 102704 50506
rect 102652 50442 102704 50448
rect 102558 49856 102614 49865
rect 102558 49791 102614 49800
rect 102664 49321 102692 50442
rect 135048 50409 135076 51326
rect 135034 50400 135090 50409
rect 135034 50335 135090 50344
rect 134852 50228 134904 50234
rect 134852 50170 134904 50176
rect 134864 49321 134892 50170
rect 135324 49865 135352 51598
rect 135402 51559 135458 51568
rect 136704 51118 136732 52375
rect 136782 51896 136838 51905
rect 136782 51831 136838 51840
rect 136796 51390 136824 51831
rect 136874 51760 136930 51769
rect 136874 51695 136930 51704
rect 136888 51662 136916 51695
rect 172032 51662 172060 52375
rect 172662 51896 172718 51905
rect 172662 51831 172664 51840
rect 172716 51831 172718 51840
rect 172664 51802 172716 51808
rect 172662 51760 172718 51769
rect 172662 51695 172664 51704
rect 172716 51695 172718 51704
rect 173768 51724 173820 51730
rect 172664 51666 172716 51672
rect 173768 51666 173820 51672
rect 136876 51656 136928 51662
rect 136876 51598 136928 51604
rect 172020 51656 172072 51662
rect 172020 51598 172072 51604
rect 136784 51384 136836 51390
rect 136784 51326 136836 51332
rect 135404 51112 135456 51118
rect 135404 51054 135456 51060
rect 136692 51112 136744 51118
rect 136692 51054 136744 51060
rect 135416 50953 135444 51054
rect 135402 50944 135458 50953
rect 135402 50879 135458 50888
rect 136782 50672 136838 50681
rect 136782 50607 136838 50616
rect 171650 50672 171706 50681
rect 171650 50607 171652 50616
rect 135404 50296 135456 50302
rect 135404 50238 135456 50244
rect 135310 49856 135366 49865
rect 135310 49791 135366 49800
rect 102650 49312 102706 49321
rect 102468 49276 102520 49282
rect 102650 49247 102706 49256
rect 134850 49312 134906 49321
rect 134850 49247 134906 49256
rect 102468 49218 102520 49224
rect 66402 48768 66458 48777
rect 66402 48703 66458 48712
rect 102374 48768 102430 48777
rect 102374 48703 102430 48712
rect 64930 48224 64986 48233
rect 64930 48159 64986 48168
rect 63734 47816 63790 47825
rect 63734 47751 63790 47760
rect 62906 47272 62962 47281
rect 62906 47207 62962 47216
rect 64944 47174 64972 48159
rect 66416 47825 66444 48703
rect 100626 48360 100682 48369
rect 100626 48295 100682 48304
rect 100640 47922 100668 48295
rect 102480 48097 102508 49218
rect 102560 49004 102612 49010
rect 102560 48946 102612 48952
rect 102466 48088 102522 48097
rect 102466 48023 102522 48032
rect 100628 47916 100680 47922
rect 100628 47858 100680 47864
rect 65022 47816 65078 47825
rect 65022 47751 65078 47760
rect 66402 47816 66458 47825
rect 66402 47751 66458 47760
rect 65036 47242 65064 47751
rect 100626 47680 100682 47689
rect 100626 47615 100628 47624
rect 100680 47615 100682 47624
rect 102376 47644 102428 47650
rect 100628 47586 100680 47592
rect 102376 47586 102428 47592
rect 66402 47544 66458 47553
rect 66402 47479 66404 47488
rect 66456 47479 66458 47488
rect 100626 47544 100682 47553
rect 100626 47479 100628 47488
rect 66404 47450 66456 47456
rect 100680 47479 100682 47488
rect 100628 47450 100680 47456
rect 65024 47236 65076 47242
rect 65024 47178 65076 47184
rect 62908 47168 62960 47174
rect 62908 47110 62960 47116
rect 64932 47168 64984 47174
rect 64932 47110 64984 47116
rect 62920 46193 62948 47110
rect 66402 47000 66458 47009
rect 66402 46935 66458 46944
rect 66416 46426 66444 46935
rect 102388 46465 102416 47586
rect 102572 47553 102600 48946
rect 135312 48868 135364 48874
rect 135312 48810 135364 48816
rect 134760 48460 134812 48466
rect 134760 48402 134812 48408
rect 102652 47916 102704 47922
rect 102652 47858 102704 47864
rect 102558 47544 102614 47553
rect 102468 47508 102520 47514
rect 102558 47479 102614 47488
rect 102468 47450 102520 47456
rect 100626 46456 100682 46465
rect 63736 46420 63788 46426
rect 63736 46362 63788 46368
rect 66404 46420 66456 46426
rect 100626 46391 100682 46400
rect 102374 46456 102430 46465
rect 102374 46391 102430 46400
rect 66404 46362 66456 46368
rect 62906 46184 62962 46193
rect 62906 46119 62962 46128
rect 62814 45640 62870 45649
rect 62814 45575 62870 45584
rect 63748 44969 63776 46362
rect 65298 46320 65354 46329
rect 100640 46290 100668 46391
rect 65298 46255 65354 46264
rect 100628 46284 100680 46290
rect 63734 44960 63790 44969
rect 63734 44895 63790 44904
rect 63736 44856 63788 44862
rect 63736 44798 63788 44804
rect 63644 44788 63696 44794
rect 63644 44730 63696 44736
rect 62816 44720 62868 44726
rect 62816 44662 62868 44668
rect 62828 44425 62856 44662
rect 62814 44416 62870 44425
rect 62814 44351 62870 44360
rect 63656 43337 63684 44730
rect 63748 43881 63776 44798
rect 65312 44726 65340 46255
rect 100628 46226 100680 46232
rect 100902 46184 100958 46193
rect 100902 46119 100904 46128
rect 100956 46119 100958 46128
rect 102376 46148 102428 46154
rect 100904 46090 100956 46096
rect 102376 46090 102428 46096
rect 66402 45776 66458 45785
rect 66402 45711 66458 45720
rect 65666 45232 65722 45241
rect 65666 45167 65722 45176
rect 65680 44794 65708 45167
rect 66416 44862 66444 45711
rect 100534 45368 100590 45377
rect 100534 45303 100590 45312
rect 100548 45270 100576 45303
rect 100536 45264 100588 45270
rect 100536 45206 100588 45212
rect 99982 45096 100038 45105
rect 99982 45031 100038 45040
rect 99996 44998 100024 45031
rect 99984 44992 100036 44998
rect 99984 44934 100036 44940
rect 66404 44856 66456 44862
rect 66404 44798 66456 44804
rect 65668 44788 65720 44794
rect 65668 44730 65720 44736
rect 65300 44720 65352 44726
rect 102388 44697 102416 46090
rect 102480 45921 102508 47450
rect 102664 47009 102692 47858
rect 134772 47553 134800 48402
rect 135324 48097 135352 48810
rect 135416 48777 135444 50238
rect 136796 50234 136824 50607
rect 171704 50607 171706 50616
rect 171652 50578 171704 50584
rect 136874 50400 136930 50409
rect 136874 50335 136930 50344
rect 136888 50302 136916 50335
rect 136876 50296 136928 50302
rect 136876 50238 136928 50244
rect 172662 50264 172718 50273
rect 136784 50228 136836 50234
rect 172718 50222 172796 50250
rect 172662 50199 172718 50208
rect 136784 50170 136836 50176
rect 136874 49448 136930 49457
rect 136874 49383 136930 49392
rect 171834 49448 171890 49457
rect 171834 49383 171890 49392
rect 136888 48942 136916 49383
rect 171848 48942 171876 49383
rect 172662 49040 172718 49049
rect 172662 48975 172664 48984
rect 172716 48975 172718 48984
rect 172664 48946 172716 48952
rect 136876 48936 136928 48942
rect 136782 48904 136838 48913
rect 136876 48878 136928 48884
rect 171836 48936 171888 48942
rect 171836 48878 171888 48884
rect 172768 48874 172796 50222
rect 173780 49865 173808 51666
rect 173872 51633 173900 53026
rect 174056 52177 174084 53162
rect 174136 52948 174188 52954
rect 174136 52890 174188 52896
rect 174148 52721 174176 52890
rect 174134 52712 174190 52721
rect 174134 52647 174190 52656
rect 174042 52168 174098 52177
rect 174042 52103 174098 52112
rect 173952 51860 174004 51866
rect 173952 51802 174004 51808
rect 173858 51624 173914 51633
rect 173858 51559 173914 51568
rect 173964 50409 173992 51802
rect 174044 51656 174096 51662
rect 174044 51598 174096 51604
rect 174056 50953 174084 51598
rect 174042 50944 174098 50953
rect 174042 50879 174098 50888
rect 174044 50636 174096 50642
rect 174044 50578 174096 50584
rect 173950 50400 174006 50409
rect 173950 50335 174006 50344
rect 173766 49856 173822 49865
rect 173766 49791 173822 49800
rect 174056 49321 174084 50578
rect 174042 49312 174098 49321
rect 174042 49247 174098 49256
rect 173952 49004 174004 49010
rect 173952 48946 174004 48952
rect 136782 48839 136838 48848
rect 172756 48868 172808 48874
rect 135402 48768 135458 48777
rect 135402 48703 135458 48712
rect 136796 48466 136824 48839
rect 172756 48810 172808 48816
rect 136784 48460 136836 48466
rect 136784 48402 136836 48408
rect 136690 48360 136746 48369
rect 136690 48295 136746 48304
rect 172110 48360 172166 48369
rect 172110 48295 172166 48304
rect 135310 48088 135366 48097
rect 135310 48023 135366 48032
rect 134758 47544 134814 47553
rect 134758 47479 134814 47488
rect 135404 47508 135456 47514
rect 135404 47450 135456 47456
rect 134852 47372 134904 47378
rect 134852 47314 134904 47320
rect 102650 47000 102706 47009
rect 102650 46935 102706 46944
rect 134864 46465 134892 47314
rect 135312 47168 135364 47174
rect 135312 47110 135364 47116
rect 135324 47009 135352 47110
rect 135310 47000 135366 47009
rect 135310 46935 135366 46944
rect 134850 46456 134906 46465
rect 134850 46391 134906 46400
rect 102560 46284 102612 46290
rect 102560 46226 102612 46232
rect 102466 45912 102522 45921
rect 102466 45847 102522 45856
rect 102468 45264 102520 45270
rect 102572 45241 102600 46226
rect 134668 46080 134720 46086
rect 134668 46022 134720 46028
rect 134680 45241 134708 46022
rect 135416 45921 135444 47450
rect 136704 47174 136732 48295
rect 136782 47680 136838 47689
rect 172124 47650 172152 48295
rect 172662 47952 172718 47961
rect 172662 47887 172718 47896
rect 172570 47680 172626 47689
rect 136782 47615 136838 47624
rect 172112 47644 172164 47650
rect 136796 47378 136824 47615
rect 172570 47615 172626 47624
rect 172112 47586 172164 47592
rect 172584 47582 172612 47615
rect 172572 47576 172624 47582
rect 136874 47544 136930 47553
rect 172572 47518 172624 47524
rect 172676 47514 172704 47887
rect 173860 47576 173912 47582
rect 173964 47553 173992 48946
rect 174044 48936 174096 48942
rect 174044 48878 174096 48884
rect 174056 48097 174084 48878
rect 174136 48868 174188 48874
rect 174136 48810 174188 48816
rect 174148 48777 174176 48810
rect 174134 48768 174190 48777
rect 174134 48703 174190 48712
rect 174042 48088 174098 48097
rect 174042 48023 174098 48032
rect 174044 47644 174096 47650
rect 174044 47586 174096 47592
rect 173860 47518 173912 47524
rect 173950 47544 174006 47553
rect 136874 47479 136876 47488
rect 136928 47479 136930 47488
rect 172664 47508 172716 47514
rect 136876 47450 136928 47456
rect 172664 47450 172716 47456
rect 136784 47372 136836 47378
rect 136784 47314 136836 47320
rect 136692 47168 136744 47174
rect 136692 47110 136744 47116
rect 136782 46456 136838 46465
rect 136782 46391 136838 46400
rect 172662 46456 172718 46465
rect 172662 46391 172664 46400
rect 136796 46086 136824 46391
rect 172716 46391 172718 46400
rect 172664 46362 172716 46368
rect 137518 46184 137574 46193
rect 137518 46119 137574 46128
rect 172662 46184 172718 46193
rect 172718 46142 172796 46170
rect 172662 46119 172718 46128
rect 136784 46080 136836 46086
rect 136784 46022 136836 46028
rect 135402 45912 135458 45921
rect 135402 45847 135458 45856
rect 136690 45368 136746 45377
rect 136690 45303 136746 45312
rect 102468 45206 102520 45212
rect 102558 45232 102614 45241
rect 65300 44662 65352 44668
rect 102374 44688 102430 44697
rect 102374 44623 102430 44632
rect 65298 44552 65354 44561
rect 65298 44487 65354 44496
rect 63734 43872 63790 43881
rect 63734 43807 63790 43816
rect 63920 43564 63972 43570
rect 63920 43506 63972 43512
rect 63736 43360 63788 43366
rect 63642 43328 63698 43337
rect 63736 43302 63788 43308
rect 63642 43263 63698 43272
rect 63748 42793 63776 43302
rect 63828 42884 63880 42890
rect 63828 42826 63880 42832
rect 63734 42784 63790 42793
rect 63734 42719 63790 42728
rect 63736 42000 63788 42006
rect 63736 41942 63788 41948
rect 63748 41025 63776 41942
rect 63840 41569 63868 42826
rect 63932 42113 63960 43506
rect 65312 43366 65340 44487
rect 102480 44153 102508 45206
rect 102558 45167 102614 45176
rect 134666 45232 134722 45241
rect 134666 45167 134722 45176
rect 102560 44992 102612 44998
rect 102560 44934 102612 44940
rect 99890 44144 99946 44153
rect 102466 44144 102522 44153
rect 99890 44079 99892 44088
rect 99944 44079 99946 44088
rect 102284 44108 102336 44114
rect 99892 44050 99944 44056
rect 102466 44079 102522 44088
rect 102284 44050 102336 44056
rect 66402 44008 66458 44017
rect 66402 43943 66458 43952
rect 66416 43570 66444 43943
rect 66404 43564 66456 43570
rect 66404 43506 66456 43512
rect 100626 43464 100682 43473
rect 100626 43399 100682 43408
rect 100640 43366 100668 43399
rect 65300 43360 65352 43366
rect 100628 43360 100680 43366
rect 65300 43302 65352 43308
rect 66402 43328 66458 43337
rect 100628 43302 100680 43308
rect 66402 43263 66458 43272
rect 66416 42890 66444 43263
rect 102296 43065 102324 44050
rect 102572 43609 102600 44934
rect 135036 44720 135088 44726
rect 135034 44688 135036 44697
rect 135088 44688 135090 44697
rect 135034 44623 135090 44632
rect 136704 44454 136732 45303
rect 136782 44960 136838 44969
rect 136782 44895 136838 44904
rect 135404 44448 135456 44454
rect 135404 44390 135456 44396
rect 136692 44448 136744 44454
rect 136692 44390 136744 44396
rect 135036 44312 135088 44318
rect 135036 44254 135088 44260
rect 135048 43609 135076 44254
rect 135416 44153 135444 44390
rect 136796 44318 136824 44895
rect 137532 44726 137560 46119
rect 172768 46034 172796 46142
rect 172768 46006 172888 46034
rect 171834 45368 171890 45377
rect 171834 45303 171890 45312
rect 171848 44794 171876 45303
rect 172662 44960 172718 44969
rect 172718 44918 172796 44946
rect 172662 44895 172718 44904
rect 171836 44788 171888 44794
rect 171836 44730 171888 44736
rect 137520 44720 137572 44726
rect 137520 44662 137572 44668
rect 172768 44318 172796 44918
rect 172860 44726 172888 46006
rect 173872 45921 173900 47518
rect 173950 47479 174006 47488
rect 174056 47009 174084 47586
rect 174228 47440 174280 47446
rect 174228 47382 174280 47388
rect 174042 47000 174098 47009
rect 174042 46935 174098 46944
rect 174240 46465 174268 47382
rect 174226 46456 174282 46465
rect 174044 46420 174096 46426
rect 174226 46391 174282 46400
rect 174044 46362 174096 46368
rect 173858 45912 173914 45921
rect 173858 45847 173914 45856
rect 174056 45241 174084 46362
rect 174042 45232 174098 45241
rect 174042 45167 174098 45176
rect 172848 44720 172900 44726
rect 174136 44720 174188 44726
rect 172848 44662 172900 44668
rect 174134 44688 174136 44697
rect 174188 44688 174190 44697
rect 174134 44623 174190 44632
rect 174688 44652 174740 44658
rect 174688 44594 174740 44600
rect 136784 44312 136836 44318
rect 136784 44254 136836 44260
rect 172756 44312 172808 44318
rect 172756 44254 172808 44260
rect 174504 44312 174556 44318
rect 174504 44254 174556 44260
rect 135402 44144 135458 44153
rect 135402 44079 135458 44088
rect 136782 44144 136838 44153
rect 136782 44079 136838 44088
rect 171834 44144 171890 44153
rect 171834 44079 171890 44088
rect 102558 43600 102614 43609
rect 102558 43535 102614 43544
rect 135034 43600 135090 43609
rect 135034 43535 135090 43544
rect 102376 43292 102428 43298
rect 102376 43234 102428 43240
rect 134944 43292 134996 43298
rect 134944 43234 134996 43240
rect 102282 43056 102338 43065
rect 102282 42991 102338 43000
rect 100626 42920 100682 42929
rect 66404 42884 66456 42890
rect 100626 42855 100682 42864
rect 66404 42826 66456 42832
rect 66402 42784 66458 42793
rect 66402 42719 66458 42728
rect 65298 42240 65354 42249
rect 65298 42175 65354 42184
rect 63918 42104 63974 42113
rect 63918 42039 63974 42048
rect 63826 41560 63882 41569
rect 63826 41495 63882 41504
rect 63734 41016 63790 41025
rect 63734 40951 63790 40960
rect 65312 40578 65340 42175
rect 66416 42006 66444 42719
rect 100640 42686 100668 42855
rect 100628 42680 100680 42686
rect 100628 42622 100680 42628
rect 102388 42385 102416 43234
rect 102560 42680 102612 42686
rect 102560 42622 102612 42628
rect 100626 42376 100682 42385
rect 100626 42311 100682 42320
rect 102374 42376 102430 42385
rect 102374 42311 102430 42320
rect 100640 42210 100668 42311
rect 100628 42204 100680 42210
rect 100628 42146 100680 42152
rect 102468 42204 102520 42210
rect 102468 42146 102520 42152
rect 100626 42104 100682 42113
rect 100626 42039 100628 42048
rect 100680 42039 100682 42048
rect 102376 42068 102428 42074
rect 100628 42010 100680 42016
rect 102376 42010 102428 42016
rect 66404 42000 66456 42006
rect 66404 41942 66456 41948
rect 71628 41926 71964 41954
rect 79080 41926 79416 41954
rect 62816 40572 62868 40578
rect 62816 40514 62868 40520
rect 65300 40572 65352 40578
rect 65300 40514 65352 40520
rect 62828 40481 62856 40514
rect 62814 40472 62870 40481
rect 62814 40407 62870 40416
rect 66402 40472 66458 40481
rect 66402 40407 66458 40416
rect 66312 39892 66364 39898
rect 66312 39834 66364 39840
rect 62814 39520 62870 39529
rect 62814 39455 62870 39464
rect 62828 39218 62856 39455
rect 62816 39212 62868 39218
rect 62816 39154 62868 39160
rect 30524 33636 30576 33642
rect 30524 33578 30576 33584
rect 66220 33636 66272 33642
rect 66220 33578 66272 33584
rect 66232 32729 66260 33578
rect 66218 32720 66274 32729
rect 66218 32655 66274 32664
rect 66324 24705 66352 39834
rect 66310 24696 66366 24705
rect 66310 24631 66366 24640
rect 13318 19664 13374 19673
rect 13318 19599 13374 19608
rect 66416 16817 66444 40407
rect 71936 39966 71964 41926
rect 71924 39960 71976 39966
rect 71924 39902 71976 39908
rect 72568 39212 72620 39218
rect 72568 39154 72620 39160
rect 72580 36786 72608 39154
rect 79388 37790 79416 41926
rect 86288 41926 86624 41954
rect 94016 41926 94076 41954
rect 82504 39960 82556 39966
rect 82504 39902 82556 39908
rect 79376 37784 79428 37790
rect 79376 37726 79428 37732
rect 82516 36786 82544 39902
rect 86288 39898 86316 41926
rect 94016 40481 94044 41926
rect 102388 40753 102416 42010
rect 102480 41297 102508 42146
rect 102572 41841 102600 42622
rect 134956 42385 134984 43234
rect 136796 43094 136824 44079
rect 171848 43570 171876 44079
rect 174516 43609 174544 44254
rect 174700 44153 174728 44594
rect 174686 44144 174742 44153
rect 174686 44079 174742 44088
rect 172662 43600 172718 43609
rect 171836 43564 171888 43570
rect 174502 43600 174558 43609
rect 172662 43535 172718 43544
rect 174044 43564 174096 43570
rect 171836 43506 171888 43512
rect 136874 43464 136930 43473
rect 136874 43399 136930 43408
rect 136888 43366 136916 43399
rect 172676 43366 172704 43535
rect 174502 43535 174558 43544
rect 174044 43506 174096 43512
rect 136876 43360 136928 43366
rect 136876 43302 136928 43308
rect 172664 43360 172716 43366
rect 172664 43302 172716 43308
rect 135404 43088 135456 43094
rect 135402 43056 135404 43065
rect 136784 43088 136836 43094
rect 135456 43056 135458 43065
rect 174056 43065 174084 43506
rect 174228 43292 174280 43298
rect 174228 43234 174280 43240
rect 136784 43030 136836 43036
rect 174042 43056 174098 43065
rect 135402 42991 135458 43000
rect 174042 42991 174098 43000
rect 136690 42920 136746 42929
rect 136690 42855 136746 42864
rect 172570 42920 172626 42929
rect 172570 42855 172626 42864
rect 134942 42376 134998 42385
rect 134942 42311 134998 42320
rect 135404 41932 135456 41938
rect 135404 41874 135456 41880
rect 135312 41864 135364 41870
rect 102558 41832 102614 41841
rect 102558 41767 102614 41776
rect 135310 41832 135312 41841
rect 135364 41832 135366 41841
rect 135310 41767 135366 41776
rect 134852 41524 134904 41530
rect 134852 41466 134904 41472
rect 102466 41288 102522 41297
rect 102466 41223 102522 41232
rect 134864 40753 134892 41466
rect 135416 41297 135444 41874
rect 136704 41870 136732 42855
rect 136874 42376 136930 42385
rect 136874 42311 136930 42320
rect 172386 42376 172442 42385
rect 172386 42311 172388 42320
rect 136782 42104 136838 42113
rect 136782 42039 136838 42048
rect 136692 41864 136744 41870
rect 136692 41806 136744 41812
rect 136796 41530 136824 42039
rect 136888 42006 136916 42311
rect 172440 42311 172442 42320
rect 172388 42282 172440 42288
rect 172584 42006 172612 42855
rect 174240 42385 174268 43234
rect 174226 42376 174282 42385
rect 173952 42340 174004 42346
rect 174226 42311 174282 42320
rect 173952 42282 174004 42288
rect 172662 42104 172718 42113
rect 172662 42039 172664 42048
rect 172716 42039 172718 42048
rect 172664 42010 172716 42016
rect 136876 42000 136928 42006
rect 136876 41942 136928 41948
rect 172572 42000 172624 42006
rect 172572 41942 172624 41948
rect 136784 41524 136836 41530
rect 136784 41466 136836 41472
rect 135402 41288 135458 41297
rect 135402 41223 135458 41232
rect 102374 40744 102430 40753
rect 102374 40679 102430 40688
rect 134850 40744 134906 40753
rect 134850 40679 134906 40688
rect 94002 40472 94058 40481
rect 94002 40407 94058 40416
rect 102374 40200 102430 40209
rect 102374 40135 102430 40144
rect 86276 39892 86328 39898
rect 86276 39834 86328 39840
rect 102388 39218 102416 40135
rect 109642 40064 109698 40073
rect 109532 40022 109642 40050
rect 109642 39999 109698 40008
rect 143604 39966 143632 41940
rect 143592 39960 143644 39966
rect 118824 39886 118884 39914
rect 93176 39212 93228 39218
rect 93176 39154 93228 39160
rect 102376 39212 102428 39218
rect 102376 39154 102428 39160
rect 93188 36786 93216 39154
rect 72580 36758 72916 36786
rect 82516 36758 82852 36786
rect 92880 36758 93216 36786
rect 118856 33642 118884 39886
rect 127780 39886 128116 39914
rect 143592 39902 143644 39908
rect 138072 39892 138124 39898
rect 127780 37790 127808 39886
rect 138072 39834 138124 39840
rect 134482 39656 134538 39665
rect 134482 39591 134538 39600
rect 134496 39218 134524 39591
rect 134484 39212 134536 39218
rect 134484 39154 134536 39160
rect 127768 37784 127820 37790
rect 127768 37726 127820 37732
rect 118844 33636 118896 33642
rect 118844 33578 118896 33584
rect 136876 33636 136928 33642
rect 136876 33578 136928 33584
rect 136888 33409 136916 33578
rect 136874 33400 136930 33409
rect 136874 33335 136930 33344
rect 138084 25113 138112 39834
rect 138162 39792 138218 39801
rect 138162 39727 138218 39736
rect 138070 25104 138126 25113
rect 138070 25039 138126 25048
rect 138176 17089 138204 39727
rect 144880 39212 144932 39218
rect 144880 39154 144932 39160
rect 144892 36772 144920 39154
rect 151056 37790 151084 41940
rect 154816 39960 154868 39966
rect 154816 39902 154868 39908
rect 151044 37784 151096 37790
rect 151044 37726 151096 37732
rect 154828 36772 154856 39902
rect 158600 39898 158628 41940
rect 158588 39892 158640 39898
rect 158588 39834 158640 39840
rect 166052 39801 166080 41940
rect 173964 41297 173992 42282
rect 174044 42068 174096 42074
rect 174044 42010 174096 42016
rect 173950 41288 174006 41297
rect 173950 41223 174006 41232
rect 174056 40753 174084 42010
rect 174136 41932 174188 41938
rect 174136 41874 174188 41880
rect 174148 41841 174176 41874
rect 174134 41832 174190 41841
rect 174134 41767 174190 41776
rect 174042 40744 174098 40753
rect 174042 40679 174098 40688
rect 181402 40064 181458 40073
rect 181458 40022 181522 40050
rect 181402 39999 181458 40008
rect 166038 39792 166094 39801
rect 166038 39727 166094 39736
rect 174134 39520 174190 39529
rect 174134 39455 174190 39464
rect 174148 39218 174176 39455
rect 164844 39212 164896 39218
rect 164844 39154 164896 39160
rect 174136 39212 174188 39218
rect 174136 39154 174188 39160
rect 164856 36772 164884 39154
rect 190800 37722 190828 39900
rect 200092 37790 200120 39900
rect 200080 37784 200132 37790
rect 200080 37726 200132 37732
rect 205152 37722 205180 68802
rect 222540 44561 222568 141902
rect 222816 127550 222844 142038
rect 222908 139761 222936 146782
rect 223552 141966 223580 149479
rect 223540 141960 223592 141966
rect 223540 141902 223592 141908
rect 222894 139752 222950 139761
rect 222894 139687 222950 139696
rect 222804 127544 222856 127550
rect 222804 127486 222856 127492
rect 222712 124824 222764 124830
rect 222712 124766 222764 124772
rect 222724 116210 222752 124766
rect 222724 116182 223028 116210
rect 222710 115952 222766 115961
rect 222710 115887 222766 115896
rect 222620 115100 222672 115106
rect 222620 115042 222672 115048
rect 222632 103290 222660 115042
rect 222724 110278 222752 115887
rect 223000 115106 223028 116182
rect 222988 115100 223040 115106
rect 222988 115042 223040 115048
rect 222712 110272 222764 110278
rect 222712 110214 222764 110220
rect 222804 107960 222856 107966
rect 222724 107908 222804 107914
rect 222724 107902 222856 107908
rect 222724 107886 222844 107902
rect 222724 103426 222752 107886
rect 224472 105761 224500 163487
rect 224458 105752 224514 105761
rect 224458 105687 224514 105696
rect 222724 103398 223028 103426
rect 222632 103262 222752 103290
rect 222724 97034 222752 103262
rect 223000 97154 223028 103398
rect 222988 97148 223040 97154
rect 222988 97090 223040 97096
rect 223540 97148 223592 97154
rect 223540 97090 223592 97096
rect 222724 97006 222844 97034
rect 222816 92598 222844 97006
rect 223552 96377 223580 97090
rect 223538 96368 223594 96377
rect 223538 96303 223594 96312
rect 222804 92592 222856 92598
rect 222804 92534 222856 92540
rect 223540 92592 223592 92598
rect 223540 92534 223592 92540
rect 223552 92161 223580 92534
rect 223538 92152 223594 92161
rect 223538 92087 223594 92096
rect 223538 85216 223594 85225
rect 223538 85151 223594 85160
rect 223552 84846 223580 85151
rect 222804 84840 222856 84846
rect 222724 84788 222804 84794
rect 222724 84782 222856 84788
rect 223540 84840 223592 84846
rect 223540 84782 223592 84788
rect 222724 84766 222844 84782
rect 222724 73642 222752 84766
rect 223538 75288 223594 75297
rect 223538 75223 223594 75232
rect 223552 75122 223580 75223
rect 222988 75116 223040 75122
rect 222988 75058 223040 75064
rect 223540 75116 223592 75122
rect 223540 75058 223592 75064
rect 222724 73626 222844 73642
rect 222724 73620 222856 73626
rect 222724 73614 222804 73620
rect 222804 73562 222856 73568
rect 223000 68066 223028 75058
rect 223080 73620 223132 73626
rect 223080 73562 223132 73568
rect 223092 68361 223120 73562
rect 223078 68352 223134 68361
rect 223078 68287 223134 68296
rect 222632 68038 223028 68066
rect 222632 63986 222660 68038
rect 222632 63958 222752 63986
rect 222526 44552 222582 44561
rect 222526 44487 222582 44496
rect 222724 40730 222752 63958
rect 222540 40702 222752 40730
rect 222540 40594 222568 40702
rect 222448 40566 222568 40594
rect 222448 40458 222476 40566
rect 222448 40430 222568 40458
rect 222540 37790 222568 40430
rect 222528 37784 222580 37790
rect 222528 37726 222580 37732
rect 190788 37716 190840 37722
rect 190788 37658 190840 37664
rect 205140 37716 205192 37722
rect 205140 37658 205192 37664
rect 222712 28196 222764 28202
rect 222712 28138 222764 28144
rect 222724 20761 222752 28138
rect 222710 20752 222766 20761
rect 222710 20687 222766 20696
rect 138162 17080 138218 17089
rect 138162 17015 138218 17024
rect 66402 16808 66458 16817
rect 66402 16743 66458 16752
rect 71292 12822 71628 12850
rect 71292 10998 71320 12822
rect 79066 12630 79094 12836
rect 86624 12822 86960 12850
rect 77996 12624 78048 12630
rect 77996 12566 78048 12572
rect 79054 12624 79106 12630
rect 79054 12566 79106 12572
rect 23532 10992 23584 10998
rect 23532 10934 23584 10940
rect 71280 10992 71332 10998
rect 71280 10934 71332 10940
rect 23544 9304 23572 10934
rect 50764 10924 50816 10930
rect 50764 10866 50816 10872
rect 50776 9304 50804 10866
rect 78008 9304 78036 12566
rect 86932 11746 86960 12822
rect 94016 12822 94076 12850
rect 86920 11740 86972 11746
rect 86920 11682 86972 11688
rect 94016 11678 94044 12822
rect 132552 11740 132604 11746
rect 132552 11682 132604 11688
rect 94004 11672 94056 11678
rect 94004 11614 94056 11620
rect 105228 10992 105280 10998
rect 105228 10934 105280 10940
rect 105240 9304 105268 10934
rect 132564 9304 132592 11682
rect 143604 10930 143632 12836
rect 151056 10998 151084 12836
rect 151044 10992 151096 10998
rect 151044 10934 151096 10940
rect 143592 10924 143644 10930
rect 143592 10866 143644 10872
rect 158600 10454 158628 12836
rect 166052 11746 166080 12836
rect 166040 11740 166092 11746
rect 166040 11682 166092 11688
rect 214248 11740 214300 11746
rect 214248 11682 214300 11688
rect 187016 11672 187068 11678
rect 187016 11614 187068 11620
rect 158588 10448 158640 10454
rect 158588 10390 158640 10396
rect 159784 10448 159836 10454
rect 159784 10390 159836 10396
rect 159796 9304 159824 10390
rect 187028 9304 187056 11614
rect 214260 9304 214288 11682
rect 23530 8824 23586 9304
rect 50762 8824 50818 9304
rect 77994 8824 78050 9304
rect 105226 8824 105282 9304
rect 132550 8824 132606 9304
rect 159782 8824 159838 9304
rect 187014 8824 187070 9304
rect 214246 8824 214302 9304
<< via2 >>
rect 98234 238704 98290 238760
rect 169994 238704 170050 238760
rect 55822 217216 55878 217272
rect 62538 215312 62594 215368
rect 62630 214632 62686 214688
rect 10466 214224 10522 214280
rect 63642 213952 63698 214008
rect 62538 213292 62594 213328
rect 62538 213272 62540 213292
rect 62540 213272 62592 213292
rect 62592 213272 62594 213292
rect 10466 213136 10522 213192
rect 98326 230680 98382 230736
rect 168522 230136 168578 230192
rect 98418 222792 98474 222848
rect 135402 215584 135458 215640
rect 102374 215312 102430 215368
rect 102374 214652 102430 214688
rect 102374 214632 102376 214652
rect 102376 214632 102428 214652
rect 102428 214632 102430 214652
rect 135402 214632 135458 214688
rect 65022 213544 65078 213600
rect 102374 213952 102430 214008
rect 135034 213952 135090 214008
rect 100994 213408 101050 213464
rect 151042 215856 151098 215912
rect 223078 234896 223134 234952
rect 170086 222812 170142 222848
rect 170086 222792 170088 222812
rect 170088 222792 170140 222812
rect 170140 222792 170142 222812
rect 174226 215720 174282 215776
rect 174042 214632 174098 214688
rect 171834 213988 171836 214008
rect 171836 213988 171888 214008
rect 171888 213988 171890 214008
rect 171834 213952 171890 213988
rect 174226 213952 174282 214008
rect 136782 213408 136838 213464
rect 62354 212592 62410 212648
rect 66218 212864 66274 212920
rect 102466 213272 102522 213328
rect 135402 213272 135458 213328
rect 174042 213272 174098 213328
rect 172662 213036 172664 213056
rect 172664 213036 172716 213056
rect 172716 213036 172718 213056
rect 100994 212864 101050 212920
rect 136782 212864 136838 212920
rect 102374 212592 102430 212648
rect 134666 212592 134722 212648
rect 65022 212184 65078 212240
rect 100534 212184 100590 212240
rect 62630 211912 62686 211968
rect 62630 211232 62686 211288
rect 66402 211640 66458 211696
rect 65022 211096 65078 211152
rect 64930 210688 64986 210744
rect 62630 210552 62686 210608
rect 172662 213000 172718 213036
rect 171742 212592 171798 212648
rect 174226 212592 174282 212648
rect 136874 212184 136930 212240
rect 102374 211932 102430 211968
rect 102374 211912 102376 211932
rect 102376 211912 102428 211932
rect 102428 211912 102430 211932
rect 134298 211912 134354 211968
rect 101086 211640 101142 211696
rect 174042 211912 174098 211968
rect 136966 211640 137022 211696
rect 172662 211504 172718 211560
rect 172570 211404 172572 211424
rect 172572 211404 172624 211424
rect 172624 211404 172626 211424
rect 172570 211368 172626 211404
rect 174134 211232 174190 211288
rect 100994 211096 101050 211152
rect 136874 211096 136930 211152
rect 66402 210688 66458 210744
rect 171834 210724 171836 210744
rect 171836 210724 171888 210744
rect 171888 210724 171890 210744
rect 171834 210688 171890 210724
rect 65482 210416 65538 210472
rect 62630 209872 62686 209928
rect 174134 209872 174190 209928
rect 65022 209464 65078 209520
rect 171926 209328 171982 209384
rect 62722 209192 62778 209248
rect 65482 209192 65538 209248
rect 135310 209192 135366 209248
rect 174594 209192 174650 209248
rect 171466 208784 171522 208840
rect 65022 208648 65078 208704
rect 137702 208648 137758 208704
rect 62538 208512 62594 208568
rect 65666 208124 65722 208160
rect 65666 208104 65668 208124
rect 65668 208104 65720 208124
rect 65720 208104 65722 208124
rect 135402 207832 135458 207888
rect 174042 207832 174098 207888
rect 136874 207424 136930 207480
rect 172570 207324 172572 207344
rect 172572 207324 172624 207344
rect 172624 207324 172626 207344
rect 172570 207288 172626 207324
rect 62630 207152 62686 207208
rect 65666 206900 65722 206936
rect 65666 206880 65668 206900
rect 65668 206880 65720 206900
rect 65720 206880 65722 206900
rect 172662 202276 172718 202312
rect 172662 202256 172664 202276
rect 172664 202256 172716 202276
rect 172716 202256 172718 202276
rect 65022 202120 65078 202176
rect 174226 201984 174282 202040
rect 62630 201712 62686 201768
rect 65022 200896 65078 200952
rect 172662 200780 172718 200816
rect 172662 200760 172664 200780
rect 172664 200760 172716 200780
rect 172716 200760 172718 200780
rect 100902 200660 100904 200680
rect 100904 200660 100956 200680
rect 100956 200660 100958 200680
rect 100902 200624 100958 200660
rect 62630 200388 62632 200408
rect 62632 200388 62684 200408
rect 62684 200388 62686 200408
rect 62630 200352 62686 200388
rect 136782 200624 136838 200680
rect 102374 200352 102430 200408
rect 135402 200352 135458 200408
rect 174134 200352 174190 200408
rect 65022 199672 65078 199728
rect 171650 199536 171706 199592
rect 136782 199400 136838 199456
rect 100902 199300 100904 199320
rect 100904 199300 100956 199320
rect 100956 199300 100958 199320
rect 100902 199264 100958 199300
rect 62354 199028 62356 199048
rect 62356 199028 62408 199048
rect 62408 199028 62410 199048
rect 62354 198992 62410 199028
rect 102374 198992 102430 199048
rect 134758 198992 134814 199048
rect 175238 198992 175294 199048
rect 65022 198448 65078 198504
rect 172662 198196 172718 198232
rect 172662 198176 172664 198196
rect 172664 198176 172716 198196
rect 172716 198176 172718 198196
rect 100810 198060 100866 198096
rect 100810 198040 100812 198060
rect 100812 198040 100864 198060
rect 100864 198040 100866 198060
rect 136782 198040 136838 198096
rect 172662 198060 172718 198096
rect 172662 198040 172664 198060
rect 172664 198040 172716 198060
rect 172716 198040 172718 198060
rect 65666 197924 65722 197960
rect 65666 197904 65668 197924
rect 65668 197904 65720 197924
rect 65720 197904 65722 197924
rect 100902 197924 100958 197960
rect 100902 197904 100904 197924
rect 100904 197904 100956 197924
rect 100956 197904 100958 197924
rect 136690 197904 136746 197960
rect 62630 197632 62686 197688
rect 102374 197632 102430 197688
rect 65022 197224 65078 197280
rect 62538 196952 62594 197008
rect 62538 196308 62540 196328
rect 62540 196308 62592 196328
rect 62592 196308 62594 196328
rect 62538 196272 62594 196308
rect 135402 197632 135458 197688
rect 174134 197632 174190 197688
rect 174226 197496 174282 197552
rect 135402 197396 135404 197416
rect 135404 197396 135456 197416
rect 135456 197396 135458 197416
rect 135402 197360 135458 197396
rect 102466 196952 102522 197008
rect 100718 196816 100774 196872
rect 136782 196816 136838 196872
rect 172570 196836 172626 196872
rect 172570 196816 172572 196836
rect 172572 196816 172624 196836
rect 172624 196816 172626 196836
rect 66218 196680 66274 196736
rect 100902 196564 100958 196600
rect 100902 196544 100904 196564
rect 100904 196544 100956 196564
rect 100956 196544 100958 196564
rect 136690 196544 136746 196600
rect 102374 196272 102430 196328
rect 65022 195728 65078 195784
rect 62630 195592 62686 195648
rect 135402 196272 135458 196328
rect 172662 196564 172718 196600
rect 172662 196544 172664 196564
rect 172664 196544 172716 196564
rect 172716 196544 172718 196564
rect 174134 196272 174190 196328
rect 135402 196172 135404 196192
rect 135404 196172 135456 196192
rect 135456 196172 135458 196192
rect 135402 196136 135458 196172
rect 174226 196136 174282 196192
rect 172386 195728 172442 195784
rect 100902 195592 100958 195648
rect 102466 195592 102522 195648
rect 136874 195592 136930 195648
rect 66402 195456 66458 195512
rect 100902 195204 100958 195240
rect 100902 195184 100904 195204
rect 100904 195184 100956 195204
rect 100956 195184 100958 195204
rect 62630 194912 62686 194968
rect 65022 194504 65078 194560
rect 62538 194232 62594 194288
rect 64930 193688 64986 193744
rect 62538 193588 62540 193608
rect 62540 193588 62592 193608
rect 62592 193588 62594 193608
rect 62538 193552 62594 193588
rect 62630 192872 62686 192928
rect 11938 192600 11994 192656
rect 62538 192228 62540 192248
rect 62540 192228 62592 192248
rect 62592 192228 62594 192248
rect 62538 192192 62594 192228
rect 62354 191512 62410 191568
rect 100626 194388 100682 194424
rect 100626 194368 100628 194388
rect 100628 194368 100680 194388
rect 100680 194368 100682 194388
rect 136782 195184 136838 195240
rect 172662 195340 172718 195376
rect 172662 195320 172664 195340
rect 172664 195320 172716 195340
rect 172716 195320 172718 195340
rect 102558 194912 102614 194968
rect 135402 194912 135458 194968
rect 135402 194812 135404 194832
rect 135404 194812 135456 194832
rect 135456 194812 135458 194832
rect 135402 194776 135458 194812
rect 174226 194912 174282 194968
rect 174134 194776 174190 194832
rect 136782 194368 136838 194424
rect 171742 194368 171798 194424
rect 66402 194232 66458 194288
rect 102374 194232 102430 194288
rect 100626 193844 100682 193880
rect 100626 193824 100628 193844
rect 100628 193824 100680 193844
rect 100680 193824 100682 193844
rect 99890 193280 99946 193336
rect 136690 193824 136746 193880
rect 102466 193552 102522 193608
rect 135402 193552 135458 193608
rect 172662 193960 172718 194016
rect 174134 193552 174190 193608
rect 135402 193452 135404 193472
rect 135404 193452 135456 193472
rect 135456 193452 135458 193472
rect 135402 193416 135458 193452
rect 174226 193416 174282 193472
rect 136782 193280 136838 193336
rect 172018 193280 172074 193336
rect 102374 192872 102430 192928
rect 65022 192736 65078 192792
rect 100626 192600 100682 192656
rect 65666 192484 65722 192520
rect 65666 192464 65668 192484
rect 65668 192464 65720 192484
rect 65720 192464 65722 192484
rect 100534 192464 100590 192520
rect 136690 192600 136746 192656
rect 102466 192192 102522 192248
rect 65022 191512 65078 191568
rect 102374 191512 102430 191568
rect 62630 190832 62686 190888
rect 100626 191376 100682 191432
rect 65206 191240 65262 191296
rect 62354 190152 62410 190208
rect 62630 189508 62632 189528
rect 62632 189508 62684 189528
rect 62684 189508 62686 189528
rect 62630 189472 62686 189508
rect 62630 188792 62686 188848
rect 65022 189608 65078 189664
rect 100902 191104 100958 191160
rect 66310 190696 66366 190752
rect 100442 190288 100498 190344
rect 66402 190152 66458 190208
rect 102282 190152 102338 190208
rect 99982 189900 100038 189936
rect 99982 189880 99984 189900
rect 99984 189880 100036 189900
rect 100036 189880 100038 189900
rect 66310 189608 66366 189664
rect 102374 188792 102430 188848
rect 135218 192092 135220 192112
rect 135220 192092 135272 192112
rect 135272 192092 135274 192112
rect 135218 192056 135274 192092
rect 102650 190832 102706 190888
rect 135402 192192 135458 192248
rect 172662 192756 172718 192792
rect 172662 192736 172664 192756
rect 172664 192736 172716 192756
rect 172716 192736 172718 192756
rect 171650 192620 171706 192656
rect 171650 192600 171652 192620
rect 171652 192600 171704 192620
rect 171704 192600 171706 192620
rect 136874 192464 136930 192520
rect 174134 192192 174190 192248
rect 174226 192056 174282 192112
rect 136782 191376 136838 191432
rect 172662 191376 172718 191432
rect 135310 190832 135366 190888
rect 137150 191104 137206 191160
rect 171834 191124 171890 191160
rect 171834 191104 171836 191124
rect 171836 191104 171888 191124
rect 171888 191104 171890 191124
rect 135402 190732 135404 190752
rect 135404 190732 135456 190752
rect 135456 190732 135458 190752
rect 135402 190696 135458 190732
rect 223538 211096 223594 211152
rect 207898 201712 207954 201768
rect 207254 192464 207310 192520
rect 207254 192328 207310 192384
rect 174318 190832 174374 190888
rect 174042 190696 174098 190752
rect 136782 190288 136838 190344
rect 171650 190288 171706 190344
rect 102558 189472 102614 189528
rect 134206 189472 134262 189528
rect 137242 189880 137298 189936
rect 171834 189880 171890 189936
rect 134758 189236 134760 189256
rect 134760 189236 134812 189256
rect 134812 189236 134814 189256
rect 134758 189200 134814 189236
rect 175330 189472 175386 189528
rect 174410 189200 174466 189256
rect 63642 188112 63698 188168
rect 102466 188112 102522 188168
rect 134942 188148 134944 188168
rect 134944 188148 134996 188168
rect 134996 188148 134998 188168
rect 134942 188112 134998 188148
rect 175422 188112 175478 188168
rect 11938 179680 11994 179736
rect 38158 184460 38214 184496
rect 38158 184440 38160 184460
rect 38160 184440 38212 184460
rect 38212 184440 38214 184460
rect 40182 184440 40238 184496
rect 54902 184168 54958 184224
rect 60146 184168 60202 184224
rect 31994 178184 32050 178240
rect 37422 178184 37478 178240
rect 59594 178184 59650 178240
rect 12030 170976 12086 171032
rect 11938 149760 11994 149816
rect 12122 169208 12178 169264
rect 105594 184712 105650 184768
rect 105594 182264 105650 182320
rect 105318 178456 105374 178512
rect 105226 177912 105282 177968
rect 105134 176688 105190 176744
rect 57386 174784 57442 174840
rect 106146 183624 106202 183680
rect 117094 185392 117150 185448
rect 116910 184712 116966 184768
rect 118198 185392 118254 185448
rect 119118 185392 119174 185448
rect 117646 184712 117702 184768
rect 118106 184712 118162 184768
rect 119486 185256 119542 185312
rect 119578 184712 119634 184768
rect 121142 185392 121198 185448
rect 121602 185256 121658 185312
rect 120682 185120 120738 185176
rect 122430 185120 122486 185176
rect 120314 184984 120370 185040
rect 122890 184984 122946 185040
rect 125098 185256 125154 185312
rect 124914 184848 124970 184904
rect 125466 185120 125522 185176
rect 126662 185392 126718 185448
rect 125834 184984 125890 185040
rect 126478 184712 126534 184768
rect 129974 185256 130030 185312
rect 130434 185120 130490 185176
rect 131446 184984 131502 185040
rect 129330 184848 129386 184904
rect 132182 185392 132238 185448
rect 131630 184712 131686 184768
rect 108538 183488 108594 183544
rect 106054 181176 106110 181232
rect 108078 181176 108134 181232
rect 105962 179816 106018 179872
rect 107894 178864 107950 178920
rect 106146 175364 106148 175384
rect 106148 175364 106200 175384
rect 106200 175364 106202 175384
rect 106146 175328 106202 175364
rect 105410 174376 105466 174432
rect 107894 176416 107950 176472
rect 106330 172880 106386 172936
rect 176986 180768 177042 180824
rect 176894 177368 176950 177424
rect 177722 184168 177778 184224
rect 177354 183080 177410 183136
rect 177170 181856 177226 181912
rect 197456 184984 197512 185040
rect 202194 184984 202250 185040
rect 198514 184440 198570 184496
rect 203390 184440 203446 184496
rect 198882 184168 198938 184224
rect 203942 184168 203998 184224
rect 180298 183488 180354 183544
rect 179654 181176 179710 181232
rect 177814 179680 177870 179736
rect 177630 178456 177686 178512
rect 177078 176144 177134 176200
rect 177170 175056 177226 175112
rect 107894 174104 107950 174160
rect 106422 172200 106478 172256
rect 108078 171792 108134 171848
rect 105962 170976 106018 171032
rect 179654 178864 179710 178920
rect 179654 176416 179710 176472
rect 225194 187296 225250 187352
rect 207254 182944 207310 183000
rect 225194 179680 225250 179736
rect 204494 178184 204550 178240
rect 201090 177640 201146 177696
rect 179654 174104 179710 174160
rect 178090 173968 178146 174024
rect 177814 172744 177870 172800
rect 179654 171792 179710 171848
rect 177722 171656 177778 171712
rect 177538 170432 177594 170488
rect 105686 169888 105742 169944
rect 178182 169344 178238 169400
rect 106606 167304 106662 167360
rect 106514 166896 106570 166952
rect 223538 169208 223594 169264
rect 177170 165944 177226 166000
rect 105226 165400 105282 165456
rect 32638 164856 32694 164912
rect 37422 164856 37478 164912
rect 59594 164856 59650 164912
rect 200998 164856 201054 164912
rect 204494 164856 204550 164912
rect 12214 159280 12270 159336
rect 12122 149352 12178 149408
rect 12122 127728 12178 127784
rect 12030 105696 12086 105752
rect 31994 151528 32050 151584
rect 107802 164720 107858 164776
rect 177538 164720 177594 164776
rect 179562 164720 179618 164776
rect 105778 164176 105834 164232
rect 105594 163516 105650 163552
rect 105594 163496 105596 163516
rect 105596 163496 105648 163516
rect 105648 163496 105650 163516
rect 176986 163632 177042 163688
rect 105686 162272 105742 162328
rect 105226 161068 105282 161104
rect 105226 161048 105228 161068
rect 105228 161048 105280 161068
rect 105280 161048 105282 161068
rect 176986 162544 177042 162600
rect 107802 162408 107858 162464
rect 107434 159960 107490 160016
rect 105594 159688 105650 159744
rect 105778 158464 105834 158520
rect 106146 157940 106202 157976
rect 106146 157920 106148 157940
rect 106148 157920 106200 157940
rect 106200 157920 106202 157940
rect 106146 156716 106202 156752
rect 106146 156696 106148 156716
rect 106148 156696 106200 156716
rect 106200 156696 106202 156716
rect 105778 155356 105834 155392
rect 105778 155336 105780 155356
rect 105780 155336 105832 155356
rect 105832 155336 105834 155356
rect 57478 154792 57534 154848
rect 106422 154112 106478 154168
rect 105226 151664 105282 151720
rect 59594 151548 59650 151584
rect 59594 151528 59596 151548
rect 59596 151528 59648 151548
rect 59648 151528 59650 151548
rect 105134 149624 105190 149680
rect 31902 141328 31958 141384
rect 62814 142008 62870 142064
rect 62814 140920 62870 140976
rect 62722 140648 62778 140704
rect 62814 139696 62870 139752
rect 62814 139424 62870 139480
rect 62722 138880 62778 138936
rect 62354 137656 62410 137712
rect 30522 137112 30578 137168
rect 30430 127728 30486 127784
rect 12214 106104 12270 106160
rect 12122 95768 12178 95824
rect 12030 75096 12086 75152
rect 11938 62856 11994 62912
rect 62814 137112 62870 137168
rect 91242 141872 91298 141928
rect 102282 142552 102338 142608
rect 101178 142416 101234 142472
rect 66218 139424 66274 139480
rect 100626 139016 100682 139072
rect 66402 138880 66458 138936
rect 100534 138608 100590 138664
rect 63458 138336 63514 138392
rect 66218 138200 66274 138256
rect 66402 137656 66458 137712
rect 100350 137248 100406 137304
rect 62906 136568 62962 136624
rect 66034 136432 66090 136488
rect 65022 136160 65078 136216
rect 62722 135616 62778 135672
rect 62630 135344 62686 135400
rect 62722 134800 62778 134856
rect 62906 134256 62962 134312
rect 66402 135888 66458 135944
rect 100994 138372 100996 138392
rect 100996 138372 101048 138392
rect 101048 138372 101050 138392
rect 100994 138336 101050 138372
rect 100718 137792 100774 137848
rect 100626 136044 100682 136080
rect 100626 136024 100628 136044
rect 100628 136024 100680 136044
rect 100680 136024 100682 136044
rect 100902 136568 100958 136624
rect 100902 135908 100958 135944
rect 100902 135888 100904 135908
rect 100904 135888 100956 135908
rect 100956 135888 100958 135908
rect 66310 135208 66366 135264
rect 100074 134800 100130 134856
rect 66402 134664 66458 134720
rect 100902 134664 100958 134720
rect 65850 134120 65906 134176
rect 62998 133576 63054 133632
rect 62814 132760 62870 132816
rect 62722 132488 62778 132544
rect 62814 130756 62816 130776
rect 62816 130756 62868 130776
rect 62868 130756 62870 130776
rect 62814 130720 62870 130756
rect 100074 133576 100130 133632
rect 66402 133440 66458 133496
rect 100902 133188 100958 133224
rect 100902 133168 100904 133188
rect 100904 133168 100956 133188
rect 100956 133168 100958 133188
rect 105410 150984 105466 151040
rect 105962 147176 106018 147232
rect 177538 161320 177594 161376
rect 177354 160232 177410 160288
rect 179562 162408 179618 162464
rect 179194 159960 179250 160016
rect 177630 159008 177686 159064
rect 107802 157648 107858 157704
rect 107710 155336 107766 155392
rect 106606 152888 106662 152944
rect 107618 152888 107674 152944
rect 106698 148264 106754 148320
rect 178182 157940 178238 157976
rect 178182 157920 178184 157940
rect 178184 157920 178236 157940
rect 178236 157920 178238 157940
rect 177354 156832 177410 156888
rect 178090 155608 178146 155664
rect 178274 154520 178330 154576
rect 132366 151528 132422 151584
rect 108722 150576 108778 150632
rect 108630 148264 108686 148320
rect 108538 145952 108594 146008
rect 176894 151120 176950 151176
rect 177170 149896 177226 149952
rect 134114 142008 134170 142064
rect 103110 141464 103166 141520
rect 102282 140920 102338 140976
rect 102374 140376 102430 140432
rect 102374 139696 102430 139752
rect 102466 139152 102522 139208
rect 102558 138608 102614 138664
rect 102374 137928 102430 137984
rect 102466 137384 102522 137440
rect 102834 136840 102890 136896
rect 102466 136296 102522 136352
rect 101178 134528 101234 134584
rect 102374 135616 102430 135672
rect 102190 133848 102246 133904
rect 102098 133304 102154 133360
rect 65022 132488 65078 132544
rect 63642 131536 63698 131592
rect 63550 131264 63606 131320
rect 100442 132352 100498 132408
rect 66402 132216 66458 132272
rect 65666 131708 65668 131728
rect 65668 131708 65720 131728
rect 65720 131708 65722 131728
rect 65666 131672 65722 131708
rect 100902 131944 100958 132000
rect 100902 131708 100904 131728
rect 100904 131708 100956 131728
rect 100956 131708 100958 131728
rect 100902 131672 100958 131708
rect 66310 131128 66366 131184
rect 100442 130604 100498 130640
rect 100442 130584 100444 130604
rect 100444 130584 100496 130604
rect 100496 130584 100498 130604
rect 66402 130448 66458 130504
rect 100902 130448 100958 130504
rect 63458 130176 63514 130232
rect 65482 129904 65538 129960
rect 63274 129496 63330 129552
rect 62722 128680 62778 128736
rect 62630 128408 62686 128464
rect 62814 127456 62870 127512
rect 100074 129360 100130 129416
rect 66402 129224 66458 129280
rect 102098 131536 102154 131592
rect 102650 135072 102706 135128
rect 102466 134528 102522 134584
rect 102282 132760 102338 132816
rect 102374 132216 102430 132272
rect 102190 130992 102246 131048
rect 102006 129224 102062 129280
rect 100902 128988 100904 129008
rect 100904 128988 100956 129008
rect 100956 128988 100958 129008
rect 100902 128952 100958 128988
rect 100350 128272 100406 128328
rect 66402 128136 66458 128192
rect 65022 127864 65078 127920
rect 62906 127184 62962 127240
rect 102374 130448 102430 130504
rect 102374 129768 102430 129824
rect 102282 128680 102338 128736
rect 102190 128136 102246 128192
rect 100534 127612 100590 127648
rect 100534 127592 100536 127612
rect 100536 127592 100588 127612
rect 100588 127592 100590 127612
rect 100442 127048 100498 127104
rect 66310 126912 66366 126968
rect 62814 126640 62870 126696
rect 65022 126504 65078 126560
rect 62630 125960 62686 126016
rect 62814 125416 62870 125472
rect 62722 124600 62778 124656
rect 66402 126232 66458 126288
rect 100902 126368 100958 126424
rect 100810 126268 100812 126288
rect 100812 126268 100864 126288
rect 100864 126268 100866 126288
rect 100810 126232 100866 126268
rect 102098 127456 102154 127512
rect 102190 126912 102246 126968
rect 102282 126368 102338 126424
rect 66310 125688 66366 125744
rect 102006 125688 102062 125744
rect 100902 125280 100958 125336
rect 66402 125144 66458 125200
rect 100810 124892 100866 124928
rect 100810 124872 100812 124892
rect 100812 124872 100864 124892
rect 100864 124872 100866 124892
rect 65022 124736 65078 124792
rect 66310 124736 66366 124792
rect 62906 124328 62962 124384
rect 100258 124056 100314 124112
rect 66402 123920 66458 123976
rect 62814 123648 62870 123704
rect 65022 123648 65078 123704
rect 62630 123104 62686 123160
rect 62814 122560 62870 122616
rect 62814 121336 62870 121392
rect 102098 123920 102154 123976
rect 100902 123376 100958 123432
rect 100166 122832 100222 122888
rect 66310 122696 66366 122752
rect 65022 122424 65078 122480
rect 63550 121608 63606 121664
rect 63458 120520 63514 120576
rect 100626 122424 100682 122480
rect 66402 122152 66458 122208
rect 100902 122172 100958 122208
rect 100902 122152 100904 122172
rect 100904 122152 100956 122172
rect 100956 122152 100958 122172
rect 101822 122968 101878 123024
rect 100074 121064 100130 121120
rect 66218 120928 66274 120984
rect 65022 120656 65078 120712
rect 63642 120248 63698 120304
rect 65482 119704 65538 119760
rect 62814 119568 62870 119624
rect 65022 119432 65078 119488
rect 62722 118752 62778 118808
rect 62814 118480 62870 118536
rect 100902 120948 100958 120984
rect 100902 120928 100904 120948
rect 100904 120928 100956 120948
rect 100956 120928 100958 120948
rect 100442 119840 100498 119896
rect 100902 119296 100958 119352
rect 66402 119160 66458 119216
rect 64930 118480 64986 118536
rect 62906 117800 62962 117856
rect 62814 117292 62816 117312
rect 62816 117292 62868 117312
rect 62868 117292 62870 117312
rect 62814 117256 62870 117292
rect 100626 118616 100682 118672
rect 65022 118208 65078 118264
rect 66402 118208 66458 118264
rect 100258 118072 100314 118128
rect 66402 117936 66458 117992
rect 100534 117936 100590 117992
rect 62814 116712 62870 116768
rect 66402 116712 66458 116768
rect 100258 116732 100314 116768
rect 100258 116712 100260 116732
rect 100260 116712 100312 116732
rect 100312 116712 100314 116732
rect 65022 116440 65078 116496
rect 62722 116168 62778 116224
rect 62814 115488 62870 115544
rect 65022 115080 65078 115136
rect 62814 114672 62870 114728
rect 100902 116848 100958 116904
rect 62814 114400 62870 114456
rect 56926 113176 56982 113232
rect 31994 104200 32050 104256
rect 37422 104200 37478 104256
rect 56834 100800 56890 100856
rect 32638 90872 32694 90928
rect 36410 90872 36466 90928
rect 72014 113176 72070 113232
rect 100902 115508 100958 115544
rect 100902 115488 100904 115508
rect 100904 115488 100956 115508
rect 100956 115488 100958 115508
rect 102374 125144 102430 125200
rect 102282 124600 102338 124656
rect 102374 123376 102430 123432
rect 102190 122832 102246 122888
rect 102282 122288 102338 122344
rect 102374 121608 102430 121664
rect 102282 121064 102338 121120
rect 102098 120520 102154 120576
rect 102006 119840 102062 119896
rect 102374 119296 102430 119352
rect 102190 118752 102246 118808
rect 102282 118208 102338 118264
rect 134298 138880 134354 138936
rect 134482 138336 134538 138392
rect 135402 140920 135458 140976
rect 135402 140684 135404 140704
rect 135404 140684 135456 140704
rect 135456 140684 135458 140704
rect 135402 140648 135458 140684
rect 135402 139696 135458 139752
rect 162174 141872 162230 141928
rect 174134 144864 174190 144920
rect 174226 140648 174282 140704
rect 135402 139460 135404 139480
rect 135404 139460 135456 139480
rect 135456 139460 135458 139480
rect 135402 139424 135458 139460
rect 174318 139424 174374 139480
rect 136874 139016 136930 139072
rect 172478 139016 172534 139072
rect 134574 137656 134630 137712
rect 136966 138880 137022 138936
rect 172662 138744 172718 138800
rect 135126 136568 135182 136624
rect 135034 134800 135090 134856
rect 136874 137792 136930 137848
rect 172202 137792 172258 137848
rect 136966 137268 137022 137304
rect 136966 137248 136968 137268
rect 136968 137248 137020 137268
rect 137020 137248 137022 137268
rect 174134 137656 174190 137712
rect 172662 137268 172718 137304
rect 172662 137248 172664 137268
rect 172664 137248 172716 137268
rect 172716 137248 172718 137268
rect 135402 136840 135458 136896
rect 136782 136568 136838 136624
rect 172018 136568 172074 136624
rect 135310 135616 135366 135672
rect 135218 135344 135274 135400
rect 136874 136024 136930 136080
rect 136966 135908 137022 135944
rect 136966 135888 136968 135908
rect 136968 135888 137020 135908
rect 137020 135888 137022 135908
rect 172570 136180 172626 136216
rect 172570 136160 172572 136180
rect 172572 136160 172624 136180
rect 172624 136160 172626 136180
rect 172662 136044 172718 136080
rect 172662 136024 172664 136044
rect 172664 136024 172716 136044
rect 172716 136024 172718 136044
rect 173950 135616 174006 135672
rect 174226 137112 174282 137168
rect 174318 136568 174374 136624
rect 174042 135344 174098 135400
rect 136874 134800 136930 134856
rect 171834 134800 171890 134856
rect 135126 134256 135182 134312
rect 134942 133576 134998 133632
rect 136966 134664 137022 134720
rect 172662 134548 172718 134584
rect 172662 134528 172664 134548
rect 172664 134528 172716 134548
rect 172716 134528 172718 134548
rect 135218 132488 135274 132544
rect 135126 131536 135182 131592
rect 134942 129496 134998 129552
rect 174318 134800 174374 134856
rect 174134 134256 174190 134312
rect 136966 133576 137022 133632
rect 172202 133596 172258 133632
rect 172202 133576 172204 133596
rect 172204 133576 172256 133596
rect 172256 133576 172258 133596
rect 172662 133168 172718 133224
rect 136874 133052 136930 133088
rect 136874 133032 136876 133052
rect 136876 133032 136928 133052
rect 136928 133032 136930 133052
rect 135402 132760 135458 132816
rect 174226 132760 174282 132816
rect 174318 132488 174374 132544
rect 136782 132352 136838 132408
rect 172386 132352 172442 132408
rect 135310 131264 135366 131320
rect 136874 131944 136930 132000
rect 172018 131944 172074 132000
rect 172662 131828 172718 131864
rect 172662 131808 172664 131828
rect 172664 131808 172716 131828
rect 172716 131808 172718 131828
rect 136966 131708 136968 131728
rect 136968 131708 137020 131728
rect 137020 131708 137022 131728
rect 136966 131672 137022 131708
rect 135310 130720 135366 130776
rect 172662 130720 172718 130776
rect 136874 130584 136930 130640
rect 136966 130448 137022 130504
rect 172662 130332 172718 130368
rect 172662 130312 172664 130332
rect 172664 130312 172716 130332
rect 172716 130312 172718 130332
rect 135218 130176 135274 130232
rect 135034 128408 135090 128464
rect 135126 127456 135182 127512
rect 134666 126640 134722 126696
rect 171834 129496 171890 129552
rect 136966 129360 137022 129416
rect 171834 129108 171890 129144
rect 171834 129088 171836 129108
rect 171836 129088 171888 129108
rect 171888 129088 171890 129108
rect 136874 128972 136930 129008
rect 136874 128952 136876 128972
rect 136876 128952 136928 128972
rect 136928 128952 136930 128972
rect 135402 128680 135458 128736
rect 136782 128272 136838 128328
rect 172570 128272 172626 128328
rect 135310 127184 135366 127240
rect 171558 127864 171614 127920
rect 136874 127612 136930 127648
rect 136874 127592 136876 127612
rect 136876 127592 136928 127612
rect 136928 127592 136930 127612
rect 174226 128680 174282 128736
rect 174318 128408 174374 128464
rect 174134 127456 174190 127512
rect 136782 127048 136838 127104
rect 172018 127048 172074 127104
rect 135218 125960 135274 126016
rect 135034 124328 135090 124384
rect 136874 126368 136930 126424
rect 136966 126252 137022 126288
rect 136966 126232 136968 126252
rect 136968 126232 137020 126252
rect 137020 126232 137022 126252
rect 172202 126640 172258 126696
rect 174226 126640 174282 126696
rect 172662 126096 172718 126152
rect 135402 125416 135458 125472
rect 174134 125416 174190 125472
rect 136782 125280 136838 125336
rect 171834 125300 171890 125336
rect 171834 125280 171836 125300
rect 171836 125280 171888 125300
rect 171888 125280 171890 125300
rect 135310 124600 135366 124656
rect 172202 125008 172258 125064
rect 136874 124872 136930 124928
rect 136782 124056 136838 124112
rect 171834 124056 171890 124112
rect 135218 123648 135274 123704
rect 135126 123104 135182 123160
rect 135310 122560 135366 122616
rect 136874 123396 136930 123432
rect 174318 124600 174374 124656
rect 172570 123648 172626 123704
rect 174226 123648 174282 123704
rect 136874 123376 136876 123396
rect 136876 123376 136928 123396
rect 136928 123376 136930 123396
rect 136874 122832 136930 122888
rect 171834 122832 171890 122888
rect 136966 122424 137022 122480
rect 174134 122560 174190 122616
rect 172018 122424 172074 122480
rect 137058 122172 137114 122208
rect 137058 122152 137060 122172
rect 137060 122152 137112 122172
rect 137112 122152 137114 122172
rect 172662 122036 172718 122072
rect 172662 122016 172664 122036
rect 172664 122016 172716 122036
rect 172716 122016 172718 122036
rect 135402 121880 135458 121936
rect 135310 121336 135366 121392
rect 136782 121064 136838 121120
rect 172110 121064 172166 121120
rect 135218 120520 135274 120576
rect 135126 120248 135182 120304
rect 172662 120812 172718 120848
rect 172662 120792 172664 120812
rect 172664 120792 172716 120812
rect 172716 120792 172718 120812
rect 136966 120656 137022 120712
rect 136782 119840 136838 119896
rect 134850 119568 134906 119624
rect 102374 117528 102430 117584
rect 102282 116984 102338 117040
rect 102466 116440 102522 116496
rect 102190 114672 102246 114728
rect 102650 115760 102706 115816
rect 102374 115216 102430 115272
rect 102282 114128 102338 114184
rect 101822 113720 101878 113776
rect 59870 104200 59926 104256
rect 105318 109132 105320 109152
rect 105320 109132 105372 109152
rect 105372 109132 105374 109152
rect 105318 109096 105374 109132
rect 105410 106784 105466 106840
rect 105226 105696 105282 105752
rect 105778 110184 105834 110240
rect 105686 107872 105742 107928
rect 134114 117256 134170 117312
rect 134666 116712 134722 116768
rect 135310 119024 135366 119080
rect 136874 119316 136930 119352
rect 136874 119296 136876 119316
rect 136876 119296 136928 119316
rect 136928 119296 136930 119316
rect 171834 119840 171890 119896
rect 171834 119568 171890 119624
rect 136966 118616 137022 118672
rect 171834 118616 171890 118672
rect 135310 118516 135312 118536
rect 135312 118516 135364 118536
rect 135364 118516 135366 118536
rect 135310 118480 135366 118516
rect 136782 118072 136838 118128
rect 135218 117528 135274 117584
rect 136874 117956 136930 117992
rect 136874 117936 136876 117956
rect 136876 117936 136928 117956
rect 136928 117936 136930 117956
rect 171650 118228 171706 118264
rect 171650 118208 171652 118228
rect 171652 118208 171704 118228
rect 171704 118208 171706 118228
rect 174318 119568 174374 119624
rect 174226 119024 174282 119080
rect 174134 118480 174190 118536
rect 172662 118092 172718 118128
rect 172662 118072 172664 118092
rect 172664 118072 172716 118092
rect 172716 118072 172718 118092
rect 136782 116848 136838 116904
rect 172662 116848 172718 116904
rect 135126 116168 135182 116224
rect 134850 115488 134906 115544
rect 136874 116712 136930 116768
rect 172570 116576 172626 116632
rect 174042 117256 174098 117312
rect 173950 116712 174006 116768
rect 136782 115488 136838 115544
rect 135310 114944 135366 115000
rect 134850 114436 134852 114456
rect 134852 114436 134904 114456
rect 134904 114436 134906 114456
rect 134850 114400 134906 114436
rect 108538 109504 108594 109560
rect 107894 107212 107950 107248
rect 107894 107192 107896 107212
rect 107896 107192 107948 107212
rect 107948 107192 107950 107212
rect 106054 104472 106110 104528
rect 105594 103384 105650 103440
rect 105134 102160 105190 102216
rect 105962 101072 106018 101128
rect 105778 98760 105834 98816
rect 108446 104880 108502 104936
rect 107894 102432 107950 102488
rect 171834 115644 171890 115680
rect 171834 115624 171836 115644
rect 171836 115624 171888 115644
rect 171888 115624 171890 115644
rect 174134 115488 174190 115544
rect 174318 116168 174374 116224
rect 174226 114944 174282 115000
rect 174042 114400 174098 114456
rect 132274 105424 132330 105480
rect 132550 105424 132606 105480
rect 107894 100120 107950 100176
rect 106422 99984 106478 100040
rect 106330 97672 106386 97728
rect 107894 97808 107950 97864
rect 106422 96448 106478 96504
rect 106238 95360 106294 95416
rect 108446 95360 108502 95416
rect 106514 94272 106570 94328
rect 105870 91708 105926 91744
rect 105870 91688 105872 91708
rect 105872 91688 105924 91708
rect 105924 91688 105926 91708
rect 59594 90872 59650 90928
rect 107802 90736 107858 90792
rect 105226 90328 105282 90384
rect 105134 89260 105190 89296
rect 105134 89240 105136 89260
rect 105136 89240 105188 89260
rect 105188 89240 105190 89260
rect 105870 87880 105926 87936
rect 106422 86656 106478 86712
rect 105594 86248 105650 86304
rect 106330 84772 106386 84808
rect 106330 84752 106332 84772
rect 106332 84752 106384 84772
rect 106384 84752 106386 84772
rect 105594 83412 105650 83448
rect 105594 83392 105596 83412
rect 105596 83392 105648 83412
rect 105648 83392 105650 83412
rect 105502 82168 105558 82224
rect 107894 88424 107950 88480
rect 107802 85976 107858 86032
rect 107710 83664 107766 83720
rect 56926 81896 56982 81952
rect 57478 81896 57534 81952
rect 107894 81352 107950 81408
rect 105226 80944 105282 81000
rect 57478 80808 57534 80864
rect 105134 79856 105190 79912
rect 106974 79312 107030 79368
rect 106330 77816 106386 77872
rect 31994 77544 32050 77600
rect 37422 77544 37478 77600
rect 59594 77580 59596 77600
rect 59596 77580 59648 77600
rect 59648 77580 59650 77600
rect 31902 68704 31958 68760
rect 48278 68976 48334 69032
rect 49474 68976 49530 69032
rect 49014 68840 49070 68896
rect 50854 68840 50910 68896
rect 59594 77544 59650 77580
rect 105410 76456 105466 76512
rect 105226 75232 105282 75288
rect 103202 73532 103258 73588
rect 102558 73328 102614 73384
rect 102558 71968 102614 72024
rect 102650 71832 102706 71888
rect 62814 66664 62870 66720
rect 62722 66120 62778 66176
rect 62906 65576 62962 65632
rect 62814 64896 62870 64952
rect 62722 64352 62778 64408
rect 63366 67208 63422 67264
rect 62998 63808 63054 63864
rect 62354 63264 62410 63320
rect 29234 62856 29290 62912
rect 12030 41232 12086 41288
rect 91242 69248 91298 69304
rect 66402 65440 66458 65496
rect 66402 64896 66458 64952
rect 63274 62720 63330 62776
rect 66402 64236 66458 64272
rect 66402 64216 66404 64236
rect 66404 64216 66456 64236
rect 66456 64216 66458 64236
rect 101362 71152 101418 71208
rect 101914 71016 101970 71072
rect 102650 70880 102706 70936
rect 102466 67480 102522 67536
rect 102374 66936 102430 66992
rect 102558 66392 102614 66448
rect 102374 65848 102430 65904
rect 100902 65460 100958 65496
rect 100902 65440 100904 65460
rect 100904 65440 100956 65460
rect 100956 65440 100958 65460
rect 100626 64488 100682 64544
rect 100902 64100 100958 64136
rect 100902 64080 100904 64100
rect 100904 64080 100956 64100
rect 100956 64080 100958 64100
rect 66310 63672 66366 63728
rect 102374 63536 102430 63592
rect 100442 63264 100498 63320
rect 66402 63128 66458 63184
rect 100902 62740 100958 62776
rect 100902 62720 100904 62740
rect 100904 62720 100956 62740
rect 100956 62720 100958 62740
rect 66310 62448 66366 62504
rect 63550 62040 63606 62096
rect 63458 61496 63514 61552
rect 100258 62040 100314 62096
rect 66402 61904 66458 61960
rect 63182 60952 63238 61008
rect 62814 60408 62870 60464
rect 100902 61380 100958 61416
rect 100902 61360 100904 61380
rect 100904 61360 100956 61380
rect 100956 61360 100958 61380
rect 66218 61224 66274 61280
rect 102650 65168 102706 65224
rect 102742 64624 102798 64680
rect 106422 74144 106478 74200
rect 108722 78904 108778 78960
rect 108814 76592 108870 76648
rect 108630 74280 108686 74336
rect 108538 71968 108594 72024
rect 117830 69112 117886 69168
rect 117094 68568 117150 68624
rect 118198 68568 118254 68624
rect 119394 69112 119450 69168
rect 119118 68432 119174 68488
rect 121142 68432 121198 68488
rect 175238 142180 175240 142200
rect 175240 142180 175292 142200
rect 175292 142180 175294 142200
rect 175238 142144 175294 142180
rect 174778 140920 174834 140976
rect 174962 139696 175018 139752
rect 177354 147584 177410 147640
rect 178550 153296 178606 153352
rect 178458 152208 178514 152264
rect 178366 148808 178422 148864
rect 179562 157648 179618 157704
rect 179470 155336 179526 155392
rect 179378 152888 179434 152944
rect 200538 151548 200594 151584
rect 200538 151528 200540 151548
rect 200540 151528 200592 151548
rect 200592 151528 200594 151548
rect 180482 150576 180538 150632
rect 180390 148264 180446 148320
rect 180298 145952 180354 146008
rect 224458 163496 224514 163552
rect 207438 163224 207494 163280
rect 223538 159144 223594 159200
rect 207438 153704 207494 153760
rect 207346 153296 207402 153352
rect 204494 151528 204550 151584
rect 175422 138880 175478 138936
rect 175146 138336 175202 138392
rect 207254 137112 207310 137168
rect 174502 133576 174558 133632
rect 174870 131264 174926 131320
rect 175330 131536 175386 131592
rect 175422 130720 175478 130776
rect 175238 130176 175294 130232
rect 175146 129496 175202 129552
rect 174502 127184 174558 127240
rect 174594 125960 174650 126016
rect 174502 124328 174558 124384
rect 174594 123104 174650 123160
rect 175054 121336 175110 121392
rect 175330 121608 175386 121664
rect 175422 120520 175478 120576
rect 175146 120248 175202 120304
rect 204678 117936 204734 117992
rect 174502 117800 174558 117856
rect 176986 106784 177042 106840
rect 177170 109096 177226 109152
rect 177262 107872 177318 107928
rect 177078 105696 177134 105752
rect 177722 110184 177778 110240
rect 180298 109504 180354 109560
rect 179654 107192 179710 107248
rect 177446 104472 177502 104528
rect 177354 103384 177410 103440
rect 176894 102160 176950 102216
rect 176986 101072 177042 101128
rect 179654 104880 179710 104936
rect 177538 99984 177594 100040
rect 177630 97672 177686 97728
rect 179654 102432 179710 102488
rect 223538 149488 223594 149544
rect 207990 127728 208046 127784
rect 207898 118480 207954 118536
rect 201090 104200 201146 104256
rect 204586 104200 204642 104256
rect 179654 100120 179710 100176
rect 177814 98760 177870 98816
rect 179654 97808 179710 97864
rect 177722 96448 177778 96504
rect 177538 95360 177594 95416
rect 179562 95360 179618 95416
rect 177446 94308 177448 94328
rect 177448 94308 177500 94328
rect 177500 94308 177502 94328
rect 177446 94272 177502 94308
rect 177538 91960 177594 92016
rect 204494 90872 204550 90928
rect 177354 90736 177410 90792
rect 179562 90736 179618 90792
rect 200998 90328 201054 90384
rect 177354 89648 177410 89704
rect 177354 88560 177410 88616
rect 178918 87336 178974 87392
rect 178090 86248 178146 86304
rect 177538 85024 177594 85080
rect 178182 83936 178238 83992
rect 177722 82848 177778 82904
rect 177354 81624 177410 81680
rect 179654 88424 179710 88480
rect 179562 85976 179618 86032
rect 179470 83664 179526 83720
rect 178918 81352 178974 81408
rect 178182 80536 178238 80592
rect 178826 79312 178882 79368
rect 178274 78224 178330 78280
rect 177722 77136 177778 77192
rect 177170 75912 177226 75968
rect 174502 72920 174558 72976
rect 135310 67480 135366 67536
rect 135034 66936 135090 66992
rect 135310 66428 135312 66448
rect 135312 66428 135364 66448
rect 135364 66428 135366 66448
rect 135310 66392 135366 66428
rect 134666 65848 134722 65904
rect 102834 64080 102890 64136
rect 134482 64080 134538 64136
rect 102558 62992 102614 63048
rect 102466 62312 102522 62368
rect 102374 61224 102430 61280
rect 63734 60136 63790 60192
rect 62722 59184 62778 59240
rect 100626 60816 100682 60872
rect 66310 60680 66366 60736
rect 100902 60272 100958 60328
rect 66402 60156 66458 60192
rect 135310 65204 135312 65224
rect 135312 65204 135364 65224
rect 135364 65204 135366 65224
rect 135310 65168 135366 65204
rect 135034 64624 135090 64680
rect 134666 62992 134722 63048
rect 102650 61768 102706 61824
rect 102558 60680 102614 60736
rect 66402 60136 66404 60156
rect 66404 60136 66456 60156
rect 66456 60136 66458 60156
rect 99706 60020 99762 60056
rect 99706 60000 99708 60020
rect 99708 60000 99760 60020
rect 99760 60000 99762 60020
rect 66310 59456 66366 59512
rect 63734 58640 63790 58696
rect 62814 58096 62870 58152
rect 62630 57552 62686 57608
rect 62630 55784 62686 55840
rect 100626 59048 100682 59104
rect 66402 58912 66458 58968
rect 100626 58660 100682 58696
rect 100626 58640 100628 58660
rect 100628 58640 100680 58660
rect 100680 58640 100682 58660
rect 102466 60136 102522 60192
rect 102374 58368 102430 58424
rect 65022 58232 65078 58288
rect 63550 57008 63606 57064
rect 100626 57824 100682 57880
rect 66402 57688 66458 57744
rect 100626 57280 100682 57336
rect 66402 57164 66458 57200
rect 66402 57144 66404 57164
rect 66404 57144 66456 57164
rect 66456 57144 66458 57164
rect 100534 57164 100590 57200
rect 100534 57144 100536 57164
rect 100536 57144 100588 57164
rect 100588 57144 100590 57164
rect 66310 56464 66366 56520
rect 62906 56328 62962 56384
rect 62814 55240 62870 55296
rect 62722 54696 62778 54752
rect 135034 62312 135090 62368
rect 136874 65460 136930 65496
rect 136874 65440 136876 65460
rect 136876 65440 136928 65460
rect 136928 65440 136930 65460
rect 136874 64488 136930 64544
rect 136966 64116 136968 64136
rect 136968 64116 137020 64136
rect 137020 64116 137022 64136
rect 136966 64080 137022 64116
rect 177354 73600 177410 73656
rect 178366 74824 178422 74880
rect 179654 76592 179710 76648
rect 180482 78904 180538 78960
rect 180390 74280 180446 74336
rect 180298 71968 180354 72024
rect 189314 69112 189370 69168
rect 190234 69112 190290 69168
rect 190418 69112 190474 69168
rect 190142 68976 190198 69032
rect 191338 69248 191394 69304
rect 191430 68976 191486 69032
rect 191982 69112 192038 69168
rect 193086 69248 193142 69304
rect 204494 77544 204550 77600
rect 201090 77000 201146 77056
rect 201090 69384 201146 69440
rect 202194 69384 202250 69440
rect 174686 67480 174742 67536
rect 174042 66936 174098 66992
rect 173950 66392 174006 66448
rect 173858 65848 173914 65904
rect 171834 65576 171890 65632
rect 169534 65168 169590 65224
rect 171650 64352 171706 64408
rect 135586 63536 135642 63592
rect 136874 63264 136930 63320
rect 136966 62740 137022 62776
rect 136966 62720 136968 62740
rect 136968 62720 137020 62740
rect 137020 62720 137022 62740
rect 171742 64080 171798 64136
rect 174134 64624 174190 64680
rect 174226 64080 174282 64136
rect 174134 63536 174190 63592
rect 172018 63400 172074 63456
rect 172662 62720 172718 62776
rect 136782 62040 136838 62096
rect 171650 62060 171706 62096
rect 171650 62040 171652 62060
rect 171652 62040 171704 62060
rect 171704 62040 171706 62060
rect 135402 61768 135458 61824
rect 134482 60680 134538 60736
rect 134850 60136 134906 60192
rect 102742 59456 102798 59512
rect 102650 58912 102706 58968
rect 134390 58912 134446 58968
rect 102558 57824 102614 57880
rect 102466 57280 102522 57336
rect 100626 56056 100682 56112
rect 102374 56056 102430 56112
rect 66402 55940 66458 55976
rect 66402 55920 66404 55940
rect 66404 55920 66456 55940
rect 66456 55920 66458 55940
rect 100902 55804 100958 55840
rect 100902 55784 100904 55804
rect 100904 55784 100956 55804
rect 100956 55784 100958 55804
rect 30522 53472 30578 53528
rect 63274 53472 63330 53528
rect 66310 55240 66366 55296
rect 100626 54852 100682 54888
rect 100626 54832 100628 54852
rect 100628 54832 100680 54852
rect 100680 54832 100682 54852
rect 66402 54716 66458 54752
rect 66402 54696 66404 54716
rect 66404 54696 66456 54716
rect 66456 54696 66458 54716
rect 100810 54580 100866 54616
rect 100810 54560 100812 54580
rect 100812 54560 100864 54580
rect 100864 54560 100866 54580
rect 102466 55512 102522 55568
rect 135310 61224 135366 61280
rect 136874 61360 136930 61416
rect 172662 61380 172718 61416
rect 172662 61360 172664 61380
rect 172664 61360 172716 61380
rect 172716 61360 172718 61380
rect 174226 62992 174282 63048
rect 173858 61224 173914 61280
rect 136782 60816 136838 60872
rect 172202 60816 172258 60872
rect 135218 59456 135274 59512
rect 134482 58368 134538 58424
rect 135034 57280 135090 57336
rect 102650 56600 102706 56656
rect 136966 60272 137022 60328
rect 136874 60000 136930 60056
rect 172662 60272 172718 60328
rect 172662 59864 172718 59920
rect 136782 59048 136838 59104
rect 172662 59048 172718 59104
rect 136874 58640 136930 58696
rect 172662 58660 172718 58696
rect 172662 58640 172664 58660
rect 172664 58640 172716 58660
rect 172716 58640 172718 58660
rect 174318 62312 174374 62368
rect 174134 61768 174190 61824
rect 174134 60680 174190 60736
rect 174042 60136 174098 60192
rect 173950 59456 174006 59512
rect 174042 58912 174098 58968
rect 135402 57824 135458 57880
rect 136782 57824 136838 57880
rect 172110 57824 172166 57880
rect 173766 57824 173822 57880
rect 135218 56600 135274 56656
rect 134574 56056 134630 56112
rect 102558 54968 102614 55024
rect 102374 54424 102430 54480
rect 63550 54152 63606 54208
rect 66310 54152 66366 54208
rect 100626 53608 100682 53664
rect 66402 53472 66458 53528
rect 102466 53200 102522 53256
rect 100626 53084 100682 53120
rect 100626 53064 100628 53084
rect 100628 53064 100680 53084
rect 100680 53064 100682 53084
rect 63458 52928 63514 52984
rect 63366 52384 63422 52440
rect 62814 51296 62870 51352
rect 62722 49528 62778 49584
rect 65666 52928 65722 52984
rect 63734 51840 63790 51896
rect 100626 52384 100682 52440
rect 66402 52248 66458 52304
rect 100626 51840 100682 51896
rect 66402 51724 66458 51760
rect 66402 51704 66404 51724
rect 66404 51704 66456 51724
rect 66456 51704 66458 51724
rect 100534 51704 100590 51760
rect 102650 53744 102706 53800
rect 102558 52656 102614 52712
rect 102374 51568 102430 51624
rect 66402 51160 66458 51216
rect 63734 50616 63790 50672
rect 100626 50616 100682 50672
rect 62906 50072 62962 50128
rect 66402 50500 66458 50536
rect 66402 50480 66404 50500
rect 66404 50480 66456 50500
rect 66456 50480 66458 50500
rect 100626 50364 100682 50400
rect 100626 50344 100628 50364
rect 100628 50344 100680 50364
rect 100680 50344 100682 50364
rect 102466 50344 102522 50400
rect 65482 49936 65538 49992
rect 63826 48984 63882 49040
rect 100626 49392 100682 49448
rect 66402 49256 66458 49312
rect 62814 48440 62870 48496
rect 62722 46672 62778 46728
rect 100626 49004 100682 49040
rect 100626 48984 100628 49004
rect 100628 48984 100680 49004
rect 100680 48984 100682 49004
rect 135310 55512 135366 55568
rect 136874 57280 136930 57336
rect 136966 57180 136968 57200
rect 136968 57180 137020 57200
rect 137020 57180 137022 57200
rect 136966 57144 137022 57180
rect 172662 57416 172718 57472
rect 172570 57280 172626 57336
rect 136782 56056 136838 56112
rect 172662 56076 172718 56112
rect 172662 56056 172664 56076
rect 172664 56056 172716 56076
rect 172716 56056 172718 56076
rect 136874 55804 136930 55840
rect 136874 55784 136876 55804
rect 136876 55784 136928 55804
rect 136928 55784 136930 55804
rect 172662 55784 172718 55840
rect 135402 54968 135458 55024
rect 136782 54832 136838 54888
rect 171742 54832 171798 54888
rect 135034 54424 135090 54480
rect 137150 54580 137206 54616
rect 137150 54560 137152 54580
rect 137152 54560 137204 54580
rect 137204 54560 137206 54580
rect 172846 54424 172902 54480
rect 134298 53744 134354 53800
rect 136782 53608 136838 53664
rect 172570 53608 172626 53664
rect 135126 53200 135182 53256
rect 134206 52656 134262 52712
rect 102742 52112 102798 52168
rect 135034 52112 135090 52168
rect 136874 53064 136930 53120
rect 172662 53084 172718 53120
rect 172662 53064 172664 53084
rect 172664 53064 172716 53084
rect 172716 53064 172718 53084
rect 174134 58368 174190 58424
rect 174042 57280 174098 57336
rect 173858 56600 173914 56656
rect 174042 56328 174098 56384
rect 173950 55512 174006 55568
rect 173766 54968 173822 55024
rect 174042 54424 174098 54480
rect 174134 53744 174190 53800
rect 174226 53200 174282 53256
rect 136690 52384 136746 52440
rect 172018 52384 172074 52440
rect 102650 50888 102706 50944
rect 102558 49800 102614 49856
rect 135034 50344 135090 50400
rect 135402 51568 135458 51624
rect 136782 51840 136838 51896
rect 136874 51704 136930 51760
rect 172662 51860 172718 51896
rect 172662 51840 172664 51860
rect 172664 51840 172716 51860
rect 172716 51840 172718 51860
rect 172662 51724 172718 51760
rect 172662 51704 172664 51724
rect 172664 51704 172716 51724
rect 172716 51704 172718 51724
rect 135402 50888 135458 50944
rect 136782 50616 136838 50672
rect 171650 50636 171706 50672
rect 171650 50616 171652 50636
rect 171652 50616 171704 50636
rect 171704 50616 171706 50636
rect 135310 49800 135366 49856
rect 102650 49256 102706 49312
rect 134850 49256 134906 49312
rect 66402 48712 66458 48768
rect 102374 48712 102430 48768
rect 64930 48168 64986 48224
rect 63734 47760 63790 47816
rect 62906 47216 62962 47272
rect 100626 48304 100682 48360
rect 102466 48032 102522 48088
rect 65022 47760 65078 47816
rect 66402 47760 66458 47816
rect 100626 47644 100682 47680
rect 100626 47624 100628 47644
rect 100628 47624 100680 47644
rect 100680 47624 100682 47644
rect 66402 47508 66458 47544
rect 66402 47488 66404 47508
rect 66404 47488 66456 47508
rect 66456 47488 66458 47508
rect 100626 47508 100682 47544
rect 100626 47488 100628 47508
rect 100628 47488 100680 47508
rect 100680 47488 100682 47508
rect 66402 46944 66458 47000
rect 102558 47488 102614 47544
rect 100626 46400 100682 46456
rect 102374 46400 102430 46456
rect 62906 46128 62962 46184
rect 62814 45584 62870 45640
rect 65298 46264 65354 46320
rect 63734 44904 63790 44960
rect 62814 44360 62870 44416
rect 100902 46148 100958 46184
rect 100902 46128 100904 46148
rect 100904 46128 100956 46148
rect 100956 46128 100958 46148
rect 66402 45720 66458 45776
rect 65666 45176 65722 45232
rect 100534 45312 100590 45368
rect 99982 45040 100038 45096
rect 136874 50344 136930 50400
rect 172662 50208 172718 50264
rect 136874 49392 136930 49448
rect 171834 49392 171890 49448
rect 172662 49004 172718 49040
rect 172662 48984 172664 49004
rect 172664 48984 172716 49004
rect 172716 48984 172718 49004
rect 136782 48848 136838 48904
rect 174134 52656 174190 52712
rect 174042 52112 174098 52168
rect 173858 51568 173914 51624
rect 174042 50888 174098 50944
rect 173950 50344 174006 50400
rect 173766 49800 173822 49856
rect 174042 49256 174098 49312
rect 135402 48712 135458 48768
rect 136690 48304 136746 48360
rect 172110 48304 172166 48360
rect 135310 48032 135366 48088
rect 134758 47488 134814 47544
rect 102650 46944 102706 47000
rect 135310 46944 135366 47000
rect 134850 46400 134906 46456
rect 102466 45856 102522 45912
rect 136782 47624 136838 47680
rect 172662 47896 172718 47952
rect 172570 47624 172626 47680
rect 136874 47508 136930 47544
rect 174134 48712 174190 48768
rect 174042 48032 174098 48088
rect 136874 47488 136876 47508
rect 136876 47488 136928 47508
rect 136928 47488 136930 47508
rect 136782 46400 136838 46456
rect 172662 46420 172718 46456
rect 172662 46400 172664 46420
rect 172664 46400 172716 46420
rect 172716 46400 172718 46420
rect 137518 46128 137574 46184
rect 172662 46128 172718 46184
rect 135402 45856 135458 45912
rect 136690 45312 136746 45368
rect 102374 44632 102430 44688
rect 65298 44496 65354 44552
rect 63734 43816 63790 43872
rect 63642 43272 63698 43328
rect 63734 42728 63790 42784
rect 102558 45176 102614 45232
rect 134666 45176 134722 45232
rect 99890 44108 99946 44144
rect 99890 44088 99892 44108
rect 99892 44088 99944 44108
rect 99944 44088 99946 44108
rect 102466 44088 102522 44144
rect 66402 43952 66458 44008
rect 100626 43408 100682 43464
rect 66402 43272 66458 43328
rect 135034 44668 135036 44688
rect 135036 44668 135088 44688
rect 135088 44668 135090 44688
rect 135034 44632 135090 44668
rect 136782 44904 136838 44960
rect 171834 45312 171890 45368
rect 172662 44904 172718 44960
rect 173950 47488 174006 47544
rect 174042 46944 174098 47000
rect 174226 46400 174282 46456
rect 173858 45856 173914 45912
rect 174042 45176 174098 45232
rect 174134 44668 174136 44688
rect 174136 44668 174188 44688
rect 174188 44668 174190 44688
rect 174134 44632 174190 44668
rect 135402 44088 135458 44144
rect 136782 44088 136838 44144
rect 171834 44088 171890 44144
rect 102558 43544 102614 43600
rect 135034 43544 135090 43600
rect 102282 43000 102338 43056
rect 100626 42864 100682 42920
rect 66402 42728 66458 42784
rect 65298 42184 65354 42240
rect 63918 42048 63974 42104
rect 63826 41504 63882 41560
rect 63734 40960 63790 41016
rect 100626 42320 100682 42376
rect 102374 42320 102430 42376
rect 100626 42068 100682 42104
rect 100626 42048 100628 42068
rect 100628 42048 100680 42068
rect 100680 42048 100682 42068
rect 62814 40416 62870 40472
rect 66402 40416 66458 40472
rect 62814 39464 62870 39520
rect 66218 32664 66274 32720
rect 66310 24640 66366 24696
rect 13318 19608 13374 19664
rect 174686 44088 174742 44144
rect 172662 43544 172718 43600
rect 136874 43408 136930 43464
rect 174502 43544 174558 43600
rect 135402 43036 135404 43056
rect 135404 43036 135456 43056
rect 135456 43036 135458 43056
rect 135402 43000 135458 43036
rect 174042 43000 174098 43056
rect 136690 42864 136746 42920
rect 172570 42864 172626 42920
rect 134942 42320 134998 42376
rect 102558 41776 102614 41832
rect 135310 41812 135312 41832
rect 135312 41812 135364 41832
rect 135364 41812 135366 41832
rect 135310 41776 135366 41812
rect 102466 41232 102522 41288
rect 136874 42320 136930 42376
rect 172386 42340 172442 42376
rect 172386 42320 172388 42340
rect 172388 42320 172440 42340
rect 172440 42320 172442 42340
rect 136782 42048 136838 42104
rect 174226 42320 174282 42376
rect 172662 42068 172718 42104
rect 172662 42048 172664 42068
rect 172664 42048 172716 42068
rect 172716 42048 172718 42068
rect 135402 41232 135458 41288
rect 102374 40688 102430 40744
rect 134850 40688 134906 40744
rect 94002 40416 94058 40472
rect 102374 40144 102430 40200
rect 109642 40008 109698 40064
rect 134482 39600 134538 39656
rect 136874 33344 136930 33400
rect 138162 39736 138218 39792
rect 138070 25048 138126 25104
rect 173950 41232 174006 41288
rect 174134 41776 174190 41832
rect 174042 40688 174098 40744
rect 181402 40008 181458 40064
rect 166038 39736 166094 39792
rect 174134 39464 174190 39520
rect 222894 139696 222950 139752
rect 222710 115896 222766 115952
rect 224458 105696 224514 105752
rect 223538 96312 223594 96368
rect 223538 92096 223594 92152
rect 223538 85160 223594 85216
rect 223538 75232 223594 75288
rect 223078 68296 223134 68352
rect 222526 44496 222582 44552
rect 222710 20696 222766 20752
rect 138162 17024 138218 17080
rect 66402 16752 66458 16808
<< metal3 >>
rect 98229 238762 98295 238765
rect 169989 238762 170055 238765
rect 96652 238760 98295 238762
rect 96652 238704 98234 238760
rect 98290 238704 98295 238760
rect 96652 238702 98295 238704
rect 168780 238760 170055 238762
rect 168780 238704 169994 238760
rect 170050 238704 170055 238760
rect 168780 238702 170055 238704
rect 98229 238699 98295 238702
rect 169989 238699 170055 238702
rect 9896 235906 10376 235936
rect 9896 235846 10570 235906
rect 9896 235816 10376 235846
rect 10510 235226 10570 235846
rect 20622 235226 20628 235228
rect 10510 235166 20628 235226
rect 20622 235164 20628 235166
rect 20692 235164 20698 235228
rect 223073 234954 223139 234957
rect 227416 234954 227896 234984
rect 223073 234952 227896 234954
rect 223073 234896 223078 234952
rect 223134 234896 227896 234952
rect 223073 234894 227896 234896
rect 223073 234891 223139 234894
rect 227416 234864 227896 234894
rect 98321 230738 98387 230741
rect 96652 230736 98387 230738
rect 96652 230680 98326 230736
rect 98382 230680 98387 230736
rect 96652 230678 98387 230680
rect 98321 230675 98387 230678
rect 168566 230197 168626 230708
rect 168517 230192 168626 230197
rect 168517 230136 168522 230192
rect 168578 230136 168626 230192
rect 168517 230134 168626 230136
rect 168517 230131 168583 230134
rect 98413 222850 98479 222853
rect 170081 222850 170147 222853
rect 96652 222848 98479 222850
rect 96652 222792 98418 222848
rect 98474 222792 98479 222848
rect 96652 222790 98479 222792
rect 168780 222848 170147 222850
rect 168780 222792 170086 222848
rect 170142 222792 170147 222848
rect 168780 222790 170147 222792
rect 98413 222787 98479 222790
rect 170081 222787 170147 222790
rect 37918 217212 37924 217276
rect 37988 217274 37994 217276
rect 55817 217274 55883 217277
rect 37988 217272 55883 217274
rect 37988 217216 55822 217272
rect 55878 217216 55883 217272
rect 37988 217214 55883 217216
rect 37988 217212 37994 217214
rect 55817 217211 55883 217214
rect 151037 215914 151103 215917
rect 204254 215914 204260 215916
rect 151037 215912 204260 215914
rect 151037 215856 151042 215912
rect 151098 215856 204260 215912
rect 151037 215854 204260 215856
rect 151037 215851 151103 215854
rect 204254 215852 204260 215854
rect 204324 215852 204330 215916
rect 174221 215778 174287 215781
rect 174221 215776 177090 215778
rect 174221 215720 174226 215776
rect 174282 215720 177090 215776
rect 174221 215718 177090 215720
rect 174221 215715 174287 215718
rect 135397 215642 135463 215645
rect 132686 215640 135463 215642
rect 132686 215584 135402 215640
rect 135458 215584 135463 215640
rect 132686 215582 135463 215584
rect 132686 215408 132746 215582
rect 135397 215579 135463 215582
rect 177030 215408 177090 215718
rect 62533 215370 62599 215373
rect 60588 215368 62599 215370
rect 60588 215312 62538 215368
rect 62594 215312 62599 215368
rect 60588 215310 62599 215312
rect 62533 215307 62599 215310
rect 102369 215370 102435 215373
rect 102369 215368 104932 215370
rect 102369 215312 102374 215368
rect 102430 215312 104932 215368
rect 102369 215310 104932 215312
rect 102369 215307 102435 215310
rect 62625 214690 62691 214693
rect 60588 214688 62691 214690
rect 60588 214632 62630 214688
rect 62686 214632 62691 214688
rect 60588 214630 62691 214632
rect 62625 214627 62691 214630
rect 102369 214690 102435 214693
rect 135397 214690 135463 214693
rect 102369 214688 104932 214690
rect 102369 214632 102374 214688
rect 102430 214632 104932 214688
rect 102369 214630 104932 214632
rect 132716 214688 135463 214690
rect 132716 214632 135402 214688
rect 135458 214632 135463 214688
rect 132716 214630 135463 214632
rect 102369 214627 102435 214630
rect 135397 214627 135463 214630
rect 174037 214690 174103 214693
rect 174037 214688 177060 214690
rect 174037 214632 174042 214688
rect 174098 214632 177060 214688
rect 174037 214630 177060 214632
rect 174037 214627 174103 214630
rect 9896 214282 10376 214312
rect 10461 214282 10527 214285
rect 9896 214280 10527 214282
rect 9896 214224 10466 214280
rect 10522 214224 10527 214280
rect 9896 214222 10527 214224
rect 9896 214192 10376 214222
rect 10461 214219 10527 214222
rect 63637 214010 63703 214013
rect 60588 214008 63703 214010
rect 60588 213952 63642 214008
rect 63698 213952 63703 214008
rect 60588 213950 63703 213952
rect 63637 213947 63703 213950
rect 102369 214010 102435 214013
rect 135029 214010 135095 214013
rect 171829 214010 171895 214013
rect 102369 214008 104932 214010
rect 102369 213952 102374 214008
rect 102430 213952 104932 214008
rect 102369 213950 104932 213952
rect 132716 214008 135095 214010
rect 132716 213952 135034 214008
rect 135090 213952 135095 214008
rect 132716 213950 135095 213952
rect 102369 213947 102435 213950
rect 135029 213947 135095 213950
rect 169670 214008 171895 214010
rect 169670 213952 171834 214008
rect 171890 213952 171895 214008
rect 169670 213950 171895 213952
rect 65017 213602 65083 213605
rect 65017 213600 67978 213602
rect 65017 213544 65022 213600
rect 65078 213544 67978 213600
rect 65017 213542 67978 213544
rect 65017 213539 65083 213542
rect 67918 213436 67978 213542
rect 100989 213466 101055 213469
rect 97756 213464 101055 213466
rect 97756 213408 100994 213464
rect 101050 213408 101055 213464
rect 97756 213406 101055 213408
rect 100989 213403 101055 213406
rect 136777 213466 136843 213469
rect 136777 213464 140076 213466
rect 136777 213408 136782 213464
rect 136838 213408 140076 213464
rect 169670 213436 169730 213950
rect 171829 213947 171895 213950
rect 174221 214010 174287 214013
rect 174221 214008 177060 214010
rect 174221 213952 174226 214008
rect 174282 213952 177060 214008
rect 174221 213950 177060 213952
rect 174221 213947 174287 213950
rect 136777 213406 140076 213408
rect 136777 213403 136843 213406
rect 62533 213330 62599 213333
rect 60588 213328 62599 213330
rect 60588 213272 62538 213328
rect 62594 213272 62599 213328
rect 60588 213270 62599 213272
rect 62533 213267 62599 213270
rect 102461 213330 102527 213333
rect 135397 213330 135463 213333
rect 102461 213328 104932 213330
rect 102461 213272 102466 213328
rect 102522 213272 104932 213328
rect 102461 213270 104932 213272
rect 132716 213328 135463 213330
rect 132716 213272 135402 213328
rect 135458 213272 135463 213328
rect 132716 213270 135463 213272
rect 102461 213267 102527 213270
rect 135397 213267 135463 213270
rect 174037 213330 174103 213333
rect 174037 213328 177060 213330
rect 174037 213272 174042 213328
rect 174098 213272 177060 213328
rect 174037 213270 177060 213272
rect 174037 213267 174103 213270
rect 10461 213194 10527 213197
rect 20806 213194 20812 213196
rect 10461 213192 20812 213194
rect 10461 213136 10466 213192
rect 10522 213136 20812 213192
rect 10461 213134 20812 213136
rect 10461 213131 10527 213134
rect 20806 213132 20812 213134
rect 20876 213132 20882 213196
rect 172657 213058 172723 213061
rect 169670 213056 172723 213058
rect 169670 213000 172662 213056
rect 172718 213000 172723 213056
rect 169670 212998 172723 213000
rect 66213 212922 66279 212925
rect 100989 212922 101055 212925
rect 66213 212920 67948 212922
rect 66213 212864 66218 212920
rect 66274 212864 67948 212920
rect 66213 212862 67948 212864
rect 97756 212920 101055 212922
rect 97756 212864 100994 212920
rect 101050 212864 101055 212920
rect 97756 212862 101055 212864
rect 66213 212859 66279 212862
rect 100989 212859 101055 212862
rect 136777 212922 136843 212925
rect 136777 212920 140076 212922
rect 136777 212864 136782 212920
rect 136838 212864 140076 212920
rect 169670 212892 169730 212998
rect 172657 212995 172723 212998
rect 136777 212862 140076 212864
rect 136777 212859 136843 212862
rect 62349 212650 62415 212653
rect 60588 212648 62415 212650
rect 60588 212592 62354 212648
rect 62410 212592 62415 212648
rect 60588 212590 62415 212592
rect 62349 212587 62415 212590
rect 102369 212650 102435 212653
rect 134661 212650 134727 212653
rect 171737 212650 171803 212653
rect 102369 212648 104932 212650
rect 102369 212592 102374 212648
rect 102430 212592 104932 212648
rect 102369 212590 104932 212592
rect 132716 212648 134727 212650
rect 132716 212592 134666 212648
rect 134722 212592 134727 212648
rect 132716 212590 134727 212592
rect 102369 212587 102435 212590
rect 134661 212587 134727 212590
rect 169670 212648 171803 212650
rect 169670 212592 171742 212648
rect 171798 212592 171803 212648
rect 169670 212590 171803 212592
rect 65017 212242 65083 212245
rect 100529 212242 100595 212245
rect 65017 212240 67948 212242
rect 65017 212184 65022 212240
rect 65078 212184 67948 212240
rect 65017 212182 67948 212184
rect 97756 212240 100595 212242
rect 97756 212184 100534 212240
rect 100590 212184 100595 212240
rect 97756 212182 100595 212184
rect 65017 212179 65083 212182
rect 100529 212179 100595 212182
rect 136869 212242 136935 212245
rect 136869 212240 140076 212242
rect 136869 212184 136874 212240
rect 136930 212184 140076 212240
rect 169670 212212 169730 212590
rect 171737 212587 171803 212590
rect 174221 212650 174287 212653
rect 174221 212648 177060 212650
rect 174221 212592 174226 212648
rect 174282 212592 177060 212648
rect 174221 212590 177060 212592
rect 174221 212587 174287 212590
rect 136869 212182 140076 212184
rect 136869 212179 136935 212182
rect 62625 211970 62691 211973
rect 60588 211968 62691 211970
rect 60588 211912 62630 211968
rect 62686 211912 62691 211968
rect 60588 211910 62691 211912
rect 62625 211907 62691 211910
rect 102369 211970 102435 211973
rect 134293 211970 134359 211973
rect 102369 211968 104932 211970
rect 102369 211912 102374 211968
rect 102430 211912 104932 211968
rect 102369 211910 104932 211912
rect 132716 211968 134359 211970
rect 132716 211912 134298 211968
rect 134354 211912 134359 211968
rect 132716 211910 134359 211912
rect 102369 211907 102435 211910
rect 134293 211907 134359 211910
rect 174037 211970 174103 211973
rect 174037 211968 177060 211970
rect 174037 211912 174042 211968
rect 174098 211912 177060 211968
rect 174037 211910 177060 211912
rect 174037 211907 174103 211910
rect 66397 211698 66463 211701
rect 101081 211698 101147 211701
rect 66397 211696 67948 211698
rect 66397 211640 66402 211696
rect 66458 211640 67948 211696
rect 66397 211638 67948 211640
rect 97756 211696 101147 211698
rect 97756 211640 101086 211696
rect 101142 211640 101147 211696
rect 97756 211638 101147 211640
rect 66397 211635 66463 211638
rect 101081 211635 101147 211638
rect 136961 211698 137027 211701
rect 136961 211696 140076 211698
rect 136961 211640 136966 211696
rect 137022 211640 140076 211696
rect 136961 211638 140076 211640
rect 136961 211635 137027 211638
rect 169854 211562 169914 211668
rect 204806 211636 204812 211700
rect 204876 211636 204882 211700
rect 172657 211562 172723 211565
rect 169854 211560 172723 211562
rect 169854 211504 172662 211560
rect 172718 211504 172723 211560
rect 169854 211502 172723 211504
rect 172657 211499 172723 211502
rect 172565 211426 172631 211429
rect 169670 211424 172631 211426
rect 169670 211368 172570 211424
rect 172626 211368 172631 211424
rect 169670 211366 172631 211368
rect 62625 211290 62691 211293
rect 60588 211288 62691 211290
rect 60588 211232 62630 211288
rect 62686 211232 62691 211288
rect 60588 211230 62691 211232
rect 62625 211227 62691 211230
rect 65017 211154 65083 211157
rect 100989 211154 101055 211157
rect 65017 211152 67948 211154
rect 65017 211096 65022 211152
rect 65078 211096 67948 211152
rect 65017 211094 67948 211096
rect 97756 211152 101055 211154
rect 97756 211096 100994 211152
rect 101050 211096 101055 211152
rect 97756 211094 101055 211096
rect 65017 211091 65083 211094
rect 100989 211091 101055 211094
rect 104902 210882 104962 211260
rect 97726 210822 104962 210882
rect 132686 210882 132746 211260
rect 136869 211154 136935 211157
rect 136869 211152 140076 211154
rect 136869 211096 136874 211152
rect 136930 211096 140076 211152
rect 169670 211124 169730 211366
rect 172565 211363 172631 211366
rect 174129 211290 174195 211293
rect 174129 211288 177060 211290
rect 174129 211232 174134 211288
rect 174190 211232 177060 211288
rect 174129 211230 177060 211232
rect 174129 211227 174195 211230
rect 204814 211124 204874 211636
rect 223533 211154 223599 211157
rect 227416 211154 227896 211184
rect 223533 211152 227896 211154
rect 136869 211094 140076 211096
rect 223533 211096 223538 211152
rect 223594 211096 227896 211152
rect 223533 211094 227896 211096
rect 136869 211091 136935 211094
rect 223533 211091 223599 211094
rect 227416 211064 227896 211094
rect 132686 210822 140106 210882
rect 64925 210746 64991 210749
rect 66397 210746 66463 210749
rect 64925 210744 66463 210746
rect 64925 210688 64930 210744
rect 64986 210688 66402 210744
rect 66458 210688 66463 210744
rect 64925 210686 66463 210688
rect 64925 210683 64991 210686
rect 66397 210683 66463 210686
rect 62625 210610 62691 210613
rect 60588 210608 62691 210610
rect 60588 210552 62630 210608
rect 62686 210552 62691 210608
rect 60588 210550 62691 210552
rect 62625 210547 62691 210550
rect 65477 210474 65543 210477
rect 65477 210472 67948 210474
rect 65477 210416 65482 210472
rect 65538 210416 67948 210472
rect 97726 210444 97786 210822
rect 65477 210414 67948 210416
rect 65477 210411 65543 210414
rect 104902 210338 104962 210580
rect 100854 210278 104962 210338
rect 132686 210338 132746 210580
rect 140046 210444 140106 210822
rect 171829 210746 171895 210749
rect 169670 210744 171895 210746
rect 169670 210688 171834 210744
rect 171890 210688 171895 210744
rect 169670 210686 171895 210688
rect 169670 210444 169730 210686
rect 171829 210683 171895 210686
rect 177030 210338 177090 210580
rect 132686 210278 136978 210338
rect 100854 210202 100914 210278
rect 97726 210142 100914 210202
rect 136918 210202 136978 210278
rect 172798 210278 177090 210338
rect 172798 210202 172858 210278
rect 136918 210142 140106 210202
rect 62625 209930 62691 209933
rect 60588 209928 62691 209930
rect 60588 209872 62630 209928
rect 62686 209872 62691 209928
rect 97726 209900 97786 210142
rect 140046 209900 140106 210142
rect 169670 210142 172858 210202
rect 169670 209900 169730 210142
rect 174129 209930 174195 209933
rect 174129 209928 177060 209930
rect 60588 209870 62691 209872
rect 62625 209867 62691 209870
rect 65017 209522 65083 209525
rect 67918 209522 67978 209900
rect 104902 209522 104962 209900
rect 132686 209658 132746 209900
rect 174129 209872 174134 209928
rect 174190 209872 177060 209928
rect 174129 209870 177060 209872
rect 174129 209867 174195 209870
rect 132686 209598 140106 209658
rect 65017 209520 67978 209522
rect 65017 209464 65022 209520
rect 65078 209464 67978 209520
rect 65017 209462 67978 209464
rect 97726 209462 104962 209522
rect 65017 209459 65083 209462
rect 62717 209250 62783 209253
rect 60588 209248 62783 209250
rect 60588 209192 62722 209248
rect 62778 209192 62783 209248
rect 60588 209190 62783 209192
rect 62717 209187 62783 209190
rect 65477 209250 65543 209253
rect 65477 209248 67948 209250
rect 65477 209192 65482 209248
rect 65538 209192 67948 209248
rect 97726 209220 97786 209462
rect 135305 209250 135371 209253
rect 132716 209248 135371 209250
rect 65477 209190 67948 209192
rect 65477 209187 65543 209190
rect 104902 208978 104962 209220
rect 132716 209192 135310 209248
rect 135366 209192 135371 209248
rect 140046 209220 140106 209598
rect 171921 209386 171987 209389
rect 169670 209384 171987 209386
rect 169670 209328 171926 209384
rect 171982 209328 171987 209384
rect 169670 209326 171987 209328
rect 169670 209220 169730 209326
rect 171921 209323 171987 209326
rect 174589 209250 174655 209253
rect 174589 209248 177060 209250
rect 132716 209190 135371 209192
rect 135305 209187 135371 209190
rect 174589 209192 174594 209248
rect 174650 209192 177060 209248
rect 174589 209190 177060 209192
rect 174589 209187 174655 209190
rect 101038 208918 104962 208978
rect 101038 208842 101098 208918
rect 171461 208842 171527 208845
rect 97726 208782 101098 208842
rect 169670 208840 171527 208842
rect 169670 208784 171466 208840
rect 171522 208784 171527 208840
rect 169670 208782 171527 208784
rect 65017 208706 65083 208709
rect 65017 208704 67948 208706
rect 65017 208648 65022 208704
rect 65078 208648 67948 208704
rect 97726 208676 97786 208782
rect 137697 208706 137763 208709
rect 137697 208704 140076 208706
rect 65017 208646 67948 208648
rect 137697 208648 137702 208704
rect 137758 208648 140076 208704
rect 169670 208676 169730 208782
rect 171461 208779 171527 208782
rect 137697 208646 140076 208648
rect 65017 208643 65083 208646
rect 137697 208643 137763 208646
rect 62533 208570 62599 208573
rect 60588 208568 62599 208570
rect 60588 208512 62538 208568
rect 62594 208512 62599 208568
rect 60588 208510 62599 208512
rect 62533 208507 62599 208510
rect 65661 208162 65727 208165
rect 104902 208162 104962 208540
rect 65661 208160 67948 208162
rect 65661 208104 65666 208160
rect 65722 208104 67948 208160
rect 65661 208102 67948 208104
rect 97756 208102 104962 208162
rect 132686 208162 132746 208540
rect 177030 208298 177090 208540
rect 169670 208238 177090 208298
rect 132686 208102 140076 208162
rect 169670 208132 169730 208238
rect 65661 208099 65727 208102
rect 135397 207890 135463 207893
rect 132716 207888 135463 207890
rect 60558 207618 60618 207860
rect 104902 207618 104962 207860
rect 132716 207832 135402 207888
rect 135458 207832 135463 207888
rect 132716 207830 135463 207832
rect 135397 207827 135463 207830
rect 174037 207890 174103 207893
rect 174037 207888 177060 207890
rect 174037 207832 174042 207888
rect 174098 207832 177060 207888
rect 174037 207830 177060 207832
rect 174037 207827 174103 207830
rect 60558 207558 63700 207618
rect 63640 207482 63700 207558
rect 102326 207558 104962 207618
rect 102326 207482 102386 207558
rect 63640 207422 67948 207482
rect 97756 207422 102386 207482
rect 136869 207482 136935 207485
rect 136869 207480 140076 207482
rect 136869 207424 136874 207480
rect 136930 207424 140076 207480
rect 136869 207422 140076 207424
rect 136869 207419 136935 207422
rect 169854 207346 169914 207452
rect 172565 207346 172631 207349
rect 169854 207344 172631 207346
rect 169854 207288 172570 207344
rect 172626 207288 172631 207344
rect 169854 207286 172631 207288
rect 172565 207283 172631 207286
rect 62625 207210 62691 207213
rect 60588 207208 62691 207210
rect 60588 207152 62630 207208
rect 62686 207152 62691 207208
rect 60588 207150 62691 207152
rect 62625 207147 62691 207150
rect 65661 206938 65727 206941
rect 104902 206938 104962 207180
rect 132716 207150 140106 207210
rect 65661 206936 67948 206938
rect 65661 206880 65666 206936
rect 65722 206880 67948 206936
rect 65661 206878 67948 206880
rect 97756 206878 104962 206938
rect 140046 206908 140106 207150
rect 65661 206875 65727 206878
rect 169854 206802 169914 206908
rect 177030 206802 177090 207180
rect 169854 206742 177090 206802
rect 60558 206258 60618 206500
rect 104902 206258 104962 206500
rect 132716 206470 140106 206530
rect 60558 206198 67948 206258
rect 97756 206198 104962 206258
rect 140046 206228 140106 206470
rect 169670 206470 177060 206530
rect 169670 206228 169730 206470
rect 60558 205714 60618 205820
rect 104902 205714 104962 205820
rect 132716 205790 140106 205850
rect 60558 205654 67948 205714
rect 97756 205654 104962 205714
rect 140046 205684 140106 205790
rect 169854 205578 169914 205684
rect 177030 205578 177090 205820
rect 169854 205518 177090 205578
rect 169670 205246 176538 205306
rect 60588 205110 67948 205170
rect 97756 205110 104932 205170
rect 132716 205110 140076 205170
rect 169670 205140 169730 205246
rect 176478 205238 176538 205246
rect 176478 205178 177060 205238
rect 60588 204430 67948 204490
rect 97756 204430 104932 204490
rect 132716 204430 140076 204490
rect 169854 204354 169914 204460
rect 177030 204354 177090 204460
rect 169854 204294 177090 204354
rect 169670 204022 177090 204082
rect 169670 203916 169730 204022
rect 60558 203538 60618 203780
rect 67918 203538 67978 203916
rect 177030 203848 177090 204022
rect 97726 203810 97786 203848
rect 140046 203810 140106 203848
rect 97726 203750 104932 203810
rect 132716 203750 140106 203810
rect 60558 203478 67978 203538
rect 60558 203206 67948 203266
rect 60558 203100 60618 203206
rect 97726 203130 97786 203168
rect 140046 203130 140106 203168
rect 97726 203070 104932 203130
rect 132716 203070 140106 203130
rect 169854 202994 169914 203236
rect 177030 202994 177090 203100
rect 169854 202934 177090 202994
rect 60558 202662 67948 202722
rect 60558 202420 60618 202662
rect 97726 202450 97786 202624
rect 140046 202450 140106 202624
rect 169854 202586 169914 202692
rect 169854 202526 176538 202586
rect 176478 202518 176538 202526
rect 176478 202458 177060 202518
rect 97726 202390 104932 202450
rect 132716 202390 140106 202450
rect 172657 202314 172723 202317
rect 169670 202312 172723 202314
rect 169670 202256 172662 202312
rect 172718 202256 172723 202312
rect 169670 202254 172723 202256
rect 65017 202178 65083 202181
rect 65017 202176 67948 202178
rect 65017 202120 65022 202176
rect 65078 202120 67948 202176
rect 65017 202118 67948 202120
rect 97756 202118 101466 202178
rect 65017 202115 65083 202118
rect 101406 202042 101466 202118
rect 136918 202118 140076 202178
rect 169670 202148 169730 202254
rect 172657 202251 172723 202254
rect 136918 202042 136978 202118
rect 101406 201982 104962 202042
rect 62625 201770 62691 201773
rect 60588 201768 62691 201770
rect 60588 201712 62630 201768
rect 62686 201712 62691 201768
rect 104902 201740 104962 201982
rect 132686 201982 136978 202042
rect 174221 202042 174287 202045
rect 174221 202040 177090 202042
rect 174221 201984 174226 202040
rect 174282 201984 177090 202040
rect 174221 201982 177090 201984
rect 132686 201808 132746 201982
rect 174221 201979 174287 201982
rect 177030 201808 177090 201982
rect 207893 201770 207959 201773
rect 204844 201768 207959 201770
rect 60588 201710 62691 201712
rect 204844 201712 207898 201768
rect 207954 201712 207959 201768
rect 204844 201710 207959 201712
rect 62625 201707 62691 201710
rect 207893 201707 207959 201710
rect 60558 201438 67948 201498
rect 60558 201060 60618 201438
rect 97726 201090 97786 201400
rect 140046 201090 140106 201400
rect 169854 201362 169914 201468
rect 169854 201302 177090 201362
rect 177030 201128 177090 201302
rect 97726 201030 104932 201090
rect 132716 201030 140106 201090
rect 65017 200954 65083 200957
rect 65017 200952 67948 200954
rect 65017 200896 65022 200952
rect 65078 200896 67948 200952
rect 65017 200894 67948 200896
rect 65017 200891 65083 200894
rect 97726 200682 97786 200856
rect 100897 200682 100963 200685
rect 97726 200680 100963 200682
rect 97726 200624 100902 200680
rect 100958 200624 100963 200680
rect 97726 200622 100963 200624
rect 100897 200619 100963 200622
rect 136777 200682 136843 200685
rect 140046 200682 140106 200856
rect 169854 200818 169914 200924
rect 172657 200818 172723 200821
rect 169854 200816 172723 200818
rect 169854 200760 172662 200816
rect 172718 200760 172723 200816
rect 169854 200758 172723 200760
rect 172657 200755 172723 200758
rect 136777 200680 140106 200682
rect 136777 200624 136782 200680
rect 136838 200624 140106 200680
rect 136777 200622 140106 200624
rect 136777 200619 136843 200622
rect 62625 200410 62691 200413
rect 60588 200408 62691 200410
rect 60588 200352 62630 200408
rect 62686 200352 62691 200408
rect 60588 200350 62691 200352
rect 62625 200347 62691 200350
rect 102369 200410 102435 200413
rect 135397 200410 135463 200413
rect 102369 200408 104932 200410
rect 102369 200352 102374 200408
rect 102430 200352 104932 200408
rect 102369 200350 104932 200352
rect 132716 200408 135463 200410
rect 132716 200352 135402 200408
rect 135458 200352 135463 200408
rect 132716 200350 135463 200352
rect 102369 200347 102435 200350
rect 135397 200347 135463 200350
rect 174129 200410 174195 200413
rect 174129 200408 177060 200410
rect 174129 200352 174134 200408
rect 174190 200352 177060 200408
rect 174129 200350 177060 200352
rect 174129 200347 174195 200350
rect 60558 200214 67948 200274
rect 60558 199700 60618 200214
rect 97726 200002 97786 200176
rect 140046 200002 140106 200176
rect 169854 200138 169914 200244
rect 169854 200078 177090 200138
rect 97726 199942 104962 200002
rect 65017 199730 65083 199733
rect 65017 199728 67948 199730
rect 65017 199672 65022 199728
rect 65078 199672 67948 199728
rect 104902 199700 104962 199942
rect 132686 199942 140106 200002
rect 132686 199768 132746 199942
rect 177030 199768 177090 200078
rect 65017 199670 67948 199672
rect 65017 199667 65083 199670
rect 97726 199322 97786 199632
rect 136777 199458 136843 199461
rect 140046 199458 140106 199632
rect 169854 199594 169914 199700
rect 171645 199594 171711 199597
rect 169854 199592 171711 199594
rect 169854 199536 171650 199592
rect 171706 199536 171711 199592
rect 169854 199534 171711 199536
rect 171645 199531 171711 199534
rect 136777 199456 140106 199458
rect 136777 199400 136782 199456
rect 136838 199400 140106 199456
rect 136777 199398 140106 199400
rect 136777 199395 136843 199398
rect 100897 199322 100963 199325
rect 97726 199320 100963 199322
rect 97726 199264 100902 199320
rect 100958 199264 100963 199320
rect 97726 199262 100963 199264
rect 100897 199259 100963 199262
rect 62349 199050 62415 199053
rect 60588 199048 62415 199050
rect 60588 198992 62354 199048
rect 62410 198992 62415 199048
rect 60588 198990 62415 198992
rect 62349 198987 62415 198990
rect 67918 198778 67978 199156
rect 60558 198718 67978 198778
rect 97726 198778 97786 199088
rect 102369 199050 102435 199053
rect 134753 199050 134819 199053
rect 102369 199048 104932 199050
rect 102369 198992 102374 199048
rect 102430 198992 104932 199048
rect 102369 198990 104932 198992
rect 132716 199048 134819 199050
rect 132716 198992 134758 199048
rect 134814 198992 134819 199048
rect 132716 198990 134819 198992
rect 102369 198987 102435 198990
rect 134753 198987 134819 198990
rect 140046 198778 140106 199088
rect 169854 198914 169914 199156
rect 175233 199050 175299 199053
rect 175233 199048 177060 199050
rect 175233 198992 175238 199048
rect 175294 198992 177060 199048
rect 175233 198990 177060 198992
rect 175233 198987 175299 198990
rect 169854 198854 177090 198914
rect 97726 198718 104962 198778
rect 60558 198340 60618 198718
rect 65017 198506 65083 198509
rect 65017 198504 67948 198506
rect 65017 198448 65022 198504
rect 65078 198448 67948 198504
rect 65017 198446 67948 198448
rect 65017 198443 65083 198446
rect 97726 198098 97786 198408
rect 104902 198340 104962 198718
rect 132686 198718 140106 198778
rect 132686 198408 132746 198718
rect 100805 198098 100871 198101
rect 97726 198096 100871 198098
rect 97726 198040 100810 198096
rect 100866 198040 100871 198096
rect 97726 198038 100871 198040
rect 100805 198035 100871 198038
rect 136777 198098 136843 198101
rect 140046 198098 140106 198408
rect 169854 198234 169914 198476
rect 177030 198408 177090 198854
rect 172657 198234 172723 198237
rect 169854 198232 172723 198234
rect 169854 198176 172662 198232
rect 172718 198176 172723 198232
rect 169854 198174 172723 198176
rect 172657 198171 172723 198174
rect 172657 198098 172723 198101
rect 136777 198096 140106 198098
rect 136777 198040 136782 198096
rect 136838 198040 140106 198096
rect 136777 198038 140106 198040
rect 169670 198096 172723 198098
rect 169670 198040 172662 198096
rect 172718 198040 172723 198096
rect 169670 198038 172723 198040
rect 136777 198035 136843 198038
rect 65661 197962 65727 197965
rect 100897 197962 100963 197965
rect 65661 197960 67948 197962
rect 65661 197904 65666 197960
rect 65722 197904 67948 197960
rect 65661 197902 67948 197904
rect 97756 197960 100963 197962
rect 97756 197904 100902 197960
rect 100958 197904 100963 197960
rect 97756 197902 100963 197904
rect 65661 197899 65727 197902
rect 100897 197899 100963 197902
rect 136685 197962 136751 197965
rect 136685 197960 140076 197962
rect 136685 197904 136690 197960
rect 136746 197904 140076 197960
rect 169670 197932 169730 198038
rect 172657 198035 172723 198038
rect 136685 197902 140076 197904
rect 136685 197899 136751 197902
rect 62625 197690 62691 197693
rect 60588 197688 62691 197690
rect 60588 197632 62630 197688
rect 62686 197632 62691 197688
rect 60588 197630 62691 197632
rect 62625 197627 62691 197630
rect 102369 197690 102435 197693
rect 135397 197690 135463 197693
rect 102369 197688 104932 197690
rect 102369 197632 102374 197688
rect 102430 197632 104932 197688
rect 102369 197630 104932 197632
rect 132716 197688 135463 197690
rect 132716 197632 135402 197688
rect 135458 197632 135463 197688
rect 132716 197630 135463 197632
rect 102369 197627 102435 197630
rect 135397 197627 135463 197630
rect 174129 197690 174195 197693
rect 174129 197688 177060 197690
rect 174129 197632 174134 197688
rect 174190 197632 177060 197688
rect 174129 197630 177060 197632
rect 174129 197627 174195 197630
rect 174221 197554 174287 197557
rect 174221 197552 177090 197554
rect 174221 197496 174226 197552
rect 174282 197496 177090 197552
rect 174221 197494 177090 197496
rect 174221 197491 174287 197494
rect 135397 197418 135463 197421
rect 132686 197416 135463 197418
rect 132686 197360 135402 197416
rect 135458 197360 135463 197416
rect 132686 197358 135463 197360
rect 65017 197282 65083 197285
rect 65017 197280 67948 197282
rect 65017 197224 65022 197280
rect 65078 197224 67948 197280
rect 65017 197222 67948 197224
rect 65017 197219 65083 197222
rect 62533 197010 62599 197013
rect 60588 197008 62599 197010
rect 60588 196952 62538 197008
rect 62594 196952 62599 197008
rect 60588 196950 62599 196952
rect 62533 196947 62599 196950
rect 97726 196874 97786 197184
rect 132686 197048 132746 197358
rect 135397 197355 135463 197358
rect 102461 197010 102527 197013
rect 102461 197008 104932 197010
rect 102461 196952 102466 197008
rect 102522 196952 104932 197008
rect 102461 196950 104932 196952
rect 102461 196947 102527 196950
rect 100713 196874 100779 196877
rect 97726 196872 100779 196874
rect 97726 196816 100718 196872
rect 100774 196816 100779 196872
rect 97726 196814 100779 196816
rect 100713 196811 100779 196814
rect 136777 196874 136843 196877
rect 140046 196874 140106 197184
rect 136777 196872 140106 196874
rect 136777 196816 136782 196872
rect 136838 196816 140106 196872
rect 136777 196814 140106 196816
rect 169854 196874 169914 197252
rect 177030 197048 177090 197494
rect 172565 196874 172631 196877
rect 169854 196872 172631 196874
rect 169854 196816 172570 196872
rect 172626 196816 172631 196872
rect 169854 196814 172631 196816
rect 136777 196811 136843 196814
rect 172565 196811 172631 196814
rect 66213 196738 66279 196741
rect 66213 196736 67948 196738
rect 66213 196680 66218 196736
rect 66274 196680 67948 196736
rect 66213 196678 67948 196680
rect 66213 196675 66279 196678
rect 97726 196602 97786 196640
rect 100897 196602 100963 196605
rect 97726 196600 100963 196602
rect 97726 196544 100902 196600
rect 100958 196544 100963 196600
rect 97726 196542 100963 196544
rect 100897 196539 100963 196542
rect 136685 196602 136751 196605
rect 140046 196602 140106 196640
rect 136685 196600 140106 196602
rect 136685 196544 136690 196600
rect 136746 196544 140106 196600
rect 136685 196542 140106 196544
rect 169854 196602 169914 196708
rect 172657 196602 172723 196605
rect 169854 196600 172723 196602
rect 169854 196544 172662 196600
rect 172718 196544 172723 196600
rect 169854 196542 172723 196544
rect 136685 196539 136751 196542
rect 172657 196539 172723 196542
rect 62533 196330 62599 196333
rect 60588 196328 62599 196330
rect 60588 196272 62538 196328
rect 62594 196272 62599 196328
rect 60588 196270 62599 196272
rect 62533 196267 62599 196270
rect 102369 196330 102435 196333
rect 135397 196330 135463 196333
rect 102369 196328 104932 196330
rect 102369 196272 102374 196328
rect 102430 196272 104932 196328
rect 102369 196270 104932 196272
rect 132716 196328 135463 196330
rect 132716 196272 135402 196328
rect 135458 196272 135463 196328
rect 132716 196270 135463 196272
rect 102369 196267 102435 196270
rect 135397 196267 135463 196270
rect 174129 196330 174195 196333
rect 174129 196328 177060 196330
rect 174129 196272 174134 196328
rect 174190 196272 177060 196328
rect 174129 196270 177060 196272
rect 174129 196267 174195 196270
rect 135397 196194 135463 196197
rect 132686 196192 135463 196194
rect 65017 195786 65083 195789
rect 67918 195786 67978 196164
rect 132686 196136 135402 196192
rect 135458 196136 135463 196192
rect 174221 196194 174287 196197
rect 174221 196192 177090 196194
rect 132686 196134 135463 196136
rect 65017 195784 67978 195786
rect 65017 195728 65022 195784
rect 65078 195728 67978 195784
rect 65017 195726 67978 195728
rect 65017 195723 65083 195726
rect 62625 195650 62691 195653
rect 60588 195648 62691 195650
rect 60588 195592 62630 195648
rect 62686 195592 62691 195648
rect 60588 195590 62691 195592
rect 97726 195650 97786 196096
rect 132686 195688 132746 196134
rect 135397 196131 135463 196134
rect 100897 195650 100963 195653
rect 97726 195648 100963 195650
rect 97726 195592 100902 195648
rect 100958 195592 100963 195648
rect 97726 195590 100963 195592
rect 62625 195587 62691 195590
rect 100897 195587 100963 195590
rect 102461 195650 102527 195653
rect 136869 195650 136935 195653
rect 140046 195650 140106 196096
rect 169854 195786 169914 196164
rect 174221 196136 174226 196192
rect 174282 196136 177090 196192
rect 174221 196134 177090 196136
rect 174221 196131 174287 196134
rect 172381 195786 172447 195789
rect 169854 195784 172447 195786
rect 169854 195728 172386 195784
rect 172442 195728 172447 195784
rect 169854 195726 172447 195728
rect 172381 195723 172447 195726
rect 177030 195688 177090 196134
rect 102461 195648 104932 195650
rect 102461 195592 102466 195648
rect 102522 195592 104932 195648
rect 102461 195590 104932 195592
rect 136869 195648 140106 195650
rect 136869 195592 136874 195648
rect 136930 195592 140106 195648
rect 136869 195590 140106 195592
rect 102461 195587 102527 195590
rect 136869 195587 136935 195590
rect 66397 195514 66463 195517
rect 66397 195512 67948 195514
rect 66397 195456 66402 195512
rect 66458 195456 67948 195512
rect 66397 195454 67948 195456
rect 66397 195451 66463 195454
rect 97726 195242 97786 195416
rect 100897 195242 100963 195245
rect 97726 195240 100963 195242
rect 97726 195184 100902 195240
rect 100958 195184 100963 195240
rect 97726 195182 100963 195184
rect 100897 195179 100963 195182
rect 136777 195242 136843 195245
rect 140046 195242 140106 195416
rect 169854 195378 169914 195484
rect 172657 195378 172723 195381
rect 169854 195376 172723 195378
rect 169854 195320 172662 195376
rect 172718 195320 172723 195376
rect 169854 195318 172723 195320
rect 172657 195315 172723 195318
rect 136777 195240 140106 195242
rect 136777 195184 136782 195240
rect 136838 195184 140106 195240
rect 136777 195182 140106 195184
rect 136777 195179 136843 195182
rect 62625 194970 62691 194973
rect 60588 194968 62691 194970
rect 60588 194912 62630 194968
rect 62686 194912 62691 194968
rect 102553 194970 102619 194973
rect 135397 194970 135463 194973
rect 102553 194968 104932 194970
rect 60588 194910 62691 194912
rect 62625 194907 62691 194910
rect 65017 194562 65083 194565
rect 67918 194562 67978 194940
rect 102553 194912 102558 194968
rect 102614 194912 104932 194968
rect 102553 194910 104932 194912
rect 132716 194968 135463 194970
rect 132716 194912 135402 194968
rect 135458 194912 135463 194968
rect 174221 194970 174287 194973
rect 174221 194968 177060 194970
rect 132716 194910 135463 194912
rect 102553 194907 102619 194910
rect 135397 194907 135463 194910
rect 65017 194560 67978 194562
rect 65017 194504 65022 194560
rect 65078 194504 67978 194560
rect 65017 194502 67978 194504
rect 65017 194499 65083 194502
rect 97726 194426 97786 194872
rect 135397 194834 135463 194837
rect 132686 194832 135463 194834
rect 132686 194776 135402 194832
rect 135458 194776 135463 194832
rect 132686 194774 135463 194776
rect 100621 194426 100687 194429
rect 97726 194424 100687 194426
rect 97726 194368 100626 194424
rect 100682 194368 100687 194424
rect 97726 194366 100687 194368
rect 100621 194363 100687 194366
rect 132686 194328 132746 194774
rect 135397 194771 135463 194774
rect 136777 194426 136843 194429
rect 140046 194426 140106 194872
rect 136777 194424 140106 194426
rect 136777 194368 136782 194424
rect 136838 194368 140106 194424
rect 136777 194366 140106 194368
rect 169854 194426 169914 194940
rect 174221 194912 174226 194968
rect 174282 194912 177060 194968
rect 174221 194910 177060 194912
rect 174221 194907 174287 194910
rect 174129 194834 174195 194837
rect 174129 194832 177090 194834
rect 174129 194776 174134 194832
rect 174190 194776 177090 194832
rect 174129 194774 177090 194776
rect 174129 194771 174195 194774
rect 171737 194426 171803 194429
rect 169854 194424 171803 194426
rect 169854 194368 171742 194424
rect 171798 194368 171803 194424
rect 169854 194366 171803 194368
rect 136777 194363 136843 194366
rect 171737 194363 171803 194366
rect 177030 194328 177090 194774
rect 62533 194290 62599 194293
rect 60588 194288 62599 194290
rect 60588 194232 62538 194288
rect 62594 194232 62599 194288
rect 60588 194230 62599 194232
rect 62533 194227 62599 194230
rect 66397 194290 66463 194293
rect 102369 194290 102435 194293
rect 66397 194288 67948 194290
rect 66397 194232 66402 194288
rect 66458 194232 67948 194288
rect 66397 194230 67948 194232
rect 102369 194288 104932 194290
rect 102369 194232 102374 194288
rect 102430 194232 104932 194288
rect 102369 194230 104932 194232
rect 66397 194227 66463 194230
rect 102369 194227 102435 194230
rect 97726 193882 97786 194192
rect 100621 193882 100687 193885
rect 97726 193880 100687 193882
rect 97726 193824 100626 193880
rect 100682 193824 100687 193880
rect 97726 193822 100687 193824
rect 100621 193819 100687 193822
rect 136685 193882 136751 193885
rect 140046 193882 140106 194192
rect 169854 194018 169914 194260
rect 172657 194018 172723 194021
rect 169854 194016 172723 194018
rect 169854 193960 172662 194016
rect 172718 193960 172723 194016
rect 169854 193958 172723 193960
rect 172657 193955 172723 193958
rect 136685 193880 140106 193882
rect 136685 193824 136690 193880
rect 136746 193824 140106 193880
rect 136685 193822 140106 193824
rect 136685 193819 136751 193822
rect 64925 193746 64991 193749
rect 64925 193744 67948 193746
rect 64925 193688 64930 193744
rect 64986 193688 67948 193744
rect 64925 193686 67948 193688
rect 64925 193683 64991 193686
rect 62533 193610 62599 193613
rect 60588 193608 62599 193610
rect 60588 193552 62538 193608
rect 62594 193552 62599 193608
rect 60588 193550 62599 193552
rect 62533 193547 62599 193550
rect 97726 193338 97786 193648
rect 102461 193610 102527 193613
rect 135397 193610 135463 193613
rect 102461 193608 104932 193610
rect 102461 193552 102466 193608
rect 102522 193552 104932 193608
rect 102461 193550 104932 193552
rect 132716 193608 135463 193610
rect 132716 193552 135402 193608
rect 135458 193552 135463 193608
rect 132716 193550 135463 193552
rect 102461 193547 102527 193550
rect 135397 193547 135463 193550
rect 135397 193474 135463 193477
rect 132686 193472 135463 193474
rect 132686 193416 135402 193472
rect 135458 193416 135463 193472
rect 132686 193414 135463 193416
rect 99885 193338 99951 193341
rect 97726 193336 99951 193338
rect 97726 193280 99890 193336
rect 99946 193280 99951 193336
rect 97726 193278 99951 193280
rect 99885 193275 99951 193278
rect 62625 192930 62691 192933
rect 60588 192928 62691 192930
rect 60588 192872 62630 192928
rect 62686 192872 62691 192928
rect 60588 192870 62691 192872
rect 62625 192867 62691 192870
rect 65017 192794 65083 192797
rect 67918 192794 67978 193172
rect 65017 192792 67978 192794
rect 65017 192736 65022 192792
rect 65078 192736 67978 192792
rect 65017 192734 67978 192736
rect 65017 192731 65083 192734
rect 9896 192658 10376 192688
rect 11933 192658 11999 192661
rect 9896 192656 11999 192658
rect 9896 192600 11938 192656
rect 11994 192600 11999 192656
rect 9896 192598 11999 192600
rect 97726 192658 97786 193104
rect 132686 192968 132746 193414
rect 135397 193411 135463 193414
rect 136777 193338 136843 193341
rect 140046 193338 140106 193648
rect 136777 193336 140106 193338
rect 136777 193280 136782 193336
rect 136838 193280 140106 193336
rect 136777 193278 140106 193280
rect 169854 193338 169914 193716
rect 174129 193610 174195 193613
rect 174129 193608 177060 193610
rect 174129 193552 174134 193608
rect 174190 193552 177060 193608
rect 174129 193550 177060 193552
rect 174129 193547 174195 193550
rect 174221 193474 174287 193477
rect 174221 193472 177090 193474
rect 174221 193416 174226 193472
rect 174282 193416 177090 193472
rect 174221 193414 177090 193416
rect 174221 193411 174287 193414
rect 172013 193338 172079 193341
rect 169854 193336 172079 193338
rect 169854 193280 172018 193336
rect 172074 193280 172079 193336
rect 169854 193278 172079 193280
rect 136777 193275 136843 193278
rect 172013 193275 172079 193278
rect 102369 192930 102435 192933
rect 102369 192928 104932 192930
rect 102369 192872 102374 192928
rect 102430 192872 104932 192928
rect 102369 192870 104932 192872
rect 102369 192867 102435 192870
rect 100621 192658 100687 192661
rect 97726 192656 100687 192658
rect 97726 192600 100626 192656
rect 100682 192600 100687 192656
rect 97726 192598 100687 192600
rect 9896 192568 10376 192598
rect 11933 192595 11999 192598
rect 100621 192595 100687 192598
rect 136685 192658 136751 192661
rect 140046 192658 140106 193104
rect 169854 192794 169914 193172
rect 177030 192968 177090 193414
rect 172657 192794 172723 192797
rect 169854 192792 172723 192794
rect 169854 192736 172662 192792
rect 172718 192736 172723 192792
rect 169854 192734 172723 192736
rect 172657 192731 172723 192734
rect 171645 192658 171711 192661
rect 136685 192656 140106 192658
rect 136685 192600 136690 192656
rect 136746 192600 140106 192656
rect 136685 192598 140106 192600
rect 169670 192656 171711 192658
rect 169670 192600 171650 192656
rect 171706 192600 171711 192656
rect 169670 192598 171711 192600
rect 136685 192595 136751 192598
rect 65661 192522 65727 192525
rect 100529 192522 100595 192525
rect 65661 192520 67948 192522
rect 65661 192464 65666 192520
rect 65722 192464 67948 192520
rect 65661 192462 67948 192464
rect 97756 192520 100595 192522
rect 97756 192464 100534 192520
rect 100590 192464 100595 192520
rect 97756 192462 100595 192464
rect 65661 192459 65727 192462
rect 100529 192459 100595 192462
rect 136869 192522 136935 192525
rect 136869 192520 140076 192522
rect 136869 192464 136874 192520
rect 136930 192464 140076 192520
rect 169670 192492 169730 192598
rect 171645 192595 171711 192598
rect 207249 192522 207315 192525
rect 207566 192522 207572 192524
rect 204844 192520 207572 192522
rect 136869 192462 140076 192464
rect 204844 192464 207254 192520
rect 207310 192464 207572 192520
rect 204844 192462 207572 192464
rect 136869 192459 136935 192462
rect 207249 192459 207315 192462
rect 207566 192460 207572 192462
rect 207636 192460 207642 192524
rect 207249 192386 207315 192389
rect 207566 192386 207572 192388
rect 207249 192384 207572 192386
rect 207249 192328 207254 192384
rect 207310 192328 207572 192384
rect 207249 192326 207572 192328
rect 207249 192323 207315 192326
rect 207566 192324 207572 192326
rect 207636 192324 207642 192388
rect 62533 192250 62599 192253
rect 60588 192248 62599 192250
rect 60588 192192 62538 192248
rect 62594 192192 62599 192248
rect 60588 192190 62599 192192
rect 62533 192187 62599 192190
rect 102461 192250 102527 192253
rect 135397 192250 135463 192253
rect 102461 192248 104932 192250
rect 102461 192192 102466 192248
rect 102522 192192 104932 192248
rect 102461 192190 104932 192192
rect 132716 192248 135463 192250
rect 132716 192192 135402 192248
rect 135458 192192 135463 192248
rect 132716 192190 135463 192192
rect 102461 192187 102527 192190
rect 135397 192187 135463 192190
rect 174129 192250 174195 192253
rect 174129 192248 177060 192250
rect 174129 192192 174134 192248
rect 174190 192192 177060 192248
rect 174129 192190 177060 192192
rect 174129 192187 174195 192190
rect 135213 192114 135279 192117
rect 132686 192112 135279 192114
rect 132686 192056 135218 192112
rect 135274 192056 135279 192112
rect 132686 192054 135279 192056
rect 62349 191570 62415 191573
rect 60588 191568 62415 191570
rect 60588 191512 62354 191568
rect 62410 191512 62415 191568
rect 60588 191510 62415 191512
rect 62349 191507 62415 191510
rect 65017 191570 65083 191573
rect 67918 191570 67978 191948
rect 65017 191568 67978 191570
rect 65017 191512 65022 191568
rect 65078 191512 67978 191568
rect 65017 191510 67978 191512
rect 65017 191507 65083 191510
rect 97726 191434 97786 191880
rect 132686 191608 132746 192054
rect 135213 192051 135279 192054
rect 174221 192114 174287 192117
rect 174221 192112 177090 192114
rect 174221 192056 174226 192112
rect 174282 192056 177090 192112
rect 174221 192054 177090 192056
rect 174221 192051 174287 192054
rect 102369 191570 102435 191573
rect 102369 191568 104932 191570
rect 102369 191512 102374 191568
rect 102430 191512 104932 191568
rect 102369 191510 104932 191512
rect 102369 191507 102435 191510
rect 100621 191434 100687 191437
rect 97726 191432 100687 191434
rect 97726 191376 100626 191432
rect 100682 191376 100687 191432
rect 97726 191374 100687 191376
rect 100621 191371 100687 191374
rect 136777 191434 136843 191437
rect 140046 191434 140106 191880
rect 136777 191432 140106 191434
rect 136777 191376 136782 191432
rect 136838 191376 140106 191432
rect 136777 191374 140106 191376
rect 169854 191434 169914 191948
rect 177030 191608 177090 192054
rect 172657 191434 172723 191437
rect 169854 191432 172723 191434
rect 169854 191376 172662 191432
rect 172718 191376 172723 191432
rect 169854 191374 172723 191376
rect 136777 191371 136843 191374
rect 172657 191371 172723 191374
rect 65201 191298 65267 191301
rect 65201 191296 67948 191298
rect 65201 191240 65206 191296
rect 65262 191240 67948 191296
rect 65201 191238 67948 191240
rect 65201 191235 65267 191238
rect 97726 191162 97786 191200
rect 100897 191162 100963 191165
rect 97726 191160 100963 191162
rect 97726 191104 100902 191160
rect 100958 191104 100963 191160
rect 97726 191102 100963 191104
rect 100897 191099 100963 191102
rect 137145 191162 137211 191165
rect 140046 191162 140106 191200
rect 137145 191160 140106 191162
rect 137145 191104 137150 191160
rect 137206 191104 140106 191160
rect 137145 191102 140106 191104
rect 169854 191162 169914 191268
rect 171829 191162 171895 191165
rect 169854 191160 171895 191162
rect 169854 191104 171834 191160
rect 171890 191104 171895 191160
rect 169854 191102 171895 191104
rect 137145 191099 137211 191102
rect 171829 191099 171895 191102
rect 62625 190890 62691 190893
rect 60588 190888 62691 190890
rect 60588 190832 62630 190888
rect 62686 190832 62691 190888
rect 60588 190830 62691 190832
rect 62625 190827 62691 190830
rect 102645 190890 102711 190893
rect 135305 190890 135371 190893
rect 102645 190888 104932 190890
rect 102645 190832 102650 190888
rect 102706 190832 104932 190888
rect 102645 190830 104932 190832
rect 132716 190888 135371 190890
rect 132716 190832 135310 190888
rect 135366 190832 135371 190888
rect 132716 190830 135371 190832
rect 102645 190827 102711 190830
rect 135305 190827 135371 190830
rect 174313 190890 174379 190893
rect 174313 190888 177060 190890
rect 174313 190832 174318 190888
rect 174374 190832 177060 190888
rect 174313 190830 177060 190832
rect 174313 190827 174379 190830
rect 66305 190754 66371 190757
rect 135397 190754 135463 190757
rect 66305 190752 67948 190754
rect 66305 190696 66310 190752
rect 66366 190696 67948 190752
rect 66305 190694 67948 190696
rect 132686 190752 135463 190754
rect 132686 190696 135402 190752
rect 135458 190696 135463 190752
rect 174037 190754 174103 190757
rect 174037 190752 177090 190754
rect 132686 190694 135463 190696
rect 66305 190691 66371 190694
rect 97726 190346 97786 190656
rect 100437 190346 100503 190349
rect 97726 190344 100503 190346
rect 97726 190288 100442 190344
rect 100498 190288 100503 190344
rect 97726 190286 100503 190288
rect 100437 190283 100503 190286
rect 132686 190248 132746 190694
rect 135397 190691 135463 190694
rect 136777 190346 136843 190349
rect 140046 190346 140106 190656
rect 136777 190344 140106 190346
rect 136777 190288 136782 190344
rect 136838 190288 140106 190344
rect 136777 190286 140106 190288
rect 169854 190346 169914 190724
rect 174037 190696 174042 190752
rect 174098 190696 177090 190752
rect 174037 190694 177090 190696
rect 174037 190691 174103 190694
rect 171645 190346 171711 190349
rect 169854 190344 171711 190346
rect 169854 190288 171650 190344
rect 171706 190288 171711 190344
rect 169854 190286 171711 190288
rect 136777 190283 136843 190286
rect 171645 190283 171711 190286
rect 177030 190248 177090 190694
rect 62349 190210 62415 190213
rect 60588 190208 62415 190210
rect 60588 190152 62354 190208
rect 62410 190152 62415 190208
rect 60588 190150 62415 190152
rect 62349 190147 62415 190150
rect 66397 190210 66463 190213
rect 102277 190210 102343 190213
rect 66397 190208 67948 190210
rect 66397 190152 66402 190208
rect 66458 190152 67948 190208
rect 66397 190150 67948 190152
rect 102277 190208 104932 190210
rect 102277 190152 102282 190208
rect 102338 190152 104932 190208
rect 102277 190150 104932 190152
rect 66397 190147 66463 190150
rect 102277 190147 102343 190150
rect 97726 189938 97786 190112
rect 99977 189938 100043 189941
rect 97726 189936 100043 189938
rect 97726 189880 99982 189936
rect 100038 189880 100043 189936
rect 97726 189878 100043 189880
rect 99977 189875 100043 189878
rect 137237 189938 137303 189941
rect 140046 189938 140106 190112
rect 137237 189936 140106 189938
rect 137237 189880 137242 189936
rect 137298 189880 140106 189936
rect 137237 189878 140106 189880
rect 169854 189938 169914 190180
rect 171829 189938 171895 189941
rect 169854 189936 171895 189938
rect 169854 189880 171834 189936
rect 171890 189880 171895 189936
rect 169854 189878 171895 189880
rect 137237 189875 137303 189878
rect 171829 189875 171895 189878
rect 65017 189666 65083 189669
rect 66305 189666 66371 189669
rect 65017 189664 66371 189666
rect 65017 189608 65022 189664
rect 65078 189608 66310 189664
rect 66366 189608 66371 189664
rect 65017 189606 66371 189608
rect 65017 189603 65083 189606
rect 66305 189603 66371 189606
rect 62625 189530 62691 189533
rect 60588 189528 62691 189530
rect 60588 189472 62630 189528
rect 62686 189472 62691 189528
rect 60588 189470 62691 189472
rect 62625 189467 62691 189470
rect 102553 189530 102619 189533
rect 134201 189530 134267 189533
rect 102553 189528 104932 189530
rect 102553 189472 102558 189528
rect 102614 189472 104932 189528
rect 102553 189470 104932 189472
rect 132716 189528 134267 189530
rect 132716 189472 134206 189528
rect 134262 189472 134267 189528
rect 132716 189470 134267 189472
rect 102553 189467 102619 189470
rect 134201 189467 134267 189470
rect 175325 189530 175391 189533
rect 175325 189528 177060 189530
rect 175325 189472 175330 189528
rect 175386 189472 177060 189528
rect 175325 189470 177060 189472
rect 175325 189467 175391 189470
rect 134753 189258 134819 189261
rect 132686 189256 134819 189258
rect 132686 189200 134758 189256
rect 134814 189200 134819 189256
rect 132686 189198 134819 189200
rect 132686 188888 132746 189198
rect 134753 189195 134819 189198
rect 174405 189258 174471 189261
rect 174405 189256 177090 189258
rect 174405 189200 174410 189256
rect 174466 189200 177090 189256
rect 174405 189198 177090 189200
rect 174405 189195 174471 189198
rect 177030 188888 177090 189198
rect 62625 188850 62691 188853
rect 60588 188848 62691 188850
rect 60588 188792 62630 188848
rect 62686 188792 62691 188848
rect 60588 188790 62691 188792
rect 62625 188787 62691 188790
rect 102369 188850 102435 188853
rect 102369 188848 104932 188850
rect 102369 188792 102374 188848
rect 102430 188792 104932 188848
rect 102369 188790 104932 188792
rect 102369 188787 102435 188790
rect 63637 188170 63703 188173
rect 60588 188168 63703 188170
rect 60588 188112 63642 188168
rect 63698 188112 63703 188168
rect 60588 188110 63703 188112
rect 63637 188107 63703 188110
rect 102461 188170 102527 188173
rect 134937 188170 135003 188173
rect 102461 188168 104932 188170
rect 102461 188112 102466 188168
rect 102522 188112 104932 188168
rect 102461 188110 104932 188112
rect 132716 188168 135003 188170
rect 132716 188112 134942 188168
rect 134998 188112 135003 188168
rect 132716 188110 135003 188112
rect 102461 188107 102527 188110
rect 134937 188107 135003 188110
rect 175417 188170 175483 188173
rect 175417 188168 177060 188170
rect 175417 188112 175422 188168
rect 175478 188112 177060 188168
rect 175417 188110 177060 188112
rect 175417 188107 175483 188110
rect 225189 187354 225255 187357
rect 227416 187354 227896 187384
rect 225189 187352 227896 187354
rect 225189 187296 225194 187352
rect 225250 187296 227896 187352
rect 225189 187294 227896 187296
rect 225189 187291 225255 187294
rect 227416 187264 227896 187294
rect 117089 185450 117155 185453
rect 118193 185450 118259 185453
rect 117089 185448 118259 185450
rect 117089 185392 117094 185448
rect 117150 185392 118198 185448
rect 118254 185392 118259 185448
rect 117089 185390 118259 185392
rect 117089 185387 117155 185390
rect 118193 185387 118259 185390
rect 119113 185450 119179 185453
rect 121137 185450 121203 185453
rect 119113 185448 121203 185450
rect 119113 185392 119118 185448
rect 119174 185392 121142 185448
rect 121198 185392 121203 185448
rect 119113 185390 121203 185392
rect 119113 185387 119179 185390
rect 121137 185387 121203 185390
rect 126657 185450 126723 185453
rect 132177 185450 132243 185453
rect 126657 185448 132243 185450
rect 126657 185392 126662 185448
rect 126718 185392 132182 185448
rect 132238 185392 132243 185448
rect 126657 185390 132243 185392
rect 126657 185387 126723 185390
rect 132177 185387 132243 185390
rect 119481 185314 119547 185317
rect 121597 185314 121663 185317
rect 119481 185312 121663 185314
rect 119481 185256 119486 185312
rect 119542 185256 121602 185312
rect 121658 185256 121663 185312
rect 119481 185254 121663 185256
rect 119481 185251 119547 185254
rect 121597 185251 121663 185254
rect 125093 185314 125159 185317
rect 129969 185314 130035 185317
rect 125093 185312 130035 185314
rect 125093 185256 125098 185312
rect 125154 185256 129974 185312
rect 130030 185256 130035 185312
rect 125093 185254 130035 185256
rect 125093 185251 125159 185254
rect 129969 185251 130035 185254
rect 120677 185178 120743 185181
rect 122425 185178 122491 185181
rect 120677 185176 122491 185178
rect 120677 185120 120682 185176
rect 120738 185120 122430 185176
rect 122486 185120 122491 185176
rect 120677 185118 122491 185120
rect 120677 185115 120743 185118
rect 122425 185115 122491 185118
rect 125461 185178 125527 185181
rect 130429 185178 130495 185181
rect 125461 185176 130495 185178
rect 125461 185120 125466 185176
rect 125522 185120 130434 185176
rect 130490 185120 130495 185176
rect 125461 185118 130495 185120
rect 125461 185115 125527 185118
rect 130429 185115 130495 185118
rect 120309 185042 120375 185045
rect 122885 185042 122951 185045
rect 120309 185040 122951 185042
rect 120309 184984 120314 185040
rect 120370 184984 122890 185040
rect 122946 184984 122951 185040
rect 120309 184982 122951 184984
rect 120309 184979 120375 184982
rect 122885 184979 122951 184982
rect 125829 185042 125895 185045
rect 131441 185042 131507 185045
rect 125829 185040 131507 185042
rect 125829 184984 125834 185040
rect 125890 184984 131446 185040
rect 131502 184984 131507 185040
rect 125829 184982 131507 184984
rect 125829 184979 125895 184982
rect 131441 184979 131507 184982
rect 197451 185042 197517 185045
rect 202189 185042 202255 185045
rect 197451 185040 202255 185042
rect 197451 184984 197456 185040
rect 197512 184984 202194 185040
rect 202250 184984 202255 185040
rect 197451 184982 202255 184984
rect 197451 184979 197517 184982
rect 202189 184979 202255 184982
rect 124909 184906 124975 184909
rect 129325 184906 129391 184909
rect 124909 184904 129391 184906
rect 124909 184848 124914 184904
rect 124970 184848 129330 184904
rect 129386 184848 129391 184904
rect 124909 184846 129391 184848
rect 124909 184843 124975 184846
rect 129325 184843 129391 184846
rect 105589 184770 105655 184773
rect 102694 184768 105655 184770
rect 102694 184712 105594 184768
rect 105650 184712 105655 184768
rect 102694 184710 105655 184712
rect 38153 184498 38219 184501
rect 40177 184498 40243 184501
rect 38153 184496 40243 184498
rect 38153 184440 38158 184496
rect 38214 184440 40182 184496
rect 40238 184440 40243 184496
rect 38153 184438 40243 184440
rect 38153 184435 38219 184438
rect 40177 184435 40243 184438
rect 54897 184226 54963 184229
rect 60141 184226 60207 184229
rect 54897 184224 60207 184226
rect 102694 184224 102754 184710
rect 105589 184707 105655 184710
rect 116905 184770 116971 184773
rect 117641 184770 117707 184773
rect 116905 184768 117707 184770
rect 116905 184712 116910 184768
rect 116966 184712 117646 184768
rect 117702 184712 117707 184768
rect 116905 184710 117707 184712
rect 116905 184707 116971 184710
rect 117641 184707 117707 184710
rect 118101 184770 118167 184773
rect 119573 184770 119639 184773
rect 118101 184768 119639 184770
rect 118101 184712 118106 184768
rect 118162 184712 119578 184768
rect 119634 184712 119639 184768
rect 118101 184710 119639 184712
rect 118101 184707 118167 184710
rect 119573 184707 119639 184710
rect 126473 184770 126539 184773
rect 131625 184770 131691 184773
rect 126473 184768 131691 184770
rect 126473 184712 126478 184768
rect 126534 184712 131630 184768
rect 131686 184712 131691 184768
rect 126473 184710 131691 184712
rect 126473 184707 126539 184710
rect 131625 184707 131691 184710
rect 198509 184498 198575 184501
rect 203385 184498 203451 184501
rect 198509 184496 203451 184498
rect 198509 184440 198514 184496
rect 198570 184440 203390 184496
rect 203446 184440 203451 184496
rect 198509 184438 203451 184440
rect 198509 184435 198575 184438
rect 203385 184435 203451 184438
rect 177717 184226 177783 184229
rect 174852 184224 177783 184226
rect 54897 184168 54902 184224
rect 54958 184168 60146 184224
rect 60202 184168 60207 184224
rect 54897 184166 60207 184168
rect 174852 184168 177722 184224
rect 177778 184168 177783 184224
rect 174852 184166 177783 184168
rect 54897 184163 54963 184166
rect 60141 184163 60207 184166
rect 177717 184163 177783 184166
rect 198877 184226 198943 184229
rect 203937 184226 204003 184229
rect 198877 184224 204003 184226
rect 198877 184168 198882 184224
rect 198938 184168 203942 184224
rect 203998 184168 204003 184224
rect 198877 184166 204003 184168
rect 198877 184163 198943 184166
rect 203937 184163 204003 184166
rect 106141 183682 106207 183685
rect 102694 183680 106207 183682
rect 102694 183624 106146 183680
rect 106202 183624 106207 183680
rect 102694 183622 106207 183624
rect 20070 183484 20076 183548
rect 20140 183546 20146 183548
rect 20622 183546 20628 183548
rect 20140 183486 20628 183546
rect 20140 183484 20146 183486
rect 20622 183484 20628 183486
rect 20692 183484 20698 183548
rect 102694 183136 102754 183622
rect 106141 183619 106207 183622
rect 108533 183546 108599 183549
rect 180293 183546 180359 183549
rect 108533 183544 111004 183546
rect 108533 183488 108538 183544
rect 108594 183488 111004 183544
rect 108533 183486 111004 183488
rect 180293 183544 182948 183546
rect 180293 183488 180298 183544
rect 180354 183488 182948 183544
rect 180293 183486 182948 183488
rect 108533 183483 108599 183486
rect 180293 183483 180359 183486
rect 177349 183138 177415 183141
rect 174852 183136 177415 183138
rect 174852 183080 177354 183136
rect 177410 183080 177415 183136
rect 174852 183078 177415 183080
rect 177349 183075 177415 183078
rect 207249 183002 207315 183005
rect 207206 183000 207315 183002
rect 207206 182944 207254 183000
rect 207310 182944 207315 183000
rect 207206 182939 207315 182944
rect 207206 182868 207266 182939
rect 207198 182804 207204 182868
rect 207268 182804 207274 182868
rect 20806 182532 20812 182596
rect 20876 182594 20882 182596
rect 28718 182594 28724 182596
rect 20876 182534 28724 182594
rect 20876 182532 20882 182534
rect 28718 182532 28724 182534
rect 28788 182532 28794 182596
rect 105589 182322 105655 182325
rect 102694 182320 105655 182322
rect 102694 182264 105594 182320
rect 105650 182264 105655 182320
rect 102694 182262 105655 182264
rect 102694 181912 102754 182262
rect 105589 182259 105655 182262
rect 177165 181914 177231 181917
rect 174852 181912 177231 181914
rect 174852 181856 177170 181912
rect 177226 181856 177231 181912
rect 174852 181854 177231 181856
rect 177165 181851 177231 181854
rect 106049 181234 106115 181237
rect 102694 181232 106115 181234
rect 102694 181176 106054 181232
rect 106110 181176 106115 181232
rect 102694 181174 106115 181176
rect 102694 180824 102754 181174
rect 106049 181171 106115 181174
rect 108073 181234 108139 181237
rect 179649 181234 179715 181237
rect 108073 181232 111004 181234
rect 108073 181176 108078 181232
rect 108134 181176 111004 181232
rect 108073 181174 111004 181176
rect 179649 181232 182948 181234
rect 179649 181176 179654 181232
rect 179710 181176 182948 181232
rect 179649 181174 182948 181176
rect 108073 181171 108139 181174
rect 179649 181171 179715 181174
rect 176981 180826 177047 180829
rect 174852 180824 177047 180826
rect 174852 180768 176986 180824
rect 177042 180768 177047 180824
rect 174852 180766 177047 180768
rect 176981 180763 177047 180766
rect 105957 179874 106023 179877
rect 103062 179872 106023 179874
rect 103062 179816 105962 179872
rect 106018 179816 106023 179872
rect 103062 179814 106023 179816
rect 103062 179766 103122 179814
rect 105957 179811 106023 179814
rect 11933 179738 11999 179741
rect 11933 179736 14036 179738
rect 11933 179680 11938 179736
rect 11994 179680 14036 179736
rect 102724 179706 103122 179766
rect 177809 179738 177875 179741
rect 225189 179738 225255 179741
rect 174852 179736 177875 179738
rect 11933 179678 14036 179680
rect 174852 179680 177814 179736
rect 177870 179680 177875 179736
rect 174852 179678 177875 179680
rect 223796 179736 225255 179738
rect 223796 179680 225194 179736
rect 225250 179680 225255 179736
rect 223796 179678 225255 179680
rect 11933 179675 11999 179678
rect 177809 179675 177875 179678
rect 225189 179675 225255 179678
rect 107889 178922 107955 178925
rect 179649 178922 179715 178925
rect 107889 178920 111004 178922
rect 107889 178864 107894 178920
rect 107950 178864 111004 178920
rect 107889 178862 111004 178864
rect 179649 178920 182948 178922
rect 179649 178864 179654 178920
rect 179710 178864 182948 178920
rect 179649 178862 182948 178864
rect 107889 178859 107955 178862
rect 179649 178859 179715 178862
rect 105313 178514 105379 178517
rect 177625 178514 177691 178517
rect 102724 178512 105379 178514
rect 102724 178456 105318 178512
rect 105374 178456 105379 178512
rect 102724 178454 105379 178456
rect 174852 178512 177691 178514
rect 174852 178456 177630 178512
rect 177686 178456 177691 178512
rect 174852 178454 177691 178456
rect 105313 178451 105379 178454
rect 177625 178451 177691 178454
rect 31989 178242 32055 178245
rect 29860 178240 32055 178242
rect 29860 178184 31994 178240
rect 32050 178184 32055 178240
rect 29860 178182 32055 178184
rect 31989 178179 32055 178182
rect 37417 178242 37483 178245
rect 59589 178242 59655 178245
rect 204489 178242 204555 178245
rect 37417 178240 39060 178242
rect 37417 178184 37422 178240
rect 37478 178184 39060 178240
rect 37417 178182 39060 178184
rect 59589 178240 62980 178242
rect 59589 178184 59594 178240
rect 59650 178184 62980 178240
rect 59589 178182 62980 178184
rect 126828 178182 134924 178242
rect 204489 178240 207972 178242
rect 204489 178184 204494 178240
rect 204550 178184 207972 178240
rect 37417 178179 37483 178182
rect 59589 178179 59655 178182
rect 105221 177970 105287 177973
rect 102694 177968 105287 177970
rect 102694 177912 105226 177968
rect 105282 177912 105287 177968
rect 102694 177910 105287 177912
rect 102694 177424 102754 177910
rect 105221 177907 105287 177910
rect 198742 177698 198802 178184
rect 204489 178182 207972 178184
rect 204489 178179 204555 178182
rect 201085 177698 201151 177701
rect 198742 177696 201151 177698
rect 198742 177640 201090 177696
rect 201146 177640 201151 177696
rect 198742 177638 201151 177640
rect 201085 177635 201151 177638
rect 176889 177426 176955 177429
rect 174852 177424 176955 177426
rect 174852 177368 176894 177424
rect 176950 177368 176955 177424
rect 174852 177366 176955 177368
rect 176889 177363 176955 177366
rect 105129 176746 105195 176749
rect 102694 176744 105195 176746
rect 102694 176688 105134 176744
rect 105190 176688 105195 176744
rect 102694 176686 105195 176688
rect 102694 176200 102754 176686
rect 105129 176683 105195 176686
rect 107889 176474 107955 176477
rect 179649 176474 179715 176477
rect 107889 176472 111004 176474
rect 107889 176416 107894 176472
rect 107950 176416 111004 176472
rect 107889 176414 111004 176416
rect 179649 176472 182948 176474
rect 179649 176416 179654 176472
rect 179710 176416 182948 176472
rect 179649 176414 182948 176416
rect 107889 176411 107955 176414
rect 179649 176411 179715 176414
rect 177073 176202 177139 176205
rect 174852 176200 177139 176202
rect 174852 176144 177078 176200
rect 177134 176144 177139 176200
rect 174852 176142 177139 176144
rect 177073 176139 177139 176142
rect 106141 175386 106207 175389
rect 102694 175384 106207 175386
rect 102694 175328 106146 175384
rect 106202 175328 106207 175384
rect 102694 175326 106207 175328
rect 102694 175112 102754 175326
rect 106141 175323 106207 175326
rect 177165 175114 177231 175117
rect 174852 175112 177231 175114
rect 174852 175056 177170 175112
rect 177226 175056 177231 175112
rect 174852 175054 177231 175056
rect 177165 175051 177231 175054
rect 57381 174842 57447 174845
rect 54884 174840 57447 174842
rect 54884 174784 57386 174840
rect 57442 174784 57447 174840
rect 54884 174782 57447 174784
rect 57381 174779 57447 174782
rect 105405 174434 105471 174437
rect 102694 174432 105471 174434
rect 102694 174376 105410 174432
rect 105466 174376 105471 174432
rect 102694 174374 105471 174376
rect 102694 174024 102754 174374
rect 105405 174371 105471 174374
rect 107889 174162 107955 174165
rect 179649 174162 179715 174165
rect 107889 174160 111004 174162
rect 107889 174104 107894 174160
rect 107950 174104 111004 174160
rect 107889 174102 111004 174104
rect 179649 174160 182948 174162
rect 179649 174104 179654 174160
rect 179710 174104 182948 174160
rect 179649 174102 182948 174104
rect 107889 174099 107955 174102
rect 179649 174099 179715 174102
rect 178085 174026 178151 174029
rect 174852 174024 178151 174026
rect 174852 173968 178090 174024
rect 178146 173968 178151 174024
rect 174852 173966 178151 173968
rect 178085 173963 178151 173966
rect 106325 172938 106391 172941
rect 103062 172936 106391 172938
rect 103062 172880 106330 172936
rect 106386 172880 106391 172936
rect 103062 172878 106391 172880
rect 103062 172830 103122 172878
rect 106325 172875 106391 172878
rect 207382 172876 207388 172940
rect 207452 172938 207458 172940
rect 207566 172938 207572 172940
rect 207452 172878 207572 172938
rect 207452 172876 207458 172878
rect 207566 172876 207572 172878
rect 207636 172876 207642 172940
rect 102724 172770 103122 172830
rect 177809 172802 177875 172805
rect 174852 172800 177875 172802
rect 174852 172744 177814 172800
rect 177870 172744 177875 172800
rect 174852 172742 177875 172744
rect 177809 172739 177875 172742
rect 106417 172258 106483 172261
rect 102694 172256 106483 172258
rect 102694 172200 106422 172256
rect 106478 172200 106483 172256
rect 102694 172198 106483 172200
rect 102694 171712 102754 172198
rect 106417 172195 106483 172198
rect 108073 171850 108139 171853
rect 179649 171850 179715 171853
rect 108073 171848 111004 171850
rect 108073 171792 108078 171848
rect 108134 171792 111004 171848
rect 108073 171790 111004 171792
rect 179649 171848 182948 171850
rect 179649 171792 179654 171848
rect 179710 171792 182948 171848
rect 179649 171790 182948 171792
rect 108073 171787 108139 171790
rect 179649 171787 179715 171790
rect 177717 171714 177783 171717
rect 174852 171712 177783 171714
rect 174852 171656 177722 171712
rect 177778 171656 177783 171712
rect 174852 171654 177783 171656
rect 177717 171651 177783 171654
rect 9896 171034 10376 171064
rect 12025 171034 12091 171037
rect 105957 171034 106023 171037
rect 9896 171032 12091 171034
rect 9896 170976 12030 171032
rect 12086 170976 12091 171032
rect 9896 170974 12091 170976
rect 9896 170944 10376 170974
rect 12025 170971 12091 170974
rect 102694 171032 106023 171034
rect 102694 170976 105962 171032
rect 106018 170976 106023 171032
rect 102694 170974 106023 170976
rect 102694 170488 102754 170974
rect 105957 170971 106023 170974
rect 177533 170490 177599 170493
rect 174852 170488 177599 170490
rect 174852 170432 177538 170488
rect 177594 170432 177599 170488
rect 174852 170430 177599 170432
rect 177533 170427 177599 170430
rect 105681 169946 105747 169949
rect 102694 169944 105747 169946
rect 102694 169888 105686 169944
rect 105742 169888 105747 169944
rect 102694 169886 105747 169888
rect 12117 169266 12183 169269
rect 14006 169266 14066 169752
rect 102694 169400 102754 169886
rect 105681 169883 105747 169886
rect 178177 169402 178243 169405
rect 174852 169400 178243 169402
rect 12117 169264 14066 169266
rect 12117 169208 12122 169264
rect 12178 169208 14066 169264
rect 12117 169206 14066 169208
rect 12117 169203 12183 169206
rect 110974 168994 111034 169372
rect 174852 169344 178182 169400
rect 178238 169344 178243 169400
rect 174852 169342 178243 169344
rect 178177 169339 178243 169342
rect 182918 168994 182978 169372
rect 223582 169269 223642 169780
rect 223533 169264 223642 169269
rect 223533 169208 223538 169264
rect 223594 169208 223642 169264
rect 223533 169206 223642 169208
rect 223533 169203 223599 169206
rect 107846 168934 111034 168994
rect 179606 168934 182978 168994
rect 107846 168858 107906 168934
rect 179606 168858 179666 168934
rect 102694 168798 107906 168858
rect 174822 168798 179666 168858
rect 102694 168312 102754 168798
rect 174822 168284 174882 168798
rect 106601 167362 106667 167365
rect 106601 167360 111218 167362
rect 106601 167304 106606 167360
rect 106662 167304 111218 167360
rect 106601 167302 111218 167304
rect 106601 167299 106667 167302
rect 102724 167002 103122 167062
rect 111158 167060 111218 167302
rect 174852 167030 182948 167090
rect 103062 166954 103122 167002
rect 106509 166954 106575 166957
rect 103062 166952 106575 166954
rect 103062 166896 106514 166952
rect 106570 166896 106575 166952
rect 103062 166894 106575 166896
rect 106509 166891 106575 166894
rect 177165 166002 177231 166005
rect 174852 166000 177231 166002
rect 174852 165944 177170 166000
rect 177226 165944 177231 166000
rect 102694 165458 102754 165944
rect 174852 165942 177231 165944
rect 177165 165939 177231 165942
rect 105221 165458 105287 165461
rect 102694 165456 105287 165458
rect 102694 165400 105226 165456
rect 105282 165400 105287 165456
rect 102694 165398 105287 165400
rect 105221 165395 105287 165398
rect 32633 164914 32699 164917
rect 29860 164912 32699 164914
rect 29860 164856 32638 164912
rect 32694 164856 32699 164912
rect 29860 164854 32699 164856
rect 32633 164851 32699 164854
rect 37417 164914 37483 164917
rect 59589 164914 59655 164917
rect 200993 164914 201059 164917
rect 37417 164912 39060 164914
rect 37417 164856 37422 164912
rect 37478 164856 39060 164912
rect 37417 164854 39060 164856
rect 59589 164912 62980 164914
rect 59589 164856 59594 164912
rect 59650 164856 62980 164912
rect 59589 164854 62980 164856
rect 126828 164854 134924 164914
rect 198772 164912 201059 164914
rect 198772 164856 200998 164912
rect 201054 164856 201059 164912
rect 198772 164854 201059 164856
rect 37417 164851 37483 164854
rect 59589 164851 59655 164854
rect 200993 164851 201059 164854
rect 204489 164914 204555 164917
rect 204489 164912 207972 164914
rect 204489 164856 204494 164912
rect 204550 164856 207972 164912
rect 204489 164854 207972 164856
rect 204489 164851 204555 164854
rect 107797 164778 107863 164781
rect 177533 164778 177599 164781
rect 107797 164776 111004 164778
rect 107797 164720 107802 164776
rect 107858 164720 111004 164776
rect 102694 164234 102754 164720
rect 107797 164718 111004 164720
rect 174852 164776 177599 164778
rect 174852 164720 177538 164776
rect 177594 164720 177599 164776
rect 174852 164718 177599 164720
rect 107797 164715 107863 164718
rect 177533 164715 177599 164718
rect 179557 164778 179623 164781
rect 179557 164776 182948 164778
rect 179557 164720 179562 164776
rect 179618 164720 182948 164776
rect 179557 164718 182948 164720
rect 179557 164715 179623 164718
rect 105773 164234 105839 164237
rect 102694 164232 105839 164234
rect 102694 164176 105778 164232
rect 105834 164176 105839 164232
rect 102694 164174 105839 164176
rect 105773 164171 105839 164174
rect 176981 163690 177047 163693
rect 174852 163688 177047 163690
rect 102724 163602 103122 163662
rect 174852 163632 176986 163688
rect 177042 163632 177047 163688
rect 174852 163630 177047 163632
rect 176981 163627 177047 163630
rect 103062 163554 103122 163602
rect 105589 163554 105655 163557
rect 103062 163552 105655 163554
rect 103062 163496 105594 163552
rect 105650 163496 105655 163552
rect 103062 163494 105655 163496
rect 105589 163491 105655 163494
rect 224453 163554 224519 163557
rect 227416 163554 227896 163584
rect 224453 163552 227896 163554
rect 224453 163496 224458 163552
rect 224514 163496 227896 163552
rect 224453 163494 227896 163496
rect 224453 163491 224519 163494
rect 227416 163464 227896 163494
rect 207433 163282 207499 163285
rect 207566 163282 207572 163284
rect 207433 163280 207572 163282
rect 207433 163224 207438 163280
rect 207494 163224 207572 163280
rect 207433 163222 207572 163224
rect 207433 163219 207499 163222
rect 207566 163220 207572 163222
rect 207636 163220 207642 163284
rect 176981 162602 177047 162605
rect 174852 162600 177047 162602
rect 174852 162544 176986 162600
rect 177042 162544 177047 162600
rect 102694 162330 102754 162544
rect 174852 162542 177047 162544
rect 176981 162539 177047 162542
rect 107797 162466 107863 162469
rect 179557 162466 179623 162469
rect 107797 162464 111004 162466
rect 107797 162408 107802 162464
rect 107858 162408 111004 162464
rect 107797 162406 111004 162408
rect 179557 162464 182948 162466
rect 179557 162408 179562 162464
rect 179618 162408 182948 162464
rect 179557 162406 182948 162408
rect 107797 162403 107863 162406
rect 179557 162403 179623 162406
rect 105681 162330 105747 162333
rect 102694 162328 105747 162330
rect 102694 162272 105686 162328
rect 105742 162272 105747 162328
rect 102694 162270 105747 162272
rect 105681 162267 105747 162270
rect 177533 161378 177599 161381
rect 174852 161376 177599 161378
rect 174852 161320 177538 161376
rect 177594 161320 177599 161376
rect 102694 161106 102754 161320
rect 174852 161318 177599 161320
rect 177533 161315 177599 161318
rect 105221 161106 105287 161109
rect 102694 161104 105287 161106
rect 102694 161048 105226 161104
rect 105282 161048 105287 161104
rect 102694 161046 105287 161048
rect 105221 161043 105287 161046
rect 177349 160290 177415 160293
rect 174852 160288 177415 160290
rect 174852 160232 177354 160288
rect 177410 160232 177415 160288
rect 102694 159746 102754 160232
rect 174852 160230 177415 160232
rect 177349 160227 177415 160230
rect 107429 160018 107495 160021
rect 179189 160018 179255 160021
rect 107429 160016 111004 160018
rect 107429 159960 107434 160016
rect 107490 159960 111004 160016
rect 107429 159958 111004 159960
rect 179189 160016 182948 160018
rect 179189 159960 179194 160016
rect 179250 159960 182948 160016
rect 179189 159958 182948 159960
rect 107429 159955 107495 159958
rect 179189 159955 179255 159958
rect 105589 159746 105655 159749
rect 102694 159744 105655 159746
rect 102694 159688 105594 159744
rect 105650 159688 105655 159744
rect 12209 159338 12275 159341
rect 14006 159338 14066 159688
rect 102694 159686 105655 159688
rect 105589 159683 105655 159686
rect 12209 159336 14066 159338
rect 12209 159280 12214 159336
rect 12270 159280 14066 159336
rect 12209 159278 14066 159280
rect 12209 159275 12275 159278
rect 223582 159205 223642 159716
rect 223533 159200 223642 159205
rect 223533 159144 223538 159200
rect 223594 159144 223642 159200
rect 223533 159142 223642 159144
rect 223533 159139 223599 159142
rect 177625 159066 177691 159069
rect 174852 159064 177691 159066
rect 174852 159008 177630 159064
rect 177686 159008 177691 159064
rect 102694 158522 102754 159008
rect 174852 159006 177691 159008
rect 177625 159003 177691 159006
rect 105773 158522 105839 158525
rect 102694 158520 105839 158522
rect 102694 158464 105778 158520
rect 105834 158464 105839 158520
rect 102694 158462 105839 158464
rect 105773 158459 105839 158462
rect 106141 157978 106207 157981
rect 178177 157978 178243 157981
rect 102724 157976 106207 157978
rect 102724 157920 106146 157976
rect 106202 157920 106207 157976
rect 102724 157918 106207 157920
rect 174852 157976 178243 157978
rect 174852 157920 178182 157976
rect 178238 157920 178243 157976
rect 174852 157918 178243 157920
rect 106141 157915 106207 157918
rect 178177 157915 178243 157918
rect 107797 157706 107863 157709
rect 179557 157706 179623 157709
rect 107797 157704 111004 157706
rect 107797 157648 107802 157704
rect 107858 157648 111004 157704
rect 107797 157646 111004 157648
rect 179557 157704 182948 157706
rect 179557 157648 179562 157704
rect 179618 157648 182948 157704
rect 179557 157646 182948 157648
rect 107797 157643 107863 157646
rect 179557 157643 179623 157646
rect 177349 156890 177415 156893
rect 174852 156888 177415 156890
rect 102724 156802 103122 156862
rect 174852 156832 177354 156888
rect 177410 156832 177415 156888
rect 174852 156830 177415 156832
rect 177349 156827 177415 156830
rect 103062 156754 103122 156802
rect 106141 156754 106207 156757
rect 103062 156752 106207 156754
rect 103062 156696 106146 156752
rect 106202 156696 106207 156752
rect 103062 156694 106207 156696
rect 106141 156691 106207 156694
rect 178085 155666 178151 155669
rect 174852 155664 178151 155666
rect 174852 155608 178090 155664
rect 178146 155608 178151 155664
rect 102694 155394 102754 155608
rect 174852 155606 178151 155608
rect 178085 155603 178151 155606
rect 105773 155394 105839 155397
rect 102694 155392 105839 155394
rect 102694 155336 105778 155392
rect 105834 155336 105839 155392
rect 102694 155334 105839 155336
rect 105773 155331 105839 155334
rect 107705 155394 107771 155397
rect 179465 155394 179531 155397
rect 107705 155392 111004 155394
rect 107705 155336 107710 155392
rect 107766 155336 111004 155392
rect 107705 155334 111004 155336
rect 179465 155392 182948 155394
rect 179465 155336 179470 155392
rect 179526 155336 182948 155392
rect 179465 155334 182948 155336
rect 107705 155331 107771 155334
rect 179465 155331 179531 155334
rect 57473 154850 57539 154853
rect 54884 154848 57539 154850
rect 54884 154792 57478 154848
rect 57534 154792 57539 154848
rect 54884 154790 57539 154792
rect 57473 154787 57539 154790
rect 178269 154578 178335 154581
rect 174852 154576 178335 154578
rect 174852 154520 178274 154576
rect 178330 154520 178335 154576
rect 102694 154170 102754 154520
rect 174852 154518 178335 154520
rect 178269 154515 178335 154518
rect 106417 154170 106483 154173
rect 102694 154168 106483 154170
rect 102694 154112 106422 154168
rect 106478 154112 106483 154168
rect 102694 154110 106483 154112
rect 106417 154107 106483 154110
rect 207433 153764 207499 153765
rect 207382 153762 207388 153764
rect 207342 153702 207388 153762
rect 207452 153760 207499 153764
rect 207494 153704 207499 153760
rect 207382 153700 207388 153702
rect 207452 153700 207499 153704
rect 207433 153699 207499 153700
rect 178545 153354 178611 153357
rect 174852 153352 178611 153354
rect 174852 153296 178550 153352
rect 178606 153296 178611 153352
rect 102694 152946 102754 153296
rect 174852 153294 178611 153296
rect 178545 153291 178611 153294
rect 207341 153356 207407 153357
rect 207341 153352 207388 153356
rect 207452 153354 207458 153356
rect 207341 153296 207346 153352
rect 207341 153292 207388 153296
rect 207452 153294 207498 153354
rect 207452 153292 207458 153294
rect 207341 153291 207407 153292
rect 106601 152946 106667 152949
rect 102694 152944 106667 152946
rect 102694 152888 106606 152944
rect 106662 152888 106667 152944
rect 102694 152886 106667 152888
rect 106601 152883 106667 152886
rect 107613 152946 107679 152949
rect 179373 152946 179439 152949
rect 107613 152944 111004 152946
rect 107613 152888 107618 152944
rect 107674 152888 111004 152944
rect 107613 152886 111004 152888
rect 179373 152944 182948 152946
rect 179373 152888 179378 152944
rect 179434 152888 182948 152944
rect 179373 152886 182948 152888
rect 107613 152883 107679 152886
rect 179373 152883 179439 152886
rect 178453 152266 178519 152269
rect 174852 152264 178519 152266
rect 174852 152208 178458 152264
rect 178514 152208 178519 152264
rect 102694 151722 102754 152208
rect 174852 152206 178519 152208
rect 178453 152203 178519 152206
rect 105221 151722 105287 151725
rect 102694 151720 105287 151722
rect 102694 151664 105226 151720
rect 105282 151664 105287 151720
rect 102694 151662 105287 151664
rect 105221 151659 105287 151662
rect 31989 151586 32055 151589
rect 29860 151584 32055 151586
rect 29860 151528 31994 151584
rect 32050 151528 32055 151584
rect 29860 151526 32055 151528
rect 31989 151523 32055 151526
rect 37918 151524 37924 151588
rect 37988 151586 37994 151588
rect 59589 151586 59655 151589
rect 132361 151586 132427 151589
rect 200533 151586 200599 151589
rect 37988 151526 39060 151586
rect 59589 151584 62980 151586
rect 59589 151528 59594 151584
rect 59650 151528 62980 151584
rect 59589 151526 62980 151528
rect 126828 151584 134924 151586
rect 126828 151528 132366 151584
rect 132422 151528 134924 151584
rect 126828 151526 134924 151528
rect 198772 151584 200599 151586
rect 198772 151528 200538 151584
rect 200594 151528 200599 151584
rect 198772 151526 200599 151528
rect 37988 151524 37994 151526
rect 59589 151523 59655 151526
rect 132361 151523 132427 151526
rect 200533 151523 200599 151526
rect 204489 151586 204555 151589
rect 204489 151584 207972 151586
rect 204489 151528 204494 151584
rect 204550 151528 207972 151584
rect 204489 151526 207972 151528
rect 204489 151523 204555 151526
rect 176889 151178 176955 151181
rect 174852 151176 176955 151178
rect 102724 151090 103122 151150
rect 174852 151120 176894 151176
rect 176950 151120 176955 151176
rect 174852 151118 176955 151120
rect 176889 151115 176955 151118
rect 103062 151042 103122 151090
rect 105405 151042 105471 151045
rect 103062 151040 105471 151042
rect 103062 150984 105410 151040
rect 105466 150984 105471 151040
rect 103062 150982 105471 150984
rect 105405 150979 105471 150982
rect 108717 150634 108783 150637
rect 180477 150634 180543 150637
rect 108717 150632 111004 150634
rect 108717 150576 108722 150632
rect 108778 150576 111004 150632
rect 108717 150574 111004 150576
rect 180477 150632 182948 150634
rect 180477 150576 180482 150632
rect 180538 150576 182948 150632
rect 180477 150574 182948 150576
rect 108717 150571 108783 150574
rect 180477 150571 180543 150574
rect 177165 149954 177231 149957
rect 174852 149952 177231 149954
rect 174852 149896 177170 149952
rect 177226 149896 177231 149952
rect 11933 149818 11999 149821
rect 11933 149816 14036 149818
rect 11933 149760 11938 149816
rect 11994 149760 14036 149816
rect 11933 149758 14036 149760
rect 11933 149755 11999 149758
rect 102694 149682 102754 149896
rect 174852 149894 177231 149896
rect 177165 149891 177231 149894
rect 105129 149682 105195 149685
rect 102694 149680 105195 149682
rect 102694 149624 105134 149680
rect 105190 149624 105195 149680
rect 102694 149622 105195 149624
rect 105129 149619 105195 149622
rect 223582 149549 223642 149788
rect 223533 149544 223642 149549
rect 223533 149488 223538 149544
rect 223594 149488 223642 149544
rect 223533 149486 223642 149488
rect 223533 149483 223599 149486
rect 9896 149410 10376 149440
rect 12117 149410 12183 149413
rect 9896 149408 12183 149410
rect 9896 149352 12122 149408
rect 12178 149352 12183 149408
rect 9896 149350 12183 149352
rect 9896 149320 10376 149350
rect 12117 149347 12183 149350
rect 178361 148866 178427 148869
rect 174852 148864 178427 148866
rect 174852 148808 178366 148864
rect 178422 148808 178427 148864
rect 102694 148322 102754 148808
rect 174852 148806 178427 148808
rect 178361 148803 178427 148806
rect 106693 148322 106759 148325
rect 102694 148320 106759 148322
rect 102694 148264 106698 148320
rect 106754 148264 106759 148320
rect 102694 148262 106759 148264
rect 106693 148259 106759 148262
rect 108625 148322 108691 148325
rect 180385 148322 180451 148325
rect 108625 148320 111004 148322
rect 108625 148264 108630 148320
rect 108686 148264 111004 148320
rect 108625 148262 111004 148264
rect 180385 148320 182948 148322
rect 180385 148264 180390 148320
rect 180446 148264 182948 148320
rect 180385 148262 182948 148264
rect 108625 148259 108691 148262
rect 180385 148259 180451 148262
rect 177349 147642 177415 147645
rect 174852 147640 177415 147642
rect 174852 147584 177354 147640
rect 177410 147584 177415 147640
rect 102694 147234 102754 147584
rect 174852 147582 177415 147584
rect 177349 147579 177415 147582
rect 105957 147234 106023 147237
rect 102694 147232 106023 147234
rect 102694 147176 105962 147232
rect 106018 147176 106023 147232
rect 102694 147174 106023 147176
rect 105957 147171 106023 147174
rect 176838 146554 176844 146556
rect 174852 146494 176844 146554
rect 176838 146492 176844 146494
rect 176908 146492 176914 146556
rect 17126 146084 17132 146148
rect 17196 146146 17202 146148
rect 20438 146146 20444 146148
rect 17196 146086 20444 146146
rect 17196 146084 17202 146086
rect 20438 146084 20444 146086
rect 20508 146084 20514 146148
rect 108533 146010 108599 146013
rect 180293 146010 180359 146013
rect 108533 146008 111004 146010
rect 108533 145952 108538 146008
rect 108594 145952 111004 146008
rect 108533 145950 111004 145952
rect 180293 146008 182948 146010
rect 180293 145952 180298 146008
rect 180354 145952 182948 146008
rect 180293 145950 182948 145952
rect 108533 145947 108599 145950
rect 180293 145947 180359 145950
rect 174129 144922 174195 144925
rect 174454 144922 174514 145436
rect 174129 144920 174514 144922
rect 174129 144864 174134 144920
rect 174190 144864 174514 144920
rect 174129 144862 174514 144864
rect 174129 144859 174195 144862
rect 20438 142548 20444 142612
rect 20508 142610 20514 142612
rect 101030 142610 101036 142612
rect 20508 142550 101036 142610
rect 20508 142548 20514 142550
rect 101030 142548 101036 142550
rect 101100 142610 101106 142612
rect 102277 142610 102343 142613
rect 101100 142608 102343 142610
rect 101100 142552 102282 142608
rect 102338 142552 102343 142608
rect 101100 142550 102343 142552
rect 101100 142548 101106 142550
rect 102277 142547 102343 142550
rect 28718 142412 28724 142476
rect 28788 142474 28794 142476
rect 101173 142474 101239 142477
rect 28788 142472 101239 142474
rect 28788 142416 101178 142472
rect 101234 142416 101239 142472
rect 28788 142414 101239 142416
rect 28788 142412 28794 142414
rect 101173 142411 101239 142414
rect 175233 142202 175299 142205
rect 175233 142200 177090 142202
rect 175233 142144 175238 142200
rect 175294 142144 177090 142200
rect 175233 142142 177090 142144
rect 175233 142139 175299 142142
rect 62809 142066 62875 142069
rect 134109 142066 134175 142069
rect 60742 142064 62875 142066
rect 60742 142008 62814 142064
rect 62870 142008 62875 142064
rect 60742 142006 62875 142008
rect 60742 141560 60802 142006
rect 62809 142003 62875 142006
rect 132686 142064 134175 142066
rect 132686 142008 134114 142064
rect 134170 142008 134175 142064
rect 132686 142006 134175 142008
rect 91237 141930 91303 141933
rect 101582 141930 101588 141932
rect 91237 141928 101588 141930
rect 91237 141872 91242 141928
rect 91298 141872 101588 141928
rect 91237 141870 101588 141872
rect 91237 141867 91303 141870
rect 101582 141868 101588 141870
rect 101652 141868 101658 141932
rect 132686 141560 132746 142006
rect 134109 142003 134175 142006
rect 162169 141930 162235 141933
rect 173342 141930 173348 141932
rect 162169 141928 173348 141930
rect 162169 141872 162174 141928
rect 162230 141872 173348 141928
rect 162169 141870 173348 141872
rect 162169 141867 162235 141870
rect 173342 141868 173348 141870
rect 173412 141868 173418 141932
rect 177030 141560 177090 142142
rect 103105 141522 103171 141525
rect 103105 141520 104932 141522
rect 103105 141464 103110 141520
rect 103166 141464 104932 141520
rect 103105 141462 104932 141464
rect 103105 141459 103171 141462
rect 31897 141388 31963 141389
rect 31846 141386 31852 141388
rect 31806 141326 31852 141386
rect 31916 141384 31963 141388
rect 31958 141328 31963 141384
rect 31846 141324 31852 141326
rect 31916 141324 31963 141328
rect 31897 141323 31963 141324
rect 62809 140978 62875 140981
rect 60772 140976 62875 140978
rect 60772 140920 62814 140976
rect 62870 140920 62875 140976
rect 60772 140918 62875 140920
rect 62809 140915 62875 140918
rect 102277 140978 102343 140981
rect 135397 140978 135463 140981
rect 102277 140976 104932 140978
rect 102277 140920 102282 140976
rect 102338 140920 104932 140976
rect 102277 140918 104932 140920
rect 132716 140976 135463 140978
rect 132716 140920 135402 140976
rect 135458 140920 135463 140976
rect 132716 140918 135463 140920
rect 102277 140915 102343 140918
rect 135397 140915 135463 140918
rect 174773 140978 174839 140981
rect 174773 140976 177060 140978
rect 174773 140920 174778 140976
rect 174834 140920 177060 140976
rect 174773 140918 177060 140920
rect 174773 140915 174839 140918
rect 62717 140706 62783 140709
rect 135397 140706 135463 140709
rect 60742 140704 62783 140706
rect 60742 140648 62722 140704
rect 62778 140648 62783 140704
rect 60742 140646 62783 140648
rect 60742 140472 60802 140646
rect 62717 140643 62783 140646
rect 132686 140704 135463 140706
rect 132686 140648 135402 140704
rect 135458 140648 135463 140704
rect 132686 140646 135463 140648
rect 132686 140472 132746 140646
rect 135397 140643 135463 140646
rect 174221 140706 174287 140709
rect 174221 140704 177090 140706
rect 174221 140648 174226 140704
rect 174282 140648 177090 140704
rect 174221 140646 177090 140648
rect 174221 140643 174287 140646
rect 177030 140472 177090 140646
rect 102369 140434 102435 140437
rect 102369 140432 104932 140434
rect 102369 140376 102374 140432
rect 102430 140376 104932 140432
rect 102369 140374 104932 140376
rect 102369 140371 102435 140374
rect 62809 139754 62875 139757
rect 60772 139752 62875 139754
rect 60772 139696 62814 139752
rect 62870 139696 62875 139752
rect 60772 139694 62875 139696
rect 62809 139691 62875 139694
rect 102369 139754 102435 139757
rect 135397 139754 135463 139757
rect 102369 139752 104932 139754
rect 102369 139696 102374 139752
rect 102430 139696 104932 139752
rect 102369 139694 104932 139696
rect 132716 139752 135463 139754
rect 132716 139696 135402 139752
rect 135458 139696 135463 139752
rect 132716 139694 135463 139696
rect 102369 139691 102435 139694
rect 135397 139691 135463 139694
rect 174957 139754 175023 139757
rect 222889 139754 222955 139757
rect 227416 139754 227896 139784
rect 174957 139752 177060 139754
rect 174957 139696 174962 139752
rect 175018 139696 177060 139752
rect 174957 139694 177060 139696
rect 222889 139752 227896 139754
rect 222889 139696 222894 139752
rect 222950 139696 227896 139752
rect 222889 139694 227896 139696
rect 174957 139691 175023 139694
rect 222889 139691 222955 139694
rect 227416 139664 227896 139694
rect 62809 139482 62875 139485
rect 60742 139480 62875 139482
rect 60742 139424 62814 139480
rect 62870 139424 62875 139480
rect 60742 139422 62875 139424
rect 60742 139248 60802 139422
rect 62809 139419 62875 139422
rect 66213 139482 66279 139485
rect 135397 139482 135463 139485
rect 66213 139480 67948 139482
rect 66213 139424 66218 139480
rect 66274 139424 67948 139480
rect 66213 139422 67948 139424
rect 132686 139480 135463 139482
rect 132686 139424 135402 139480
rect 135458 139424 135463 139480
rect 174313 139482 174379 139485
rect 174313 139480 177090 139482
rect 132686 139422 135463 139424
rect 66213 139419 66279 139422
rect 97726 139074 97786 139384
rect 132686 139248 132746 139422
rect 135397 139419 135463 139422
rect 102461 139210 102527 139213
rect 102461 139208 104932 139210
rect 102461 139152 102466 139208
rect 102522 139152 104932 139208
rect 102461 139150 104932 139152
rect 102461 139147 102527 139150
rect 100621 139074 100687 139077
rect 97726 139072 100687 139074
rect 97726 139016 100626 139072
rect 100682 139016 100687 139072
rect 97726 139014 100687 139016
rect 100621 139011 100687 139014
rect 136869 139074 136935 139077
rect 140046 139074 140106 139384
rect 136869 139072 140106 139074
rect 136869 139016 136874 139072
rect 136930 139016 140106 139072
rect 136869 139014 140106 139016
rect 169854 139074 169914 139452
rect 174313 139424 174318 139480
rect 174374 139424 177090 139480
rect 174313 139422 177090 139424
rect 174313 139419 174379 139422
rect 177030 139248 177090 139422
rect 172473 139074 172539 139077
rect 169854 139072 172539 139074
rect 169854 139016 172478 139072
rect 172534 139016 172539 139072
rect 169854 139014 172539 139016
rect 136869 139011 136935 139014
rect 172473 139011 172539 139014
rect 62717 138938 62783 138941
rect 60742 138936 62783 138938
rect 60742 138880 62722 138936
rect 62778 138880 62783 138936
rect 60742 138878 62783 138880
rect 60742 138704 60802 138878
rect 62717 138875 62783 138878
rect 66397 138938 66463 138941
rect 134293 138938 134359 138941
rect 66397 138936 67948 138938
rect 66397 138880 66402 138936
rect 66458 138880 67948 138936
rect 66397 138878 67948 138880
rect 132686 138936 134359 138938
rect 132686 138880 134298 138936
rect 134354 138880 134359 138936
rect 132686 138878 134359 138880
rect 66397 138875 66463 138878
rect 97726 138666 97786 138840
rect 132686 138704 132746 138878
rect 134293 138875 134359 138878
rect 136961 138938 137027 138941
rect 175417 138938 175483 138941
rect 136961 138936 140076 138938
rect 136961 138880 136966 138936
rect 137022 138880 140076 138936
rect 175417 138936 177090 138938
rect 136961 138878 140076 138880
rect 136961 138875 137027 138878
rect 169854 138802 169914 138908
rect 175417 138880 175422 138936
rect 175478 138880 177090 138936
rect 175417 138878 177090 138880
rect 175417 138875 175483 138878
rect 172657 138802 172723 138805
rect 169854 138800 172723 138802
rect 169854 138744 172662 138800
rect 172718 138744 172723 138800
rect 169854 138742 172723 138744
rect 172657 138739 172723 138742
rect 177030 138704 177090 138878
rect 100529 138666 100595 138669
rect 97726 138664 100595 138666
rect 97726 138608 100534 138664
rect 100590 138608 100595 138664
rect 97726 138606 100595 138608
rect 100529 138603 100595 138606
rect 102553 138666 102619 138669
rect 102553 138664 104932 138666
rect 102553 138608 102558 138664
rect 102614 138608 104932 138664
rect 102553 138606 104932 138608
rect 102553 138603 102619 138606
rect 63453 138394 63519 138397
rect 60742 138392 63519 138394
rect 60742 138336 63458 138392
rect 63514 138336 63519 138392
rect 60742 138334 63519 138336
rect 60742 138024 60802 138334
rect 63453 138331 63519 138334
rect 100989 138394 101055 138397
rect 102134 138394 102140 138396
rect 100989 138392 102140 138394
rect 100989 138336 100994 138392
rect 101050 138336 102140 138392
rect 100989 138334 102140 138336
rect 100989 138331 101055 138334
rect 102134 138332 102140 138334
rect 102204 138332 102210 138396
rect 134477 138394 134543 138397
rect 132686 138392 134543 138394
rect 132686 138336 134482 138392
rect 134538 138336 134543 138392
rect 132686 138334 134543 138336
rect 66213 138258 66279 138261
rect 66213 138256 67948 138258
rect 66213 138200 66218 138256
rect 66274 138200 67948 138256
rect 66213 138198 67948 138200
rect 66213 138195 66279 138198
rect 97726 137850 97786 138160
rect 132686 138024 132746 138334
rect 134477 138331 134543 138334
rect 175141 138394 175207 138397
rect 175141 138392 177090 138394
rect 175141 138336 175146 138392
rect 175202 138336 177090 138392
rect 175141 138334 177090 138336
rect 175141 138331 175207 138334
rect 102369 137986 102435 137989
rect 102369 137984 104932 137986
rect 102369 137928 102374 137984
rect 102430 137928 104932 137984
rect 102369 137926 104932 137928
rect 102369 137923 102435 137926
rect 100713 137850 100779 137853
rect 97726 137848 100779 137850
rect 97726 137792 100718 137848
rect 100774 137792 100779 137848
rect 97726 137790 100779 137792
rect 100713 137787 100779 137790
rect 136869 137850 136935 137853
rect 140046 137850 140106 138160
rect 136869 137848 140106 137850
rect 136869 137792 136874 137848
rect 136930 137792 140106 137848
rect 136869 137790 140106 137792
rect 169854 137850 169914 138228
rect 177030 138024 177090 138334
rect 172197 137850 172263 137853
rect 169854 137848 172263 137850
rect 169854 137792 172202 137848
rect 172258 137792 172263 137848
rect 169854 137790 172263 137792
rect 136869 137787 136935 137790
rect 172197 137787 172263 137790
rect 62349 137714 62415 137717
rect 60742 137712 62415 137714
rect 60742 137656 62354 137712
rect 62410 137656 62415 137712
rect 60742 137654 62415 137656
rect 60742 137480 60802 137654
rect 62349 137651 62415 137654
rect 66397 137714 66463 137717
rect 134569 137714 134635 137717
rect 66397 137712 67948 137714
rect 66397 137656 66402 137712
rect 66458 137656 67948 137712
rect 66397 137654 67948 137656
rect 132686 137712 134635 137714
rect 132686 137656 134574 137712
rect 134630 137656 134635 137712
rect 174129 137714 174195 137717
rect 174129 137712 177090 137714
rect 132686 137654 134635 137656
rect 66397 137651 66463 137654
rect 97726 137306 97786 137616
rect 132686 137480 132746 137654
rect 134569 137651 134635 137654
rect 102461 137442 102527 137445
rect 102461 137440 104932 137442
rect 102461 137384 102466 137440
rect 102522 137384 104932 137440
rect 102461 137382 104932 137384
rect 102461 137379 102527 137382
rect 100345 137306 100411 137309
rect 97726 137304 100411 137306
rect 97726 137248 100350 137304
rect 100406 137248 100411 137304
rect 97726 137246 100411 137248
rect 100345 137243 100411 137246
rect 136961 137306 137027 137309
rect 140046 137306 140106 137616
rect 136961 137304 140106 137306
rect 136961 137248 136966 137304
rect 137022 137248 140106 137304
rect 136961 137246 140106 137248
rect 169854 137306 169914 137684
rect 174129 137656 174134 137712
rect 174190 137656 177090 137712
rect 174129 137654 177090 137656
rect 174129 137651 174195 137654
rect 177030 137480 177090 137654
rect 172657 137306 172723 137309
rect 169854 137304 172723 137306
rect 169854 137248 172662 137304
rect 172718 137248 172723 137304
rect 169854 137246 172723 137248
rect 136961 137243 137027 137246
rect 172657 137243 172723 137246
rect 30517 137170 30583 137173
rect 62809 137170 62875 137173
rect 30517 137168 32988 137170
rect 30517 137112 30522 137168
rect 30578 137112 32988 137168
rect 30517 137110 32988 137112
rect 60742 137168 62875 137170
rect 60742 137112 62814 137168
rect 62870 137112 62875 137168
rect 174221 137170 174287 137173
rect 207249 137170 207315 137173
rect 174221 137168 177090 137170
rect 60742 137110 62875 137112
rect 30517 137107 30583 137110
rect 60742 136936 60802 137110
rect 62809 137107 62875 137110
rect 62901 136626 62967 136629
rect 67918 136626 67978 137140
rect 60742 136624 62967 136626
rect 60742 136568 62906 136624
rect 62962 136568 62967 136624
rect 60742 136566 62967 136568
rect 60742 136392 60802 136566
rect 62901 136563 62967 136566
rect 65894 136566 67978 136626
rect 97726 136626 97786 137072
rect 102829 136898 102895 136901
rect 135397 136898 135463 136901
rect 102829 136896 104932 136898
rect 102829 136840 102834 136896
rect 102890 136840 104932 136896
rect 102829 136838 104932 136840
rect 132716 136896 135463 136898
rect 132716 136840 135402 136896
rect 135458 136840 135463 136896
rect 132716 136838 135463 136840
rect 102829 136835 102895 136838
rect 135397 136835 135463 136838
rect 100897 136626 100963 136629
rect 135121 136626 135187 136629
rect 97726 136624 100963 136626
rect 97726 136568 100902 136624
rect 100958 136568 100963 136624
rect 97726 136566 100963 136568
rect 65017 136218 65083 136221
rect 65894 136218 65954 136566
rect 100897 136563 100963 136566
rect 132686 136624 135187 136626
rect 132686 136568 135126 136624
rect 135182 136568 135187 136624
rect 132686 136566 135187 136568
rect 66029 136490 66095 136493
rect 66029 136488 67948 136490
rect 66029 136432 66034 136488
rect 66090 136432 67948 136488
rect 66029 136430 67948 136432
rect 66029 136427 66095 136430
rect 132686 136392 132746 136566
rect 135121 136563 135187 136566
rect 136777 136626 136843 136629
rect 140046 136626 140106 137072
rect 136777 136624 140106 136626
rect 136777 136568 136782 136624
rect 136838 136568 140106 136624
rect 136777 136566 140106 136568
rect 169854 136626 169914 137140
rect 174221 137112 174226 137168
rect 174282 137112 177090 137168
rect 174221 137110 177090 137112
rect 204844 137168 207315 137170
rect 204844 137112 207254 137168
rect 207310 137112 207315 137168
rect 204844 137110 207315 137112
rect 174221 137107 174287 137110
rect 177030 136936 177090 137110
rect 207249 137107 207315 137110
rect 172013 136626 172079 136629
rect 169854 136624 172079 136626
rect 169854 136568 172018 136624
rect 172074 136568 172079 136624
rect 169854 136566 172079 136568
rect 136777 136563 136843 136566
rect 172013 136563 172079 136566
rect 174313 136626 174379 136629
rect 174313 136624 177090 136626
rect 174313 136568 174318 136624
rect 174374 136568 177090 136624
rect 174313 136566 177090 136568
rect 174313 136563 174379 136566
rect 65017 136216 65954 136218
rect 65017 136160 65022 136216
rect 65078 136160 65954 136216
rect 65017 136158 65954 136160
rect 65017 136155 65083 136158
rect 97726 136082 97786 136392
rect 102461 136354 102527 136357
rect 102461 136352 104932 136354
rect 102461 136296 102466 136352
rect 102522 136296 104932 136352
rect 102461 136294 104932 136296
rect 102461 136291 102527 136294
rect 100621 136082 100687 136085
rect 97726 136080 100687 136082
rect 97726 136024 100626 136080
rect 100682 136024 100687 136080
rect 97726 136022 100687 136024
rect 100621 136019 100687 136022
rect 136869 136082 136935 136085
rect 140046 136082 140106 136392
rect 169854 136218 169914 136460
rect 177030 136392 177090 136566
rect 172565 136218 172631 136221
rect 169854 136216 172631 136218
rect 169854 136160 172570 136216
rect 172626 136160 172631 136216
rect 169854 136158 172631 136160
rect 172565 136155 172631 136158
rect 172657 136082 172723 136085
rect 136869 136080 140106 136082
rect 136869 136024 136874 136080
rect 136930 136024 140106 136080
rect 136869 136022 140106 136024
rect 169670 136080 172723 136082
rect 169670 136024 172662 136080
rect 172718 136024 172723 136080
rect 169670 136022 172723 136024
rect 136869 136019 136935 136022
rect 66397 135946 66463 135949
rect 100897 135946 100963 135949
rect 66397 135944 67948 135946
rect 66397 135888 66402 135944
rect 66458 135888 67948 135944
rect 66397 135886 67948 135888
rect 97756 135944 100963 135946
rect 97756 135888 100902 135944
rect 100958 135888 100963 135944
rect 97756 135886 100963 135888
rect 66397 135883 66463 135886
rect 100897 135883 100963 135886
rect 136961 135946 137027 135949
rect 136961 135944 140076 135946
rect 136961 135888 136966 135944
rect 137022 135888 140076 135944
rect 169670 135916 169730 136022
rect 172657 136019 172723 136022
rect 136961 135886 140076 135888
rect 136961 135883 137027 135886
rect 62717 135674 62783 135677
rect 60772 135672 62783 135674
rect 60772 135616 62722 135672
rect 62778 135616 62783 135672
rect 60772 135614 62783 135616
rect 62717 135611 62783 135614
rect 102369 135674 102435 135677
rect 135305 135674 135371 135677
rect 102369 135672 104932 135674
rect 102369 135616 102374 135672
rect 102430 135616 104932 135672
rect 102369 135614 104932 135616
rect 132716 135672 135371 135674
rect 132716 135616 135310 135672
rect 135366 135616 135371 135672
rect 132716 135614 135371 135616
rect 102369 135611 102435 135614
rect 135305 135611 135371 135614
rect 173945 135674 174011 135677
rect 173945 135672 177060 135674
rect 173945 135616 173950 135672
rect 174006 135616 177060 135672
rect 173945 135614 177060 135616
rect 173945 135611 174011 135614
rect 62625 135402 62691 135405
rect 135213 135402 135279 135405
rect 60742 135400 62691 135402
rect 60742 135344 62630 135400
rect 62686 135344 62691 135400
rect 60742 135342 62691 135344
rect 60742 135168 60802 135342
rect 62625 135339 62691 135342
rect 132686 135400 135279 135402
rect 132686 135344 135218 135400
rect 135274 135344 135279 135400
rect 132686 135342 135279 135344
rect 66305 135266 66371 135269
rect 66305 135264 67948 135266
rect 66305 135208 66310 135264
rect 66366 135208 67948 135264
rect 66305 135206 67948 135208
rect 66305 135203 66371 135206
rect 132686 135168 132746 135342
rect 135213 135339 135279 135342
rect 174037 135402 174103 135405
rect 174037 135400 177090 135402
rect 174037 135344 174042 135400
rect 174098 135344 177090 135400
rect 174037 135342 177090 135344
rect 174037 135339 174103 135342
rect 62717 134858 62783 134861
rect 60742 134856 62783 134858
rect 60742 134800 62722 134856
rect 62778 134800 62783 134856
rect 60742 134798 62783 134800
rect 97726 134858 97786 135168
rect 102645 135130 102711 135133
rect 102645 135128 104932 135130
rect 102645 135072 102650 135128
rect 102706 135072 104932 135128
rect 102645 135070 104932 135072
rect 102645 135067 102711 135070
rect 100069 134858 100135 134861
rect 135029 134858 135095 134861
rect 97726 134856 100135 134858
rect 97726 134800 100074 134856
rect 100130 134800 100135 134856
rect 97726 134798 100135 134800
rect 60742 134624 60802 134798
rect 62717 134795 62783 134798
rect 100069 134795 100135 134798
rect 132686 134856 135095 134858
rect 132686 134800 135034 134856
rect 135090 134800 135095 134856
rect 132686 134798 135095 134800
rect 66397 134722 66463 134725
rect 100897 134722 100963 134725
rect 66397 134720 67948 134722
rect 66397 134664 66402 134720
rect 66458 134664 67948 134720
rect 66397 134662 67948 134664
rect 97756 134720 100963 134722
rect 97756 134664 100902 134720
rect 100958 134664 100963 134720
rect 97756 134662 100963 134664
rect 66397 134659 66463 134662
rect 100897 134659 100963 134662
rect 132686 134624 132746 134798
rect 135029 134795 135095 134798
rect 136869 134858 136935 134861
rect 140046 134858 140106 135168
rect 136869 134856 140106 134858
rect 136869 134800 136874 134856
rect 136930 134800 140106 134856
rect 136869 134798 140106 134800
rect 169854 134858 169914 135236
rect 177030 135168 177090 135342
rect 171829 134858 171895 134861
rect 169854 134856 171895 134858
rect 169854 134800 171834 134856
rect 171890 134800 171895 134856
rect 169854 134798 171895 134800
rect 136869 134795 136935 134798
rect 171829 134795 171895 134798
rect 174313 134858 174379 134861
rect 174313 134856 177090 134858
rect 174313 134800 174318 134856
rect 174374 134800 177090 134856
rect 174313 134798 177090 134800
rect 174313 134795 174379 134798
rect 136961 134722 137027 134725
rect 136961 134720 140076 134722
rect 136961 134664 136966 134720
rect 137022 134664 140076 134720
rect 136961 134662 140076 134664
rect 136961 134659 137027 134662
rect 101173 134586 101239 134589
rect 102461 134586 102527 134589
rect 169854 134586 169914 134692
rect 177030 134624 177090 134798
rect 172657 134586 172723 134589
rect 101173 134584 101834 134586
rect 101173 134528 101178 134584
rect 101234 134528 101834 134584
rect 101173 134526 101834 134528
rect 101173 134523 101239 134526
rect 101774 134452 101834 134526
rect 102461 134584 104932 134586
rect 102461 134528 102466 134584
rect 102522 134528 104932 134584
rect 102461 134526 104932 134528
rect 169854 134584 172723 134586
rect 169854 134528 172662 134584
rect 172718 134528 172723 134584
rect 169854 134526 172723 134528
rect 102461 134523 102527 134526
rect 172657 134523 172723 134526
rect 101766 134388 101772 134452
rect 101836 134388 101842 134452
rect 62901 134314 62967 134317
rect 135121 134314 135187 134317
rect 60742 134312 62967 134314
rect 60742 134256 62906 134312
rect 62962 134256 62967 134312
rect 60742 134254 62967 134256
rect 60742 133944 60802 134254
rect 62901 134251 62967 134254
rect 132686 134312 135187 134314
rect 132686 134256 135126 134312
rect 135182 134256 135187 134312
rect 132686 134254 135187 134256
rect 65845 134178 65911 134181
rect 65845 134176 67948 134178
rect 65845 134120 65850 134176
rect 65906 134120 67948 134176
rect 65845 134118 67948 134120
rect 65845 134115 65911 134118
rect 62993 133634 63059 133637
rect 60742 133632 63059 133634
rect 60742 133576 62998 133632
rect 63054 133576 63059 133632
rect 60742 133574 63059 133576
rect 97726 133634 97786 134080
rect 132686 133944 132746 134254
rect 135121 134251 135187 134254
rect 174129 134314 174195 134317
rect 174129 134312 177090 134314
rect 174129 134256 174134 134312
rect 174190 134256 177090 134312
rect 174129 134254 177090 134256
rect 174129 134251 174195 134254
rect 102185 133906 102251 133909
rect 102185 133904 104932 133906
rect 102185 133848 102190 133904
rect 102246 133848 104932 133904
rect 102185 133846 104932 133848
rect 102185 133843 102251 133846
rect 100069 133634 100135 133637
rect 134937 133634 135003 133637
rect 97726 133632 100135 133634
rect 97726 133576 100074 133632
rect 100130 133576 100135 133632
rect 97726 133574 100135 133576
rect 60742 133400 60802 133574
rect 62993 133571 63059 133574
rect 100069 133571 100135 133574
rect 132686 133632 135003 133634
rect 132686 133576 134942 133632
rect 134998 133576 135003 133632
rect 132686 133574 135003 133576
rect 66397 133498 66463 133501
rect 66397 133496 67948 133498
rect 66397 133440 66402 133496
rect 66458 133440 67948 133496
rect 66397 133438 67948 133440
rect 66397 133435 66463 133438
rect 132686 133400 132746 133574
rect 134937 133571 135003 133574
rect 136961 133634 137027 133637
rect 140046 133634 140106 134080
rect 136961 133632 140106 133634
rect 136961 133576 136966 133632
rect 137022 133576 140106 133632
rect 136961 133574 140106 133576
rect 169854 133634 169914 134148
rect 177030 133944 177090 134254
rect 172197 133634 172263 133637
rect 169854 133632 172263 133634
rect 169854 133576 172202 133632
rect 172258 133576 172263 133632
rect 169854 133574 172263 133576
rect 136961 133571 137027 133574
rect 172197 133571 172263 133574
rect 174497 133634 174563 133637
rect 174497 133632 177090 133634
rect 174497 133576 174502 133632
rect 174558 133576 177090 133632
rect 174497 133574 177090 133576
rect 174497 133571 174563 133574
rect 97726 133226 97786 133400
rect 102093 133362 102159 133365
rect 102093 133360 104932 133362
rect 102093 133304 102098 133360
rect 102154 133304 104932 133360
rect 102093 133302 104932 133304
rect 102093 133299 102159 133302
rect 100897 133226 100963 133229
rect 97726 133224 100963 133226
rect 97726 133168 100902 133224
rect 100958 133168 100963 133224
rect 97726 133166 100963 133168
rect 100897 133163 100963 133166
rect 136869 133090 136935 133093
rect 140046 133090 140106 133400
rect 169854 133226 169914 133468
rect 177030 133400 177090 133574
rect 172657 133226 172723 133229
rect 169854 133224 172723 133226
rect 169854 133168 172662 133224
rect 172718 133168 172723 133224
rect 169854 133166 172723 133168
rect 172657 133163 172723 133166
rect 136869 133088 140106 133090
rect 136869 133032 136874 133088
rect 136930 133032 140106 133088
rect 136869 133030 140106 133032
rect 136869 133027 136935 133030
rect 62809 132818 62875 132821
rect 60772 132816 62875 132818
rect 60772 132760 62814 132816
rect 62870 132760 62875 132816
rect 60772 132758 62875 132760
rect 62809 132755 62875 132758
rect 62717 132546 62783 132549
rect 60742 132544 62783 132546
rect 60742 132488 62722 132544
rect 62778 132488 62783 132544
rect 60742 132486 62783 132488
rect 60742 132312 60802 132486
rect 62717 132483 62783 132486
rect 65017 132546 65083 132549
rect 67918 132546 67978 132924
rect 65017 132544 67978 132546
rect 65017 132488 65022 132544
rect 65078 132488 67978 132544
rect 65017 132486 67978 132488
rect 65017 132483 65083 132486
rect 97726 132410 97786 132856
rect 102277 132818 102343 132821
rect 135397 132818 135463 132821
rect 102277 132816 104932 132818
rect 102277 132760 102282 132816
rect 102338 132760 104932 132816
rect 102277 132758 104932 132760
rect 132716 132816 135463 132818
rect 132716 132760 135402 132816
rect 135458 132760 135463 132816
rect 132716 132758 135463 132760
rect 102277 132755 102343 132758
rect 135397 132755 135463 132758
rect 135213 132546 135279 132549
rect 132686 132544 135279 132546
rect 132686 132488 135218 132544
rect 135274 132488 135279 132544
rect 132686 132486 135279 132488
rect 100437 132410 100503 132413
rect 97726 132408 100503 132410
rect 97726 132352 100442 132408
rect 100498 132352 100503 132408
rect 97726 132350 100503 132352
rect 100437 132347 100503 132350
rect 132686 132312 132746 132486
rect 135213 132483 135279 132486
rect 136777 132410 136843 132413
rect 140046 132410 140106 132856
rect 136777 132408 140106 132410
rect 136777 132352 136782 132408
rect 136838 132352 140106 132408
rect 136777 132350 140106 132352
rect 169854 132410 169914 132924
rect 174221 132818 174287 132821
rect 174221 132816 177060 132818
rect 174221 132760 174226 132816
rect 174282 132760 177060 132816
rect 174221 132758 177060 132760
rect 174221 132755 174287 132758
rect 174313 132546 174379 132549
rect 174313 132544 177090 132546
rect 174313 132488 174318 132544
rect 174374 132488 177090 132544
rect 174313 132486 177090 132488
rect 174313 132483 174379 132486
rect 172381 132410 172447 132413
rect 169854 132408 172447 132410
rect 169854 132352 172386 132408
rect 172442 132352 172447 132408
rect 169854 132350 172447 132352
rect 136777 132347 136843 132350
rect 172381 132347 172447 132350
rect 177030 132312 177090 132486
rect 66397 132274 66463 132277
rect 102369 132274 102435 132277
rect 66397 132272 67948 132274
rect 66397 132216 66402 132272
rect 66458 132216 67948 132272
rect 66397 132214 67948 132216
rect 102369 132272 104932 132274
rect 102369 132216 102374 132272
rect 102430 132216 104932 132272
rect 102369 132214 104932 132216
rect 66397 132211 66463 132214
rect 102369 132211 102435 132214
rect 97726 132002 97786 132176
rect 100897 132002 100963 132005
rect 97726 132000 100963 132002
rect 97726 131944 100902 132000
rect 100958 131944 100963 132000
rect 97726 131942 100963 131944
rect 100897 131939 100963 131942
rect 136869 132002 136935 132005
rect 140046 132002 140106 132176
rect 136869 132000 140106 132002
rect 136869 131944 136874 132000
rect 136930 131944 140106 132000
rect 136869 131942 140106 131944
rect 169854 132002 169914 132244
rect 172013 132002 172079 132005
rect 169854 132000 172079 132002
rect 169854 131944 172018 132000
rect 172074 131944 172079 132000
rect 169854 131942 172079 131944
rect 136869 131939 136935 131942
rect 172013 131939 172079 131942
rect 172657 131866 172723 131869
rect 169670 131864 172723 131866
rect 169670 131808 172662 131864
rect 172718 131808 172723 131864
rect 169670 131806 172723 131808
rect 65661 131730 65727 131733
rect 100897 131730 100963 131733
rect 65661 131728 67948 131730
rect 65661 131672 65666 131728
rect 65722 131672 67948 131728
rect 65661 131670 67948 131672
rect 97756 131728 100963 131730
rect 97756 131672 100902 131728
rect 100958 131672 100963 131728
rect 97756 131670 100963 131672
rect 65661 131667 65727 131670
rect 100897 131667 100963 131670
rect 136961 131730 137027 131733
rect 136961 131728 140076 131730
rect 136961 131672 136966 131728
rect 137022 131672 140076 131728
rect 169670 131700 169730 131806
rect 172657 131803 172723 131806
rect 136961 131670 140076 131672
rect 136961 131667 137027 131670
rect 63637 131594 63703 131597
rect 60772 131592 63703 131594
rect 60772 131536 63642 131592
rect 63698 131536 63703 131592
rect 60772 131534 63703 131536
rect 63637 131531 63703 131534
rect 102093 131594 102159 131597
rect 135121 131594 135187 131597
rect 102093 131592 104932 131594
rect 102093 131536 102098 131592
rect 102154 131536 104932 131592
rect 102093 131534 104932 131536
rect 132716 131592 135187 131594
rect 132716 131536 135126 131592
rect 135182 131536 135187 131592
rect 132716 131534 135187 131536
rect 102093 131531 102159 131534
rect 135121 131531 135187 131534
rect 175325 131594 175391 131597
rect 175325 131592 177060 131594
rect 175325 131536 175330 131592
rect 175386 131536 177060 131592
rect 175325 131534 177060 131536
rect 175325 131531 175391 131534
rect 63545 131322 63611 131325
rect 135305 131322 135371 131325
rect 60742 131320 63611 131322
rect 60742 131264 63550 131320
rect 63606 131264 63611 131320
rect 60742 131262 63611 131264
rect 60742 131088 60802 131262
rect 63545 131259 63611 131262
rect 132686 131320 135371 131322
rect 132686 131264 135310 131320
rect 135366 131264 135371 131320
rect 132686 131262 135371 131264
rect 66305 131186 66371 131189
rect 66305 131184 67948 131186
rect 66305 131128 66310 131184
rect 66366 131128 67948 131184
rect 66305 131126 67948 131128
rect 66305 131123 66371 131126
rect 132686 131088 132746 131262
rect 135305 131259 135371 131262
rect 174865 131322 174931 131325
rect 174865 131320 177090 131322
rect 174865 131264 174870 131320
rect 174926 131264 177090 131320
rect 174865 131262 177090 131264
rect 174865 131259 174931 131262
rect 62809 130778 62875 130781
rect 60742 130776 62875 130778
rect 60742 130720 62814 130776
rect 62870 130720 62875 130776
rect 60742 130718 62875 130720
rect 60742 130544 60802 130718
rect 62809 130715 62875 130718
rect 97726 130642 97786 131088
rect 102185 131050 102251 131053
rect 102185 131048 104932 131050
rect 102185 130992 102190 131048
rect 102246 130992 104932 131048
rect 102185 130990 104932 130992
rect 102185 130987 102251 130990
rect 135305 130778 135371 130781
rect 132686 130776 135371 130778
rect 132686 130720 135310 130776
rect 135366 130720 135371 130776
rect 132686 130718 135371 130720
rect 100437 130642 100503 130645
rect 97726 130640 100503 130642
rect 97726 130584 100442 130640
rect 100498 130584 100503 130640
rect 97726 130582 100503 130584
rect 100437 130579 100503 130582
rect 132686 130544 132746 130718
rect 135305 130715 135371 130718
rect 136869 130642 136935 130645
rect 140046 130642 140106 131088
rect 169854 130778 169914 131156
rect 177030 131088 177090 131262
rect 172657 130778 172723 130781
rect 169854 130776 172723 130778
rect 169854 130720 172662 130776
rect 172718 130720 172723 130776
rect 169854 130718 172723 130720
rect 172657 130715 172723 130718
rect 175417 130778 175483 130781
rect 175417 130776 177090 130778
rect 175417 130720 175422 130776
rect 175478 130720 177090 130776
rect 175417 130718 177090 130720
rect 175417 130715 175483 130718
rect 136869 130640 140106 130642
rect 136869 130584 136874 130640
rect 136930 130584 140106 130640
rect 136869 130582 140106 130584
rect 136869 130579 136935 130582
rect 177030 130544 177090 130718
rect 66397 130506 66463 130509
rect 100897 130506 100963 130509
rect 66397 130504 67948 130506
rect 66397 130448 66402 130504
rect 66458 130448 67948 130504
rect 66397 130446 67948 130448
rect 97756 130504 100963 130506
rect 97756 130448 100902 130504
rect 100958 130448 100963 130504
rect 97756 130446 100963 130448
rect 66397 130443 66463 130446
rect 100897 130443 100963 130446
rect 102369 130506 102435 130509
rect 136961 130506 137027 130509
rect 102369 130504 104932 130506
rect 102369 130448 102374 130504
rect 102430 130448 104932 130504
rect 102369 130446 104932 130448
rect 136961 130504 140076 130506
rect 136961 130448 136966 130504
rect 137022 130448 140076 130504
rect 136961 130446 140076 130448
rect 102369 130443 102435 130446
rect 136961 130443 137027 130446
rect 169854 130370 169914 130476
rect 172657 130370 172723 130373
rect 169854 130368 172723 130370
rect 169854 130312 172662 130368
rect 172718 130312 172723 130368
rect 169854 130310 172723 130312
rect 172657 130307 172723 130310
rect 63453 130234 63519 130237
rect 135213 130234 135279 130237
rect 60742 130232 63519 130234
rect 60742 130176 63458 130232
rect 63514 130176 63519 130232
rect 60742 130174 63519 130176
rect 60742 129864 60802 130174
rect 63453 130171 63519 130174
rect 132686 130232 135279 130234
rect 132686 130176 135218 130232
rect 135274 130176 135279 130232
rect 132686 130174 135279 130176
rect 65477 129962 65543 129965
rect 65477 129960 67948 129962
rect 65477 129904 65482 129960
rect 65538 129904 67948 129960
rect 65477 129902 67948 129904
rect 65477 129899 65543 129902
rect 132686 129864 132746 130174
rect 135213 130171 135279 130174
rect 175233 130234 175299 130237
rect 175233 130232 177090 130234
rect 175233 130176 175238 130232
rect 175294 130176 177090 130232
rect 175233 130174 177090 130176
rect 175233 130171 175299 130174
rect 63269 129554 63335 129557
rect 60742 129552 63335 129554
rect 60742 129496 63274 129552
rect 63330 129496 63335 129552
rect 60742 129494 63335 129496
rect 60742 129320 60802 129494
rect 63269 129491 63335 129494
rect 97726 129418 97786 129864
rect 102369 129826 102435 129829
rect 102369 129824 104932 129826
rect 102369 129768 102374 129824
rect 102430 129768 104932 129824
rect 102369 129766 104932 129768
rect 102369 129763 102435 129766
rect 134937 129554 135003 129557
rect 132686 129552 135003 129554
rect 132686 129496 134942 129552
rect 134998 129496 135003 129552
rect 132686 129494 135003 129496
rect 100069 129418 100135 129421
rect 97726 129416 100135 129418
rect 97726 129360 100074 129416
rect 100130 129360 100135 129416
rect 97726 129358 100135 129360
rect 100069 129355 100135 129358
rect 132686 129320 132746 129494
rect 134937 129491 135003 129494
rect 136961 129418 137027 129421
rect 140046 129418 140106 129864
rect 169854 129554 169914 129932
rect 177030 129864 177090 130174
rect 171829 129554 171895 129557
rect 169854 129552 171895 129554
rect 169854 129496 171834 129552
rect 171890 129496 171895 129552
rect 169854 129494 171895 129496
rect 171829 129491 171895 129494
rect 175141 129554 175207 129557
rect 175141 129552 177090 129554
rect 175141 129496 175146 129552
rect 175202 129496 177090 129552
rect 175141 129494 177090 129496
rect 175141 129491 175207 129494
rect 136961 129416 140106 129418
rect 136961 129360 136966 129416
rect 137022 129360 140106 129416
rect 136961 129358 140106 129360
rect 136961 129355 137027 129358
rect 177030 129320 177090 129494
rect 66397 129282 66463 129285
rect 102001 129282 102067 129285
rect 66397 129280 67948 129282
rect 66397 129224 66402 129280
rect 66458 129224 67948 129280
rect 66397 129222 67948 129224
rect 102001 129280 104932 129282
rect 102001 129224 102006 129280
rect 102062 129224 104932 129280
rect 102001 129222 104932 129224
rect 66397 129219 66463 129222
rect 102001 129219 102067 129222
rect 97726 129010 97786 129184
rect 100897 129010 100963 129013
rect 97726 129008 100963 129010
rect 97726 128952 100902 129008
rect 100958 128952 100963 129008
rect 97726 128950 100963 128952
rect 100897 128947 100963 128950
rect 136869 129010 136935 129013
rect 140046 129010 140106 129184
rect 169854 129146 169914 129252
rect 171829 129146 171895 129149
rect 169854 129144 171895 129146
rect 169854 129088 171834 129144
rect 171890 129088 171895 129144
rect 169854 129086 171895 129088
rect 171829 129083 171895 129086
rect 136869 129008 140106 129010
rect 136869 128952 136874 129008
rect 136930 128952 140106 129008
rect 136869 128950 140106 128952
rect 136869 128947 136935 128950
rect 62717 128738 62783 128741
rect 60772 128736 62783 128738
rect 60772 128680 62722 128736
rect 62778 128680 62783 128736
rect 102277 128738 102343 128741
rect 135397 128738 135463 128741
rect 102277 128736 104932 128738
rect 60772 128678 62783 128680
rect 62717 128675 62783 128678
rect 62625 128466 62691 128469
rect 60742 128464 62691 128466
rect 60742 128408 62630 128464
rect 62686 128408 62691 128464
rect 60742 128406 62691 128408
rect 60742 128232 60802 128406
rect 62625 128403 62691 128406
rect 67918 128330 67978 128708
rect 102277 128680 102282 128736
rect 102338 128680 104932 128736
rect 102277 128678 104932 128680
rect 132716 128736 135463 128738
rect 132716 128680 135402 128736
rect 135458 128680 135463 128736
rect 174221 128738 174287 128741
rect 174221 128736 177060 128738
rect 132716 128678 135463 128680
rect 102277 128675 102343 128678
rect 135397 128675 135463 128678
rect 66262 128270 67978 128330
rect 97726 128330 97786 128640
rect 135029 128466 135095 128469
rect 132686 128464 135095 128466
rect 132686 128408 135034 128464
rect 135090 128408 135095 128464
rect 132686 128406 135095 128408
rect 100345 128330 100411 128333
rect 97726 128328 100411 128330
rect 97726 128272 100350 128328
rect 100406 128272 100411 128328
rect 97726 128270 100411 128272
rect 65017 127922 65083 127925
rect 66262 127922 66322 128270
rect 100345 128267 100411 128270
rect 132686 128232 132746 128406
rect 135029 128403 135095 128406
rect 136777 128330 136843 128333
rect 140046 128330 140106 128640
rect 136777 128328 140106 128330
rect 136777 128272 136782 128328
rect 136838 128272 140106 128328
rect 136777 128270 140106 128272
rect 169854 128330 169914 128708
rect 174221 128680 174226 128736
rect 174282 128680 177060 128736
rect 174221 128678 177060 128680
rect 174221 128675 174287 128678
rect 174313 128466 174379 128469
rect 174313 128464 177090 128466
rect 174313 128408 174318 128464
rect 174374 128408 177090 128464
rect 174313 128406 177090 128408
rect 174313 128403 174379 128406
rect 172565 128330 172631 128333
rect 169854 128328 172631 128330
rect 169854 128272 172570 128328
rect 172626 128272 172631 128328
rect 169854 128270 172631 128272
rect 136777 128267 136843 128270
rect 172565 128267 172631 128270
rect 177030 128232 177090 128406
rect 66397 128194 66463 128197
rect 102185 128194 102251 128197
rect 66397 128192 67948 128194
rect 66397 128136 66402 128192
rect 66458 128136 67948 128192
rect 66397 128134 67948 128136
rect 102185 128192 104932 128194
rect 102185 128136 102190 128192
rect 102246 128136 104932 128192
rect 102185 128134 104932 128136
rect 66397 128131 66463 128134
rect 102185 128131 102251 128134
rect 65017 127920 66322 127922
rect 65017 127864 65022 127920
rect 65078 127864 66322 127920
rect 65017 127862 66322 127864
rect 65017 127859 65083 127862
rect 9896 127786 10376 127816
rect 12117 127786 12183 127789
rect 9896 127784 12183 127786
rect 9896 127728 12122 127784
rect 12178 127728 12183 127784
rect 9896 127726 12183 127728
rect 9896 127696 10376 127726
rect 12117 127723 12183 127726
rect 30425 127786 30491 127789
rect 30425 127784 32988 127786
rect 30425 127728 30430 127784
rect 30486 127728 32988 127784
rect 30425 127726 32988 127728
rect 30425 127723 30491 127726
rect 97726 127650 97786 128096
rect 100529 127650 100595 127653
rect 97726 127648 100595 127650
rect 97726 127592 100534 127648
rect 100590 127592 100595 127648
rect 97726 127590 100595 127592
rect 100529 127587 100595 127590
rect 136869 127650 136935 127653
rect 140046 127650 140106 128096
rect 169854 127922 169914 128164
rect 171553 127922 171619 127925
rect 169854 127920 171619 127922
rect 169854 127864 171558 127920
rect 171614 127864 171619 127920
rect 169854 127862 171619 127864
rect 171553 127859 171619 127862
rect 207985 127786 208051 127789
rect 204844 127784 208051 127786
rect 204844 127728 207990 127784
rect 208046 127728 208051 127784
rect 204844 127726 208051 127728
rect 207985 127723 208051 127726
rect 136869 127648 140106 127650
rect 136869 127592 136874 127648
rect 136930 127592 140106 127648
rect 136869 127590 140106 127592
rect 136869 127587 136935 127590
rect 62809 127514 62875 127517
rect 60772 127512 62875 127514
rect 60772 127456 62814 127512
rect 62870 127456 62875 127512
rect 102093 127514 102159 127517
rect 135121 127514 135187 127517
rect 102093 127512 104932 127514
rect 60772 127454 62875 127456
rect 62809 127451 62875 127454
rect 62901 127242 62967 127245
rect 60742 127240 62967 127242
rect 60742 127184 62906 127240
rect 62962 127184 62967 127240
rect 60742 127182 62967 127184
rect 60742 127008 60802 127182
rect 62901 127179 62967 127182
rect 67918 127106 67978 127484
rect 102093 127456 102098 127512
rect 102154 127456 104932 127512
rect 102093 127454 104932 127456
rect 132716 127512 135187 127514
rect 132716 127456 135126 127512
rect 135182 127456 135187 127512
rect 174129 127514 174195 127517
rect 174129 127512 177060 127514
rect 132716 127454 135187 127456
rect 102093 127451 102159 127454
rect 135121 127451 135187 127454
rect 66078 127046 67978 127106
rect 97726 127106 97786 127416
rect 135305 127242 135371 127245
rect 132686 127240 135371 127242
rect 132686 127184 135310 127240
rect 135366 127184 135371 127240
rect 132686 127182 135371 127184
rect 100437 127106 100503 127109
rect 97726 127104 100503 127106
rect 97726 127048 100442 127104
rect 100498 127048 100503 127104
rect 97726 127046 100503 127048
rect 62809 126698 62875 126701
rect 60742 126696 62875 126698
rect 60742 126640 62814 126696
rect 62870 126640 62875 126696
rect 60742 126638 62875 126640
rect 60742 126464 60802 126638
rect 62809 126635 62875 126638
rect 65017 126562 65083 126565
rect 66078 126562 66138 127046
rect 100437 127043 100503 127046
rect 132686 127008 132746 127182
rect 135305 127179 135371 127182
rect 136777 127106 136843 127109
rect 140046 127106 140106 127416
rect 136777 127104 140106 127106
rect 136777 127048 136782 127104
rect 136838 127048 140106 127104
rect 136777 127046 140106 127048
rect 169854 127106 169914 127484
rect 174129 127456 174134 127512
rect 174190 127456 177060 127512
rect 174129 127454 177060 127456
rect 174129 127451 174195 127454
rect 174497 127242 174563 127245
rect 174497 127240 177090 127242
rect 174497 127184 174502 127240
rect 174558 127184 177090 127240
rect 174497 127182 177090 127184
rect 174497 127179 174563 127182
rect 172013 127106 172079 127109
rect 169854 127104 172079 127106
rect 169854 127048 172018 127104
rect 172074 127048 172079 127104
rect 169854 127046 172079 127048
rect 136777 127043 136843 127046
rect 172013 127043 172079 127046
rect 177030 127008 177090 127182
rect 66305 126970 66371 126973
rect 102185 126970 102251 126973
rect 66305 126968 67948 126970
rect 66305 126912 66310 126968
rect 66366 126912 67948 126968
rect 66305 126910 67948 126912
rect 102185 126968 104932 126970
rect 102185 126912 102190 126968
rect 102246 126912 104932 126968
rect 102185 126910 104932 126912
rect 66305 126907 66371 126910
rect 102185 126907 102251 126910
rect 65017 126560 66138 126562
rect 65017 126504 65022 126560
rect 65078 126504 66138 126560
rect 65017 126502 66138 126504
rect 65017 126499 65083 126502
rect 97726 126426 97786 126872
rect 134661 126698 134727 126701
rect 132686 126696 134727 126698
rect 132686 126640 134666 126696
rect 134722 126640 134727 126696
rect 132686 126638 134727 126640
rect 132686 126464 132746 126638
rect 134661 126635 134727 126638
rect 100897 126426 100963 126429
rect 97726 126424 100963 126426
rect 97726 126368 100902 126424
rect 100958 126368 100963 126424
rect 97726 126366 100963 126368
rect 100897 126363 100963 126366
rect 102277 126426 102343 126429
rect 136869 126426 136935 126429
rect 140046 126426 140106 126872
rect 169854 126698 169914 126940
rect 172197 126698 172263 126701
rect 169854 126696 172263 126698
rect 169854 126640 172202 126696
rect 172258 126640 172263 126696
rect 169854 126638 172263 126640
rect 172197 126635 172263 126638
rect 174221 126698 174287 126701
rect 174221 126696 177090 126698
rect 174221 126640 174226 126696
rect 174282 126640 177090 126696
rect 174221 126638 177090 126640
rect 174221 126635 174287 126638
rect 177030 126464 177090 126638
rect 102277 126424 104932 126426
rect 102277 126368 102282 126424
rect 102338 126368 104932 126424
rect 102277 126366 104932 126368
rect 136869 126424 140106 126426
rect 136869 126368 136874 126424
rect 136930 126368 140106 126424
rect 136869 126366 140106 126368
rect 102277 126363 102343 126366
rect 136869 126363 136935 126366
rect 66397 126290 66463 126293
rect 100805 126290 100871 126293
rect 66397 126288 67948 126290
rect 66397 126232 66402 126288
rect 66458 126232 67948 126288
rect 66397 126230 67948 126232
rect 97756 126288 100871 126290
rect 97756 126232 100810 126288
rect 100866 126232 100871 126288
rect 97756 126230 100871 126232
rect 66397 126227 66463 126230
rect 100805 126227 100871 126230
rect 136961 126290 137027 126293
rect 136961 126288 140076 126290
rect 136961 126232 136966 126288
rect 137022 126232 140076 126288
rect 136961 126230 140076 126232
rect 136961 126227 137027 126230
rect 169854 126154 169914 126260
rect 172657 126154 172723 126157
rect 169854 126152 172723 126154
rect 169854 126096 172662 126152
rect 172718 126096 172723 126152
rect 169854 126094 172723 126096
rect 172657 126091 172723 126094
rect 62625 126018 62691 126021
rect 135213 126018 135279 126021
rect 60742 126016 62691 126018
rect 60742 125960 62630 126016
rect 62686 125960 62691 126016
rect 60742 125958 62691 125960
rect 60742 125784 60802 125958
rect 62625 125955 62691 125958
rect 132686 126016 135279 126018
rect 132686 125960 135218 126016
rect 135274 125960 135279 126016
rect 132686 125958 135279 125960
rect 132686 125784 132746 125958
rect 135213 125955 135279 125958
rect 174589 126018 174655 126021
rect 174589 126016 177090 126018
rect 174589 125960 174594 126016
rect 174650 125960 177090 126016
rect 174589 125958 177090 125960
rect 174589 125955 174655 125958
rect 177030 125784 177090 125958
rect 66305 125746 66371 125749
rect 102001 125746 102067 125749
rect 66305 125744 67948 125746
rect 66305 125688 66310 125744
rect 66366 125688 67948 125744
rect 66305 125686 67948 125688
rect 102001 125744 104932 125746
rect 102001 125688 102006 125744
rect 102062 125688 104932 125744
rect 102001 125686 104932 125688
rect 66305 125683 66371 125686
rect 102001 125683 102067 125686
rect 62809 125474 62875 125477
rect 60742 125472 62875 125474
rect 60742 125416 62814 125472
rect 62870 125416 62875 125472
rect 60742 125414 62875 125416
rect 60742 125240 60802 125414
rect 62809 125411 62875 125414
rect 97726 125338 97786 125648
rect 135397 125474 135463 125477
rect 132686 125472 135463 125474
rect 132686 125416 135402 125472
rect 135458 125416 135463 125472
rect 132686 125414 135463 125416
rect 100897 125338 100963 125341
rect 97726 125336 100963 125338
rect 97726 125280 100902 125336
rect 100958 125280 100963 125336
rect 97726 125278 100963 125280
rect 100897 125275 100963 125278
rect 132686 125240 132746 125414
rect 135397 125411 135463 125414
rect 136777 125338 136843 125341
rect 140046 125338 140106 125648
rect 136777 125336 140106 125338
rect 136777 125280 136782 125336
rect 136838 125280 140106 125336
rect 136777 125278 140106 125280
rect 169854 125338 169914 125716
rect 174129 125474 174195 125477
rect 174129 125472 177090 125474
rect 174129 125416 174134 125472
rect 174190 125416 177090 125472
rect 174129 125414 177090 125416
rect 174129 125411 174195 125414
rect 171829 125338 171895 125341
rect 169854 125336 171895 125338
rect 169854 125280 171834 125336
rect 171890 125280 171895 125336
rect 169854 125278 171895 125280
rect 136777 125275 136843 125278
rect 171829 125275 171895 125278
rect 177030 125240 177090 125414
rect 66397 125202 66463 125205
rect 102369 125202 102435 125205
rect 66397 125200 67948 125202
rect 66397 125144 66402 125200
rect 66458 125144 67948 125200
rect 66397 125142 67948 125144
rect 102369 125200 104932 125202
rect 102369 125144 102374 125200
rect 102430 125144 104932 125200
rect 102369 125142 104932 125144
rect 66397 125139 66463 125142
rect 102369 125139 102435 125142
rect 97726 124930 97786 125104
rect 100805 124930 100871 124933
rect 97726 124928 100871 124930
rect 97726 124872 100810 124928
rect 100866 124872 100871 124928
rect 97726 124870 100871 124872
rect 100805 124867 100871 124870
rect 136869 124930 136935 124933
rect 140046 124930 140106 125104
rect 169854 125066 169914 125172
rect 172197 125066 172263 125069
rect 169854 125064 172263 125066
rect 169854 125008 172202 125064
rect 172258 125008 172263 125064
rect 169854 125006 172263 125008
rect 172197 125003 172263 125006
rect 136869 124928 140106 124930
rect 136869 124872 136874 124928
rect 136930 124872 140106 124928
rect 136869 124870 140106 124872
rect 136869 124867 136935 124870
rect 65017 124794 65083 124797
rect 66305 124794 66371 124797
rect 65017 124792 66371 124794
rect 65017 124736 65022 124792
rect 65078 124736 66310 124792
rect 66366 124736 66371 124792
rect 65017 124734 66371 124736
rect 65017 124731 65083 124734
rect 66305 124731 66371 124734
rect 62717 124658 62783 124661
rect 60772 124656 62783 124658
rect 60772 124600 62722 124656
rect 62778 124600 62783 124656
rect 60772 124598 62783 124600
rect 62717 124595 62783 124598
rect 102277 124658 102343 124661
rect 135305 124658 135371 124661
rect 102277 124656 104932 124658
rect 102277 124600 102282 124656
rect 102338 124600 104932 124656
rect 102277 124598 104932 124600
rect 132716 124656 135371 124658
rect 132716 124600 135310 124656
rect 135366 124600 135371 124656
rect 132716 124598 135371 124600
rect 102277 124595 102343 124598
rect 135305 124595 135371 124598
rect 174313 124658 174379 124661
rect 174313 124656 177060 124658
rect 174313 124600 174318 124656
rect 174374 124600 177060 124656
rect 174313 124598 177060 124600
rect 174313 124595 174379 124598
rect 62901 124386 62967 124389
rect 60742 124384 62967 124386
rect 60742 124328 62906 124384
rect 62962 124328 62967 124384
rect 60742 124326 62967 124328
rect 60742 124016 60802 124326
rect 62901 124323 62967 124326
rect 67918 124114 67978 124492
rect 66262 124054 67978 124114
rect 97726 124114 97786 124424
rect 135029 124386 135095 124389
rect 132686 124384 135095 124386
rect 132686 124328 135034 124384
rect 135090 124328 135095 124384
rect 132686 124326 135095 124328
rect 100253 124114 100319 124117
rect 97726 124112 100319 124114
rect 97726 124056 100258 124112
rect 100314 124056 100319 124112
rect 97726 124054 100319 124056
rect 62809 123706 62875 123709
rect 60742 123704 62875 123706
rect 60742 123648 62814 123704
rect 62870 123648 62875 123704
rect 60742 123646 62875 123648
rect 60742 123472 60802 123646
rect 62809 123643 62875 123646
rect 65017 123706 65083 123709
rect 66262 123706 66322 124054
rect 100253 124051 100319 124054
rect 132686 124016 132746 124326
rect 135029 124323 135095 124326
rect 136777 124114 136843 124117
rect 140046 124114 140106 124424
rect 136777 124112 140106 124114
rect 136777 124056 136782 124112
rect 136838 124056 140106 124112
rect 136777 124054 140106 124056
rect 169854 124114 169914 124492
rect 174497 124386 174563 124389
rect 174497 124384 177090 124386
rect 174497 124328 174502 124384
rect 174558 124328 177090 124384
rect 174497 124326 177090 124328
rect 174497 124323 174563 124326
rect 171829 124114 171895 124117
rect 169854 124112 171895 124114
rect 169854 124056 171834 124112
rect 171890 124056 171895 124112
rect 169854 124054 171895 124056
rect 136777 124051 136843 124054
rect 171829 124051 171895 124054
rect 177030 124016 177090 124326
rect 66397 123978 66463 123981
rect 102093 123978 102159 123981
rect 66397 123976 67948 123978
rect 66397 123920 66402 123976
rect 66458 123920 67948 123976
rect 66397 123918 67948 123920
rect 102093 123976 104932 123978
rect 102093 123920 102098 123976
rect 102154 123920 104932 123976
rect 102093 123918 104932 123920
rect 66397 123915 66463 123918
rect 102093 123915 102159 123918
rect 65017 123704 66322 123706
rect 65017 123648 65022 123704
rect 65078 123648 66322 123704
rect 65017 123646 66322 123648
rect 65017 123643 65083 123646
rect 97726 123434 97786 123880
rect 135213 123706 135279 123709
rect 132686 123704 135279 123706
rect 132686 123648 135218 123704
rect 135274 123648 135279 123704
rect 132686 123646 135279 123648
rect 101950 123570 101956 123572
rect 101774 123510 101956 123570
rect 100897 123434 100963 123437
rect 101774 123436 101834 123510
rect 101950 123508 101956 123510
rect 102020 123508 102026 123572
rect 132686 123472 132746 123646
rect 135213 123643 135279 123646
rect 97726 123432 100963 123434
rect 97726 123376 100902 123432
rect 100958 123376 100963 123432
rect 97726 123374 100963 123376
rect 100897 123371 100963 123374
rect 101766 123372 101772 123436
rect 101836 123372 101842 123436
rect 102369 123434 102435 123437
rect 136869 123434 136935 123437
rect 140046 123434 140106 123880
rect 169854 123706 169914 123948
rect 172565 123706 172631 123709
rect 169854 123704 172631 123706
rect 169854 123648 172570 123704
rect 172626 123648 172631 123704
rect 169854 123646 172631 123648
rect 172565 123643 172631 123646
rect 174221 123706 174287 123709
rect 174221 123704 177090 123706
rect 174221 123648 174226 123704
rect 174282 123648 177090 123704
rect 174221 123646 177090 123648
rect 174221 123643 174287 123646
rect 177030 123472 177090 123646
rect 102369 123432 104932 123434
rect 102369 123376 102374 123432
rect 102430 123376 104932 123432
rect 102369 123374 104932 123376
rect 136869 123432 140106 123434
rect 136869 123376 136874 123432
rect 136930 123376 140106 123432
rect 136869 123374 140106 123376
rect 102369 123371 102435 123374
rect 136869 123371 136935 123374
rect 62625 123162 62691 123165
rect 60742 123160 62691 123162
rect 60742 123104 62630 123160
rect 62686 123104 62691 123160
rect 60742 123102 62691 123104
rect 60742 122928 60802 123102
rect 62625 123099 62691 123102
rect 67918 122890 67978 123268
rect 66078 122830 67978 122890
rect 97726 122890 97786 123200
rect 101766 123168 101772 123232
rect 101836 123168 101842 123232
rect 101774 123029 101834 123168
rect 135121 123162 135187 123165
rect 132686 123160 135187 123162
rect 132686 123104 135126 123160
rect 135182 123104 135187 123160
rect 132686 123102 135187 123104
rect 101774 123024 101883 123029
rect 101774 122968 101822 123024
rect 101878 122968 101883 123024
rect 101774 122966 101883 122968
rect 101817 122963 101883 122966
rect 132686 122928 132746 123102
rect 135121 123099 135187 123102
rect 100161 122890 100227 122893
rect 97726 122888 100227 122890
rect 97726 122832 100166 122888
rect 100222 122832 100227 122888
rect 97726 122830 100227 122832
rect 62809 122618 62875 122621
rect 60742 122616 62875 122618
rect 60742 122560 62814 122616
rect 62870 122560 62875 122616
rect 60742 122558 62875 122560
rect 60742 122384 60802 122558
rect 62809 122555 62875 122558
rect 65017 122482 65083 122485
rect 66078 122482 66138 122830
rect 100161 122827 100227 122830
rect 102185 122890 102251 122893
rect 136869 122890 136935 122893
rect 140046 122890 140106 123200
rect 102185 122888 104932 122890
rect 102185 122832 102190 122888
rect 102246 122832 104932 122888
rect 102185 122830 104932 122832
rect 136869 122888 140106 122890
rect 136869 122832 136874 122888
rect 136930 122832 140106 122888
rect 136869 122830 140106 122832
rect 169854 122890 169914 123268
rect 174589 123162 174655 123165
rect 174589 123160 177090 123162
rect 174589 123104 174594 123160
rect 174650 123104 177090 123160
rect 174589 123102 177090 123104
rect 174589 123099 174655 123102
rect 177030 122928 177090 123102
rect 171829 122890 171895 122893
rect 169854 122888 171895 122890
rect 169854 122832 171834 122888
rect 171890 122832 171895 122888
rect 169854 122830 171895 122832
rect 102185 122827 102251 122830
rect 136869 122827 136935 122830
rect 171829 122827 171895 122830
rect 66305 122754 66371 122757
rect 66305 122752 67948 122754
rect 66305 122696 66310 122752
rect 66366 122696 67948 122752
rect 66305 122694 67948 122696
rect 66305 122691 66371 122694
rect 65017 122480 66138 122482
rect 65017 122424 65022 122480
rect 65078 122424 66138 122480
rect 65017 122422 66138 122424
rect 97726 122482 97786 122656
rect 135305 122618 135371 122621
rect 132686 122616 135371 122618
rect 132686 122560 135310 122616
rect 135366 122560 135371 122616
rect 132686 122558 135371 122560
rect 100621 122482 100687 122485
rect 97726 122480 100687 122482
rect 97726 122424 100626 122480
rect 100682 122424 100687 122480
rect 97726 122422 100687 122424
rect 65017 122419 65083 122422
rect 100621 122419 100687 122422
rect 132686 122384 132746 122558
rect 135305 122555 135371 122558
rect 136961 122482 137027 122485
rect 140046 122482 140106 122656
rect 136961 122480 140106 122482
rect 136961 122424 136966 122480
rect 137022 122424 140106 122480
rect 136961 122422 140106 122424
rect 169854 122482 169914 122724
rect 174129 122618 174195 122621
rect 174129 122616 177090 122618
rect 174129 122560 174134 122616
rect 174190 122560 177090 122616
rect 174129 122558 177090 122560
rect 174129 122555 174195 122558
rect 172013 122482 172079 122485
rect 169854 122480 172079 122482
rect 169854 122424 172018 122480
rect 172074 122424 172079 122480
rect 169854 122422 172079 122424
rect 136961 122419 137027 122422
rect 172013 122419 172079 122422
rect 177030 122384 177090 122558
rect 102277 122346 102343 122349
rect 102277 122344 104932 122346
rect 102277 122288 102282 122344
rect 102338 122288 104932 122344
rect 102277 122286 104932 122288
rect 102277 122283 102343 122286
rect 66397 122210 66463 122213
rect 100897 122210 100963 122213
rect 66397 122208 67948 122210
rect 66397 122152 66402 122208
rect 66458 122152 67948 122208
rect 66397 122150 67948 122152
rect 97756 122208 100963 122210
rect 97756 122152 100902 122208
rect 100958 122152 100963 122208
rect 97756 122150 100963 122152
rect 66397 122147 66463 122150
rect 100897 122147 100963 122150
rect 137053 122210 137119 122213
rect 137053 122208 140076 122210
rect 137053 122152 137058 122208
rect 137114 122152 140076 122208
rect 137053 122150 140076 122152
rect 137053 122147 137119 122150
rect 169854 122074 169914 122180
rect 172657 122074 172723 122077
rect 169854 122072 172723 122074
rect 169854 122016 172662 122072
rect 172718 122016 172723 122072
rect 169854 122014 172723 122016
rect 172657 122011 172723 122014
rect 135397 121938 135463 121941
rect 132686 121936 135463 121938
rect 132686 121880 135402 121936
rect 135458 121880 135463 121936
rect 132686 121878 135463 121880
rect 132686 121704 132746 121878
rect 135397 121875 135463 121878
rect 63545 121666 63611 121669
rect 60772 121664 63611 121666
rect 60772 121608 63550 121664
rect 63606 121608 63611 121664
rect 60772 121606 63611 121608
rect 63545 121603 63611 121606
rect 102369 121666 102435 121669
rect 175325 121666 175391 121669
rect 102369 121664 104932 121666
rect 102369 121608 102374 121664
rect 102430 121608 104932 121664
rect 102369 121606 104932 121608
rect 175325 121664 177060 121666
rect 175325 121608 175330 121664
rect 175386 121608 177060 121664
rect 175325 121606 177060 121608
rect 102369 121603 102435 121606
rect 175325 121603 175391 121606
rect 62809 121394 62875 121397
rect 60742 121392 62875 121394
rect 60742 121336 62814 121392
rect 62870 121336 62875 121392
rect 60742 121334 62875 121336
rect 60742 121160 60802 121334
rect 62809 121331 62875 121334
rect 67918 121122 67978 121500
rect 66078 121062 67978 121122
rect 97726 121122 97786 121432
rect 135305 121394 135371 121397
rect 132686 121392 135371 121394
rect 132686 121336 135310 121392
rect 135366 121336 135371 121392
rect 132686 121334 135371 121336
rect 132686 121160 132746 121334
rect 135305 121331 135371 121334
rect 100069 121122 100135 121125
rect 97726 121120 100135 121122
rect 97726 121064 100074 121120
rect 100130 121064 100135 121120
rect 97726 121062 100135 121064
rect 65017 120714 65083 120717
rect 66078 120714 66138 121062
rect 100069 121059 100135 121062
rect 102277 121122 102343 121125
rect 136777 121122 136843 121125
rect 140046 121122 140106 121432
rect 102277 121120 104932 121122
rect 102277 121064 102282 121120
rect 102338 121064 104932 121120
rect 102277 121062 104932 121064
rect 136777 121120 140106 121122
rect 136777 121064 136782 121120
rect 136838 121064 140106 121120
rect 136777 121062 140106 121064
rect 169854 121122 169914 121500
rect 175049 121394 175115 121397
rect 175049 121392 177090 121394
rect 175049 121336 175054 121392
rect 175110 121336 177090 121392
rect 175049 121334 177090 121336
rect 175049 121331 175115 121334
rect 177030 121160 177090 121334
rect 172105 121122 172171 121125
rect 169854 121120 172171 121122
rect 169854 121064 172110 121120
rect 172166 121064 172171 121120
rect 169854 121062 172171 121064
rect 102277 121059 102343 121062
rect 136777 121059 136843 121062
rect 172105 121059 172171 121062
rect 66213 120986 66279 120989
rect 100897 120986 100963 120989
rect 66213 120984 67948 120986
rect 66213 120928 66218 120984
rect 66274 120928 67948 120984
rect 66213 120926 67948 120928
rect 97756 120984 100963 120986
rect 97756 120928 100902 120984
rect 100958 120928 100963 120984
rect 97756 120926 100963 120928
rect 66213 120923 66279 120926
rect 100897 120923 100963 120926
rect 65017 120712 66138 120714
rect 65017 120656 65022 120712
rect 65078 120656 66138 120712
rect 65017 120654 66138 120656
rect 136961 120714 137027 120717
rect 140046 120714 140106 120888
rect 169854 120850 169914 120956
rect 172657 120850 172723 120853
rect 169854 120848 172723 120850
rect 169854 120792 172662 120848
rect 172718 120792 172723 120848
rect 169854 120790 172723 120792
rect 172657 120787 172723 120790
rect 136961 120712 140106 120714
rect 136961 120656 136966 120712
rect 137022 120656 140106 120712
rect 136961 120654 140106 120656
rect 65017 120651 65083 120654
rect 136961 120651 137027 120654
rect 63453 120578 63519 120581
rect 60772 120576 63519 120578
rect 60772 120520 63458 120576
rect 63514 120520 63519 120576
rect 60772 120518 63519 120520
rect 63453 120515 63519 120518
rect 102093 120578 102159 120581
rect 135213 120578 135279 120581
rect 102093 120576 104932 120578
rect 102093 120520 102098 120576
rect 102154 120520 104932 120576
rect 102093 120518 104932 120520
rect 132716 120576 135279 120578
rect 132716 120520 135218 120576
rect 135274 120520 135279 120576
rect 132716 120518 135279 120520
rect 102093 120515 102159 120518
rect 135213 120515 135279 120518
rect 175417 120578 175483 120581
rect 175417 120576 177060 120578
rect 175417 120520 175422 120576
rect 175478 120520 177060 120576
rect 175417 120518 177060 120520
rect 175417 120515 175483 120518
rect 63637 120306 63703 120309
rect 135121 120306 135187 120309
rect 60742 120304 63703 120306
rect 60742 120248 63642 120304
rect 63698 120248 63703 120304
rect 132686 120304 135187 120306
rect 60742 120246 63703 120248
rect 60742 119936 60802 120246
rect 63637 120243 63703 120246
rect 67918 119898 67978 120276
rect 132686 120248 135126 120304
rect 135182 120248 135187 120304
rect 175141 120306 175207 120309
rect 175141 120304 177090 120306
rect 132686 120246 135187 120248
rect 65342 119838 67978 119898
rect 97726 119898 97786 120208
rect 132686 119936 132746 120246
rect 135121 120243 135187 120246
rect 100437 119898 100503 119901
rect 97726 119896 100503 119898
rect 97726 119840 100442 119896
rect 100498 119840 100503 119896
rect 97726 119838 100503 119840
rect 62809 119626 62875 119629
rect 60742 119624 62875 119626
rect 60742 119568 62814 119624
rect 62870 119568 62875 119624
rect 60742 119566 62875 119568
rect 60742 119392 60802 119566
rect 62809 119563 62875 119566
rect 65017 119490 65083 119493
rect 65342 119490 65402 119838
rect 100437 119835 100503 119838
rect 102001 119898 102067 119901
rect 136777 119898 136843 119901
rect 140046 119898 140106 120208
rect 102001 119896 104932 119898
rect 102001 119840 102006 119896
rect 102062 119840 104932 119896
rect 102001 119838 104932 119840
rect 136777 119896 140106 119898
rect 136777 119840 136782 119896
rect 136838 119840 140106 119896
rect 136777 119838 140106 119840
rect 169854 119898 169914 120276
rect 175141 120248 175146 120304
rect 175202 120248 177090 120304
rect 175141 120246 177090 120248
rect 175141 120243 175207 120246
rect 177030 119936 177090 120246
rect 171829 119898 171895 119901
rect 169854 119896 171895 119898
rect 169854 119840 171834 119896
rect 171890 119840 171895 119896
rect 169854 119838 171895 119840
rect 102001 119835 102067 119838
rect 136777 119835 136843 119838
rect 171829 119835 171895 119838
rect 65477 119762 65543 119765
rect 65477 119760 67948 119762
rect 65477 119704 65482 119760
rect 65538 119704 67948 119760
rect 65477 119702 67948 119704
rect 65477 119699 65543 119702
rect 65017 119488 65402 119490
rect 65017 119432 65022 119488
rect 65078 119432 65402 119488
rect 65017 119430 65402 119432
rect 65017 119427 65083 119430
rect 97726 119354 97786 119664
rect 134845 119626 134911 119629
rect 132686 119624 134911 119626
rect 132686 119568 134850 119624
rect 134906 119568 134911 119624
rect 132686 119566 134911 119568
rect 132686 119392 132746 119566
rect 134845 119563 134911 119566
rect 100897 119354 100963 119357
rect 97726 119352 100963 119354
rect 97726 119296 100902 119352
rect 100958 119296 100963 119352
rect 97726 119294 100963 119296
rect 100897 119291 100963 119294
rect 102369 119354 102435 119357
rect 136869 119354 136935 119357
rect 140046 119354 140106 119664
rect 169854 119626 169914 119732
rect 171829 119626 171895 119629
rect 169854 119624 171895 119626
rect 169854 119568 171834 119624
rect 171890 119568 171895 119624
rect 169854 119566 171895 119568
rect 171829 119563 171895 119566
rect 174313 119626 174379 119629
rect 174313 119624 177090 119626
rect 174313 119568 174318 119624
rect 174374 119568 177090 119624
rect 174313 119566 177090 119568
rect 174313 119563 174379 119566
rect 177030 119392 177090 119566
rect 102369 119352 104932 119354
rect 102369 119296 102374 119352
rect 102430 119296 104932 119352
rect 102369 119294 104932 119296
rect 136869 119352 140106 119354
rect 136869 119296 136874 119352
rect 136930 119296 140106 119352
rect 136869 119294 140106 119296
rect 102369 119291 102435 119294
rect 136869 119291 136935 119294
rect 66397 119218 66463 119221
rect 66397 119216 67948 119218
rect 66397 119160 66402 119216
rect 66458 119160 67948 119216
rect 66397 119158 67948 119160
rect 66397 119155 66463 119158
rect 62717 118810 62783 118813
rect 60772 118808 62783 118810
rect 60772 118752 62722 118808
rect 62778 118752 62783 118808
rect 60772 118750 62783 118752
rect 62717 118747 62783 118750
rect 97726 118674 97786 119120
rect 135305 119082 135371 119085
rect 132686 119080 135371 119082
rect 132686 119024 135310 119080
rect 135366 119024 135371 119080
rect 132686 119022 135371 119024
rect 132686 118848 132746 119022
rect 135305 119019 135371 119022
rect 102185 118810 102251 118813
rect 102185 118808 104932 118810
rect 102185 118752 102190 118808
rect 102246 118752 104932 118808
rect 102185 118750 104932 118752
rect 102185 118747 102251 118750
rect 100621 118674 100687 118677
rect 97726 118672 100687 118674
rect 97726 118616 100626 118672
rect 100682 118616 100687 118672
rect 97726 118614 100687 118616
rect 100621 118611 100687 118614
rect 136961 118674 137027 118677
rect 140046 118674 140106 119120
rect 136961 118672 140106 118674
rect 136961 118616 136966 118672
rect 137022 118616 140106 118672
rect 136961 118614 140106 118616
rect 169854 118674 169914 119188
rect 174221 119082 174287 119085
rect 174221 119080 177090 119082
rect 174221 119024 174226 119080
rect 174282 119024 177090 119080
rect 174221 119022 177090 119024
rect 174221 119019 174287 119022
rect 177030 118848 177090 119022
rect 171829 118674 171895 118677
rect 169854 118672 171895 118674
rect 169854 118616 171834 118672
rect 171890 118616 171895 118672
rect 169854 118614 171895 118616
rect 136961 118611 137027 118614
rect 171829 118611 171895 118614
rect 31846 118476 31852 118540
rect 31916 118538 31922 118540
rect 62809 118538 62875 118541
rect 31916 118478 32988 118538
rect 60742 118536 62875 118538
rect 60742 118480 62814 118536
rect 62870 118480 62875 118536
rect 60742 118478 62875 118480
rect 31916 118476 31922 118478
rect 60742 118304 60802 118478
rect 62809 118475 62875 118478
rect 64925 118538 64991 118541
rect 135305 118538 135371 118541
rect 64925 118536 67948 118538
rect 64925 118480 64930 118536
rect 64986 118480 67948 118536
rect 64925 118478 67948 118480
rect 132686 118536 135371 118538
rect 132686 118480 135310 118536
rect 135366 118480 135371 118536
rect 174129 118538 174195 118541
rect 207893 118538 207959 118541
rect 174129 118536 177090 118538
rect 132686 118478 135371 118480
rect 64925 118475 64991 118478
rect 65017 118266 65083 118269
rect 66397 118266 66463 118269
rect 65017 118264 66463 118266
rect 65017 118208 65022 118264
rect 65078 118208 66402 118264
rect 66458 118208 66463 118264
rect 65017 118206 66463 118208
rect 65017 118203 65083 118206
rect 66397 118203 66463 118206
rect 97726 118130 97786 118440
rect 132686 118304 132746 118478
rect 135305 118475 135371 118478
rect 102277 118266 102343 118269
rect 102277 118264 104932 118266
rect 102277 118208 102282 118264
rect 102338 118208 104932 118264
rect 102277 118206 104932 118208
rect 102277 118203 102343 118206
rect 100253 118130 100319 118133
rect 97726 118128 100319 118130
rect 97726 118072 100258 118128
rect 100314 118072 100319 118128
rect 97726 118070 100319 118072
rect 100253 118067 100319 118070
rect 136777 118130 136843 118133
rect 140046 118130 140106 118440
rect 169854 118266 169914 118508
rect 174129 118480 174134 118536
rect 174190 118480 177090 118536
rect 204844 118536 207959 118538
rect 204844 118508 207898 118536
rect 174129 118478 177090 118480
rect 174129 118475 174195 118478
rect 177030 118304 177090 118478
rect 204814 118480 207898 118508
rect 207954 118480 207959 118536
rect 204814 118478 207959 118480
rect 171645 118266 171711 118269
rect 169854 118264 171711 118266
rect 169854 118208 171650 118264
rect 171706 118208 171711 118264
rect 169854 118206 171711 118208
rect 171645 118203 171711 118206
rect 172657 118130 172723 118133
rect 136777 118128 140106 118130
rect 136777 118072 136782 118128
rect 136838 118072 140106 118128
rect 136777 118070 140106 118072
rect 169670 118128 172723 118130
rect 169670 118072 172662 118128
rect 172718 118072 172723 118128
rect 169670 118070 172723 118072
rect 136777 118067 136843 118070
rect 66397 117994 66463 117997
rect 100529 117994 100595 117997
rect 66397 117992 67948 117994
rect 66397 117936 66402 117992
rect 66458 117936 67948 117992
rect 66397 117934 67948 117936
rect 97756 117992 100595 117994
rect 97756 117936 100534 117992
rect 100590 117936 100595 117992
rect 97756 117934 100595 117936
rect 66397 117931 66463 117934
rect 100529 117931 100595 117934
rect 136869 117994 136935 117997
rect 136869 117992 140076 117994
rect 136869 117936 136874 117992
rect 136930 117936 140076 117992
rect 169670 117964 169730 118070
rect 172657 118067 172723 118070
rect 204673 117994 204739 117997
rect 204814 117994 204874 118478
rect 207893 118475 207959 118478
rect 204673 117992 204874 117994
rect 136869 117934 140076 117936
rect 204673 117936 204678 117992
rect 204734 117936 204874 117992
rect 204673 117934 204874 117936
rect 136869 117931 136935 117934
rect 204673 117931 204739 117934
rect 62901 117858 62967 117861
rect 60742 117856 62967 117858
rect 60742 117800 62906 117856
rect 62962 117800 62967 117856
rect 60742 117798 62967 117800
rect 60742 117624 60802 117798
rect 62901 117795 62967 117798
rect 174497 117858 174563 117861
rect 174497 117856 177090 117858
rect 174497 117800 174502 117856
rect 174558 117800 177090 117856
rect 174497 117798 177090 117800
rect 174497 117795 174563 117798
rect 177030 117624 177090 117798
rect 102369 117586 102435 117589
rect 135213 117586 135279 117589
rect 102369 117584 104932 117586
rect 102369 117528 102374 117584
rect 102430 117528 104932 117584
rect 102369 117526 104932 117528
rect 132716 117584 135279 117586
rect 132716 117528 135218 117584
rect 135274 117528 135279 117584
rect 132716 117526 135279 117528
rect 102369 117523 102435 117526
rect 135213 117523 135279 117526
rect 62809 117314 62875 117317
rect 134109 117314 134175 117317
rect 60742 117312 62875 117314
rect 60742 117256 62814 117312
rect 62870 117256 62875 117312
rect 132686 117312 134175 117314
rect 60742 117254 62875 117256
rect 60742 117080 60802 117254
rect 62809 117251 62875 117254
rect 67918 116906 67978 117284
rect 132686 117256 134114 117312
rect 134170 117256 134175 117312
rect 174037 117314 174103 117317
rect 174037 117312 177090 117314
rect 132686 117254 134175 117256
rect 66262 116846 67978 116906
rect 97726 116906 97786 117216
rect 132686 117080 132746 117254
rect 134109 117251 134175 117254
rect 102277 117042 102343 117045
rect 102277 117040 104932 117042
rect 102277 116984 102282 117040
rect 102338 116984 104932 117040
rect 102277 116982 104932 116984
rect 102277 116979 102343 116982
rect 100897 116906 100963 116909
rect 97726 116904 100963 116906
rect 97726 116848 100902 116904
rect 100958 116848 100963 116904
rect 97726 116846 100963 116848
rect 62809 116770 62875 116773
rect 60742 116768 62875 116770
rect 60742 116712 62814 116768
rect 62870 116712 62875 116768
rect 60742 116710 62875 116712
rect 60742 116536 60802 116710
rect 62809 116707 62875 116710
rect 65017 116498 65083 116501
rect 66262 116498 66322 116846
rect 100897 116843 100963 116846
rect 136777 116906 136843 116909
rect 140046 116906 140106 117216
rect 136777 116904 140106 116906
rect 136777 116848 136782 116904
rect 136838 116848 140106 116904
rect 136777 116846 140106 116848
rect 169854 116906 169914 117284
rect 174037 117256 174042 117312
rect 174098 117256 177090 117312
rect 174037 117254 177090 117256
rect 174037 117251 174103 117254
rect 177030 117080 177090 117254
rect 172657 116906 172723 116909
rect 169854 116904 172723 116906
rect 169854 116848 172662 116904
rect 172718 116848 172723 116904
rect 169854 116846 172723 116848
rect 136777 116843 136843 116846
rect 172657 116843 172723 116846
rect 66397 116770 66463 116773
rect 100253 116770 100319 116773
rect 134661 116770 134727 116773
rect 66397 116768 67948 116770
rect 66397 116712 66402 116768
rect 66458 116712 67948 116768
rect 66397 116710 67948 116712
rect 97756 116768 100319 116770
rect 97756 116712 100258 116768
rect 100314 116712 100319 116768
rect 97756 116710 100319 116712
rect 66397 116707 66463 116710
rect 100253 116707 100319 116710
rect 132686 116768 134727 116770
rect 132686 116712 134666 116768
rect 134722 116712 134727 116768
rect 132686 116710 134727 116712
rect 132686 116536 132746 116710
rect 134661 116707 134727 116710
rect 136869 116770 136935 116773
rect 173945 116770 174011 116773
rect 136869 116768 140076 116770
rect 136869 116712 136874 116768
rect 136930 116712 140076 116768
rect 173945 116768 177090 116770
rect 136869 116710 140076 116712
rect 136869 116707 136935 116710
rect 169854 116634 169914 116740
rect 173945 116712 173950 116768
rect 174006 116712 177090 116768
rect 173945 116710 177090 116712
rect 173945 116707 174011 116710
rect 172565 116634 172631 116637
rect 169854 116632 172631 116634
rect 169854 116576 172570 116632
rect 172626 116576 172631 116632
rect 169854 116574 172631 116576
rect 172565 116571 172631 116574
rect 177030 116536 177090 116710
rect 65017 116496 66322 116498
rect 65017 116440 65022 116496
rect 65078 116440 66322 116496
rect 65017 116438 66322 116440
rect 102461 116498 102527 116501
rect 102461 116496 104932 116498
rect 102461 116440 102466 116496
rect 102522 116440 104932 116496
rect 102461 116438 104932 116440
rect 65017 116435 65083 116438
rect 102461 116435 102527 116438
rect 62717 116226 62783 116229
rect 135121 116226 135187 116229
rect 60742 116224 62783 116226
rect 60742 116168 62722 116224
rect 62778 116168 62783 116224
rect 132686 116224 135187 116226
rect 60742 116166 62783 116168
rect 60742 115856 60802 116166
rect 62717 116163 62783 116166
rect 62809 115546 62875 115549
rect 60742 115544 62875 115546
rect 60742 115488 62814 115544
rect 62870 115488 62875 115544
rect 60742 115486 62875 115488
rect 60742 115312 60802 115486
rect 62809 115483 62875 115486
rect 65017 115138 65083 115141
rect 67918 115138 67978 116196
rect 132686 116168 135126 116224
rect 135182 116168 135187 116224
rect 174313 116226 174379 116229
rect 174313 116224 177090 116226
rect 132686 116166 135187 116168
rect 97726 115546 97786 116128
rect 132686 115856 132746 116166
rect 135121 116163 135187 116166
rect 102645 115818 102711 115821
rect 102645 115816 104932 115818
rect 102645 115760 102650 115816
rect 102706 115760 104932 115816
rect 102645 115758 104932 115760
rect 102645 115755 102711 115758
rect 100897 115546 100963 115549
rect 134845 115546 134911 115549
rect 97726 115544 100963 115546
rect 97726 115488 100902 115544
rect 100958 115488 100963 115544
rect 97726 115486 100963 115488
rect 100897 115483 100963 115486
rect 132686 115544 134911 115546
rect 132686 115488 134850 115544
rect 134906 115488 134911 115544
rect 132686 115486 134911 115488
rect 132686 115312 132746 115486
rect 134845 115483 134911 115486
rect 136777 115546 136843 115549
rect 140046 115546 140106 116128
rect 169854 115682 169914 116196
rect 174313 116168 174318 116224
rect 174374 116168 177090 116224
rect 174313 116166 177090 116168
rect 174313 116163 174379 116166
rect 177030 115856 177090 116166
rect 222705 115954 222771 115957
rect 227416 115954 227896 115984
rect 222705 115952 227896 115954
rect 222705 115896 222710 115952
rect 222766 115896 227896 115952
rect 222705 115894 227896 115896
rect 222705 115891 222771 115894
rect 227416 115864 227896 115894
rect 171829 115682 171895 115685
rect 169854 115680 171895 115682
rect 169854 115624 171834 115680
rect 171890 115624 171895 115680
rect 169854 115622 171895 115624
rect 171829 115619 171895 115622
rect 136777 115544 140106 115546
rect 136777 115488 136782 115544
rect 136838 115488 140106 115544
rect 136777 115486 140106 115488
rect 174129 115546 174195 115549
rect 174129 115544 177090 115546
rect 174129 115488 174134 115544
rect 174190 115488 177090 115544
rect 174129 115486 177090 115488
rect 136777 115483 136843 115486
rect 174129 115483 174195 115486
rect 177030 115312 177090 115486
rect 102369 115274 102435 115277
rect 102369 115272 104932 115274
rect 102369 115216 102374 115272
rect 102430 115216 104932 115272
rect 102369 115214 104932 115216
rect 102369 115211 102435 115214
rect 65017 115136 67978 115138
rect 65017 115080 65022 115136
rect 65078 115080 67978 115136
rect 65017 115078 67978 115080
rect 65017 115075 65083 115078
rect 135305 115002 135371 115005
rect 132686 115000 135371 115002
rect 132686 114944 135310 115000
rect 135366 114944 135371 115000
rect 132686 114942 135371 114944
rect 132686 114768 132746 114942
rect 135305 114939 135371 114942
rect 174221 115002 174287 115005
rect 174221 115000 177090 115002
rect 174221 114944 174226 115000
rect 174282 114944 177090 115000
rect 174221 114942 177090 114944
rect 174221 114939 174287 114942
rect 177030 114768 177090 114942
rect 62809 114730 62875 114733
rect 60772 114728 62875 114730
rect 60772 114672 62814 114728
rect 62870 114672 62875 114728
rect 60772 114670 62875 114672
rect 62809 114667 62875 114670
rect 102185 114730 102251 114733
rect 102185 114728 104932 114730
rect 102185 114672 102190 114728
rect 102246 114672 104932 114728
rect 102185 114670 104932 114672
rect 102185 114667 102251 114670
rect 62809 114458 62875 114461
rect 134845 114458 134911 114461
rect 60742 114456 62875 114458
rect 60742 114400 62814 114456
rect 62870 114400 62875 114456
rect 60742 114398 62875 114400
rect 60742 114224 60802 114398
rect 62809 114395 62875 114398
rect 132686 114456 134911 114458
rect 132686 114400 134850 114456
rect 134906 114400 134911 114456
rect 132686 114398 134911 114400
rect 132686 114224 132746 114398
rect 134845 114395 134911 114398
rect 174037 114458 174103 114461
rect 174037 114456 177090 114458
rect 174037 114400 174042 114456
rect 174098 114400 177090 114456
rect 174037 114398 177090 114400
rect 174037 114395 174103 114398
rect 177030 114224 177090 114398
rect 102277 114186 102343 114189
rect 102277 114184 104932 114186
rect 102277 114128 102282 114184
rect 102338 114128 104932 114184
rect 102277 114126 104932 114128
rect 102277 114123 102343 114126
rect 101817 113780 101883 113781
rect 101766 113778 101772 113780
rect 101726 113718 101772 113778
rect 101836 113776 101883 113780
rect 101878 113720 101883 113776
rect 101766 113716 101772 113718
rect 101836 113716 101883 113720
rect 101817 113715 101883 113716
rect 56921 113236 56987 113237
rect 72009 113236 72075 113237
rect 56870 113172 56876 113236
rect 56940 113234 56987 113236
rect 56940 113232 57032 113234
rect 56982 113176 57032 113232
rect 56940 113174 57032 113176
rect 56940 113172 56987 113174
rect 71958 113172 71964 113236
rect 72028 113234 72075 113236
rect 72028 113232 72120 113234
rect 72070 113176 72120 113232
rect 72028 113174 72120 113176
rect 72028 113172 72075 113174
rect 56921 113171 56987 113172
rect 72009 113171 72075 113172
rect 105773 110242 105839 110245
rect 177717 110242 177783 110245
rect 102724 110240 105839 110242
rect 102724 110184 105778 110240
rect 105834 110184 105839 110240
rect 102724 110182 105839 110184
rect 174852 110240 177783 110242
rect 174852 110184 177722 110240
rect 177778 110184 177783 110240
rect 174852 110182 177783 110184
rect 105773 110179 105839 110182
rect 177717 110179 177783 110182
rect 108533 109562 108599 109565
rect 180293 109562 180359 109565
rect 108533 109560 111004 109562
rect 108533 109504 108538 109560
rect 108594 109504 111004 109560
rect 108533 109502 111004 109504
rect 180293 109560 182948 109562
rect 180293 109504 180298 109560
rect 180354 109504 182948 109560
rect 180293 109502 182948 109504
rect 108533 109499 108599 109502
rect 180293 109499 180359 109502
rect 105313 109154 105379 109157
rect 177165 109154 177231 109157
rect 102724 109152 105379 109154
rect 102724 109096 105318 109152
rect 105374 109096 105379 109152
rect 102724 109094 105379 109096
rect 174852 109152 177231 109154
rect 174852 109096 177170 109152
rect 177226 109096 177231 109152
rect 174852 109094 177231 109096
rect 105313 109091 105379 109094
rect 177165 109091 177231 109094
rect 105681 107930 105747 107933
rect 177257 107930 177323 107933
rect 102724 107928 105747 107930
rect 102724 107872 105686 107928
rect 105742 107872 105747 107928
rect 102724 107870 105747 107872
rect 174852 107928 177323 107930
rect 174852 107872 177262 107928
rect 177318 107872 177323 107928
rect 174852 107870 177323 107872
rect 105681 107867 105747 107870
rect 177257 107867 177323 107870
rect 107889 107250 107955 107253
rect 179649 107250 179715 107253
rect 107889 107248 111004 107250
rect 107889 107192 107894 107248
rect 107950 107192 111004 107248
rect 107889 107190 111004 107192
rect 179649 107248 182948 107250
rect 179649 107192 179654 107248
rect 179710 107192 182948 107248
rect 179649 107190 182948 107192
rect 107889 107187 107955 107190
rect 179649 107187 179715 107190
rect 105405 106842 105471 106845
rect 176981 106842 177047 106845
rect 102724 106840 105471 106842
rect 102724 106784 105410 106840
rect 105466 106784 105471 106840
rect 102724 106782 105471 106784
rect 174852 106840 177047 106842
rect 174852 106784 176986 106840
rect 177042 106784 177047 106840
rect 174852 106782 177047 106784
rect 105405 106779 105471 106782
rect 176981 106779 177047 106782
rect 9896 106162 10376 106192
rect 12209 106162 12275 106165
rect 9896 106160 12275 106162
rect 9896 106104 12214 106160
rect 12270 106104 12275 106160
rect 9896 106102 12275 106104
rect 9896 106072 10376 106102
rect 12209 106099 12275 106102
rect 12025 105754 12091 105757
rect 105221 105754 105287 105757
rect 177073 105754 177139 105757
rect 224453 105754 224519 105757
rect 12025 105752 14036 105754
rect 12025 105696 12030 105752
rect 12086 105696 14036 105752
rect 12025 105694 14036 105696
rect 102724 105752 105287 105754
rect 102724 105696 105226 105752
rect 105282 105696 105287 105752
rect 102724 105694 105287 105696
rect 174852 105752 177139 105754
rect 174852 105696 177078 105752
rect 177134 105696 177139 105752
rect 174852 105694 177139 105696
rect 223796 105752 224519 105754
rect 223796 105696 224458 105752
rect 224514 105696 224519 105752
rect 223796 105694 224519 105696
rect 12025 105691 12091 105694
rect 105221 105691 105287 105694
rect 177073 105691 177139 105694
rect 224453 105691 224519 105694
rect 132269 105482 132335 105485
rect 132545 105482 132611 105485
rect 132269 105480 132611 105482
rect 132269 105424 132274 105480
rect 132330 105424 132550 105480
rect 132606 105424 132611 105480
rect 132269 105422 132611 105424
rect 132269 105419 132335 105422
rect 132545 105419 132611 105422
rect 108441 104938 108507 104941
rect 179649 104938 179715 104941
rect 108441 104936 111004 104938
rect 108441 104880 108446 104936
rect 108502 104880 111004 104936
rect 108441 104878 111004 104880
rect 179649 104936 182948 104938
rect 179649 104880 179654 104936
rect 179710 104880 182948 104936
rect 179649 104878 182948 104880
rect 108441 104875 108507 104878
rect 179649 104875 179715 104878
rect 106049 104530 106115 104533
rect 177441 104530 177507 104533
rect 102724 104528 106115 104530
rect 102724 104472 106054 104528
rect 106110 104472 106115 104528
rect 102724 104470 106115 104472
rect 174852 104528 177507 104530
rect 174852 104472 177446 104528
rect 177502 104472 177507 104528
rect 174852 104470 177507 104472
rect 106049 104467 106115 104470
rect 177441 104467 177507 104470
rect 31989 104258 32055 104261
rect 29860 104256 32055 104258
rect 29860 104200 31994 104256
rect 32050 104200 32055 104256
rect 29860 104198 32055 104200
rect 31989 104195 32055 104198
rect 37417 104258 37483 104261
rect 59865 104258 59931 104261
rect 201085 104258 201151 104261
rect 37417 104256 39060 104258
rect 37417 104200 37422 104256
rect 37478 104200 39060 104256
rect 37417 104198 39060 104200
rect 59865 104256 62980 104258
rect 59865 104200 59870 104256
rect 59926 104200 62980 104256
rect 59865 104198 62980 104200
rect 126828 104198 134924 104258
rect 198772 104256 201151 104258
rect 198772 104200 201090 104256
rect 201146 104200 201151 104256
rect 198772 104198 201151 104200
rect 37417 104195 37483 104198
rect 59865 104195 59931 104198
rect 201085 104195 201151 104198
rect 204581 104258 204647 104261
rect 204581 104256 207972 104258
rect 204581 104200 204586 104256
rect 204642 104200 207972 104256
rect 204581 104198 207972 104200
rect 204581 104195 204647 104198
rect 105589 103442 105655 103445
rect 177349 103442 177415 103445
rect 102724 103440 105655 103442
rect 102724 103384 105594 103440
rect 105650 103384 105655 103440
rect 102724 103382 105655 103384
rect 174852 103440 177415 103442
rect 174852 103384 177354 103440
rect 177410 103384 177415 103440
rect 174852 103382 177415 103384
rect 105589 103379 105655 103382
rect 177349 103379 177415 103382
rect 107889 102490 107955 102493
rect 179649 102490 179715 102493
rect 107889 102488 111004 102490
rect 107889 102432 107894 102488
rect 107950 102432 111004 102488
rect 107889 102430 111004 102432
rect 179649 102488 182948 102490
rect 179649 102432 179654 102488
rect 179710 102432 182948 102488
rect 179649 102430 182948 102432
rect 107889 102427 107955 102430
rect 179649 102427 179715 102430
rect 105129 102218 105195 102221
rect 176889 102218 176955 102221
rect 102724 102216 105195 102218
rect 102724 102160 105134 102216
rect 105190 102160 105195 102216
rect 102724 102158 105195 102160
rect 174852 102216 176955 102218
rect 174852 102160 176894 102216
rect 176950 102160 176955 102216
rect 174852 102158 176955 102160
rect 105129 102155 105195 102158
rect 176889 102155 176955 102158
rect 105957 101130 106023 101133
rect 176981 101130 177047 101133
rect 102724 101128 106023 101130
rect 102724 101072 105962 101128
rect 106018 101072 106023 101128
rect 102724 101070 106023 101072
rect 174852 101128 177047 101130
rect 174852 101072 176986 101128
rect 177042 101072 177047 101128
rect 174852 101070 177047 101072
rect 105957 101067 106023 101070
rect 176981 101067 177047 101070
rect 56829 100858 56895 100861
rect 54884 100856 56895 100858
rect 54884 100800 56834 100856
rect 56890 100800 56895 100856
rect 54884 100798 56895 100800
rect 56829 100795 56895 100798
rect 107889 100178 107955 100181
rect 179649 100178 179715 100181
rect 107889 100176 111004 100178
rect 107889 100120 107894 100176
rect 107950 100120 111004 100176
rect 107889 100118 111004 100120
rect 179649 100176 182948 100178
rect 179649 100120 179654 100176
rect 179710 100120 182948 100176
rect 179649 100118 182948 100120
rect 107889 100115 107955 100118
rect 179649 100115 179715 100118
rect 106417 100042 106483 100045
rect 177533 100042 177599 100045
rect 102724 100040 106483 100042
rect 102724 99984 106422 100040
rect 106478 99984 106483 100040
rect 102724 99982 106483 99984
rect 174852 100040 177599 100042
rect 174852 99984 177538 100040
rect 177594 99984 177599 100040
rect 174852 99982 177599 99984
rect 106417 99979 106483 99982
rect 177533 99979 177599 99982
rect 105773 98818 105839 98821
rect 177809 98818 177875 98821
rect 102724 98816 105839 98818
rect 102724 98760 105778 98816
rect 105834 98760 105839 98816
rect 102724 98758 105839 98760
rect 174852 98816 177875 98818
rect 174852 98760 177814 98816
rect 177870 98760 177875 98816
rect 174852 98758 177875 98760
rect 105773 98755 105839 98758
rect 177809 98755 177875 98758
rect 107889 97866 107955 97869
rect 179649 97866 179715 97869
rect 107889 97864 111004 97866
rect 107889 97808 107894 97864
rect 107950 97808 111004 97864
rect 107889 97806 111004 97808
rect 179649 97864 182948 97866
rect 179649 97808 179654 97864
rect 179710 97808 182948 97864
rect 179649 97806 182948 97808
rect 107889 97803 107955 97806
rect 179649 97803 179715 97806
rect 106325 97730 106391 97733
rect 177625 97730 177691 97733
rect 102724 97728 106391 97730
rect 102724 97672 106330 97728
rect 106386 97672 106391 97728
rect 102724 97670 106391 97672
rect 174852 97728 177691 97730
rect 174852 97672 177630 97728
rect 177686 97672 177691 97728
rect 174852 97670 177691 97672
rect 106325 97667 106391 97670
rect 177625 97667 177691 97670
rect 106417 96506 106483 96509
rect 177717 96506 177783 96509
rect 102724 96504 106483 96506
rect 102724 96448 106422 96504
rect 106478 96448 106483 96504
rect 102724 96446 106483 96448
rect 174852 96504 177783 96506
rect 174852 96448 177722 96504
rect 177778 96448 177783 96504
rect 174852 96446 177783 96448
rect 106417 96443 106483 96446
rect 177717 96443 177783 96446
rect 223533 96370 223599 96373
rect 223533 96368 223642 96370
rect 223533 96312 223538 96368
rect 223594 96312 223642 96368
rect 223533 96307 223642 96312
rect 12117 95826 12183 95829
rect 12117 95824 14036 95826
rect 12117 95768 12122 95824
rect 12178 95768 14036 95824
rect 223582 95796 223642 96307
rect 12117 95766 14036 95768
rect 12117 95763 12183 95766
rect 106233 95418 106299 95421
rect 102724 95416 106299 95418
rect 102724 95360 106238 95416
rect 106294 95360 106299 95416
rect 102724 95358 106299 95360
rect 106233 95355 106299 95358
rect 108441 95418 108507 95421
rect 177533 95418 177599 95421
rect 108441 95416 111004 95418
rect 108441 95360 108446 95416
rect 108502 95360 111004 95416
rect 108441 95358 111004 95360
rect 174852 95416 177599 95418
rect 174852 95360 177538 95416
rect 177594 95360 177599 95416
rect 174852 95358 177599 95360
rect 108441 95355 108507 95358
rect 177533 95355 177599 95358
rect 179557 95418 179623 95421
rect 179557 95416 182948 95418
rect 179557 95360 179562 95416
rect 179618 95360 182948 95416
rect 179557 95358 182948 95360
rect 179557 95355 179623 95358
rect 106509 94330 106575 94333
rect 177441 94330 177507 94333
rect 102724 94328 106575 94330
rect 102724 94272 106514 94328
rect 106570 94272 106575 94328
rect 102724 94270 106575 94272
rect 174852 94328 177507 94330
rect 174852 94272 177446 94328
rect 177502 94272 177507 94328
rect 174852 94270 177507 94272
rect 106509 94267 106575 94270
rect 177441 94267 177507 94270
rect 102724 93046 111004 93106
rect 174852 93046 182948 93106
rect 223533 92154 223599 92157
rect 227416 92154 227896 92184
rect 223533 92152 227896 92154
rect 223533 92096 223538 92152
rect 223594 92096 227896 92152
rect 223533 92094 227896 92096
rect 223533 92091 223599 92094
rect 227416 92064 227896 92094
rect 177533 92018 177599 92021
rect 174852 92016 177599 92018
rect 174852 91960 177538 92016
rect 177594 91960 177599 92016
rect 174852 91958 177599 91960
rect 177533 91955 177599 91958
rect 102694 91746 102754 91920
rect 105865 91746 105931 91749
rect 102694 91744 105931 91746
rect 102694 91688 105870 91744
rect 105926 91688 105931 91744
rect 102694 91686 105931 91688
rect 105865 91683 105931 91686
rect 32633 90930 32699 90933
rect 29860 90928 32699 90930
rect 29860 90872 32638 90928
rect 32694 90872 32699 90928
rect 29860 90870 32699 90872
rect 32633 90867 32699 90870
rect 36405 90930 36471 90933
rect 59589 90930 59655 90933
rect 204489 90930 204555 90933
rect 36405 90928 39060 90930
rect 36405 90872 36410 90928
rect 36466 90872 39060 90928
rect 36405 90870 39060 90872
rect 59589 90928 62980 90930
rect 59589 90872 59594 90928
rect 59650 90872 62980 90928
rect 59589 90870 62980 90872
rect 126828 90870 134924 90930
rect 204489 90928 207972 90930
rect 204489 90872 204494 90928
rect 204550 90872 207972 90928
rect 204489 90870 207972 90872
rect 36405 90867 36471 90870
rect 59589 90867 59655 90870
rect 204489 90867 204555 90870
rect 107797 90794 107863 90797
rect 177349 90794 177415 90797
rect 107797 90792 111004 90794
rect 107797 90736 107802 90792
rect 107858 90736 111004 90792
rect 107797 90734 111004 90736
rect 174852 90792 177415 90794
rect 174852 90736 177354 90792
rect 177410 90736 177415 90792
rect 174852 90734 177415 90736
rect 107797 90731 107863 90734
rect 177349 90731 177415 90734
rect 179557 90794 179623 90797
rect 179557 90792 182948 90794
rect 179557 90736 179562 90792
rect 179618 90736 182948 90792
rect 179557 90734 182948 90736
rect 179557 90731 179623 90734
rect 102694 90386 102754 90696
rect 105221 90386 105287 90389
rect 102694 90384 105287 90386
rect 102694 90328 105226 90384
rect 105282 90328 105287 90384
rect 102694 90326 105287 90328
rect 198742 90386 198802 90832
rect 200993 90386 201059 90389
rect 198742 90384 201059 90386
rect 198742 90328 200998 90384
rect 201054 90328 201059 90384
rect 198742 90326 201059 90328
rect 105221 90323 105287 90326
rect 200993 90323 201059 90326
rect 177349 89706 177415 89709
rect 174852 89704 177415 89706
rect 174852 89648 177354 89704
rect 177410 89648 177415 89704
rect 174852 89646 177415 89648
rect 177349 89643 177415 89646
rect 102694 89298 102754 89608
rect 105129 89298 105195 89301
rect 102694 89296 105195 89298
rect 102694 89240 105134 89296
rect 105190 89240 105195 89296
rect 102694 89238 105195 89240
rect 105129 89235 105195 89238
rect 177349 88618 177415 88621
rect 174852 88616 177415 88618
rect 174852 88560 177354 88616
rect 177410 88560 177415 88616
rect 174852 88558 177415 88560
rect 177349 88555 177415 88558
rect 102694 87938 102754 88520
rect 107889 88482 107955 88485
rect 179649 88482 179715 88485
rect 107889 88480 111004 88482
rect 107889 88424 107894 88480
rect 107950 88424 111004 88480
rect 107889 88422 111004 88424
rect 179649 88480 182948 88482
rect 179649 88424 179654 88480
rect 179710 88424 182948 88480
rect 179649 88422 182948 88424
rect 107889 88419 107955 88422
rect 179649 88419 179715 88422
rect 105865 87938 105931 87941
rect 102694 87936 105931 87938
rect 102694 87880 105870 87936
rect 105926 87880 105931 87936
rect 102694 87878 105931 87880
rect 105865 87875 105931 87878
rect 178913 87394 178979 87397
rect 174852 87392 178979 87394
rect 174852 87336 178918 87392
rect 178974 87336 178979 87392
rect 174852 87334 178979 87336
rect 178913 87331 178979 87334
rect 102694 86714 102754 87296
rect 106417 86714 106483 86717
rect 102694 86712 106483 86714
rect 102694 86656 106422 86712
rect 106478 86656 106483 86712
rect 102694 86654 106483 86656
rect 106417 86651 106483 86654
rect 105589 86306 105655 86309
rect 178085 86306 178151 86309
rect 102724 86304 105655 86306
rect 102724 86248 105594 86304
rect 105650 86248 105655 86304
rect 102724 86246 105655 86248
rect 174852 86304 178151 86306
rect 174852 86248 178090 86304
rect 178146 86248 178151 86304
rect 174852 86246 178151 86248
rect 105589 86243 105655 86246
rect 178085 86243 178151 86246
rect 107797 86034 107863 86037
rect 179557 86034 179623 86037
rect 107797 86032 111004 86034
rect 107797 85976 107802 86032
rect 107858 85976 111004 86032
rect 107797 85974 111004 85976
rect 179557 86032 182948 86034
rect 179557 85976 179562 86032
rect 179618 85976 182948 86032
rect 179557 85974 182948 85976
rect 107797 85971 107863 85974
rect 179557 85971 179623 85974
rect 14006 84810 14066 85664
rect 223582 85221 223642 85732
rect 223533 85216 223642 85221
rect 223533 85160 223538 85216
rect 223594 85160 223642 85216
rect 223533 85158 223642 85160
rect 223533 85155 223599 85158
rect 177533 85082 177599 85085
rect 174852 85080 177599 85082
rect 174852 85024 177538 85080
rect 177594 85024 177599 85080
rect 174852 85022 177599 85024
rect 177533 85019 177599 85022
rect 11982 84750 14066 84810
rect 102694 84810 102754 84984
rect 106325 84810 106391 84813
rect 102694 84808 106391 84810
rect 102694 84752 106330 84808
rect 106386 84752 106391 84808
rect 102694 84750 106391 84752
rect 9896 84538 10376 84568
rect 11982 84538 12042 84750
rect 106325 84747 106391 84750
rect 9896 84478 12042 84538
rect 9896 84448 10376 84478
rect 178177 83994 178243 83997
rect 174852 83992 178243 83994
rect 174852 83936 178182 83992
rect 178238 83936 178243 83992
rect 174852 83934 178243 83936
rect 178177 83931 178243 83934
rect 102694 83450 102754 83896
rect 107705 83722 107771 83725
rect 179465 83722 179531 83725
rect 107705 83720 111004 83722
rect 107705 83664 107710 83720
rect 107766 83664 111004 83720
rect 107705 83662 111004 83664
rect 179465 83720 182948 83722
rect 179465 83664 179470 83720
rect 179526 83664 182948 83720
rect 179465 83662 182948 83664
rect 107705 83659 107771 83662
rect 179465 83659 179531 83662
rect 105589 83450 105655 83453
rect 102694 83448 105655 83450
rect 102694 83392 105594 83448
rect 105650 83392 105655 83448
rect 102694 83390 105655 83392
rect 105589 83387 105655 83390
rect 177717 82906 177783 82909
rect 174852 82904 177783 82906
rect 174852 82848 177722 82904
rect 177778 82848 177783 82904
rect 174852 82846 177783 82848
rect 177717 82843 177783 82846
rect 102694 82226 102754 82808
rect 105497 82226 105563 82229
rect 102694 82224 105563 82226
rect 102694 82168 105502 82224
rect 105558 82168 105563 82224
rect 102694 82166 105563 82168
rect 105497 82163 105563 82166
rect 56921 81954 56987 81957
rect 57473 81954 57539 81957
rect 56921 81952 57539 81954
rect 56921 81896 56926 81952
rect 56982 81896 57478 81952
rect 57534 81896 57539 81952
rect 56921 81894 57539 81896
rect 56921 81891 56987 81894
rect 57473 81891 57539 81894
rect 177349 81682 177415 81685
rect 174852 81680 177415 81682
rect 174852 81624 177354 81680
rect 177410 81624 177415 81680
rect 174852 81622 177415 81624
rect 177349 81619 177415 81622
rect 102694 81002 102754 81584
rect 107889 81410 107955 81413
rect 178913 81410 178979 81413
rect 107889 81408 111004 81410
rect 107889 81352 107894 81408
rect 107950 81352 111004 81408
rect 107889 81350 111004 81352
rect 178913 81408 182948 81410
rect 178913 81352 178918 81408
rect 178974 81352 182948 81408
rect 178913 81350 182948 81352
rect 107889 81347 107955 81350
rect 178913 81347 178979 81350
rect 105221 81002 105287 81005
rect 102694 81000 105287 81002
rect 102694 80944 105226 81000
rect 105282 80944 105287 81000
rect 102694 80942 105287 80944
rect 105221 80939 105287 80942
rect 57473 80866 57539 80869
rect 54884 80864 57539 80866
rect 54884 80808 57478 80864
rect 57534 80808 57539 80864
rect 54884 80806 57539 80808
rect 57473 80803 57539 80806
rect 178177 80594 178243 80597
rect 174852 80592 178243 80594
rect 174852 80536 178182 80592
rect 178238 80536 178243 80592
rect 174852 80534 178243 80536
rect 178177 80531 178243 80534
rect 102694 79914 102754 80496
rect 105129 79914 105195 79917
rect 102694 79912 105195 79914
rect 102694 79856 105134 79912
rect 105190 79856 105195 79912
rect 102694 79854 105195 79856
rect 105129 79851 105195 79854
rect 106969 79370 107035 79373
rect 178821 79370 178887 79373
rect 102724 79368 107035 79370
rect 102724 79312 106974 79368
rect 107030 79312 107035 79368
rect 102724 79310 107035 79312
rect 174852 79368 178887 79370
rect 174852 79312 178826 79368
rect 178882 79312 178887 79368
rect 174852 79310 178887 79312
rect 106969 79307 107035 79310
rect 178821 79307 178887 79310
rect 108717 78962 108783 78965
rect 180477 78962 180543 78965
rect 108717 78960 111004 78962
rect 108717 78904 108722 78960
rect 108778 78904 111004 78960
rect 108717 78902 111004 78904
rect 180477 78960 182948 78962
rect 180477 78904 180482 78960
rect 180538 78904 182948 78960
rect 180477 78902 182948 78904
rect 108717 78899 108783 78902
rect 180477 78899 180543 78902
rect 178269 78282 178335 78285
rect 174852 78280 178335 78282
rect 174852 78224 178274 78280
rect 178330 78224 178335 78280
rect 174852 78222 178335 78224
rect 178269 78219 178335 78222
rect 102694 77874 102754 78184
rect 106325 77874 106391 77877
rect 102694 77872 106391 77874
rect 102694 77816 106330 77872
rect 106386 77816 106391 77872
rect 102694 77814 106391 77816
rect 106325 77811 106391 77814
rect 31989 77602 32055 77605
rect 29860 77600 32055 77602
rect 29860 77544 31994 77600
rect 32050 77544 32055 77600
rect 29860 77542 32055 77544
rect 31989 77539 32055 77542
rect 37417 77602 37483 77605
rect 59589 77602 59655 77605
rect 129734 77602 129740 77604
rect 37417 77600 39060 77602
rect 37417 77544 37422 77600
rect 37478 77544 39060 77600
rect 37417 77542 39060 77544
rect 59589 77600 62980 77602
rect 59589 77544 59594 77600
rect 59650 77544 62980 77600
rect 59589 77542 62980 77544
rect 126828 77542 129740 77602
rect 37417 77539 37483 77542
rect 59589 77539 59655 77542
rect 129734 77540 129740 77542
rect 129804 77602 129810 77604
rect 204489 77602 204555 77605
rect 129804 77542 134924 77602
rect 204489 77600 207972 77602
rect 204489 77544 204494 77600
rect 204550 77544 207972 77600
rect 204489 77542 207972 77544
rect 129804 77540 129810 77542
rect 204489 77539 204555 77542
rect 177717 77194 177783 77197
rect 174852 77192 177783 77194
rect 174852 77136 177722 77192
rect 177778 77136 177783 77192
rect 174852 77134 177783 77136
rect 177717 77131 177783 77134
rect 102694 76514 102754 77096
rect 198742 77058 198802 77504
rect 201085 77058 201151 77061
rect 198742 77056 201151 77058
rect 198742 77000 201090 77056
rect 201146 77000 201151 77056
rect 198742 76998 201151 77000
rect 201085 76995 201151 76998
rect 108809 76650 108875 76653
rect 179649 76650 179715 76653
rect 108809 76648 111004 76650
rect 108809 76592 108814 76648
rect 108870 76592 111004 76648
rect 108809 76590 111004 76592
rect 179649 76648 182948 76650
rect 179649 76592 179654 76648
rect 179710 76592 182948 76648
rect 179649 76590 182948 76592
rect 108809 76587 108875 76590
rect 179649 76587 179715 76590
rect 105405 76514 105471 76517
rect 102694 76512 105471 76514
rect 102694 76456 105410 76512
rect 105466 76456 105471 76512
rect 102694 76454 105471 76456
rect 105405 76451 105471 76454
rect 177165 75970 177231 75973
rect 174852 75968 177231 75970
rect 174852 75912 177170 75968
rect 177226 75912 177231 75968
rect 174852 75910 177231 75912
rect 177165 75907 177231 75910
rect 12025 75154 12091 75157
rect 14006 75154 14066 75736
rect 102694 75290 102754 75872
rect 223582 75293 223642 75804
rect 105221 75290 105287 75293
rect 102694 75288 105287 75290
rect 102694 75232 105226 75288
rect 105282 75232 105287 75288
rect 102694 75230 105287 75232
rect 105221 75227 105287 75230
rect 223533 75288 223642 75293
rect 223533 75232 223538 75288
rect 223594 75232 223642 75288
rect 223533 75230 223642 75232
rect 223533 75227 223599 75230
rect 12025 75152 14066 75154
rect 12025 75096 12030 75152
rect 12086 75096 14066 75152
rect 12025 75094 14066 75096
rect 12025 75091 12091 75094
rect 178361 74882 178427 74885
rect 174852 74880 178427 74882
rect 174852 74824 178366 74880
rect 178422 74824 178427 74880
rect 174852 74822 178427 74824
rect 178361 74819 178427 74822
rect 102694 74202 102754 74784
rect 108625 74338 108691 74341
rect 180385 74338 180451 74341
rect 108625 74336 111004 74338
rect 108625 74280 108630 74336
rect 108686 74280 111004 74336
rect 108625 74278 111004 74280
rect 180385 74336 182948 74338
rect 180385 74280 180390 74336
rect 180446 74280 182948 74336
rect 180385 74278 182948 74280
rect 108625 74275 108691 74278
rect 180385 74275 180451 74278
rect 106417 74202 106483 74205
rect 102694 74200 106483 74202
rect 102694 74144 106422 74200
rect 106478 74144 106483 74200
rect 102694 74142 106483 74144
rect 106417 74139 106483 74142
rect 177349 73658 177415 73661
rect 174852 73656 177415 73658
rect 174852 73600 177354 73656
rect 177410 73600 177415 73656
rect 174852 73598 177415 73600
rect 177349 73595 177415 73598
rect 103197 73590 103263 73593
rect 102724 73588 103263 73590
rect 102724 73532 103202 73588
rect 103258 73532 103263 73588
rect 102724 73530 103263 73532
rect 103197 73527 103263 73530
rect 102553 73388 102619 73389
rect 102502 73324 102508 73388
rect 102572 73386 102619 73388
rect 102572 73384 102664 73386
rect 102614 73328 102664 73384
rect 102572 73326 102664 73328
rect 102572 73324 102619 73326
rect 102553 73323 102619 73324
rect 174497 72978 174563 72981
rect 174497 72976 174698 72978
rect 174497 72920 174502 72976
rect 174558 72920 174698 72976
rect 174497 72918 174698 72920
rect 174497 72915 174563 72918
rect 174638 72540 174698 72918
rect 102553 72026 102619 72029
rect 102510 72024 102619 72026
rect 102510 71968 102558 72024
rect 102614 71968 102619 72024
rect 102510 71963 102619 71968
rect 102510 71452 102570 71963
rect 102694 71893 102754 72472
rect 108533 72026 108599 72029
rect 180293 72026 180359 72029
rect 108533 72024 111004 72026
rect 108533 71968 108538 72024
rect 108594 71968 111004 72024
rect 108533 71966 111004 71968
rect 180293 72024 182948 72026
rect 180293 71968 180298 72024
rect 180354 71968 182948 72024
rect 180293 71966 182948 71968
rect 108533 71963 108599 71966
rect 180293 71963 180359 71966
rect 102645 71888 102754 71893
rect 102645 71832 102650 71888
rect 102706 71832 102754 71888
rect 102645 71830 102754 71832
rect 102645 71827 102711 71830
rect 101357 71212 101423 71213
rect 101357 71210 101404 71212
rect 101312 71208 101404 71210
rect 101312 71152 101362 71208
rect 101312 71150 101404 71152
rect 101357 71148 101404 71150
rect 101468 71148 101474 71212
rect 173342 71148 173348 71212
rect 173412 71210 173418 71212
rect 174454 71210 174514 71452
rect 173412 71150 174514 71210
rect 173412 71148 173418 71150
rect 101357 71147 101423 71148
rect 100846 71012 100852 71076
rect 100916 71074 100922 71076
rect 101909 71074 101975 71077
rect 100916 71072 101975 71074
rect 100916 71016 101914 71072
rect 101970 71016 101975 71072
rect 100916 71014 101975 71016
rect 100916 71012 100922 71014
rect 101909 71011 101975 71014
rect 101214 70876 101220 70940
rect 101284 70938 101290 70940
rect 102645 70938 102711 70941
rect 101284 70936 102711 70938
rect 101284 70880 102650 70936
rect 102706 70880 102711 70936
rect 101284 70878 102711 70880
rect 101284 70876 101290 70878
rect 102645 70875 102711 70878
rect 201085 69442 201151 69445
rect 201494 69442 201500 69444
rect 201085 69440 201500 69442
rect 201085 69384 201090 69440
rect 201146 69384 201500 69440
rect 201085 69382 201500 69384
rect 201085 69379 201151 69382
rect 201494 69380 201500 69382
rect 201564 69442 201570 69444
rect 202189 69442 202255 69445
rect 201564 69440 202255 69442
rect 201564 69384 202194 69440
rect 202250 69384 202255 69440
rect 201564 69382 202255 69384
rect 201564 69380 201570 69382
rect 202189 69379 202255 69382
rect 91237 69306 91303 69309
rect 176838 69306 176844 69308
rect 91237 69304 176844 69306
rect 91237 69248 91242 69304
rect 91298 69248 176844 69304
rect 91237 69246 176844 69248
rect 91237 69243 91303 69246
rect 176838 69244 176844 69246
rect 176908 69244 176914 69308
rect 191333 69306 191399 69309
rect 193081 69306 193147 69309
rect 191333 69304 193147 69306
rect 191333 69248 191338 69304
rect 191394 69248 193086 69304
rect 193142 69248 193147 69304
rect 191333 69246 193147 69248
rect 191333 69243 191399 69246
rect 193081 69243 193147 69246
rect 117825 69170 117891 69173
rect 119389 69170 119455 69173
rect 117825 69168 119455 69170
rect 117825 69112 117830 69168
rect 117886 69112 119394 69168
rect 119450 69112 119455 69168
rect 117825 69110 119455 69112
rect 117825 69107 117891 69110
rect 119389 69107 119455 69110
rect 189309 69170 189375 69173
rect 190229 69170 190295 69173
rect 189309 69168 190295 69170
rect 189309 69112 189314 69168
rect 189370 69112 190234 69168
rect 190290 69112 190295 69168
rect 189309 69110 190295 69112
rect 189309 69107 189375 69110
rect 190229 69107 190295 69110
rect 190413 69170 190479 69173
rect 191977 69170 192043 69173
rect 190413 69168 192043 69170
rect 190413 69112 190418 69168
rect 190474 69112 191982 69168
rect 192038 69112 192043 69168
rect 190413 69110 192043 69112
rect 190413 69107 190479 69110
rect 191977 69107 192043 69110
rect 48273 69034 48339 69037
rect 49469 69034 49535 69037
rect 48273 69032 49535 69034
rect 48273 68976 48278 69032
rect 48334 68976 49474 69032
rect 49530 68976 49535 69032
rect 48273 68974 49535 68976
rect 48273 68971 48339 68974
rect 49469 68971 49535 68974
rect 190137 69034 190203 69037
rect 191425 69034 191491 69037
rect 190137 69032 191491 69034
rect 190137 68976 190142 69032
rect 190198 68976 191430 69032
rect 191486 68976 191491 69032
rect 190137 68974 191491 68976
rect 190137 68971 190203 68974
rect 191425 68971 191491 68974
rect 49009 68898 49075 68901
rect 50849 68898 50915 68901
rect 49009 68896 50915 68898
rect 49009 68840 49014 68896
rect 49070 68840 50854 68896
rect 50910 68840 50915 68896
rect 49009 68838 50915 68840
rect 49009 68835 49075 68838
rect 50849 68835 50915 68838
rect 31897 68764 31963 68765
rect 31846 68762 31852 68764
rect 31806 68702 31852 68762
rect 31916 68760 31963 68764
rect 31958 68704 31963 68760
rect 31846 68700 31852 68702
rect 31916 68700 31963 68704
rect 31897 68699 31963 68700
rect 117089 68626 117155 68629
rect 118193 68626 118259 68629
rect 117089 68624 118259 68626
rect 117089 68568 117094 68624
rect 117150 68568 118198 68624
rect 118254 68568 118259 68624
rect 117089 68566 118259 68568
rect 117089 68563 117155 68566
rect 118193 68563 118259 68566
rect 119113 68490 119179 68493
rect 121137 68490 121203 68493
rect 119113 68488 121203 68490
rect 119113 68432 119118 68488
rect 119174 68432 121142 68488
rect 121198 68432 121203 68488
rect 119113 68430 121203 68432
rect 119113 68427 119179 68430
rect 121137 68427 121203 68430
rect 223073 68354 223139 68357
rect 227416 68354 227896 68384
rect 223073 68352 227896 68354
rect 223073 68296 223078 68352
rect 223134 68296 227896 68352
rect 223073 68294 227896 68296
rect 223073 68291 223139 68294
rect 227416 68264 227896 68294
rect 102461 67538 102527 67541
rect 135305 67538 135371 67541
rect 102461 67536 104932 67538
rect 102461 67480 102466 67536
rect 102522 67480 104932 67536
rect 102461 67478 104932 67480
rect 132716 67536 135371 67538
rect 132716 67480 135310 67536
rect 135366 67480 135371 67536
rect 132716 67478 135371 67480
rect 102461 67475 102527 67478
rect 135305 67475 135371 67478
rect 174681 67538 174747 67541
rect 174681 67536 177060 67538
rect 174681 67480 174686 67536
rect 174742 67480 177060 67536
rect 174681 67478 177060 67480
rect 174681 67475 174747 67478
rect 63361 67266 63427 67269
rect 60772 67264 63427 67266
rect 60772 67208 63366 67264
rect 63422 67208 63427 67264
rect 60772 67206 63427 67208
rect 63361 67203 63427 67206
rect 102369 66994 102435 66997
rect 135029 66994 135095 66997
rect 102369 66992 104932 66994
rect 102369 66936 102374 66992
rect 102430 66936 104932 66992
rect 102369 66934 104932 66936
rect 132716 66992 135095 66994
rect 132716 66936 135034 66992
rect 135090 66936 135095 66992
rect 132716 66934 135095 66936
rect 102369 66931 102435 66934
rect 135029 66931 135095 66934
rect 174037 66994 174103 66997
rect 174037 66992 177060 66994
rect 174037 66936 174042 66992
rect 174098 66936 177060 66992
rect 174037 66934 177060 66936
rect 174037 66931 174103 66934
rect 62809 66722 62875 66725
rect 60772 66720 62875 66722
rect 60772 66664 62814 66720
rect 62870 66664 62875 66720
rect 60772 66662 62875 66664
rect 62809 66659 62875 66662
rect 102553 66450 102619 66453
rect 135305 66450 135371 66453
rect 102553 66448 104932 66450
rect 102553 66392 102558 66448
rect 102614 66392 104932 66448
rect 102553 66390 104932 66392
rect 132716 66448 135371 66450
rect 132716 66392 135310 66448
rect 135366 66392 135371 66448
rect 132716 66390 135371 66392
rect 102553 66387 102619 66390
rect 135305 66387 135371 66390
rect 173945 66450 174011 66453
rect 173945 66448 177060 66450
rect 173945 66392 173950 66448
rect 174006 66392 177060 66448
rect 173945 66390 177060 66392
rect 173945 66387 174011 66390
rect 62717 66178 62783 66181
rect 60772 66176 62783 66178
rect 60772 66120 62722 66176
rect 62778 66120 62783 66176
rect 60772 66118 62783 66120
rect 62717 66115 62783 66118
rect 102369 65906 102435 65909
rect 134661 65906 134727 65909
rect 102369 65904 104932 65906
rect 102369 65848 102374 65904
rect 102430 65848 104932 65904
rect 102369 65846 104932 65848
rect 132716 65904 134727 65906
rect 132716 65848 134666 65904
rect 134722 65848 134727 65904
rect 132716 65846 134727 65848
rect 102369 65843 102435 65846
rect 134661 65843 134727 65846
rect 173853 65906 173919 65909
rect 173853 65904 177060 65906
rect 173853 65848 173858 65904
rect 173914 65848 177060 65904
rect 173853 65846 177060 65848
rect 173853 65843 173919 65846
rect 62901 65634 62967 65637
rect 171829 65634 171895 65637
rect 60772 65632 62967 65634
rect 60772 65576 62906 65632
rect 62962 65576 62967 65632
rect 60772 65574 62967 65576
rect 62901 65571 62967 65574
rect 169670 65632 171895 65634
rect 169670 65576 171834 65632
rect 171890 65576 171895 65632
rect 169670 65574 171895 65576
rect 66397 65498 66463 65501
rect 100897 65498 100963 65501
rect 66397 65496 67948 65498
rect 66397 65440 66402 65496
rect 66458 65440 67948 65496
rect 66397 65438 67948 65440
rect 97756 65496 100963 65498
rect 97756 65440 100902 65496
rect 100958 65440 100963 65496
rect 97756 65438 100963 65440
rect 66397 65435 66463 65438
rect 100897 65435 100963 65438
rect 136869 65498 136935 65501
rect 136869 65496 140076 65498
rect 136869 65440 136874 65496
rect 136930 65440 140076 65496
rect 169670 65468 169730 65574
rect 171829 65571 171895 65574
rect 136869 65438 140076 65440
rect 136869 65435 136935 65438
rect 102645 65226 102711 65229
rect 135305 65226 135371 65229
rect 102645 65224 104932 65226
rect 102645 65168 102650 65224
rect 102706 65168 104932 65224
rect 102645 65166 104932 65168
rect 132716 65224 135371 65226
rect 132716 65168 135310 65224
rect 135366 65168 135371 65224
rect 132716 65166 135371 65168
rect 102645 65163 102711 65166
rect 135305 65163 135371 65166
rect 169529 65226 169595 65229
rect 169529 65224 170466 65226
rect 169529 65168 169534 65224
rect 169590 65168 170466 65224
rect 169529 65166 170466 65168
rect 169529 65163 169595 65166
rect 62809 64954 62875 64957
rect 60772 64952 62875 64954
rect 60772 64896 62814 64952
rect 62870 64896 62875 64952
rect 60772 64894 62875 64896
rect 62809 64891 62875 64894
rect 66397 64954 66463 64957
rect 170406 64954 170466 65166
rect 177030 64954 177090 65128
rect 66397 64952 67948 64954
rect 66397 64896 66402 64952
rect 66458 64896 67948 64952
rect 66397 64894 67948 64896
rect 66397 64891 66463 64894
rect 97726 64546 97786 64856
rect 102737 64682 102803 64685
rect 135029 64682 135095 64685
rect 102737 64680 104932 64682
rect 102737 64624 102742 64680
rect 102798 64624 104932 64680
rect 102737 64622 104932 64624
rect 132716 64680 135095 64682
rect 132716 64624 135034 64680
rect 135090 64624 135095 64680
rect 132716 64622 135095 64624
rect 102737 64619 102803 64622
rect 135029 64619 135095 64622
rect 100621 64546 100687 64549
rect 97726 64544 100687 64546
rect 97726 64488 100626 64544
rect 100682 64488 100687 64544
rect 97726 64486 100687 64488
rect 100621 64483 100687 64486
rect 136869 64546 136935 64549
rect 140046 64546 140106 64856
rect 136869 64544 140106 64546
rect 136869 64488 136874 64544
rect 136930 64488 140106 64544
rect 136869 64486 140106 64488
rect 136869 64483 136935 64486
rect 62717 64410 62783 64413
rect 60772 64408 62783 64410
rect 60772 64352 62722 64408
rect 62778 64352 62783 64408
rect 60772 64350 62783 64352
rect 169854 64410 169914 64924
rect 170406 64894 177090 64954
rect 174129 64682 174195 64685
rect 174129 64680 177060 64682
rect 174129 64624 174134 64680
rect 174190 64624 177060 64680
rect 174129 64622 177060 64624
rect 174129 64619 174195 64622
rect 171645 64410 171711 64413
rect 169854 64408 171711 64410
rect 169854 64352 171650 64408
rect 171706 64352 171711 64408
rect 169854 64350 171711 64352
rect 62717 64347 62783 64350
rect 171645 64347 171711 64350
rect 66397 64274 66463 64277
rect 66397 64272 67948 64274
rect 66397 64216 66402 64272
rect 66458 64216 67948 64272
rect 66397 64214 67948 64216
rect 66397 64211 66463 64214
rect 97726 64138 97786 64176
rect 100897 64138 100963 64141
rect 97726 64136 100963 64138
rect 97726 64080 100902 64136
rect 100958 64080 100963 64136
rect 97726 64078 100963 64080
rect 100897 64075 100963 64078
rect 102829 64138 102895 64141
rect 134477 64138 134543 64141
rect 102829 64136 104932 64138
rect 102829 64080 102834 64136
rect 102890 64080 104932 64136
rect 102829 64078 104932 64080
rect 132716 64136 134543 64138
rect 132716 64080 134482 64136
rect 134538 64080 134543 64136
rect 132716 64078 134543 64080
rect 102829 64075 102895 64078
rect 134477 64075 134543 64078
rect 136961 64138 137027 64141
rect 140046 64138 140106 64176
rect 136961 64136 140106 64138
rect 136961 64080 136966 64136
rect 137022 64080 140106 64136
rect 136961 64078 140106 64080
rect 169854 64138 169914 64244
rect 171737 64138 171803 64141
rect 169854 64136 171803 64138
rect 169854 64080 171742 64136
rect 171798 64080 171803 64136
rect 169854 64078 171803 64080
rect 136961 64075 137027 64078
rect 171737 64075 171803 64078
rect 174221 64138 174287 64141
rect 174221 64136 177060 64138
rect 174221 64080 174226 64136
rect 174282 64080 177060 64136
rect 174221 64078 177060 64080
rect 174221 64075 174287 64078
rect 62993 63866 63059 63869
rect 60772 63864 63059 63866
rect 60772 63808 62998 63864
rect 63054 63808 63059 63864
rect 60772 63806 63059 63808
rect 62993 63803 63059 63806
rect 66305 63730 66371 63733
rect 66305 63728 67948 63730
rect 66305 63672 66310 63728
rect 66366 63672 67948 63728
rect 66305 63670 67948 63672
rect 66305 63667 66371 63670
rect 62349 63322 62415 63325
rect 60772 63320 62415 63322
rect 60772 63264 62354 63320
rect 62410 63264 62415 63320
rect 60772 63262 62415 63264
rect 97726 63322 97786 63632
rect 102369 63594 102435 63597
rect 135581 63594 135647 63597
rect 102369 63592 104932 63594
rect 102369 63536 102374 63592
rect 102430 63536 104932 63592
rect 102369 63534 104932 63536
rect 132716 63592 135647 63594
rect 132716 63536 135586 63592
rect 135642 63536 135647 63592
rect 132716 63534 135647 63536
rect 102369 63531 102435 63534
rect 135581 63531 135647 63534
rect 100437 63322 100503 63325
rect 97726 63320 100503 63322
rect 97726 63264 100442 63320
rect 100498 63264 100503 63320
rect 97726 63262 100503 63264
rect 62349 63259 62415 63262
rect 100437 63259 100503 63262
rect 136869 63322 136935 63325
rect 140046 63322 140106 63632
rect 169854 63458 169914 63700
rect 174129 63594 174195 63597
rect 174129 63592 177060 63594
rect 174129 63536 174134 63592
rect 174190 63536 177060 63592
rect 174129 63534 177060 63536
rect 174129 63531 174195 63534
rect 172013 63458 172079 63461
rect 169854 63456 172079 63458
rect 169854 63400 172018 63456
rect 172074 63400 172079 63456
rect 169854 63398 172079 63400
rect 172013 63395 172079 63398
rect 136869 63320 140106 63322
rect 136869 63264 136874 63320
rect 136930 63264 140106 63320
rect 136869 63262 140106 63264
rect 136869 63259 136935 63262
rect 66397 63186 66463 63189
rect 66397 63184 67948 63186
rect 66397 63128 66402 63184
rect 66458 63128 67948 63184
rect 66397 63126 67948 63128
rect 66397 63123 66463 63126
rect 9896 62914 10376 62944
rect 11933 62914 11999 62917
rect 9896 62912 11999 62914
rect 9896 62856 11938 62912
rect 11994 62856 11999 62912
rect 9896 62854 11999 62856
rect 9896 62824 10376 62854
rect 11933 62851 11999 62854
rect 29229 62914 29295 62917
rect 29229 62912 32988 62914
rect 29229 62856 29234 62912
rect 29290 62856 32988 62912
rect 29229 62854 32988 62856
rect 29229 62851 29295 62854
rect 63269 62778 63335 62781
rect 60772 62776 63335 62778
rect 60772 62720 63274 62776
rect 63330 62720 63335 62776
rect 60772 62718 63335 62720
rect 97726 62778 97786 63088
rect 102553 63050 102619 63053
rect 134661 63050 134727 63053
rect 102553 63048 104932 63050
rect 102553 62992 102558 63048
rect 102614 62992 104932 63048
rect 102553 62990 104932 62992
rect 132716 63048 134727 63050
rect 132716 62992 134666 63048
rect 134722 62992 134727 63048
rect 132716 62990 134727 62992
rect 102553 62987 102619 62990
rect 134661 62987 134727 62990
rect 100897 62778 100963 62781
rect 97726 62776 100963 62778
rect 97726 62720 100902 62776
rect 100958 62720 100963 62776
rect 97726 62718 100963 62720
rect 63269 62715 63335 62718
rect 100897 62715 100963 62718
rect 136961 62778 137027 62781
rect 140046 62778 140106 63088
rect 136961 62776 140106 62778
rect 136961 62720 136966 62776
rect 137022 62720 140106 62776
rect 136961 62718 140106 62720
rect 169854 62778 169914 63156
rect 174221 63050 174287 63053
rect 174221 63048 177060 63050
rect 174221 62992 174226 63048
rect 174282 62992 177060 63048
rect 174221 62990 177060 62992
rect 174221 62987 174287 62990
rect 172657 62778 172723 62781
rect 169854 62776 172723 62778
rect 169854 62720 172662 62776
rect 172718 62720 172723 62776
rect 169854 62718 172723 62720
rect 136961 62715 137027 62718
rect 172657 62715 172723 62718
rect 66305 62506 66371 62509
rect 66305 62504 67948 62506
rect 66305 62448 66310 62504
rect 66366 62448 67948 62504
rect 66305 62446 67948 62448
rect 66305 62443 66371 62446
rect 63545 62098 63611 62101
rect 60772 62096 63611 62098
rect 60772 62040 63550 62096
rect 63606 62040 63611 62096
rect 60772 62038 63611 62040
rect 97726 62098 97786 62408
rect 102461 62370 102527 62373
rect 135029 62370 135095 62373
rect 102461 62368 104932 62370
rect 102461 62312 102466 62368
rect 102522 62312 104932 62368
rect 102461 62310 104932 62312
rect 132716 62368 135095 62370
rect 132716 62312 135034 62368
rect 135090 62312 135095 62368
rect 132716 62310 135095 62312
rect 102461 62307 102527 62310
rect 135029 62307 135095 62310
rect 100253 62098 100319 62101
rect 97726 62096 100319 62098
rect 97726 62040 100258 62096
rect 100314 62040 100319 62096
rect 97726 62038 100319 62040
rect 63545 62035 63611 62038
rect 100253 62035 100319 62038
rect 136777 62098 136843 62101
rect 140046 62098 140106 62408
rect 136777 62096 140106 62098
rect 136777 62040 136782 62096
rect 136838 62040 140106 62096
rect 136777 62038 140106 62040
rect 169854 62098 169914 62476
rect 174313 62370 174379 62373
rect 174313 62368 177060 62370
rect 174313 62312 174318 62368
rect 174374 62312 177060 62368
rect 174313 62310 177060 62312
rect 174313 62307 174379 62310
rect 171645 62098 171711 62101
rect 169854 62096 171711 62098
rect 169854 62040 171650 62096
rect 171706 62040 171711 62096
rect 169854 62038 171711 62040
rect 136777 62035 136843 62038
rect 171645 62035 171711 62038
rect 66397 61962 66463 61965
rect 66397 61960 67948 61962
rect 66397 61904 66402 61960
rect 66458 61904 67948 61960
rect 66397 61902 67948 61904
rect 66397 61899 66463 61902
rect 63453 61554 63519 61557
rect 60772 61552 63519 61554
rect 60772 61496 63458 61552
rect 63514 61496 63519 61552
rect 60772 61494 63519 61496
rect 63453 61491 63519 61494
rect 97726 61418 97786 61864
rect 102645 61826 102711 61829
rect 135397 61826 135463 61829
rect 102645 61824 104932 61826
rect 102645 61768 102650 61824
rect 102706 61768 104932 61824
rect 102645 61766 104932 61768
rect 132716 61824 135463 61826
rect 132716 61768 135402 61824
rect 135458 61768 135463 61824
rect 132716 61766 135463 61768
rect 102645 61763 102711 61766
rect 135397 61763 135463 61766
rect 100897 61418 100963 61421
rect 97726 61416 100963 61418
rect 97726 61360 100902 61416
rect 100958 61360 100963 61416
rect 97726 61358 100963 61360
rect 100897 61355 100963 61358
rect 136869 61418 136935 61421
rect 140046 61418 140106 61864
rect 136869 61416 140106 61418
rect 136869 61360 136874 61416
rect 136930 61360 140106 61416
rect 136869 61358 140106 61360
rect 169854 61418 169914 61932
rect 174129 61826 174195 61829
rect 174129 61824 177060 61826
rect 174129 61768 174134 61824
rect 174190 61768 177060 61824
rect 174129 61766 177060 61768
rect 174129 61763 174195 61766
rect 172657 61418 172723 61421
rect 169854 61416 172723 61418
rect 169854 61360 172662 61416
rect 172718 61360 172723 61416
rect 169854 61358 172723 61360
rect 136869 61355 136935 61358
rect 172657 61355 172723 61358
rect 66213 61282 66279 61285
rect 102369 61282 102435 61285
rect 135305 61282 135371 61285
rect 66213 61280 67948 61282
rect 66213 61224 66218 61280
rect 66274 61224 67948 61280
rect 66213 61222 67948 61224
rect 102369 61280 104932 61282
rect 102369 61224 102374 61280
rect 102430 61224 104932 61280
rect 102369 61222 104932 61224
rect 132716 61280 135371 61282
rect 132716 61224 135310 61280
rect 135366 61224 135371 61280
rect 173853 61282 173919 61285
rect 173853 61280 177060 61282
rect 132716 61222 135371 61224
rect 66213 61219 66279 61222
rect 102369 61219 102435 61222
rect 135305 61219 135371 61222
rect 63177 61010 63243 61013
rect 60772 61008 63243 61010
rect 60772 60952 63182 61008
rect 63238 60952 63243 61008
rect 60772 60950 63243 60952
rect 63177 60947 63243 60950
rect 97726 60874 97786 61184
rect 100621 60874 100687 60877
rect 97726 60872 100687 60874
rect 97726 60816 100626 60872
rect 100682 60816 100687 60872
rect 97726 60814 100687 60816
rect 100621 60811 100687 60814
rect 136777 60874 136843 60877
rect 140046 60874 140106 61184
rect 136777 60872 140106 60874
rect 136777 60816 136782 60872
rect 136838 60816 140106 60872
rect 136777 60814 140106 60816
rect 169854 60874 169914 61252
rect 173853 61224 173858 61280
rect 173914 61224 177060 61280
rect 173853 61222 177060 61224
rect 173853 61219 173919 61222
rect 172197 60874 172263 60877
rect 169854 60872 172263 60874
rect 169854 60816 172202 60872
rect 172258 60816 172263 60872
rect 169854 60814 172263 60816
rect 136777 60811 136843 60814
rect 172197 60811 172263 60814
rect 66305 60738 66371 60741
rect 102553 60738 102619 60741
rect 134477 60738 134543 60741
rect 66305 60736 67948 60738
rect 66305 60680 66310 60736
rect 66366 60680 67948 60736
rect 66305 60678 67948 60680
rect 102553 60736 104932 60738
rect 102553 60680 102558 60736
rect 102614 60680 104932 60736
rect 102553 60678 104932 60680
rect 132716 60736 134543 60738
rect 132716 60680 134482 60736
rect 134538 60680 134543 60736
rect 174129 60738 174195 60741
rect 174129 60736 177060 60738
rect 132716 60678 134543 60680
rect 66305 60675 66371 60678
rect 102553 60675 102619 60678
rect 134477 60675 134543 60678
rect 62809 60466 62875 60469
rect 60772 60464 62875 60466
rect 60772 60408 62814 60464
rect 62870 60408 62875 60464
rect 60772 60406 62875 60408
rect 62809 60403 62875 60406
rect 97726 60330 97786 60640
rect 100897 60330 100963 60333
rect 97726 60328 100963 60330
rect 97726 60272 100902 60328
rect 100958 60272 100963 60328
rect 97726 60270 100963 60272
rect 100897 60267 100963 60270
rect 136961 60330 137027 60333
rect 140046 60330 140106 60640
rect 136961 60328 140106 60330
rect 136961 60272 136966 60328
rect 137022 60272 140106 60328
rect 136961 60270 140106 60272
rect 169854 60330 169914 60708
rect 174129 60680 174134 60736
rect 174190 60680 177060 60736
rect 174129 60678 177060 60680
rect 174129 60675 174195 60678
rect 172657 60330 172723 60333
rect 169854 60328 172723 60330
rect 169854 60272 172662 60328
rect 172718 60272 172723 60328
rect 169854 60270 172723 60272
rect 136961 60267 137027 60270
rect 172657 60267 172723 60270
rect 63729 60194 63795 60197
rect 60742 60192 63795 60194
rect 60742 60136 63734 60192
rect 63790 60136 63795 60192
rect 60742 60134 63795 60136
rect 60742 59892 60802 60134
rect 63729 60131 63795 60134
rect 66397 60194 66463 60197
rect 102461 60194 102527 60197
rect 134845 60194 134911 60197
rect 66397 60192 67948 60194
rect 66397 60136 66402 60192
rect 66458 60136 67948 60192
rect 66397 60134 67948 60136
rect 102461 60192 104932 60194
rect 102461 60136 102466 60192
rect 102522 60136 104932 60192
rect 102461 60134 104932 60136
rect 132716 60192 134911 60194
rect 132716 60136 134850 60192
rect 134906 60136 134911 60192
rect 174037 60194 174103 60197
rect 174037 60192 177060 60194
rect 132716 60134 134911 60136
rect 66397 60131 66463 60134
rect 102461 60131 102527 60134
rect 134845 60131 134911 60134
rect 97726 60058 97786 60096
rect 99701 60058 99767 60061
rect 97726 60056 99767 60058
rect 97726 60000 99706 60056
rect 99762 60000 99767 60056
rect 97726 59998 99767 60000
rect 99701 59995 99767 59998
rect 136869 60058 136935 60061
rect 140046 60058 140106 60096
rect 136869 60056 140106 60058
rect 136869 60000 136874 60056
rect 136930 60000 140106 60056
rect 136869 59998 140106 60000
rect 136869 59995 136935 59998
rect 169854 59922 169914 60164
rect 174037 60136 174042 60192
rect 174098 60136 177060 60192
rect 174037 60134 177060 60136
rect 174037 60131 174103 60134
rect 172657 59922 172723 59925
rect 169854 59920 172723 59922
rect 169854 59864 172662 59920
rect 172718 59864 172723 59920
rect 169854 59862 172723 59864
rect 172657 59859 172723 59862
rect 66305 59514 66371 59517
rect 102737 59514 102803 59517
rect 135213 59514 135279 59517
rect 66305 59512 67948 59514
rect 66305 59456 66310 59512
rect 66366 59456 67948 59512
rect 66305 59454 67948 59456
rect 102737 59512 104932 59514
rect 102737 59456 102742 59512
rect 102798 59456 104932 59512
rect 102737 59454 104932 59456
rect 132716 59512 135279 59514
rect 132716 59456 135218 59512
rect 135274 59456 135279 59512
rect 173945 59514 174011 59517
rect 173945 59512 177060 59514
rect 132716 59454 135279 59456
rect 66305 59451 66371 59454
rect 102737 59451 102803 59454
rect 135213 59451 135279 59454
rect 62717 59242 62783 59245
rect 60772 59240 62783 59242
rect 60772 59184 62722 59240
rect 62778 59184 62783 59240
rect 60772 59182 62783 59184
rect 62717 59179 62783 59182
rect 97726 59106 97786 59416
rect 100621 59106 100687 59109
rect 97726 59104 100687 59106
rect 97726 59048 100626 59104
rect 100682 59048 100687 59104
rect 97726 59046 100687 59048
rect 100621 59043 100687 59046
rect 136777 59106 136843 59109
rect 140046 59106 140106 59416
rect 136777 59104 140106 59106
rect 136777 59048 136782 59104
rect 136838 59048 140106 59104
rect 136777 59046 140106 59048
rect 169854 59106 169914 59484
rect 173945 59456 173950 59512
rect 174006 59456 177060 59512
rect 173945 59454 177060 59456
rect 173945 59451 174011 59454
rect 172657 59106 172723 59109
rect 169854 59104 172723 59106
rect 169854 59048 172662 59104
rect 172718 59048 172723 59104
rect 169854 59046 172723 59048
rect 136777 59043 136843 59046
rect 172657 59043 172723 59046
rect 66397 58970 66463 58973
rect 102645 58970 102711 58973
rect 134385 58970 134451 58973
rect 66397 58968 67948 58970
rect 66397 58912 66402 58968
rect 66458 58912 67948 58968
rect 66397 58910 67948 58912
rect 102645 58968 104932 58970
rect 102645 58912 102650 58968
rect 102706 58912 104932 58968
rect 102645 58910 104932 58912
rect 132716 58968 134451 58970
rect 132716 58912 134390 58968
rect 134446 58912 134451 58968
rect 174037 58970 174103 58973
rect 174037 58968 177060 58970
rect 132716 58910 134451 58912
rect 66397 58907 66463 58910
rect 102645 58907 102711 58910
rect 134385 58907 134451 58910
rect 63729 58698 63795 58701
rect 60772 58696 63795 58698
rect 60772 58640 63734 58696
rect 63790 58640 63795 58696
rect 60772 58638 63795 58640
rect 97726 58698 97786 58872
rect 100621 58698 100687 58701
rect 97726 58696 100687 58698
rect 97726 58640 100626 58696
rect 100682 58640 100687 58696
rect 97726 58638 100687 58640
rect 63729 58635 63795 58638
rect 100621 58635 100687 58638
rect 136869 58698 136935 58701
rect 140046 58698 140106 58872
rect 136869 58696 140106 58698
rect 136869 58640 136874 58696
rect 136930 58640 140106 58696
rect 136869 58638 140106 58640
rect 169854 58698 169914 58940
rect 174037 58912 174042 58968
rect 174098 58912 177060 58968
rect 174037 58910 177060 58912
rect 174037 58907 174103 58910
rect 172657 58698 172723 58701
rect 169854 58696 172723 58698
rect 169854 58640 172662 58696
rect 172718 58640 172723 58696
rect 169854 58638 172723 58640
rect 136869 58635 136935 58638
rect 172657 58635 172723 58638
rect 102369 58426 102435 58429
rect 134477 58426 134543 58429
rect 102369 58424 104932 58426
rect 102369 58368 102374 58424
rect 102430 58368 104932 58424
rect 102369 58366 104932 58368
rect 132716 58424 134543 58426
rect 132716 58368 134482 58424
rect 134538 58368 134543 58424
rect 132716 58366 134543 58368
rect 102369 58363 102435 58366
rect 134477 58363 134543 58366
rect 174129 58426 174195 58429
rect 174129 58424 177060 58426
rect 174129 58368 174134 58424
rect 174190 58368 177060 58424
rect 174129 58366 177060 58368
rect 174129 58363 174195 58366
rect 65017 58290 65083 58293
rect 65017 58288 67948 58290
rect 65017 58232 65022 58288
rect 65078 58232 67948 58288
rect 65017 58230 67948 58232
rect 65017 58227 65083 58230
rect 62809 58154 62875 58157
rect 60772 58152 62875 58154
rect 60772 58096 62814 58152
rect 62870 58096 62875 58152
rect 60772 58094 62875 58096
rect 62809 58091 62875 58094
rect 97726 57882 97786 58192
rect 100621 57882 100687 57885
rect 97726 57880 100687 57882
rect 97726 57824 100626 57880
rect 100682 57824 100687 57880
rect 97726 57822 100687 57824
rect 100621 57819 100687 57822
rect 102553 57882 102619 57885
rect 135397 57882 135463 57885
rect 102553 57880 104932 57882
rect 102553 57824 102558 57880
rect 102614 57824 104932 57880
rect 102553 57822 104932 57824
rect 132716 57880 135463 57882
rect 132716 57824 135402 57880
rect 135458 57824 135463 57880
rect 132716 57822 135463 57824
rect 102553 57819 102619 57822
rect 135397 57819 135463 57822
rect 136777 57882 136843 57885
rect 140046 57882 140106 58192
rect 136777 57880 140106 57882
rect 136777 57824 136782 57880
rect 136838 57824 140106 57880
rect 136777 57822 140106 57824
rect 169854 57882 169914 58260
rect 172105 57882 172171 57885
rect 169854 57880 172171 57882
rect 169854 57824 172110 57880
rect 172166 57824 172171 57880
rect 169854 57822 172171 57824
rect 136777 57819 136843 57822
rect 172105 57819 172171 57822
rect 173761 57882 173827 57885
rect 173761 57880 177060 57882
rect 173761 57824 173766 57880
rect 173822 57824 177060 57880
rect 173761 57822 177060 57824
rect 173761 57819 173827 57822
rect 66397 57746 66463 57749
rect 66397 57744 67948 57746
rect 66397 57688 66402 57744
rect 66458 57688 67948 57744
rect 66397 57686 67948 57688
rect 66397 57683 66463 57686
rect 62625 57610 62691 57613
rect 60772 57608 62691 57610
rect 60772 57552 62630 57608
rect 62686 57552 62691 57608
rect 60772 57550 62691 57552
rect 62625 57547 62691 57550
rect 97726 57338 97786 57648
rect 100621 57338 100687 57341
rect 97726 57336 100687 57338
rect 97726 57280 100626 57336
rect 100682 57280 100687 57336
rect 97726 57278 100687 57280
rect 100621 57275 100687 57278
rect 102461 57338 102527 57341
rect 135029 57338 135095 57341
rect 102461 57336 104932 57338
rect 102461 57280 102466 57336
rect 102522 57280 104932 57336
rect 102461 57278 104932 57280
rect 132716 57336 135095 57338
rect 132716 57280 135034 57336
rect 135090 57280 135095 57336
rect 132716 57278 135095 57280
rect 102461 57275 102527 57278
rect 135029 57275 135095 57278
rect 136869 57338 136935 57341
rect 140046 57338 140106 57648
rect 169854 57474 169914 57716
rect 172657 57474 172723 57477
rect 169854 57472 172723 57474
rect 169854 57416 172662 57472
rect 172718 57416 172723 57472
rect 169854 57414 172723 57416
rect 172657 57411 172723 57414
rect 172565 57338 172631 57341
rect 136869 57336 140106 57338
rect 136869 57280 136874 57336
rect 136930 57280 140106 57336
rect 136869 57278 140106 57280
rect 169670 57336 172631 57338
rect 169670 57280 172570 57336
rect 172626 57280 172631 57336
rect 169670 57278 172631 57280
rect 136869 57275 136935 57278
rect 66397 57202 66463 57205
rect 100529 57202 100595 57205
rect 66397 57200 67948 57202
rect 66397 57144 66402 57200
rect 66458 57144 67948 57200
rect 66397 57142 67948 57144
rect 97756 57200 100595 57202
rect 97756 57144 100534 57200
rect 100590 57144 100595 57200
rect 97756 57142 100595 57144
rect 66397 57139 66463 57142
rect 100529 57139 100595 57142
rect 136961 57202 137027 57205
rect 136961 57200 140076 57202
rect 136961 57144 136966 57200
rect 137022 57144 140076 57200
rect 169670 57172 169730 57278
rect 172565 57275 172631 57278
rect 174037 57338 174103 57341
rect 174037 57336 177060 57338
rect 174037 57280 174042 57336
rect 174098 57280 177060 57336
rect 174037 57278 177060 57280
rect 174037 57275 174103 57278
rect 136961 57142 140076 57144
rect 136961 57139 137027 57142
rect 63545 57066 63611 57069
rect 60772 57064 63611 57066
rect 60772 57008 63550 57064
rect 63606 57008 63611 57064
rect 60772 57006 63611 57008
rect 63545 57003 63611 57006
rect 102645 56658 102711 56661
rect 135213 56658 135279 56661
rect 102645 56656 104932 56658
rect 102645 56600 102650 56656
rect 102706 56600 104932 56656
rect 102645 56598 104932 56600
rect 132716 56656 135279 56658
rect 132716 56600 135218 56656
rect 135274 56600 135279 56656
rect 132716 56598 135279 56600
rect 102645 56595 102711 56598
rect 135213 56595 135279 56598
rect 173853 56658 173919 56661
rect 173853 56656 177060 56658
rect 173853 56600 173858 56656
rect 173914 56600 177060 56656
rect 173853 56598 177060 56600
rect 173853 56595 173919 56598
rect 66305 56522 66371 56525
rect 66305 56520 67948 56522
rect 66305 56464 66310 56520
rect 66366 56464 67948 56520
rect 66305 56462 67948 56464
rect 66305 56459 66371 56462
rect 62901 56386 62967 56389
rect 60772 56384 62967 56386
rect 60772 56328 62906 56384
rect 62962 56328 62967 56384
rect 60772 56326 62967 56328
rect 62901 56323 62967 56326
rect 97726 56114 97786 56424
rect 100621 56114 100687 56117
rect 97726 56112 100687 56114
rect 97726 56056 100626 56112
rect 100682 56056 100687 56112
rect 97726 56054 100687 56056
rect 100621 56051 100687 56054
rect 102369 56114 102435 56117
rect 134569 56114 134635 56117
rect 102369 56112 104932 56114
rect 102369 56056 102374 56112
rect 102430 56056 104932 56112
rect 102369 56054 104932 56056
rect 132716 56112 134635 56114
rect 132716 56056 134574 56112
rect 134630 56056 134635 56112
rect 132716 56054 134635 56056
rect 102369 56051 102435 56054
rect 134569 56051 134635 56054
rect 136777 56114 136843 56117
rect 140046 56114 140106 56424
rect 136777 56112 140106 56114
rect 136777 56056 136782 56112
rect 136838 56056 140106 56112
rect 136777 56054 140106 56056
rect 169854 56114 169914 56492
rect 174037 56386 174103 56389
rect 174037 56384 177090 56386
rect 174037 56328 174042 56384
rect 174098 56328 177090 56384
rect 174037 56326 177090 56328
rect 174037 56323 174103 56326
rect 172657 56114 172723 56117
rect 169854 56112 172723 56114
rect 169854 56056 172662 56112
rect 172718 56056 172723 56112
rect 177030 56084 177090 56326
rect 169854 56054 172723 56056
rect 136777 56051 136843 56054
rect 172657 56051 172723 56054
rect 66397 55978 66463 55981
rect 66397 55976 67948 55978
rect 66397 55920 66402 55976
rect 66458 55920 67948 55976
rect 66397 55918 67948 55920
rect 66397 55915 66463 55918
rect 62625 55842 62691 55845
rect 60772 55840 62691 55842
rect 60772 55784 62630 55840
rect 62686 55784 62691 55840
rect 60772 55782 62691 55784
rect 97726 55842 97786 55880
rect 100897 55842 100963 55845
rect 97726 55840 100963 55842
rect 97726 55784 100902 55840
rect 100958 55784 100963 55840
rect 97726 55782 100963 55784
rect 62625 55779 62691 55782
rect 100897 55779 100963 55782
rect 136869 55842 136935 55845
rect 140046 55842 140106 55880
rect 136869 55840 140106 55842
rect 136869 55784 136874 55840
rect 136930 55784 140106 55840
rect 136869 55782 140106 55784
rect 169854 55842 169914 55948
rect 172657 55842 172723 55845
rect 169854 55840 172723 55842
rect 169854 55784 172662 55840
rect 172718 55784 172723 55840
rect 169854 55782 172723 55784
rect 136869 55779 136935 55782
rect 172657 55779 172723 55782
rect 102461 55570 102527 55573
rect 135305 55570 135371 55573
rect 102461 55568 104932 55570
rect 102461 55512 102466 55568
rect 102522 55512 104932 55568
rect 102461 55510 104932 55512
rect 132716 55568 135371 55570
rect 132716 55512 135310 55568
rect 135366 55512 135371 55568
rect 132716 55510 135371 55512
rect 102461 55507 102527 55510
rect 135305 55507 135371 55510
rect 173945 55570 174011 55573
rect 173945 55568 177060 55570
rect 173945 55512 173950 55568
rect 174006 55512 177060 55568
rect 173945 55510 177060 55512
rect 173945 55507 174011 55510
rect 62809 55298 62875 55301
rect 60772 55296 62875 55298
rect 60772 55240 62814 55296
rect 62870 55240 62875 55296
rect 60772 55238 62875 55240
rect 62809 55235 62875 55238
rect 66305 55298 66371 55301
rect 66305 55296 67948 55298
rect 66305 55240 66310 55296
rect 66366 55240 67948 55296
rect 66305 55238 67948 55240
rect 66305 55235 66371 55238
rect 97726 54890 97786 55200
rect 102553 55026 102619 55029
rect 135397 55026 135463 55029
rect 102553 55024 104932 55026
rect 102553 54968 102558 55024
rect 102614 54968 104932 55024
rect 102553 54966 104932 54968
rect 132716 55024 135463 55026
rect 132716 54968 135402 55024
rect 135458 54968 135463 55024
rect 132716 54966 135463 54968
rect 102553 54963 102619 54966
rect 135397 54963 135463 54966
rect 100621 54890 100687 54893
rect 97726 54888 100687 54890
rect 97726 54832 100626 54888
rect 100682 54832 100687 54888
rect 97726 54830 100687 54832
rect 100621 54827 100687 54830
rect 136777 54890 136843 54893
rect 140046 54890 140106 55200
rect 136777 54888 140106 54890
rect 136777 54832 136782 54888
rect 136838 54832 140106 54888
rect 136777 54830 140106 54832
rect 169854 54890 169914 55268
rect 173761 55026 173827 55029
rect 173761 55024 177060 55026
rect 173761 54968 173766 55024
rect 173822 54968 177060 55024
rect 173761 54966 177060 54968
rect 173761 54963 173827 54966
rect 171737 54890 171803 54893
rect 169854 54888 171803 54890
rect 169854 54832 171742 54888
rect 171798 54832 171803 54888
rect 169854 54830 171803 54832
rect 136777 54827 136843 54830
rect 171737 54827 171803 54830
rect 62717 54754 62783 54757
rect 60772 54752 62783 54754
rect 60772 54696 62722 54752
rect 62778 54696 62783 54752
rect 60772 54694 62783 54696
rect 62717 54691 62783 54694
rect 66397 54754 66463 54757
rect 66397 54752 67948 54754
rect 66397 54696 66402 54752
rect 66458 54696 67948 54752
rect 66397 54694 67948 54696
rect 66397 54691 66463 54694
rect 97726 54618 97786 54656
rect 100805 54618 100871 54621
rect 97726 54616 100871 54618
rect 97726 54560 100810 54616
rect 100866 54560 100871 54616
rect 97726 54558 100871 54560
rect 100805 54555 100871 54558
rect 137145 54618 137211 54621
rect 140046 54618 140106 54656
rect 137145 54616 140106 54618
rect 137145 54560 137150 54616
rect 137206 54560 140106 54616
rect 137145 54558 140106 54560
rect 137145 54555 137211 54558
rect 102369 54482 102435 54485
rect 135029 54482 135095 54485
rect 102369 54480 104932 54482
rect 102369 54424 102374 54480
rect 102430 54424 104932 54480
rect 102369 54422 104932 54424
rect 132716 54480 135095 54482
rect 132716 54424 135034 54480
rect 135090 54424 135095 54480
rect 132716 54422 135095 54424
rect 169854 54482 169914 54724
rect 172841 54482 172907 54485
rect 169854 54480 172907 54482
rect 169854 54424 172846 54480
rect 172902 54424 172907 54480
rect 169854 54422 172907 54424
rect 102369 54419 102435 54422
rect 135029 54419 135095 54422
rect 172841 54419 172907 54422
rect 174037 54482 174103 54485
rect 174037 54480 177060 54482
rect 174037 54424 174042 54480
rect 174098 54424 177060 54480
rect 174037 54422 177060 54424
rect 174037 54419 174103 54422
rect 63545 54210 63611 54213
rect 60772 54208 63611 54210
rect 60772 54152 63550 54208
rect 63606 54152 63611 54208
rect 60772 54150 63611 54152
rect 63545 54147 63611 54150
rect 66305 54210 66371 54213
rect 66305 54208 67948 54210
rect 66305 54152 66310 54208
rect 66366 54152 67948 54208
rect 66305 54150 67948 54152
rect 66305 54147 66371 54150
rect 97726 53666 97786 54112
rect 102645 53802 102711 53805
rect 134293 53802 134359 53805
rect 102645 53800 104932 53802
rect 102645 53744 102650 53800
rect 102706 53744 104932 53800
rect 102645 53742 104932 53744
rect 132716 53800 134359 53802
rect 132716 53744 134298 53800
rect 134354 53744 134359 53800
rect 132716 53742 134359 53744
rect 102645 53739 102711 53742
rect 134293 53739 134359 53742
rect 100621 53666 100687 53669
rect 97726 53664 100687 53666
rect 97726 53608 100626 53664
rect 100682 53608 100687 53664
rect 97726 53606 100687 53608
rect 100621 53603 100687 53606
rect 136777 53666 136843 53669
rect 140046 53666 140106 54112
rect 136777 53664 140106 53666
rect 136777 53608 136782 53664
rect 136838 53608 140106 53664
rect 136777 53606 140106 53608
rect 169854 53666 169914 54180
rect 174129 53802 174195 53805
rect 174129 53800 177060 53802
rect 174129 53744 174134 53800
rect 174190 53744 177060 53800
rect 174129 53742 177060 53744
rect 174129 53739 174195 53742
rect 172565 53666 172631 53669
rect 169854 53664 172631 53666
rect 169854 53608 172570 53664
rect 172626 53608 172631 53664
rect 169854 53606 172631 53608
rect 136777 53603 136843 53606
rect 172565 53603 172631 53606
rect 30517 53530 30583 53533
rect 63269 53530 63335 53533
rect 30517 53528 32988 53530
rect 30517 53472 30522 53528
rect 30578 53472 32988 53528
rect 30517 53470 32988 53472
rect 60772 53528 63335 53530
rect 60772 53472 63274 53528
rect 63330 53472 63335 53528
rect 60772 53470 63335 53472
rect 30517 53467 30583 53470
rect 63269 53467 63335 53470
rect 66397 53530 66463 53533
rect 66397 53528 67948 53530
rect 66397 53472 66402 53528
rect 66458 53472 67948 53528
rect 66397 53470 67948 53472
rect 66397 53467 66463 53470
rect 97726 53122 97786 53432
rect 102461 53258 102527 53261
rect 135121 53258 135187 53261
rect 102461 53256 104932 53258
rect 102461 53200 102466 53256
rect 102522 53200 104932 53256
rect 102461 53198 104932 53200
rect 132716 53256 135187 53258
rect 132716 53200 135126 53256
rect 135182 53200 135187 53256
rect 132716 53198 135187 53200
rect 102461 53195 102527 53198
rect 135121 53195 135187 53198
rect 100621 53122 100687 53125
rect 97726 53120 100687 53122
rect 97726 53064 100626 53120
rect 100682 53064 100687 53120
rect 97726 53062 100687 53064
rect 100621 53059 100687 53062
rect 136869 53122 136935 53125
rect 140046 53122 140106 53432
rect 136869 53120 140106 53122
rect 136869 53064 136874 53120
rect 136930 53064 140106 53120
rect 136869 53062 140106 53064
rect 169854 53122 169914 53500
rect 174221 53258 174287 53261
rect 174221 53256 177060 53258
rect 174221 53200 174226 53256
rect 174282 53200 177060 53256
rect 174221 53198 177060 53200
rect 174221 53195 174287 53198
rect 172657 53122 172723 53125
rect 169854 53120 172723 53122
rect 169854 53064 172662 53120
rect 172718 53064 172723 53120
rect 169854 53062 172723 53064
rect 136869 53059 136935 53062
rect 172657 53059 172723 53062
rect 63453 52986 63519 52989
rect 60772 52984 63519 52986
rect 60772 52928 63458 52984
rect 63514 52928 63519 52984
rect 60772 52926 63519 52928
rect 63453 52923 63519 52926
rect 65661 52986 65727 52989
rect 65661 52984 67948 52986
rect 65661 52928 65666 52984
rect 65722 52928 67948 52984
rect 65661 52926 67948 52928
rect 65661 52923 65727 52926
rect 63361 52442 63427 52445
rect 60772 52440 63427 52442
rect 60772 52384 63366 52440
rect 63422 52384 63427 52440
rect 60772 52382 63427 52384
rect 97726 52442 97786 52888
rect 102553 52714 102619 52717
rect 134201 52714 134267 52717
rect 102553 52712 104932 52714
rect 102553 52656 102558 52712
rect 102614 52656 104932 52712
rect 102553 52654 104932 52656
rect 132716 52712 134267 52714
rect 132716 52656 134206 52712
rect 134262 52656 134267 52712
rect 132716 52654 134267 52656
rect 102553 52651 102619 52654
rect 134201 52651 134267 52654
rect 100621 52442 100687 52445
rect 97726 52440 100687 52442
rect 97726 52384 100626 52440
rect 100682 52384 100687 52440
rect 97726 52382 100687 52384
rect 63361 52379 63427 52382
rect 100621 52379 100687 52382
rect 136685 52442 136751 52445
rect 140046 52442 140106 52888
rect 136685 52440 140106 52442
rect 136685 52384 136690 52440
rect 136746 52384 140106 52440
rect 136685 52382 140106 52384
rect 169854 52442 169914 52956
rect 174129 52714 174195 52717
rect 174129 52712 177060 52714
rect 174129 52656 174134 52712
rect 174190 52656 177060 52712
rect 174129 52654 177060 52656
rect 174129 52651 174195 52654
rect 172013 52442 172079 52445
rect 169854 52440 172079 52442
rect 169854 52384 172018 52440
rect 172074 52384 172079 52440
rect 169854 52382 172079 52384
rect 136685 52379 136751 52382
rect 172013 52379 172079 52382
rect 66397 52306 66463 52309
rect 66397 52304 67948 52306
rect 66397 52248 66402 52304
rect 66458 52248 67948 52304
rect 66397 52246 67948 52248
rect 66397 52243 66463 52246
rect 63729 51898 63795 51901
rect 60772 51896 63795 51898
rect 60772 51840 63734 51896
rect 63790 51840 63795 51896
rect 60772 51838 63795 51840
rect 97726 51898 97786 52208
rect 102737 52170 102803 52173
rect 135029 52170 135095 52173
rect 102737 52168 104932 52170
rect 102737 52112 102742 52168
rect 102798 52112 104932 52168
rect 102737 52110 104932 52112
rect 132716 52168 135095 52170
rect 132716 52112 135034 52168
rect 135090 52112 135095 52168
rect 132716 52110 135095 52112
rect 102737 52107 102803 52110
rect 135029 52107 135095 52110
rect 100621 51898 100687 51901
rect 97726 51896 100687 51898
rect 97726 51840 100626 51896
rect 100682 51840 100687 51896
rect 97726 51838 100687 51840
rect 63729 51835 63795 51838
rect 100621 51835 100687 51838
rect 136777 51898 136843 51901
rect 140046 51898 140106 52208
rect 169854 52170 169914 52276
rect 174037 52170 174103 52173
rect 169854 52110 170282 52170
rect 170222 51898 170282 52110
rect 174037 52168 177060 52170
rect 174037 52112 174042 52168
rect 174098 52112 177060 52168
rect 174037 52110 177060 52112
rect 174037 52107 174103 52110
rect 172657 51898 172723 51901
rect 136777 51896 140106 51898
rect 136777 51840 136782 51896
rect 136838 51840 140106 51896
rect 136777 51838 140106 51840
rect 169670 51838 170098 51898
rect 170222 51896 172723 51898
rect 170222 51840 172662 51896
rect 172718 51840 172723 51896
rect 170222 51838 172723 51840
rect 136777 51835 136843 51838
rect 66397 51762 66463 51765
rect 100529 51762 100595 51765
rect 66397 51760 67948 51762
rect 66397 51704 66402 51760
rect 66458 51704 67948 51760
rect 66397 51702 67948 51704
rect 97756 51760 100595 51762
rect 97756 51704 100534 51760
rect 100590 51704 100595 51760
rect 97756 51702 100595 51704
rect 66397 51699 66463 51702
rect 100529 51699 100595 51702
rect 136869 51762 136935 51765
rect 136869 51760 140076 51762
rect 136869 51704 136874 51760
rect 136930 51704 140076 51760
rect 169670 51732 169730 51838
rect 170038 51762 170098 51838
rect 172657 51835 172723 51838
rect 172657 51762 172723 51765
rect 170038 51760 172723 51762
rect 136869 51702 140076 51704
rect 170038 51704 172662 51760
rect 172718 51704 172723 51760
rect 170038 51702 172723 51704
rect 136869 51699 136935 51702
rect 172657 51699 172723 51702
rect 102369 51626 102435 51629
rect 135397 51626 135463 51629
rect 102369 51624 104932 51626
rect 102369 51568 102374 51624
rect 102430 51568 104932 51624
rect 102369 51566 104932 51568
rect 132716 51624 135463 51626
rect 132716 51568 135402 51624
rect 135458 51568 135463 51624
rect 132716 51566 135463 51568
rect 102369 51563 102435 51566
rect 135397 51563 135463 51566
rect 173853 51626 173919 51629
rect 173853 51624 177060 51626
rect 173853 51568 173858 51624
rect 173914 51568 177060 51624
rect 173853 51566 177060 51568
rect 173853 51563 173919 51566
rect 62809 51354 62875 51357
rect 60772 51352 62875 51354
rect 60772 51296 62814 51352
rect 62870 51296 62875 51352
rect 60772 51294 62875 51296
rect 62809 51291 62875 51294
rect 66397 51218 66463 51221
rect 66397 51216 67948 51218
rect 66397 51160 66402 51216
rect 66458 51160 67948 51216
rect 66397 51158 67948 51160
rect 66397 51155 66463 51158
rect 63729 50674 63795 50677
rect 60772 50672 63795 50674
rect 60772 50616 63734 50672
rect 63790 50616 63795 50672
rect 60772 50614 63795 50616
rect 97726 50674 97786 51120
rect 102645 50946 102711 50949
rect 135397 50946 135463 50949
rect 102645 50944 104932 50946
rect 102645 50888 102650 50944
rect 102706 50888 104932 50944
rect 102645 50886 104932 50888
rect 132716 50944 135463 50946
rect 132716 50888 135402 50944
rect 135458 50888 135463 50944
rect 132716 50886 135463 50888
rect 102645 50883 102711 50886
rect 135397 50883 135463 50886
rect 100621 50674 100687 50677
rect 97726 50672 100687 50674
rect 97726 50616 100626 50672
rect 100682 50616 100687 50672
rect 97726 50614 100687 50616
rect 63729 50611 63795 50614
rect 100621 50611 100687 50614
rect 136777 50674 136843 50677
rect 140046 50674 140106 51120
rect 136777 50672 140106 50674
rect 136777 50616 136782 50672
rect 136838 50616 140106 50672
rect 136777 50614 140106 50616
rect 169854 50674 169914 51188
rect 174037 50946 174103 50949
rect 174037 50944 177060 50946
rect 174037 50888 174042 50944
rect 174098 50888 177060 50944
rect 174037 50886 177060 50888
rect 174037 50883 174103 50886
rect 171645 50674 171711 50677
rect 169854 50672 171711 50674
rect 169854 50616 171650 50672
rect 171706 50616 171711 50672
rect 169854 50614 171711 50616
rect 136777 50611 136843 50614
rect 171645 50611 171711 50614
rect 66397 50538 66463 50541
rect 66397 50536 67948 50538
rect 66397 50480 66402 50536
rect 66458 50480 67948 50536
rect 66397 50478 67948 50480
rect 66397 50475 66463 50478
rect 97726 50402 97786 50440
rect 100621 50402 100687 50405
rect 97726 50400 100687 50402
rect 97726 50344 100626 50400
rect 100682 50344 100687 50400
rect 97726 50342 100687 50344
rect 100621 50339 100687 50342
rect 102461 50402 102527 50405
rect 135029 50402 135095 50405
rect 102461 50400 104932 50402
rect 102461 50344 102466 50400
rect 102522 50344 104932 50400
rect 102461 50342 104932 50344
rect 132716 50400 135095 50402
rect 132716 50344 135034 50400
rect 135090 50344 135095 50400
rect 132716 50342 135095 50344
rect 102461 50339 102527 50342
rect 135029 50339 135095 50342
rect 136869 50402 136935 50405
rect 140046 50402 140106 50440
rect 136869 50400 140106 50402
rect 136869 50344 136874 50400
rect 136930 50344 140106 50400
rect 136869 50342 140106 50344
rect 136869 50339 136935 50342
rect 169854 50266 169914 50508
rect 173945 50402 174011 50405
rect 173945 50400 177060 50402
rect 173945 50344 173950 50400
rect 174006 50344 177060 50400
rect 173945 50342 177060 50344
rect 173945 50339 174011 50342
rect 172657 50266 172723 50269
rect 169854 50264 172723 50266
rect 169854 50208 172662 50264
rect 172718 50208 172723 50264
rect 169854 50206 172723 50208
rect 172657 50203 172723 50206
rect 62901 50130 62967 50133
rect 60772 50128 62967 50130
rect 60772 50072 62906 50128
rect 62962 50072 62967 50128
rect 60772 50070 62967 50072
rect 62901 50067 62967 50070
rect 65477 49994 65543 49997
rect 65477 49992 67948 49994
rect 65477 49936 65482 49992
rect 65538 49936 67948 49992
rect 65477 49934 67948 49936
rect 65477 49931 65543 49934
rect 62717 49586 62783 49589
rect 60772 49584 62783 49586
rect 60772 49528 62722 49584
rect 62778 49528 62783 49584
rect 60772 49526 62783 49528
rect 62717 49523 62783 49526
rect 97726 49450 97786 49896
rect 102553 49858 102619 49861
rect 135305 49858 135371 49861
rect 102553 49856 104932 49858
rect 102553 49800 102558 49856
rect 102614 49800 104932 49856
rect 102553 49798 104932 49800
rect 132716 49856 135371 49858
rect 132716 49800 135310 49856
rect 135366 49800 135371 49856
rect 132716 49798 135371 49800
rect 102553 49795 102619 49798
rect 135305 49795 135371 49798
rect 100621 49450 100687 49453
rect 97726 49448 100687 49450
rect 97726 49392 100626 49448
rect 100682 49392 100687 49448
rect 97726 49390 100687 49392
rect 100621 49387 100687 49390
rect 136869 49450 136935 49453
rect 140046 49450 140106 49896
rect 136869 49448 140106 49450
rect 136869 49392 136874 49448
rect 136930 49392 140106 49448
rect 136869 49390 140106 49392
rect 169854 49450 169914 49964
rect 173761 49858 173827 49861
rect 173761 49856 177060 49858
rect 173761 49800 173766 49856
rect 173822 49800 177060 49856
rect 173761 49798 177060 49800
rect 173761 49795 173827 49798
rect 171829 49450 171895 49453
rect 169854 49448 171895 49450
rect 169854 49392 171834 49448
rect 171890 49392 171895 49448
rect 169854 49390 171895 49392
rect 136869 49387 136935 49390
rect 171829 49387 171895 49390
rect 66397 49314 66463 49317
rect 102645 49314 102711 49317
rect 134845 49314 134911 49317
rect 66397 49312 67948 49314
rect 66397 49256 66402 49312
rect 66458 49256 67948 49312
rect 66397 49254 67948 49256
rect 102645 49312 104932 49314
rect 102645 49256 102650 49312
rect 102706 49256 104932 49312
rect 102645 49254 104932 49256
rect 132716 49312 134911 49314
rect 132716 49256 134850 49312
rect 134906 49256 134911 49312
rect 174037 49314 174103 49317
rect 174037 49312 177060 49314
rect 132716 49254 134911 49256
rect 66397 49251 66463 49254
rect 102645 49251 102711 49254
rect 134845 49251 134911 49254
rect 63821 49042 63887 49045
rect 60772 49040 63887 49042
rect 60772 48984 63826 49040
rect 63882 48984 63887 49040
rect 60772 48982 63887 48984
rect 97726 49042 97786 49216
rect 100621 49042 100687 49045
rect 97726 49040 100687 49042
rect 97726 48984 100626 49040
rect 100682 48984 100687 49040
rect 97726 48982 100687 48984
rect 63821 48979 63887 48982
rect 100621 48979 100687 48982
rect 136777 48906 136843 48909
rect 140046 48906 140106 49216
rect 169854 49042 169914 49284
rect 174037 49256 174042 49312
rect 174098 49256 177060 49312
rect 174037 49254 177060 49256
rect 174037 49251 174103 49254
rect 172657 49042 172723 49045
rect 169854 49040 172723 49042
rect 169854 48984 172662 49040
rect 172718 48984 172723 49040
rect 169854 48982 172723 48984
rect 172657 48979 172723 48982
rect 136777 48904 140106 48906
rect 136777 48848 136782 48904
rect 136838 48848 140106 48904
rect 136777 48846 140106 48848
rect 136777 48843 136843 48846
rect 66397 48770 66463 48773
rect 102369 48770 102435 48773
rect 135397 48770 135463 48773
rect 66397 48768 67948 48770
rect 66397 48712 66402 48768
rect 66458 48712 67948 48768
rect 66397 48710 67948 48712
rect 102369 48768 104932 48770
rect 102369 48712 102374 48768
rect 102430 48712 104932 48768
rect 102369 48710 104932 48712
rect 132716 48768 135463 48770
rect 132716 48712 135402 48768
rect 135458 48712 135463 48768
rect 174129 48770 174195 48773
rect 174129 48768 177060 48770
rect 132716 48710 135463 48712
rect 66397 48707 66463 48710
rect 102369 48707 102435 48710
rect 135397 48707 135463 48710
rect 62809 48498 62875 48501
rect 60772 48496 62875 48498
rect 60772 48440 62814 48496
rect 62870 48440 62875 48496
rect 60772 48438 62875 48440
rect 62809 48435 62875 48438
rect 97726 48362 97786 48672
rect 100621 48362 100687 48365
rect 97726 48360 100687 48362
rect 97726 48304 100626 48360
rect 100682 48304 100687 48360
rect 97726 48302 100687 48304
rect 100621 48299 100687 48302
rect 136685 48362 136751 48365
rect 140046 48362 140106 48672
rect 136685 48360 140106 48362
rect 136685 48304 136690 48360
rect 136746 48304 140106 48360
rect 136685 48302 140106 48304
rect 169854 48362 169914 48740
rect 174129 48712 174134 48768
rect 174190 48712 177060 48768
rect 174129 48710 177060 48712
rect 174129 48707 174195 48710
rect 172105 48362 172171 48365
rect 169854 48360 172171 48362
rect 169854 48304 172110 48360
rect 172166 48304 172171 48360
rect 169854 48302 172171 48304
rect 136685 48299 136751 48302
rect 172105 48299 172171 48302
rect 64925 48226 64991 48229
rect 64925 48224 67948 48226
rect 64925 48168 64930 48224
rect 64986 48168 67948 48224
rect 64925 48166 67948 48168
rect 64925 48163 64991 48166
rect 63729 47818 63795 47821
rect 60772 47816 63795 47818
rect 60772 47760 63734 47816
rect 63790 47760 63795 47816
rect 60772 47758 63795 47760
rect 63729 47755 63795 47758
rect 65017 47818 65083 47821
rect 66397 47818 66463 47821
rect 65017 47816 66463 47818
rect 65017 47760 65022 47816
rect 65078 47760 66402 47816
rect 66458 47760 66463 47816
rect 65017 47758 66463 47760
rect 65017 47755 65083 47758
rect 66397 47755 66463 47758
rect 97726 47682 97786 48128
rect 102461 48090 102527 48093
rect 135305 48090 135371 48093
rect 102461 48088 104932 48090
rect 102461 48032 102466 48088
rect 102522 48032 104932 48088
rect 102461 48030 104932 48032
rect 132716 48088 135371 48090
rect 132716 48032 135310 48088
rect 135366 48032 135371 48088
rect 132716 48030 135371 48032
rect 102461 48027 102527 48030
rect 135305 48027 135371 48030
rect 100621 47682 100687 47685
rect 97726 47680 100687 47682
rect 97726 47624 100626 47680
rect 100682 47624 100687 47680
rect 97726 47622 100687 47624
rect 100621 47619 100687 47622
rect 136777 47682 136843 47685
rect 140046 47682 140106 48128
rect 169854 47954 169914 48196
rect 174037 48090 174103 48093
rect 174037 48088 177060 48090
rect 174037 48032 174042 48088
rect 174098 48032 177060 48088
rect 174037 48030 177060 48032
rect 174037 48027 174103 48030
rect 172657 47954 172723 47957
rect 169854 47952 172723 47954
rect 169854 47896 172662 47952
rect 172718 47896 172723 47952
rect 169854 47894 172723 47896
rect 172657 47891 172723 47894
rect 172565 47682 172631 47685
rect 136777 47680 140106 47682
rect 136777 47624 136782 47680
rect 136838 47624 140106 47680
rect 136777 47622 140106 47624
rect 169670 47680 172631 47682
rect 169670 47624 172570 47680
rect 172626 47624 172631 47680
rect 169670 47622 172631 47624
rect 136777 47619 136843 47622
rect 66397 47546 66463 47549
rect 100621 47546 100687 47549
rect 66397 47544 67948 47546
rect 66397 47488 66402 47544
rect 66458 47488 67948 47544
rect 66397 47486 67948 47488
rect 97756 47544 100687 47546
rect 97756 47488 100626 47544
rect 100682 47488 100687 47544
rect 97756 47486 100687 47488
rect 66397 47483 66463 47486
rect 100621 47483 100687 47486
rect 102553 47546 102619 47549
rect 134753 47546 134819 47549
rect 102553 47544 104932 47546
rect 102553 47488 102558 47544
rect 102614 47488 104932 47544
rect 102553 47486 104932 47488
rect 132716 47544 134819 47546
rect 132716 47488 134758 47544
rect 134814 47488 134819 47544
rect 132716 47486 134819 47488
rect 102553 47483 102619 47486
rect 134753 47483 134819 47486
rect 136869 47546 136935 47549
rect 136869 47544 140076 47546
rect 136869 47488 136874 47544
rect 136930 47488 140076 47544
rect 169670 47516 169730 47622
rect 172565 47619 172631 47622
rect 173945 47546 174011 47549
rect 173945 47544 177060 47546
rect 136869 47486 140076 47488
rect 173945 47488 173950 47544
rect 174006 47488 177060 47544
rect 173945 47486 177060 47488
rect 136869 47483 136935 47486
rect 173945 47483 174011 47486
rect 62901 47274 62967 47277
rect 60772 47272 62967 47274
rect 60772 47216 62906 47272
rect 62962 47216 62967 47272
rect 60772 47214 62967 47216
rect 62901 47211 62967 47214
rect 66397 47002 66463 47005
rect 102645 47002 102711 47005
rect 135305 47002 135371 47005
rect 66397 47000 67948 47002
rect 66397 46944 66402 47000
rect 66458 46944 67948 47000
rect 66397 46942 67948 46944
rect 102645 47000 104932 47002
rect 102645 46944 102650 47000
rect 102706 46944 104932 47000
rect 102645 46942 104932 46944
rect 132716 47000 135371 47002
rect 132716 46944 135310 47000
rect 135366 46944 135371 47000
rect 174037 47002 174103 47005
rect 174037 47000 177060 47002
rect 132716 46942 135371 46944
rect 66397 46939 66463 46942
rect 102645 46939 102711 46942
rect 135305 46939 135371 46942
rect 62717 46730 62783 46733
rect 60772 46728 62783 46730
rect 60772 46672 62722 46728
rect 62778 46672 62783 46728
rect 60772 46670 62783 46672
rect 62717 46667 62783 46670
rect 97726 46458 97786 46904
rect 100621 46458 100687 46461
rect 97726 46456 100687 46458
rect 97726 46400 100626 46456
rect 100682 46400 100687 46456
rect 97726 46398 100687 46400
rect 100621 46395 100687 46398
rect 102369 46458 102435 46461
rect 134845 46458 134911 46461
rect 102369 46456 104932 46458
rect 102369 46400 102374 46456
rect 102430 46400 104932 46456
rect 102369 46398 104932 46400
rect 132716 46456 134911 46458
rect 132716 46400 134850 46456
rect 134906 46400 134911 46456
rect 132716 46398 134911 46400
rect 102369 46395 102435 46398
rect 134845 46395 134911 46398
rect 136777 46458 136843 46461
rect 140046 46458 140106 46904
rect 136777 46456 140106 46458
rect 136777 46400 136782 46456
rect 136838 46400 140106 46456
rect 136777 46398 140106 46400
rect 169854 46458 169914 46972
rect 174037 46944 174042 47000
rect 174098 46944 177060 47000
rect 174037 46942 177060 46944
rect 174037 46939 174103 46942
rect 172657 46458 172723 46461
rect 169854 46456 172723 46458
rect 169854 46400 172662 46456
rect 172718 46400 172723 46456
rect 169854 46398 172723 46400
rect 136777 46395 136843 46398
rect 172657 46395 172723 46398
rect 174221 46458 174287 46461
rect 174221 46456 177060 46458
rect 174221 46400 174226 46456
rect 174282 46400 177060 46456
rect 174221 46398 177060 46400
rect 174221 46395 174287 46398
rect 65293 46322 65359 46325
rect 65293 46320 67948 46322
rect 65293 46264 65298 46320
rect 65354 46264 67948 46320
rect 65293 46262 67948 46264
rect 65293 46259 65359 46262
rect 62901 46186 62967 46189
rect 60772 46184 62967 46186
rect 60772 46128 62906 46184
rect 62962 46128 62967 46184
rect 60772 46126 62967 46128
rect 97726 46186 97786 46224
rect 100897 46186 100963 46189
rect 97726 46184 100963 46186
rect 97726 46128 100902 46184
rect 100958 46128 100963 46184
rect 97726 46126 100963 46128
rect 62901 46123 62967 46126
rect 100897 46123 100963 46126
rect 137513 46186 137579 46189
rect 140046 46186 140106 46224
rect 137513 46184 140106 46186
rect 137513 46128 137518 46184
rect 137574 46128 140106 46184
rect 137513 46126 140106 46128
rect 169854 46186 169914 46292
rect 172657 46186 172723 46189
rect 169854 46184 172723 46186
rect 169854 46128 172662 46184
rect 172718 46128 172723 46184
rect 169854 46126 172723 46128
rect 137513 46123 137579 46126
rect 172657 46123 172723 46126
rect 102461 45914 102527 45917
rect 135397 45914 135463 45917
rect 102461 45912 104932 45914
rect 102461 45856 102466 45912
rect 102522 45856 104932 45912
rect 102461 45854 104932 45856
rect 132716 45912 135463 45914
rect 132716 45856 135402 45912
rect 135458 45856 135463 45912
rect 132716 45854 135463 45856
rect 102461 45851 102527 45854
rect 135397 45851 135463 45854
rect 173853 45914 173919 45917
rect 173853 45912 177060 45914
rect 173853 45856 173858 45912
rect 173914 45856 177060 45912
rect 173853 45854 177060 45856
rect 173853 45851 173919 45854
rect 66397 45778 66463 45781
rect 66397 45776 67948 45778
rect 66397 45720 66402 45776
rect 66458 45720 67948 45776
rect 66397 45718 67948 45720
rect 66397 45715 66463 45718
rect 62809 45642 62875 45645
rect 60772 45640 62875 45642
rect 60772 45584 62814 45640
rect 62870 45584 62875 45640
rect 60772 45582 62875 45584
rect 62809 45579 62875 45582
rect 97726 45370 97786 45680
rect 100529 45370 100595 45373
rect 97726 45368 100595 45370
rect 97726 45312 100534 45368
rect 100590 45312 100595 45368
rect 97726 45310 100595 45312
rect 100529 45307 100595 45310
rect 136685 45370 136751 45373
rect 140046 45370 140106 45680
rect 136685 45368 140106 45370
rect 136685 45312 136690 45368
rect 136746 45312 140106 45368
rect 136685 45310 140106 45312
rect 169854 45370 169914 45748
rect 171829 45370 171895 45373
rect 169854 45368 171895 45370
rect 169854 45312 171834 45368
rect 171890 45312 171895 45368
rect 169854 45310 171895 45312
rect 136685 45307 136751 45310
rect 171829 45307 171895 45310
rect 65661 45234 65727 45237
rect 102553 45234 102619 45237
rect 134661 45234 134727 45237
rect 65661 45232 67948 45234
rect 65661 45176 65666 45232
rect 65722 45176 67948 45232
rect 65661 45174 67948 45176
rect 102553 45232 104932 45234
rect 102553 45176 102558 45232
rect 102614 45176 104932 45232
rect 102553 45174 104932 45176
rect 132716 45232 134727 45234
rect 132716 45176 134666 45232
rect 134722 45176 134727 45232
rect 174037 45234 174103 45237
rect 174037 45232 177060 45234
rect 132716 45174 134727 45176
rect 65661 45171 65727 45174
rect 102553 45171 102619 45174
rect 134661 45171 134727 45174
rect 97726 45098 97786 45136
rect 99977 45098 100043 45101
rect 97726 45096 100043 45098
rect 97726 45040 99982 45096
rect 100038 45040 100043 45096
rect 97726 45038 100043 45040
rect 99977 45035 100043 45038
rect 63729 44962 63795 44965
rect 60772 44960 63795 44962
rect 60772 44904 63734 44960
rect 63790 44904 63795 44960
rect 60772 44902 63795 44904
rect 63729 44899 63795 44902
rect 136777 44962 136843 44965
rect 140046 44962 140106 45136
rect 136777 44960 140106 44962
rect 136777 44904 136782 44960
rect 136838 44904 140106 44960
rect 136777 44902 140106 44904
rect 169854 44962 169914 45204
rect 174037 45176 174042 45232
rect 174098 45176 177060 45232
rect 174037 45174 177060 45176
rect 174037 45171 174103 45174
rect 172657 44962 172723 44965
rect 169854 44960 172723 44962
rect 169854 44904 172662 44960
rect 172718 44904 172723 44960
rect 169854 44902 172723 44904
rect 136777 44899 136843 44902
rect 172657 44899 172723 44902
rect 102369 44690 102435 44693
rect 135029 44690 135095 44693
rect 102369 44688 104932 44690
rect 102369 44632 102374 44688
rect 102430 44632 104932 44688
rect 102369 44630 104932 44632
rect 132716 44688 135095 44690
rect 132716 44632 135034 44688
rect 135090 44632 135095 44688
rect 132716 44630 135095 44632
rect 102369 44627 102435 44630
rect 135029 44627 135095 44630
rect 174129 44690 174195 44693
rect 174129 44688 177060 44690
rect 174129 44632 174134 44688
rect 174190 44632 177060 44688
rect 174129 44630 177060 44632
rect 174129 44627 174195 44630
rect 65293 44554 65359 44557
rect 222521 44554 222587 44557
rect 227416 44554 227896 44584
rect 65293 44552 67948 44554
rect 65293 44496 65298 44552
rect 65354 44496 67948 44552
rect 222521 44552 227896 44554
rect 65293 44494 67948 44496
rect 65293 44491 65359 44494
rect 62809 44418 62875 44421
rect 60772 44416 62875 44418
rect 60772 44360 62814 44416
rect 62870 44360 62875 44416
rect 60772 44358 62875 44360
rect 62809 44355 62875 44358
rect 31846 44220 31852 44284
rect 31916 44282 31922 44284
rect 31916 44222 32988 44282
rect 31916 44220 31922 44222
rect 97726 44146 97786 44456
rect 99885 44146 99951 44149
rect 97726 44144 99951 44146
rect 97726 44088 99890 44144
rect 99946 44088 99951 44144
rect 97726 44086 99951 44088
rect 99885 44083 99951 44086
rect 102461 44146 102527 44149
rect 135397 44146 135463 44149
rect 102461 44144 104932 44146
rect 102461 44088 102466 44144
rect 102522 44088 104932 44144
rect 102461 44086 104932 44088
rect 132716 44144 135463 44146
rect 132716 44088 135402 44144
rect 135458 44088 135463 44144
rect 132716 44086 135463 44088
rect 102461 44083 102527 44086
rect 135397 44083 135463 44086
rect 136777 44146 136843 44149
rect 140046 44146 140106 44456
rect 136777 44144 140106 44146
rect 136777 44088 136782 44144
rect 136838 44088 140106 44144
rect 136777 44086 140106 44088
rect 169854 44146 169914 44524
rect 222521 44496 222526 44552
rect 222582 44496 227896 44552
rect 222521 44494 227896 44496
rect 222521 44491 222587 44494
rect 227416 44464 227896 44494
rect 171829 44146 171895 44149
rect 169854 44144 171895 44146
rect 169854 44088 171834 44144
rect 171890 44088 171895 44144
rect 169854 44086 171895 44088
rect 136777 44083 136843 44086
rect 171829 44083 171895 44086
rect 174681 44146 174747 44149
rect 174681 44144 177060 44146
rect 174681 44088 174686 44144
rect 174742 44088 177060 44144
rect 174681 44086 177060 44088
rect 174681 44083 174747 44086
rect 66397 44010 66463 44013
rect 66397 44008 67948 44010
rect 66397 43952 66402 44008
rect 66458 43952 67948 44008
rect 66397 43950 67948 43952
rect 66397 43947 66463 43950
rect 63729 43874 63795 43877
rect 60772 43872 63795 43874
rect 60772 43816 63734 43872
rect 63790 43816 63795 43872
rect 60772 43814 63795 43816
rect 63729 43811 63795 43814
rect 97726 43466 97786 43912
rect 102553 43602 102619 43605
rect 135029 43602 135095 43605
rect 102553 43600 104932 43602
rect 102553 43544 102558 43600
rect 102614 43544 104932 43600
rect 102553 43542 104932 43544
rect 132716 43600 135095 43602
rect 132716 43544 135034 43600
rect 135090 43544 135095 43600
rect 132716 43542 135095 43544
rect 102553 43539 102619 43542
rect 135029 43539 135095 43542
rect 100621 43466 100687 43469
rect 97726 43464 100687 43466
rect 97726 43408 100626 43464
rect 100682 43408 100687 43464
rect 97726 43406 100687 43408
rect 100621 43403 100687 43406
rect 136869 43466 136935 43469
rect 140046 43466 140106 43912
rect 169854 43602 169914 43980
rect 172657 43602 172723 43605
rect 169854 43600 172723 43602
rect 169854 43544 172662 43600
rect 172718 43544 172723 43600
rect 169854 43542 172723 43544
rect 172657 43539 172723 43542
rect 174497 43602 174563 43605
rect 174497 43600 177060 43602
rect 174497 43544 174502 43600
rect 174558 43544 177060 43600
rect 174497 43542 177060 43544
rect 174497 43539 174563 43542
rect 136869 43464 140106 43466
rect 136869 43408 136874 43464
rect 136930 43408 140106 43464
rect 136869 43406 140106 43408
rect 136869 43403 136935 43406
rect 63637 43330 63703 43333
rect 60772 43328 63703 43330
rect 60772 43272 63642 43328
rect 63698 43272 63703 43328
rect 60772 43270 63703 43272
rect 63637 43267 63703 43270
rect 66397 43330 66463 43333
rect 66397 43328 67948 43330
rect 66397 43272 66402 43328
rect 66458 43272 67948 43328
rect 66397 43270 67948 43272
rect 66397 43267 66463 43270
rect 97726 42922 97786 43232
rect 102277 43058 102343 43061
rect 135397 43058 135463 43061
rect 102277 43056 104932 43058
rect 102277 43000 102282 43056
rect 102338 43000 104932 43056
rect 102277 42998 104932 43000
rect 132716 43056 135463 43058
rect 132716 43000 135402 43056
rect 135458 43000 135463 43056
rect 132716 42998 135463 43000
rect 102277 42995 102343 42998
rect 135397 42995 135463 42998
rect 100621 42922 100687 42925
rect 97726 42920 100687 42922
rect 97726 42864 100626 42920
rect 100682 42864 100687 42920
rect 97726 42862 100687 42864
rect 100621 42859 100687 42862
rect 136685 42922 136751 42925
rect 140046 42922 140106 43232
rect 136685 42920 140106 42922
rect 136685 42864 136690 42920
rect 136746 42864 140106 42920
rect 136685 42862 140106 42864
rect 169854 42922 169914 43300
rect 174037 43058 174103 43061
rect 174037 43056 177060 43058
rect 174037 43000 174042 43056
rect 174098 43000 177060 43056
rect 174037 42998 177060 43000
rect 174037 42995 174103 42998
rect 172565 42922 172631 42925
rect 169854 42920 172631 42922
rect 169854 42864 172570 42920
rect 172626 42864 172631 42920
rect 169854 42862 172631 42864
rect 136685 42859 136751 42862
rect 172565 42859 172631 42862
rect 63729 42786 63795 42789
rect 60772 42784 63795 42786
rect 60772 42728 63734 42784
rect 63790 42728 63795 42784
rect 60772 42726 63795 42728
rect 63729 42723 63795 42726
rect 66397 42786 66463 42789
rect 66397 42784 67948 42786
rect 66397 42728 66402 42784
rect 66458 42728 67948 42784
rect 66397 42726 67948 42728
rect 66397 42723 66463 42726
rect 97726 42378 97786 42688
rect 100621 42378 100687 42381
rect 97726 42376 100687 42378
rect 97726 42320 100626 42376
rect 100682 42320 100687 42376
rect 97726 42318 100687 42320
rect 100621 42315 100687 42318
rect 102369 42378 102435 42381
rect 134937 42378 135003 42381
rect 102369 42376 104932 42378
rect 102369 42320 102374 42376
rect 102430 42320 104932 42376
rect 102369 42318 104932 42320
rect 132716 42376 135003 42378
rect 132716 42320 134942 42376
rect 134998 42320 135003 42376
rect 132716 42318 135003 42320
rect 102369 42315 102435 42318
rect 134937 42315 135003 42318
rect 136869 42378 136935 42381
rect 140046 42378 140106 42688
rect 136869 42376 140106 42378
rect 136869 42320 136874 42376
rect 136930 42320 140106 42376
rect 136869 42318 140106 42320
rect 169854 42378 169914 42756
rect 172381 42378 172447 42381
rect 169854 42376 172447 42378
rect 169854 42320 172386 42376
rect 172442 42320 172447 42376
rect 169854 42318 172447 42320
rect 136869 42315 136935 42318
rect 172381 42315 172447 42318
rect 174221 42378 174287 42381
rect 174221 42376 177060 42378
rect 174221 42320 174226 42376
rect 174282 42320 177060 42376
rect 174221 42318 177060 42320
rect 174221 42315 174287 42318
rect 65293 42242 65359 42245
rect 65293 42240 67948 42242
rect 65293 42184 65298 42240
rect 65354 42184 67948 42240
rect 65293 42182 67948 42184
rect 65293 42179 65359 42182
rect 63913 42106 63979 42109
rect 60772 42104 63979 42106
rect 60772 42048 63918 42104
rect 63974 42048 63979 42104
rect 60772 42046 63979 42048
rect 97726 42106 97786 42144
rect 100621 42106 100687 42109
rect 97726 42104 100687 42106
rect 97726 42048 100626 42104
rect 100682 42048 100687 42104
rect 97726 42046 100687 42048
rect 63913 42043 63979 42046
rect 100621 42043 100687 42046
rect 136777 42106 136843 42109
rect 140046 42106 140106 42144
rect 136777 42104 140106 42106
rect 136777 42048 136782 42104
rect 136838 42048 140106 42104
rect 136777 42046 140106 42048
rect 169854 42106 169914 42212
rect 172657 42106 172723 42109
rect 169854 42104 172723 42106
rect 169854 42048 172662 42104
rect 172718 42048 172723 42104
rect 169854 42046 172723 42048
rect 136777 42043 136843 42046
rect 172657 42043 172723 42046
rect 102553 41834 102619 41837
rect 135305 41834 135371 41837
rect 102553 41832 104932 41834
rect 102553 41776 102558 41832
rect 102614 41776 104932 41832
rect 102553 41774 104932 41776
rect 132716 41832 135371 41834
rect 132716 41776 135310 41832
rect 135366 41776 135371 41832
rect 132716 41774 135371 41776
rect 102553 41771 102619 41774
rect 135305 41771 135371 41774
rect 174129 41834 174195 41837
rect 174129 41832 177060 41834
rect 174129 41776 174134 41832
rect 174190 41776 177060 41832
rect 174129 41774 177060 41776
rect 174129 41771 174195 41774
rect 63821 41562 63887 41565
rect 60772 41560 63887 41562
rect 60772 41504 63826 41560
rect 63882 41504 63887 41560
rect 60772 41502 63887 41504
rect 63821 41499 63887 41502
rect 9896 41290 10376 41320
rect 12025 41290 12091 41293
rect 9896 41288 12091 41290
rect 9896 41232 12030 41288
rect 12086 41232 12091 41288
rect 9896 41230 12091 41232
rect 9896 41200 10376 41230
rect 12025 41227 12091 41230
rect 102461 41290 102527 41293
rect 135397 41290 135463 41293
rect 102461 41288 104932 41290
rect 102461 41232 102466 41288
rect 102522 41232 104932 41288
rect 102461 41230 104932 41232
rect 132716 41288 135463 41290
rect 132716 41232 135402 41288
rect 135458 41232 135463 41288
rect 132716 41230 135463 41232
rect 102461 41227 102527 41230
rect 135397 41227 135463 41230
rect 173945 41290 174011 41293
rect 173945 41288 177060 41290
rect 173945 41232 173950 41288
rect 174006 41232 177060 41288
rect 173945 41230 177060 41232
rect 173945 41227 174011 41230
rect 63729 41018 63795 41021
rect 60772 41016 63795 41018
rect 60772 40960 63734 41016
rect 63790 40960 63795 41016
rect 60772 40958 63795 40960
rect 63729 40955 63795 40958
rect 102369 40746 102435 40749
rect 134845 40746 134911 40749
rect 102369 40744 104932 40746
rect 102369 40688 102374 40744
rect 102430 40688 104932 40744
rect 102369 40686 104932 40688
rect 132716 40744 134911 40746
rect 132716 40688 134850 40744
rect 134906 40688 134911 40744
rect 132716 40686 134911 40688
rect 102369 40683 102435 40686
rect 134845 40683 134911 40686
rect 174037 40746 174103 40749
rect 174037 40744 177060 40746
rect 174037 40688 174042 40744
rect 174098 40688 177060 40744
rect 174037 40686 177060 40688
rect 174037 40683 174103 40686
rect 62809 40474 62875 40477
rect 60772 40472 62875 40474
rect 60772 40416 62814 40472
rect 62870 40416 62875 40472
rect 60772 40414 62875 40416
rect 62809 40411 62875 40414
rect 66254 40412 66260 40476
rect 66324 40474 66330 40476
rect 66397 40474 66463 40477
rect 93854 40474 93860 40476
rect 66324 40472 93860 40474
rect 66324 40416 66402 40472
rect 66458 40416 93860 40472
rect 66324 40414 93860 40416
rect 66324 40412 66330 40414
rect 66397 40411 66463 40414
rect 93854 40412 93860 40414
rect 93924 40474 93930 40476
rect 93997 40474 94063 40477
rect 93924 40472 94063 40474
rect 93924 40416 94002 40472
rect 94058 40416 94063 40472
rect 93924 40414 94063 40416
rect 93924 40412 93930 40414
rect 93997 40411 94063 40414
rect 102369 40202 102435 40205
rect 102369 40200 104932 40202
rect 102369 40144 102374 40200
rect 102430 40144 104932 40200
rect 102369 40142 104932 40144
rect 102369 40139 102435 40142
rect 109637 40068 109703 40069
rect 109637 40066 109684 40068
rect 109592 40064 109684 40066
rect 109592 40008 109642 40064
rect 109592 40006 109684 40008
rect 109637 40004 109684 40006
rect 109748 40004 109754 40068
rect 109637 40003 109703 40004
rect 60742 39522 60802 39832
rect 132686 39658 132746 40104
rect 136910 39732 136916 39796
rect 136980 39794 136986 39796
rect 138157 39794 138223 39797
rect 166033 39794 166099 39797
rect 166166 39794 166172 39796
rect 136980 39792 166172 39794
rect 136980 39736 138162 39792
rect 138218 39736 166038 39792
rect 166094 39736 166172 39792
rect 136980 39734 166172 39736
rect 136980 39732 136986 39734
rect 138157 39731 138223 39734
rect 166033 39731 166099 39734
rect 166166 39732 166172 39734
rect 166236 39732 166242 39796
rect 134477 39658 134543 39661
rect 132686 39656 134543 39658
rect 132686 39600 134482 39656
rect 134538 39600 134543 39656
rect 132686 39598 134543 39600
rect 134477 39595 134543 39598
rect 62809 39522 62875 39525
rect 60742 39520 62875 39522
rect 60742 39464 62814 39520
rect 62870 39464 62875 39520
rect 60742 39462 62875 39464
rect 62809 39459 62875 39462
rect 174129 39522 174195 39525
rect 177030 39522 177090 40104
rect 181397 40068 181463 40069
rect 181397 40066 181444 40068
rect 181352 40064 181444 40066
rect 181352 40008 181402 40064
rect 181352 40006 181444 40008
rect 181397 40004 181444 40006
rect 181508 40004 181514 40068
rect 181397 40003 181463 40004
rect 174129 39520 177090 39522
rect 174129 39464 174134 39520
rect 174190 39464 177090 39520
rect 174129 39462 177090 39464
rect 174129 39459 174195 39462
rect 136869 33402 136935 33405
rect 136869 33400 140106 33402
rect 136869 33344 136874 33400
rect 136930 33344 140106 33400
rect 136869 33342 140106 33344
rect 136869 33339 136935 33342
rect 140046 32760 140106 33342
rect 66213 32722 66279 32725
rect 66213 32720 67948 32722
rect 66213 32664 66218 32720
rect 66274 32664 67948 32720
rect 66213 32662 67948 32664
rect 66213 32659 66279 32662
rect 138065 25106 138131 25109
rect 138065 25104 140106 25106
rect 138065 25048 138070 25104
rect 138126 25048 140106 25104
rect 138065 25046 140106 25048
rect 138065 25043 138131 25046
rect 140046 24736 140106 25046
rect 66305 24698 66371 24701
rect 66305 24696 67948 24698
rect 66305 24640 66310 24696
rect 66366 24640 67948 24696
rect 66305 24638 67948 24640
rect 66305 24635 66371 24638
rect 222705 20754 222771 20757
rect 227416 20754 227896 20784
rect 222705 20752 227896 20754
rect 222705 20696 222710 20752
rect 222766 20696 227896 20752
rect 222705 20694 227896 20696
rect 222705 20691 222771 20694
rect 227416 20664 227896 20694
rect 9896 19666 10376 19696
rect 13313 19666 13379 19669
rect 9896 19664 13379 19666
rect 9896 19608 13318 19664
rect 13374 19608 13379 19664
rect 9896 19606 13379 19608
rect 9896 19576 10376 19606
rect 13313 19603 13379 19606
rect 138157 17082 138223 17085
rect 138157 17080 140106 17082
rect 138157 17024 138162 17080
rect 138218 17024 140106 17080
rect 138157 17022 140106 17024
rect 138157 17019 138223 17022
rect 140046 16848 140106 17022
rect 66397 16810 66463 16813
rect 66397 16808 67948 16810
rect 66397 16752 66402 16808
rect 66458 16752 67948 16808
rect 66397 16750 67948 16752
rect 66397 16747 66463 16750
<< via3 >>
rect 20628 235164 20692 235228
rect 37924 217212 37988 217276
rect 204260 215852 204324 215916
rect 20812 213132 20876 213196
rect 204812 211636 204876 211700
rect 207572 192460 207636 192524
rect 207572 192324 207636 192388
rect 20076 183484 20140 183548
rect 20628 183484 20692 183548
rect 207204 182804 207268 182868
rect 20812 182532 20876 182596
rect 28724 182532 28788 182596
rect 207388 172876 207452 172940
rect 207572 172876 207636 172940
rect 207572 163220 207636 163284
rect 207388 153760 207452 153764
rect 207388 153704 207438 153760
rect 207438 153704 207452 153760
rect 207388 153700 207452 153704
rect 207388 153352 207452 153356
rect 207388 153296 207402 153352
rect 207402 153296 207452 153352
rect 207388 153292 207452 153296
rect 37924 151524 37988 151588
rect 176844 146492 176908 146556
rect 17132 146084 17196 146148
rect 20444 146084 20508 146148
rect 20444 142548 20508 142612
rect 101036 142548 101100 142612
rect 28724 142412 28788 142476
rect 101588 141868 101652 141932
rect 173348 141868 173412 141932
rect 31852 141384 31916 141388
rect 31852 141328 31902 141384
rect 31902 141328 31916 141384
rect 31852 141324 31916 141328
rect 102140 138332 102204 138396
rect 101772 134388 101836 134452
rect 101956 123508 102020 123572
rect 101772 123372 101836 123436
rect 101772 123168 101836 123232
rect 31852 118476 31916 118540
rect 101772 113776 101836 113780
rect 101772 113720 101822 113776
rect 101822 113720 101836 113776
rect 101772 113716 101836 113720
rect 56876 113232 56940 113236
rect 56876 113176 56926 113232
rect 56926 113176 56940 113232
rect 56876 113172 56940 113176
rect 71964 113232 72028 113236
rect 71964 113176 72014 113232
rect 72014 113176 72028 113232
rect 71964 113172 72028 113176
rect 129740 77540 129804 77604
rect 102508 73384 102572 73388
rect 102508 73328 102558 73384
rect 102558 73328 102572 73384
rect 102508 73324 102572 73328
rect 101404 71208 101468 71212
rect 101404 71152 101418 71208
rect 101418 71152 101468 71208
rect 101404 71148 101468 71152
rect 173348 71148 173412 71212
rect 100852 71012 100916 71076
rect 101220 70876 101284 70940
rect 201500 69380 201564 69444
rect 176844 69244 176908 69308
rect 31852 68760 31916 68764
rect 31852 68704 31902 68760
rect 31902 68704 31916 68760
rect 31852 68700 31916 68704
rect 31852 44220 31916 44284
rect 66260 40412 66324 40476
rect 93860 40412 93924 40476
rect 109684 40064 109748 40068
rect 109684 40008 109698 40064
rect 109698 40008 109748 40064
rect 109684 40004 109748 40008
rect 136916 39732 136980 39796
rect 166172 39732 166236 39796
rect 181444 40064 181508 40068
rect 181444 40008 181458 40064
rect 181458 40008 181508 40064
rect 181444 40004 181508 40008
<< metal4 >>
rect 0 255254 4000 255376
rect 0 255018 122 255254
rect 358 255018 442 255254
rect 678 255018 762 255254
rect 998 255018 1082 255254
rect 1318 255018 1402 255254
rect 1638 255018 1722 255254
rect 1958 255018 2042 255254
rect 2278 255018 2362 255254
rect 2598 255018 2682 255254
rect 2918 255018 3002 255254
rect 3238 255018 3322 255254
rect 3558 255018 3642 255254
rect 3878 255018 4000 255254
rect 0 254934 4000 255018
rect 0 254698 122 254934
rect 358 254698 442 254934
rect 678 254698 762 254934
rect 998 254698 1082 254934
rect 1318 254698 1402 254934
rect 1638 254698 1722 254934
rect 1958 254698 2042 254934
rect 2278 254698 2362 254934
rect 2598 254698 2682 254934
rect 2918 254698 3002 254934
rect 3238 254698 3322 254934
rect 3558 254698 3642 254934
rect 3878 254698 4000 254934
rect 0 254614 4000 254698
rect 0 254378 122 254614
rect 358 254378 442 254614
rect 678 254378 762 254614
rect 998 254378 1082 254614
rect 1318 254378 1402 254614
rect 1638 254378 1722 254614
rect 1958 254378 2042 254614
rect 2278 254378 2362 254614
rect 2598 254378 2682 254614
rect 2918 254378 3002 254614
rect 3238 254378 3322 254614
rect 3558 254378 3642 254614
rect 3878 254378 4000 254614
rect 0 254294 4000 254378
rect 0 254058 122 254294
rect 358 254058 442 254294
rect 678 254058 762 254294
rect 998 254058 1082 254294
rect 1318 254058 1402 254294
rect 1638 254058 1722 254294
rect 1958 254058 2042 254294
rect 2278 254058 2362 254294
rect 2598 254058 2682 254294
rect 2918 254058 3002 254294
rect 3238 254058 3322 254294
rect 3558 254058 3642 254294
rect 3878 254058 4000 254294
rect 0 253974 4000 254058
rect 0 253738 122 253974
rect 358 253738 442 253974
rect 678 253738 762 253974
rect 998 253738 1082 253974
rect 1318 253738 1402 253974
rect 1638 253738 1722 253974
rect 1958 253738 2042 253974
rect 2278 253738 2362 253974
rect 2598 253738 2682 253974
rect 2918 253738 3002 253974
rect 3238 253738 3322 253974
rect 3558 253738 3642 253974
rect 3878 253738 4000 253974
rect 0 253654 4000 253738
rect 0 253418 122 253654
rect 358 253418 442 253654
rect 678 253418 762 253654
rect 998 253418 1082 253654
rect 1318 253418 1402 253654
rect 1638 253418 1722 253654
rect 1958 253418 2042 253654
rect 2278 253418 2362 253654
rect 2598 253418 2682 253654
rect 2918 253418 3002 253654
rect 3238 253418 3322 253654
rect 3558 253418 3642 253654
rect 3878 253418 4000 253654
rect 0 253334 4000 253418
rect 0 253098 122 253334
rect 358 253098 442 253334
rect 678 253098 762 253334
rect 998 253098 1082 253334
rect 1318 253098 1402 253334
rect 1638 253098 1722 253334
rect 1958 253098 2042 253334
rect 2278 253098 2362 253334
rect 2598 253098 2682 253334
rect 2918 253098 3002 253334
rect 3238 253098 3322 253334
rect 3558 253098 3642 253334
rect 3878 253098 4000 253334
rect 0 253014 4000 253098
rect 0 252778 122 253014
rect 358 252778 442 253014
rect 678 252778 762 253014
rect 998 252778 1082 253014
rect 1318 252778 1402 253014
rect 1638 252778 1722 253014
rect 1958 252778 2042 253014
rect 2278 252778 2362 253014
rect 2598 252778 2682 253014
rect 2918 252778 3002 253014
rect 3238 252778 3322 253014
rect 3558 252778 3642 253014
rect 3878 252778 4000 253014
rect 0 252694 4000 252778
rect 0 252458 122 252694
rect 358 252458 442 252694
rect 678 252458 762 252694
rect 998 252458 1082 252694
rect 1318 252458 1402 252694
rect 1638 252458 1722 252694
rect 1958 252458 2042 252694
rect 2278 252458 2362 252694
rect 2598 252458 2682 252694
rect 2918 252458 3002 252694
rect 3238 252458 3322 252694
rect 3558 252458 3642 252694
rect 3878 252458 4000 252694
rect 0 252374 4000 252458
rect 0 252138 122 252374
rect 358 252138 442 252374
rect 678 252138 762 252374
rect 998 252138 1082 252374
rect 1318 252138 1402 252374
rect 1638 252138 1722 252374
rect 1958 252138 2042 252374
rect 2278 252138 2362 252374
rect 2598 252138 2682 252374
rect 2918 252138 3002 252374
rect 3238 252138 3322 252374
rect 3558 252138 3642 252374
rect 3878 252138 4000 252374
rect 0 252054 4000 252138
rect 0 251818 122 252054
rect 358 251818 442 252054
rect 678 251818 762 252054
rect 998 251818 1082 252054
rect 1318 251818 1402 252054
rect 1638 251818 1722 252054
rect 1958 251818 2042 252054
rect 2278 251818 2362 252054
rect 2598 251818 2682 252054
rect 2918 251818 3002 252054
rect 3238 251818 3322 252054
rect 3558 251818 3642 252054
rect 3878 251818 4000 252054
rect 0 251734 4000 251818
rect 0 251498 122 251734
rect 358 251498 442 251734
rect 678 251498 762 251734
rect 998 251498 1082 251734
rect 1318 251498 1402 251734
rect 1638 251498 1722 251734
rect 1958 251498 2042 251734
rect 2278 251498 2362 251734
rect 2598 251498 2682 251734
rect 2918 251498 3002 251734
rect 3238 251498 3322 251734
rect 3558 251498 3642 251734
rect 3878 251498 4000 251734
rect 0 228918 4000 251498
rect 233740 255254 237740 255376
rect 233740 255018 233862 255254
rect 234098 255018 234182 255254
rect 234418 255018 234502 255254
rect 234738 255018 234822 255254
rect 235058 255018 235142 255254
rect 235378 255018 235462 255254
rect 235698 255018 235782 255254
rect 236018 255018 236102 255254
rect 236338 255018 236422 255254
rect 236658 255018 236742 255254
rect 236978 255018 237062 255254
rect 237298 255018 237382 255254
rect 237618 255018 237740 255254
rect 233740 254934 237740 255018
rect 233740 254698 233862 254934
rect 234098 254698 234182 254934
rect 234418 254698 234502 254934
rect 234738 254698 234822 254934
rect 235058 254698 235142 254934
rect 235378 254698 235462 254934
rect 235698 254698 235782 254934
rect 236018 254698 236102 254934
rect 236338 254698 236422 254934
rect 236658 254698 236742 254934
rect 236978 254698 237062 254934
rect 237298 254698 237382 254934
rect 237618 254698 237740 254934
rect 233740 254614 237740 254698
rect 233740 254378 233862 254614
rect 234098 254378 234182 254614
rect 234418 254378 234502 254614
rect 234738 254378 234822 254614
rect 235058 254378 235142 254614
rect 235378 254378 235462 254614
rect 235698 254378 235782 254614
rect 236018 254378 236102 254614
rect 236338 254378 236422 254614
rect 236658 254378 236742 254614
rect 236978 254378 237062 254614
rect 237298 254378 237382 254614
rect 237618 254378 237740 254614
rect 233740 254294 237740 254378
rect 233740 254058 233862 254294
rect 234098 254058 234182 254294
rect 234418 254058 234502 254294
rect 234738 254058 234822 254294
rect 235058 254058 235142 254294
rect 235378 254058 235462 254294
rect 235698 254058 235782 254294
rect 236018 254058 236102 254294
rect 236338 254058 236422 254294
rect 236658 254058 236742 254294
rect 236978 254058 237062 254294
rect 237298 254058 237382 254294
rect 237618 254058 237740 254294
rect 233740 253974 237740 254058
rect 233740 253738 233862 253974
rect 234098 253738 234182 253974
rect 234418 253738 234502 253974
rect 234738 253738 234822 253974
rect 235058 253738 235142 253974
rect 235378 253738 235462 253974
rect 235698 253738 235782 253974
rect 236018 253738 236102 253974
rect 236338 253738 236422 253974
rect 236658 253738 236742 253974
rect 236978 253738 237062 253974
rect 237298 253738 237382 253974
rect 237618 253738 237740 253974
rect 233740 253654 237740 253738
rect 233740 253418 233862 253654
rect 234098 253418 234182 253654
rect 234418 253418 234502 253654
rect 234738 253418 234822 253654
rect 235058 253418 235142 253654
rect 235378 253418 235462 253654
rect 235698 253418 235782 253654
rect 236018 253418 236102 253654
rect 236338 253418 236422 253654
rect 236658 253418 236742 253654
rect 236978 253418 237062 253654
rect 237298 253418 237382 253654
rect 237618 253418 237740 253654
rect 233740 253334 237740 253418
rect 233740 253098 233862 253334
rect 234098 253098 234182 253334
rect 234418 253098 234502 253334
rect 234738 253098 234822 253334
rect 235058 253098 235142 253334
rect 235378 253098 235462 253334
rect 235698 253098 235782 253334
rect 236018 253098 236102 253334
rect 236338 253098 236422 253334
rect 236658 253098 236742 253334
rect 236978 253098 237062 253334
rect 237298 253098 237382 253334
rect 237618 253098 237740 253334
rect 233740 253014 237740 253098
rect 233740 252778 233862 253014
rect 234098 252778 234182 253014
rect 234418 252778 234502 253014
rect 234738 252778 234822 253014
rect 235058 252778 235142 253014
rect 235378 252778 235462 253014
rect 235698 252778 235782 253014
rect 236018 252778 236102 253014
rect 236338 252778 236422 253014
rect 236658 252778 236742 253014
rect 236978 252778 237062 253014
rect 237298 252778 237382 253014
rect 237618 252778 237740 253014
rect 233740 252694 237740 252778
rect 233740 252458 233862 252694
rect 234098 252458 234182 252694
rect 234418 252458 234502 252694
rect 234738 252458 234822 252694
rect 235058 252458 235142 252694
rect 235378 252458 235462 252694
rect 235698 252458 235782 252694
rect 236018 252458 236102 252694
rect 236338 252458 236422 252694
rect 236658 252458 236742 252694
rect 236978 252458 237062 252694
rect 237298 252458 237382 252694
rect 237618 252458 237740 252694
rect 233740 252374 237740 252458
rect 233740 252138 233862 252374
rect 234098 252138 234182 252374
rect 234418 252138 234502 252374
rect 234738 252138 234822 252374
rect 235058 252138 235142 252374
rect 235378 252138 235462 252374
rect 235698 252138 235782 252374
rect 236018 252138 236102 252374
rect 236338 252138 236422 252374
rect 236658 252138 236742 252374
rect 236978 252138 237062 252374
rect 237298 252138 237382 252374
rect 237618 252138 237740 252374
rect 233740 252054 237740 252138
rect 233740 251818 233862 252054
rect 234098 251818 234182 252054
rect 234418 251818 234502 252054
rect 234738 251818 234822 252054
rect 235058 251818 235142 252054
rect 235378 251818 235462 252054
rect 235698 251818 235782 252054
rect 236018 251818 236102 252054
rect 236338 251818 236422 252054
rect 236658 251818 236742 252054
rect 236978 251818 237062 252054
rect 237298 251818 237382 252054
rect 237618 251818 237740 252054
rect 233740 251734 237740 251818
rect 233740 251498 233862 251734
rect 234098 251498 234182 251734
rect 234418 251498 234502 251734
rect 234738 251498 234822 251734
rect 235058 251498 235142 251734
rect 235378 251498 235462 251734
rect 235698 251498 235782 251734
rect 236018 251498 236102 251734
rect 236338 251498 236422 251734
rect 236658 251498 236742 251734
rect 236978 251498 237062 251734
rect 237298 251498 237382 251734
rect 237618 251498 237740 251734
rect 0 228682 122 228918
rect 358 228682 442 228918
rect 678 228682 762 228918
rect 998 228682 1082 228918
rect 1318 228682 1402 228918
rect 1638 228682 1722 228918
rect 1958 228682 2042 228918
rect 2278 228682 2362 228918
rect 2598 228682 2682 228918
rect 2918 228682 3002 228918
rect 3238 228682 3322 228918
rect 3558 228682 3642 228918
rect 3878 228682 4000 228918
rect 0 206518 4000 228682
rect 0 206282 122 206518
rect 358 206282 442 206518
rect 678 206282 762 206518
rect 998 206282 1082 206518
rect 1318 206282 1402 206518
rect 1638 206282 1722 206518
rect 1958 206282 2042 206518
rect 2278 206282 2362 206518
rect 2598 206282 2682 206518
rect 2918 206282 3002 206518
rect 3238 206282 3322 206518
rect 3558 206282 3642 206518
rect 3878 206282 4000 206518
rect 0 184118 4000 206282
rect 0 183882 122 184118
rect 358 183882 442 184118
rect 678 183882 762 184118
rect 998 183882 1082 184118
rect 1318 183882 1402 184118
rect 1638 183882 1722 184118
rect 1958 183882 2042 184118
rect 2278 183882 2362 184118
rect 2598 183882 2682 184118
rect 2918 183882 3002 184118
rect 3238 183882 3322 184118
rect 3558 183882 3642 184118
rect 3878 183882 4000 184118
rect 0 161718 4000 183882
rect 0 161482 122 161718
rect 358 161482 442 161718
rect 678 161482 762 161718
rect 998 161482 1082 161718
rect 1318 161482 1402 161718
rect 1638 161482 1722 161718
rect 1958 161482 2042 161718
rect 2278 161482 2362 161718
rect 2598 161482 2682 161718
rect 2918 161482 3002 161718
rect 3238 161482 3322 161718
rect 3558 161482 3642 161718
rect 3878 161482 4000 161718
rect 0 139318 4000 161482
rect 0 139082 122 139318
rect 358 139082 442 139318
rect 678 139082 762 139318
rect 998 139082 1082 139318
rect 1318 139082 1402 139318
rect 1638 139082 1722 139318
rect 1958 139082 2042 139318
rect 2278 139082 2362 139318
rect 2598 139082 2682 139318
rect 2918 139082 3002 139318
rect 3238 139082 3322 139318
rect 3558 139082 3642 139318
rect 3878 139082 4000 139318
rect 0 116918 4000 139082
rect 0 116682 122 116918
rect 358 116682 442 116918
rect 678 116682 762 116918
rect 998 116682 1082 116918
rect 1318 116682 1402 116918
rect 1638 116682 1722 116918
rect 1958 116682 2042 116918
rect 2278 116682 2362 116918
rect 2598 116682 2682 116918
rect 2918 116682 3002 116918
rect 3238 116682 3322 116918
rect 3558 116682 3642 116918
rect 3878 116682 4000 116918
rect 0 94518 4000 116682
rect 0 94282 122 94518
rect 358 94282 442 94518
rect 678 94282 762 94518
rect 998 94282 1082 94518
rect 1318 94282 1402 94518
rect 1638 94282 1722 94518
rect 1958 94282 2042 94518
rect 2278 94282 2362 94518
rect 2598 94282 2682 94518
rect 2918 94282 3002 94518
rect 3238 94282 3322 94518
rect 3558 94282 3642 94518
rect 3878 94282 4000 94518
rect 0 72118 4000 94282
rect 0 71882 122 72118
rect 358 71882 442 72118
rect 678 71882 762 72118
rect 998 71882 1082 72118
rect 1318 71882 1402 72118
rect 1638 71882 1722 72118
rect 1958 71882 2042 72118
rect 2278 71882 2362 72118
rect 2598 71882 2682 72118
rect 2918 71882 3002 72118
rect 3238 71882 3322 72118
rect 3558 71882 3642 72118
rect 3878 71882 4000 72118
rect 0 49718 4000 71882
rect 0 49482 122 49718
rect 358 49482 442 49718
rect 678 49482 762 49718
rect 998 49482 1082 49718
rect 1318 49482 1402 49718
rect 1638 49482 1722 49718
rect 1958 49482 2042 49718
rect 2278 49482 2362 49718
rect 2598 49482 2682 49718
rect 2918 49482 3002 49718
rect 3238 49482 3322 49718
rect 3558 49482 3642 49718
rect 3878 49482 4000 49718
rect 0 27318 4000 49482
rect 0 27082 122 27318
rect 358 27082 442 27318
rect 678 27082 762 27318
rect 998 27082 1082 27318
rect 1318 27082 1402 27318
rect 1638 27082 1722 27318
rect 1958 27082 2042 27318
rect 2278 27082 2362 27318
rect 2598 27082 2682 27318
rect 2918 27082 3002 27318
rect 3238 27082 3322 27318
rect 3558 27082 3642 27318
rect 3878 27082 4000 27318
rect 0 3878 4000 27082
rect 5000 250254 9000 250376
rect 5000 250018 5122 250254
rect 5358 250018 5442 250254
rect 5678 250018 5762 250254
rect 5998 250018 6082 250254
rect 6318 250018 6402 250254
rect 6638 250018 6722 250254
rect 6958 250018 7042 250254
rect 7278 250018 7362 250254
rect 7598 250018 7682 250254
rect 7918 250018 8002 250254
rect 8238 250018 8322 250254
rect 8558 250018 8642 250254
rect 8878 250018 9000 250254
rect 5000 249934 9000 250018
rect 5000 249698 5122 249934
rect 5358 249698 5442 249934
rect 5678 249698 5762 249934
rect 5998 249698 6082 249934
rect 6318 249698 6402 249934
rect 6638 249698 6722 249934
rect 6958 249698 7042 249934
rect 7278 249698 7362 249934
rect 7598 249698 7682 249934
rect 7918 249698 8002 249934
rect 8238 249698 8322 249934
rect 8558 249698 8642 249934
rect 8878 249698 9000 249934
rect 5000 249614 9000 249698
rect 5000 249378 5122 249614
rect 5358 249378 5442 249614
rect 5678 249378 5762 249614
rect 5998 249378 6082 249614
rect 6318 249378 6402 249614
rect 6638 249378 6722 249614
rect 6958 249378 7042 249614
rect 7278 249378 7362 249614
rect 7598 249378 7682 249614
rect 7918 249378 8002 249614
rect 8238 249378 8322 249614
rect 8558 249378 8642 249614
rect 8878 249378 9000 249614
rect 5000 249294 9000 249378
rect 5000 249058 5122 249294
rect 5358 249058 5442 249294
rect 5678 249058 5762 249294
rect 5998 249058 6082 249294
rect 6318 249058 6402 249294
rect 6638 249058 6722 249294
rect 6958 249058 7042 249294
rect 7278 249058 7362 249294
rect 7598 249058 7682 249294
rect 7918 249058 8002 249294
rect 8238 249058 8322 249294
rect 8558 249058 8642 249294
rect 8878 249058 9000 249294
rect 5000 248974 9000 249058
rect 5000 248738 5122 248974
rect 5358 248738 5442 248974
rect 5678 248738 5762 248974
rect 5998 248738 6082 248974
rect 6318 248738 6402 248974
rect 6638 248738 6722 248974
rect 6958 248738 7042 248974
rect 7278 248738 7362 248974
rect 7598 248738 7682 248974
rect 7918 248738 8002 248974
rect 8238 248738 8322 248974
rect 8558 248738 8642 248974
rect 8878 248738 9000 248974
rect 5000 248654 9000 248738
rect 5000 248418 5122 248654
rect 5358 248418 5442 248654
rect 5678 248418 5762 248654
rect 5998 248418 6082 248654
rect 6318 248418 6402 248654
rect 6638 248418 6722 248654
rect 6958 248418 7042 248654
rect 7278 248418 7362 248654
rect 7598 248418 7682 248654
rect 7918 248418 8002 248654
rect 8238 248418 8322 248654
rect 8558 248418 8642 248654
rect 8878 248418 9000 248654
rect 5000 248334 9000 248418
rect 5000 248098 5122 248334
rect 5358 248098 5442 248334
rect 5678 248098 5762 248334
rect 5998 248098 6082 248334
rect 6318 248098 6402 248334
rect 6638 248098 6722 248334
rect 6958 248098 7042 248334
rect 7278 248098 7362 248334
rect 7598 248098 7682 248334
rect 7918 248098 8002 248334
rect 8238 248098 8322 248334
rect 8558 248098 8642 248334
rect 8878 248098 9000 248334
rect 5000 248014 9000 248098
rect 5000 247778 5122 248014
rect 5358 247778 5442 248014
rect 5678 247778 5762 248014
rect 5998 247778 6082 248014
rect 6318 247778 6402 248014
rect 6638 247778 6722 248014
rect 6958 247778 7042 248014
rect 7278 247778 7362 248014
rect 7598 247778 7682 248014
rect 7918 247778 8002 248014
rect 8238 247778 8322 248014
rect 8558 247778 8642 248014
rect 8878 247778 9000 248014
rect 5000 247694 9000 247778
rect 5000 247458 5122 247694
rect 5358 247458 5442 247694
rect 5678 247458 5762 247694
rect 5998 247458 6082 247694
rect 6318 247458 6402 247694
rect 6638 247458 6722 247694
rect 6958 247458 7042 247694
rect 7278 247458 7362 247694
rect 7598 247458 7682 247694
rect 7918 247458 8002 247694
rect 8238 247458 8322 247694
rect 8558 247458 8642 247694
rect 8878 247458 9000 247694
rect 5000 247374 9000 247458
rect 5000 247138 5122 247374
rect 5358 247138 5442 247374
rect 5678 247138 5762 247374
rect 5998 247138 6082 247374
rect 6318 247138 6402 247374
rect 6638 247138 6722 247374
rect 6958 247138 7042 247374
rect 7278 247138 7362 247374
rect 7598 247138 7682 247374
rect 7918 247138 8002 247374
rect 8238 247138 8322 247374
rect 8558 247138 8642 247374
rect 8878 247138 9000 247374
rect 5000 247054 9000 247138
rect 5000 246818 5122 247054
rect 5358 246818 5442 247054
rect 5678 246818 5762 247054
rect 5998 246818 6082 247054
rect 6318 246818 6402 247054
rect 6638 246818 6722 247054
rect 6958 246818 7042 247054
rect 7278 246818 7362 247054
rect 7598 246818 7682 247054
rect 7918 246818 8002 247054
rect 8238 246818 8322 247054
rect 8558 246818 8642 247054
rect 8878 246818 9000 247054
rect 5000 246734 9000 246818
rect 5000 246498 5122 246734
rect 5358 246498 5442 246734
rect 5678 246498 5762 246734
rect 5998 246498 6082 246734
rect 6318 246498 6402 246734
rect 6638 246498 6722 246734
rect 6958 246498 7042 246734
rect 7278 246498 7362 246734
rect 7598 246498 7682 246734
rect 7918 246498 8002 246734
rect 8238 246498 8322 246734
rect 8558 246498 8642 246734
rect 8878 246498 9000 246734
rect 5000 240118 9000 246498
rect 228740 250254 232740 250376
rect 228740 250018 228862 250254
rect 229098 250018 229182 250254
rect 229418 250018 229502 250254
rect 229738 250018 229822 250254
rect 230058 250018 230142 250254
rect 230378 250018 230462 250254
rect 230698 250018 230782 250254
rect 231018 250018 231102 250254
rect 231338 250018 231422 250254
rect 231658 250018 231742 250254
rect 231978 250018 232062 250254
rect 232298 250018 232382 250254
rect 232618 250018 232740 250254
rect 228740 249934 232740 250018
rect 228740 249698 228862 249934
rect 229098 249698 229182 249934
rect 229418 249698 229502 249934
rect 229738 249698 229822 249934
rect 230058 249698 230142 249934
rect 230378 249698 230462 249934
rect 230698 249698 230782 249934
rect 231018 249698 231102 249934
rect 231338 249698 231422 249934
rect 231658 249698 231742 249934
rect 231978 249698 232062 249934
rect 232298 249698 232382 249934
rect 232618 249698 232740 249934
rect 228740 249614 232740 249698
rect 228740 249378 228862 249614
rect 229098 249378 229182 249614
rect 229418 249378 229502 249614
rect 229738 249378 229822 249614
rect 230058 249378 230142 249614
rect 230378 249378 230462 249614
rect 230698 249378 230782 249614
rect 231018 249378 231102 249614
rect 231338 249378 231422 249614
rect 231658 249378 231742 249614
rect 231978 249378 232062 249614
rect 232298 249378 232382 249614
rect 232618 249378 232740 249614
rect 228740 249294 232740 249378
rect 228740 249058 228862 249294
rect 229098 249058 229182 249294
rect 229418 249058 229502 249294
rect 229738 249058 229822 249294
rect 230058 249058 230142 249294
rect 230378 249058 230462 249294
rect 230698 249058 230782 249294
rect 231018 249058 231102 249294
rect 231338 249058 231422 249294
rect 231658 249058 231742 249294
rect 231978 249058 232062 249294
rect 232298 249058 232382 249294
rect 232618 249058 232740 249294
rect 228740 248974 232740 249058
rect 228740 248738 228862 248974
rect 229098 248738 229182 248974
rect 229418 248738 229502 248974
rect 229738 248738 229822 248974
rect 230058 248738 230142 248974
rect 230378 248738 230462 248974
rect 230698 248738 230782 248974
rect 231018 248738 231102 248974
rect 231338 248738 231422 248974
rect 231658 248738 231742 248974
rect 231978 248738 232062 248974
rect 232298 248738 232382 248974
rect 232618 248738 232740 248974
rect 228740 248654 232740 248738
rect 228740 248418 228862 248654
rect 229098 248418 229182 248654
rect 229418 248418 229502 248654
rect 229738 248418 229822 248654
rect 230058 248418 230142 248654
rect 230378 248418 230462 248654
rect 230698 248418 230782 248654
rect 231018 248418 231102 248654
rect 231338 248418 231422 248654
rect 231658 248418 231742 248654
rect 231978 248418 232062 248654
rect 232298 248418 232382 248654
rect 232618 248418 232740 248654
rect 228740 248334 232740 248418
rect 228740 248098 228862 248334
rect 229098 248098 229182 248334
rect 229418 248098 229502 248334
rect 229738 248098 229822 248334
rect 230058 248098 230142 248334
rect 230378 248098 230462 248334
rect 230698 248098 230782 248334
rect 231018 248098 231102 248334
rect 231338 248098 231422 248334
rect 231658 248098 231742 248334
rect 231978 248098 232062 248334
rect 232298 248098 232382 248334
rect 232618 248098 232740 248334
rect 228740 248014 232740 248098
rect 228740 247778 228862 248014
rect 229098 247778 229182 248014
rect 229418 247778 229502 248014
rect 229738 247778 229822 248014
rect 230058 247778 230142 248014
rect 230378 247778 230462 248014
rect 230698 247778 230782 248014
rect 231018 247778 231102 248014
rect 231338 247778 231422 248014
rect 231658 247778 231742 248014
rect 231978 247778 232062 248014
rect 232298 247778 232382 248014
rect 232618 247778 232740 248014
rect 228740 247694 232740 247778
rect 228740 247458 228862 247694
rect 229098 247458 229182 247694
rect 229418 247458 229502 247694
rect 229738 247458 229822 247694
rect 230058 247458 230142 247694
rect 230378 247458 230462 247694
rect 230698 247458 230782 247694
rect 231018 247458 231102 247694
rect 231338 247458 231422 247694
rect 231658 247458 231742 247694
rect 231978 247458 232062 247694
rect 232298 247458 232382 247694
rect 232618 247458 232740 247694
rect 228740 247374 232740 247458
rect 228740 247138 228862 247374
rect 229098 247138 229182 247374
rect 229418 247138 229502 247374
rect 229738 247138 229822 247374
rect 230058 247138 230142 247374
rect 230378 247138 230462 247374
rect 230698 247138 230782 247374
rect 231018 247138 231102 247374
rect 231338 247138 231422 247374
rect 231658 247138 231742 247374
rect 231978 247138 232062 247374
rect 232298 247138 232382 247374
rect 232618 247138 232740 247374
rect 228740 247054 232740 247138
rect 228740 246818 228862 247054
rect 229098 246818 229182 247054
rect 229418 246818 229502 247054
rect 229738 246818 229822 247054
rect 230058 246818 230142 247054
rect 230378 246818 230462 247054
rect 230698 246818 230782 247054
rect 231018 246818 231102 247054
rect 231338 246818 231422 247054
rect 231658 246818 231742 247054
rect 231978 246818 232062 247054
rect 232298 246818 232382 247054
rect 232618 246818 232740 247054
rect 228740 246734 232740 246818
rect 228740 246498 228862 246734
rect 229098 246498 229182 246734
rect 229418 246498 229502 246734
rect 229738 246498 229822 246734
rect 230058 246498 230142 246734
rect 230378 246498 230462 246734
rect 230698 246498 230782 246734
rect 231018 246498 231102 246734
rect 231338 246498 231422 246734
rect 231658 246498 231742 246734
rect 231978 246498 232062 246734
rect 232298 246498 232382 246734
rect 232618 246498 232740 246734
rect 5000 239882 5122 240118
rect 5358 239882 5442 240118
rect 5678 239882 5762 240118
rect 5998 239882 6082 240118
rect 6318 239882 6402 240118
rect 6638 239882 6722 240118
rect 6958 239882 7042 240118
rect 7278 239882 7362 240118
rect 7598 239882 7682 240118
rect 7918 239882 8002 240118
rect 8238 239882 8322 240118
rect 8558 239882 8642 240118
rect 8878 239882 9000 240118
rect 5000 217718 9000 239882
rect 72774 240118 73094 240160
rect 72774 239882 72816 240118
rect 73052 239882 73094 240118
rect 72774 239840 73094 239882
rect 144774 240118 145094 240160
rect 144774 239882 144816 240118
rect 145052 239882 145094 240118
rect 144774 239840 145094 239882
rect 228740 240118 232740 246498
rect 228740 239882 228862 240118
rect 229098 239882 229182 240118
rect 229418 239882 229502 240118
rect 229738 239882 229822 240118
rect 230058 239882 230142 240118
rect 230378 239882 230462 240118
rect 230698 239882 230782 240118
rect 231018 239882 231102 240118
rect 231338 239882 231422 240118
rect 231658 239882 231742 240118
rect 231978 239882 232062 240118
rect 232298 239882 232382 240118
rect 232618 239882 232740 240118
rect 20627 235228 20693 235229
rect 20627 235164 20628 235228
rect 20692 235164 20693 235228
rect 20627 235163 20693 235164
rect 5000 217482 5122 217718
rect 5358 217482 5442 217718
rect 5678 217482 5762 217718
rect 5998 217482 6082 217718
rect 6318 217482 6402 217718
rect 6638 217482 6722 217718
rect 6958 217482 7042 217718
rect 7278 217482 7362 217718
rect 7598 217482 7682 217718
rect 7918 217482 8002 217718
rect 8238 217482 8322 217718
rect 8558 217482 8642 217718
rect 8878 217482 9000 217718
rect 5000 195318 9000 217482
rect 5000 195082 5122 195318
rect 5358 195082 5442 195318
rect 5678 195082 5762 195318
rect 5998 195082 6082 195318
rect 6318 195082 6402 195318
rect 6638 195082 6722 195318
rect 6958 195082 7042 195318
rect 7278 195082 7362 195318
rect 7598 195082 7682 195318
rect 7918 195082 8002 195318
rect 8238 195082 8322 195318
rect 8558 195082 8642 195318
rect 8878 195082 9000 195318
rect 5000 172918 9000 195082
rect 20630 183549 20690 235163
rect 77774 228918 78094 228960
rect 77774 228682 77816 228918
rect 78052 228682 78094 228918
rect 77774 228640 78094 228682
rect 149774 228918 150094 228960
rect 149774 228682 149816 228918
rect 150052 228682 150094 228918
rect 149774 228640 150094 228682
rect 228740 217718 232740 239882
rect 228740 217482 228862 217718
rect 229098 217482 229182 217718
rect 229418 217482 229502 217718
rect 229738 217482 229822 217718
rect 230058 217482 230142 217718
rect 230378 217482 230462 217718
rect 230698 217482 230782 217718
rect 231018 217482 231102 217718
rect 231338 217482 231422 217718
rect 231658 217482 231742 217718
rect 231978 217482 232062 217718
rect 232298 217482 232382 217718
rect 232618 217482 232740 217718
rect 37923 217276 37989 217277
rect 37923 217212 37924 217276
rect 37988 217212 37989 217276
rect 37923 217211 37989 217212
rect 20811 213196 20877 213197
rect 20811 213132 20812 213196
rect 20876 213132 20877 213196
rect 20811 213131 20877 213132
rect 20075 183548 20141 183549
rect 20075 183484 20076 183548
rect 20140 183484 20141 183548
rect 20075 183483 20141 183484
rect 20627 183548 20693 183549
rect 20627 183484 20628 183548
rect 20692 183484 20693 183548
rect 20627 183483 20693 183484
rect 20078 183362 20138 183483
rect 20814 182597 20874 213131
rect 20811 182596 20877 182597
rect 20811 182532 20812 182596
rect 20876 182532 20877 182596
rect 20811 182531 20877 182532
rect 28723 182596 28789 182597
rect 28723 182532 28724 182596
rect 28788 182532 28789 182596
rect 28723 182531 28789 182532
rect 5000 172682 5122 172918
rect 5358 172682 5442 172918
rect 5678 172682 5762 172918
rect 5998 172682 6082 172918
rect 6318 172682 6402 172918
rect 6638 172682 6722 172918
rect 6958 172682 7042 172918
rect 7278 172682 7362 172918
rect 7598 172682 7682 172918
rect 7918 172682 8002 172918
rect 8238 172682 8322 172918
rect 8558 172682 8642 172918
rect 8878 172682 9000 172918
rect 5000 150518 9000 172682
rect 16398 166274 16458 173606
rect 17134 166362 17194 175646
rect 28726 173842 28786 182531
rect 17507 172918 17827 172960
rect 17507 172682 17549 172918
rect 17785 172682 17827 172918
rect 17507 172640 17827 172682
rect 16398 166214 16826 166274
rect 16766 156074 16826 166214
rect 20173 161718 20493 161760
rect 20173 161482 20215 161718
rect 20451 161482 20493 161718
rect 20173 161440 20493 161482
rect 16582 156014 16826 156074
rect 16582 152082 16642 156014
rect 28726 154122 28786 162726
rect 5000 150282 5122 150518
rect 5358 150282 5442 150518
rect 5678 150282 5762 150518
rect 5998 150282 6082 150518
rect 6318 150282 6402 150518
rect 6638 150282 6722 150518
rect 6958 150282 7042 150518
rect 7278 150282 7362 150518
rect 7598 150282 7682 150518
rect 7918 150282 8002 150518
rect 8238 150282 8322 150518
rect 8558 150282 8642 150518
rect 8878 150282 9000 150518
rect 5000 128118 9000 150282
rect 17134 146149 17194 153886
rect 17507 150518 17827 150560
rect 17507 150282 17549 150518
rect 17785 150282 17827 150518
rect 17507 150240 17827 150282
rect 17131 146148 17197 146149
rect 17131 146084 17132 146148
rect 17196 146084 17197 146148
rect 17131 146083 17197 146084
rect 20443 146148 20509 146149
rect 20443 146084 20444 146148
rect 20508 146084 20509 146148
rect 20443 146083 20509 146084
rect 20446 142613 20506 146083
rect 20443 142612 20509 142613
rect 20443 142548 20444 142612
rect 20508 142548 20509 142612
rect 20443 142547 20509 142548
rect 28726 142477 28786 153206
rect 37926 151589 37986 217211
rect 204259 215916 204325 215917
rect 204259 215852 204260 215916
rect 204324 215852 204325 215916
rect 204259 215851 204325 215852
rect 204262 211834 204322 215851
rect 204262 211774 204874 211834
rect 204814 211701 204874 211774
rect 204811 211700 204877 211701
rect 204811 211636 204812 211700
rect 204876 211636 204877 211700
rect 204811 211635 204877 211636
rect 42885 206518 43205 206560
rect 42885 206282 42927 206518
rect 43163 206282 43205 206518
rect 42885 206240 43205 206282
rect 78840 206518 79160 206560
rect 78840 206282 78882 206518
rect 79118 206282 79160 206518
rect 78840 206240 79160 206282
rect 150840 206518 151160 206560
rect 150840 206282 150882 206518
rect 151118 206282 151160 206518
rect 150840 206240 151160 206282
rect 187173 206518 187493 206560
rect 187173 206282 187215 206518
rect 187451 206282 187493 206518
rect 187173 206240 187493 206282
rect 38219 195318 38539 195360
rect 38219 195082 38261 195318
rect 38497 195082 38539 195318
rect 38219 195040 38539 195082
rect 73840 195318 74160 195360
rect 73840 195082 73882 195318
rect 74118 195082 74160 195318
rect 73840 195040 74160 195082
rect 145840 195318 146160 195360
rect 145840 195082 145882 195318
rect 146118 195082 146160 195318
rect 145840 195040 146160 195082
rect 182507 195318 182827 195360
rect 182507 195082 182549 195318
rect 182785 195082 182827 195318
rect 182507 195040 182827 195082
rect 228740 195318 232740 217482
rect 228740 195082 228862 195318
rect 229098 195082 229182 195318
rect 229418 195082 229502 195318
rect 229738 195082 229822 195318
rect 230058 195082 230142 195318
rect 230378 195082 230462 195318
rect 230698 195082 230782 195318
rect 231018 195082 231102 195318
rect 231338 195082 231422 195318
rect 231658 195082 231742 195318
rect 231978 195082 232062 195318
rect 232298 195082 232382 195318
rect 232618 195082 232740 195318
rect 207571 192524 207637 192525
rect 207571 192460 207572 192524
rect 207636 192460 207637 192524
rect 207571 192459 207637 192460
rect 207574 192389 207634 192459
rect 207571 192388 207637 192389
rect 207571 192324 207572 192388
rect 207636 192324 207637 192388
rect 207571 192323 207637 192324
rect 207203 182868 207269 182869
rect 207203 182804 207204 182868
rect 207268 182804 207269 182868
rect 207203 182803 207269 182804
rect 207206 175794 207266 182803
rect 207206 175734 207450 175794
rect 42507 172918 42827 172960
rect 42507 172682 42549 172918
rect 42785 172682 42827 172918
rect 42507 172640 42827 172682
rect 67104 172918 67424 172960
rect 67104 172682 67146 172918
rect 67382 172682 67424 172918
rect 67104 172640 67424 172682
rect 114507 172918 114827 172960
rect 114507 172682 114549 172918
rect 114785 172682 114827 172918
rect 114507 172640 114827 172682
rect 139104 172918 139424 172960
rect 139104 172682 139146 172918
rect 139382 172682 139424 172918
rect 139104 172640 139424 172682
rect 186507 172918 186827 172960
rect 207390 172941 207450 175734
rect 186507 172682 186549 172918
rect 186785 172682 186827 172918
rect 207387 172940 207453 172941
rect 207387 172876 207388 172940
rect 207452 172876 207453 172940
rect 207387 172875 207453 172876
rect 207571 172940 207637 172941
rect 207571 172876 207572 172940
rect 207636 172876 207637 172940
rect 207571 172875 207637 172876
rect 211507 172918 211827 172960
rect 186507 172640 186827 172682
rect 207574 163285 207634 172875
rect 211507 172682 211549 172918
rect 211785 172682 211827 172918
rect 211507 172640 211827 172682
rect 228740 172918 232740 195082
rect 228740 172682 228862 172918
rect 229098 172682 229182 172918
rect 229418 172682 229502 172918
rect 229738 172682 229822 172918
rect 230058 172682 230142 172918
rect 230378 172682 230462 172918
rect 230698 172682 230782 172918
rect 231018 172682 231102 172918
rect 231338 172682 231422 172918
rect 231658 172682 231742 172918
rect 231978 172682 232062 172918
rect 232298 172682 232382 172918
rect 232618 172682 232740 172918
rect 207571 163284 207637 163285
rect 207571 163220 207572 163284
rect 207636 163220 207637 163284
rect 207571 163219 207637 163220
rect 45173 161718 45493 161760
rect 45173 161482 45215 161718
rect 45451 161482 45493 161718
rect 45173 161440 45493 161482
rect 82464 161718 82784 161760
rect 82464 161482 82506 161718
rect 82742 161482 82784 161718
rect 82464 161440 82784 161482
rect 117173 161718 117493 161760
rect 117173 161482 117215 161718
rect 117451 161482 117493 161718
rect 117173 161440 117493 161482
rect 154464 161718 154784 161760
rect 154464 161482 154506 161718
rect 154742 161482 154784 161718
rect 154464 161440 154784 161482
rect 189173 161718 189493 161760
rect 189173 161482 189215 161718
rect 189451 161482 189493 161718
rect 189173 161440 189493 161482
rect 214173 161718 214493 161760
rect 214173 161482 214215 161718
rect 214451 161482 214493 161718
rect 214173 161440 214493 161482
rect 207387 153764 207453 153765
rect 207387 153700 207388 153764
rect 207452 153700 207453 153764
rect 207387 153699 207453 153700
rect 207390 153357 207450 153699
rect 207387 153356 207453 153357
rect 207387 153292 207388 153356
rect 207452 153292 207453 153356
rect 207387 153291 207453 153292
rect 37923 151588 37989 151589
rect 37923 151524 37924 151588
rect 37988 151524 37989 151588
rect 37923 151523 37989 151524
rect 42507 150518 42827 150560
rect 42507 150282 42549 150518
rect 42785 150282 42827 150518
rect 42507 150240 42827 150282
rect 67104 150518 67424 150560
rect 67104 150282 67146 150518
rect 67382 150282 67424 150518
rect 67104 150240 67424 150282
rect 114507 150518 114827 150560
rect 114507 150282 114549 150518
rect 114785 150282 114827 150518
rect 114507 150240 114827 150282
rect 139104 150518 139424 150560
rect 139104 150282 139146 150518
rect 139382 150282 139424 150518
rect 139104 150240 139424 150282
rect 186507 150518 186827 150560
rect 186507 150282 186549 150518
rect 186785 150282 186827 150518
rect 186507 150240 186827 150282
rect 211507 150518 211827 150560
rect 211507 150282 211549 150518
rect 211785 150282 211827 150518
rect 211507 150240 211827 150282
rect 228740 150518 232740 172682
rect 228740 150282 228862 150518
rect 229098 150282 229182 150518
rect 229418 150282 229502 150518
rect 229738 150282 229822 150518
rect 230058 150282 230142 150518
rect 230378 150282 230462 150518
rect 230698 150282 230782 150518
rect 231018 150282 231102 150518
rect 231338 150282 231422 150518
rect 231658 150282 231742 150518
rect 231978 150282 232062 150518
rect 232298 150282 232382 150518
rect 232618 150282 232740 150518
rect 176843 146556 176909 146557
rect 176843 146492 176844 146556
rect 176908 146492 176909 146556
rect 176843 146491 176909 146492
rect 101035 142612 101101 142613
rect 101035 142548 101036 142612
rect 101100 142548 101101 142612
rect 101035 142547 101101 142548
rect 28723 142476 28789 142477
rect 28723 142412 28724 142476
rect 28788 142412 28789 142476
rect 28723 142411 28789 142412
rect 31851 141388 31917 141389
rect 31851 141324 31852 141388
rect 31916 141324 31917 141388
rect 31851 141323 31917 141324
rect 5000 127882 5122 128118
rect 5358 127882 5442 128118
rect 5678 127882 5762 128118
rect 5998 127882 6082 128118
rect 6318 127882 6402 128118
rect 6638 127882 6722 128118
rect 6958 127882 7042 128118
rect 7278 127882 7362 128118
rect 7598 127882 7682 128118
rect 7918 127882 8002 128118
rect 8238 127882 8322 128118
rect 8558 127882 8642 128118
rect 8878 127882 9000 128118
rect 5000 105718 9000 127882
rect 31854 118541 31914 141323
rect 43173 139318 43493 139360
rect 43173 139082 43215 139318
rect 43451 139082 43493 139318
rect 43173 139040 43493 139082
rect 38507 128118 38827 128160
rect 38507 127882 38549 128118
rect 38785 127882 38827 128118
rect 38507 127840 38827 127882
rect 73840 128118 74160 128160
rect 73840 127882 73882 128118
rect 74118 127882 74160 128118
rect 73840 127840 74160 127882
rect 31851 118540 31917 118541
rect 31851 118476 31852 118540
rect 31916 118476 31917 118540
rect 31851 118475 31917 118476
rect 31854 114002 31914 118475
rect 43173 116918 43493 116960
rect 43173 116682 43215 116918
rect 43451 116682 43493 116918
rect 43173 116640 43493 116682
rect 56878 113237 56938 113766
rect 56875 113236 56941 113237
rect 56875 113172 56876 113236
rect 56940 113172 56941 113236
rect 56875 113171 56941 113172
rect 5000 105482 5122 105718
rect 5358 105482 5442 105718
rect 5678 105482 5762 105718
rect 5998 105482 6082 105718
rect 6318 105482 6402 105718
rect 6638 105482 6722 105718
rect 6958 105482 7042 105718
rect 7278 105482 7362 105718
rect 7598 105482 7682 105718
rect 7918 105482 8002 105718
rect 8238 105482 8322 105718
rect 8558 105482 8642 105718
rect 8878 105482 9000 105718
rect 5000 83318 9000 105482
rect 17507 105718 17827 105760
rect 17507 105482 17549 105718
rect 17785 105482 17827 105718
rect 17507 105440 17827 105482
rect 42507 105718 42827 105760
rect 42507 105482 42549 105718
rect 42785 105482 42827 105718
rect 42507 105440 42827 105482
rect 67104 105718 67424 105760
rect 67104 105482 67146 105718
rect 67382 105482 67424 105718
rect 67104 105440 67424 105482
rect 20173 94518 20493 94560
rect 20173 94282 20215 94518
rect 20451 94282 20493 94518
rect 20173 94240 20493 94282
rect 45173 94518 45493 94560
rect 45173 94282 45215 94518
rect 45451 94282 45493 94518
rect 45173 94240 45493 94282
rect 82464 94518 82784 94560
rect 82464 94282 82506 94518
rect 82742 94282 82784 94518
rect 82464 94240 82784 94282
rect 5000 83082 5122 83318
rect 5358 83082 5442 83318
rect 5678 83082 5762 83318
rect 5998 83082 6082 83318
rect 6318 83082 6402 83318
rect 6638 83082 6722 83318
rect 6958 83082 7042 83318
rect 7278 83082 7362 83318
rect 7598 83082 7682 83318
rect 7918 83082 8002 83318
rect 8238 83082 8322 83318
rect 8558 83082 8642 83318
rect 8878 83082 9000 83318
rect 5000 60918 9000 83082
rect 17507 83318 17827 83360
rect 17507 83082 17549 83318
rect 17785 83082 17827 83318
rect 17507 83040 17827 83082
rect 42507 83318 42827 83360
rect 42507 83082 42549 83318
rect 42785 83082 42827 83318
rect 42507 83040 42827 83082
rect 67104 83318 67424 83360
rect 67104 83082 67146 83318
rect 67382 83082 67424 83318
rect 67104 83040 67424 83082
rect 101038 78554 101098 142547
rect 101587 141932 101653 141933
rect 101587 141868 101588 141932
rect 101652 141868 101653 141932
rect 101587 141867 101653 141868
rect 173347 141932 173413 141933
rect 173347 141868 173348 141932
rect 173412 141868 173413 141932
rect 173347 141867 173413 141868
rect 100854 78494 101098 78554
rect 100854 71077 100914 78494
rect 101590 75834 101650 141867
rect 115173 139318 115493 139360
rect 115173 139082 115215 139318
rect 115451 139082 115493 139318
rect 115173 139040 115493 139082
rect 102139 138396 102205 138397
rect 102139 138332 102140 138396
rect 102204 138332 102205 138396
rect 102139 138331 102205 138332
rect 101771 134452 101837 134453
rect 101771 134388 101772 134452
rect 101836 134388 101837 134452
rect 101771 134387 101837 134388
rect 101774 132954 101834 134387
rect 101774 132894 102018 132954
rect 101958 123573 102018 132894
rect 101955 123572 102021 123573
rect 101955 123508 101956 123572
rect 102020 123508 102021 123572
rect 101955 123507 102021 123508
rect 101771 123436 101837 123437
rect 101771 123372 101772 123436
rect 101836 123372 101837 123436
rect 101771 123371 101837 123372
rect 101774 123233 101834 123371
rect 101771 123232 101837 123233
rect 101771 123168 101772 123232
rect 101836 123168 101837 123232
rect 101771 123167 101837 123168
rect 101771 113780 101837 113781
rect 101771 113716 101772 113780
rect 101836 113716 101837 113780
rect 101771 113715 101837 113716
rect 101774 107794 101834 113715
rect 101774 107734 102018 107794
rect 101958 94194 102018 107734
rect 101222 75774 101650 75834
rect 101774 94134 102018 94194
rect 100851 71076 100917 71077
rect 100851 71012 100852 71076
rect 100916 71012 100917 71076
rect 100851 71011 100917 71012
rect 101222 70941 101282 75774
rect 101774 74474 101834 94134
rect 101406 74414 101834 74474
rect 101406 71213 101466 74414
rect 102142 73794 102202 138331
rect 110507 128118 110827 128160
rect 110507 127882 110549 128118
rect 110785 127882 110827 128118
rect 110507 127840 110827 127882
rect 145840 128118 146160 128160
rect 145840 127882 145882 128118
rect 146118 127882 146160 128118
rect 145840 127840 146160 127882
rect 115173 116918 115493 116960
rect 115173 116682 115215 116918
rect 115451 116682 115493 116918
rect 115173 116640 115493 116682
rect 114507 105718 114827 105760
rect 114507 105482 114549 105718
rect 114785 105482 114827 105718
rect 114507 105440 114827 105482
rect 139104 105718 139424 105760
rect 139104 105482 139146 105718
rect 139382 105482 139424 105718
rect 139104 105440 139424 105482
rect 117173 94518 117493 94560
rect 117173 94282 117215 94518
rect 117451 94282 117493 94518
rect 117173 94240 117493 94282
rect 154464 94518 154784 94560
rect 154464 94282 154506 94518
rect 154742 94282 154784 94518
rect 154464 94240 154784 94282
rect 114507 83318 114827 83360
rect 114507 83082 114549 83318
rect 114785 83082 114827 83318
rect 114507 83040 114827 83082
rect 139104 83318 139424 83360
rect 139104 83082 139146 83318
rect 139382 83082 139424 83318
rect 139104 83040 139424 83082
rect 129739 77604 129805 77605
rect 129739 77540 129740 77604
rect 129804 77540 129805 77604
rect 129739 77539 129805 77540
rect 102142 73734 102570 73794
rect 102510 73389 102570 73734
rect 102507 73388 102573 73389
rect 102507 73324 102508 73388
rect 102572 73324 102573 73388
rect 102507 73323 102573 73324
rect 101403 71212 101469 71213
rect 101403 71148 101404 71212
rect 101468 71148 101469 71212
rect 101403 71147 101469 71148
rect 101219 70940 101285 70941
rect 101219 70876 101220 70940
rect 101284 70876 101285 70940
rect 101219 70875 101285 70876
rect 31851 68764 31917 68765
rect 31851 68700 31852 68764
rect 31916 68700 31917 68764
rect 31851 68699 31917 68700
rect 5000 60682 5122 60918
rect 5358 60682 5442 60918
rect 5678 60682 5762 60918
rect 5998 60682 6082 60918
rect 6318 60682 6402 60918
rect 6638 60682 6722 60918
rect 6958 60682 7042 60918
rect 7278 60682 7362 60918
rect 7598 60682 7682 60918
rect 7918 60682 8002 60918
rect 8238 60682 8322 60918
rect 8558 60682 8642 60918
rect 8878 60682 9000 60918
rect 5000 38518 9000 60682
rect 31854 44285 31914 68699
rect 38507 60918 38827 60960
rect 38507 60682 38549 60918
rect 38785 60682 38827 60918
rect 38507 60640 38827 60682
rect 73840 60918 74160 60960
rect 73840 60682 73882 60918
rect 74118 60682 74160 60918
rect 73840 60640 74160 60682
rect 110507 60918 110827 60960
rect 110507 60682 110549 60918
rect 110785 60682 110827 60918
rect 110507 60640 110827 60682
rect 43173 49718 43493 49760
rect 43173 49482 43215 49718
rect 43451 49482 43493 49718
rect 43173 49440 43493 49482
rect 78840 49718 79160 49760
rect 78840 49482 78882 49718
rect 79118 49482 79160 49718
rect 78840 49440 79160 49482
rect 115173 49718 115493 49760
rect 115173 49482 115215 49718
rect 115451 49482 115493 49718
rect 115173 49440 115493 49482
rect 31851 44284 31917 44285
rect 31851 44220 31852 44284
rect 31916 44220 31917 44284
rect 31851 44219 31917 44220
rect 31854 41242 31914 44219
rect 66262 40477 66322 41006
rect 129742 40562 129802 77539
rect 173350 71213 173410 141867
rect 173347 71212 173413 71213
rect 173347 71148 173348 71212
rect 173412 71148 173413 71212
rect 173347 71147 173413 71148
rect 176846 69309 176906 146491
rect 187173 139318 187493 139360
rect 187173 139082 187215 139318
rect 187451 139082 187493 139318
rect 187173 139040 187493 139082
rect 182507 128118 182827 128160
rect 182507 127882 182549 128118
rect 182785 127882 182827 128118
rect 182507 127840 182827 127882
rect 228740 128118 232740 150282
rect 228740 127882 228862 128118
rect 229098 127882 229182 128118
rect 229418 127882 229502 128118
rect 229738 127882 229822 128118
rect 230058 127882 230142 128118
rect 230378 127882 230462 128118
rect 230698 127882 230782 128118
rect 231018 127882 231102 128118
rect 231338 127882 231422 128118
rect 231658 127882 231742 128118
rect 231978 127882 232062 128118
rect 232298 127882 232382 128118
rect 232618 127882 232740 128118
rect 187173 116918 187493 116960
rect 187173 116682 187215 116918
rect 187451 116682 187493 116918
rect 187173 116640 187493 116682
rect 186507 105718 186827 105760
rect 186507 105482 186549 105718
rect 186785 105482 186827 105718
rect 186507 105440 186827 105482
rect 211507 105718 211827 105760
rect 211507 105482 211549 105718
rect 211785 105482 211827 105718
rect 211507 105440 211827 105482
rect 228740 105718 232740 127882
rect 228740 105482 228862 105718
rect 229098 105482 229182 105718
rect 229418 105482 229502 105718
rect 229738 105482 229822 105718
rect 230058 105482 230142 105718
rect 230378 105482 230462 105718
rect 230698 105482 230782 105718
rect 231018 105482 231102 105718
rect 231338 105482 231422 105718
rect 231658 105482 231742 105718
rect 231978 105482 232062 105718
rect 232298 105482 232382 105718
rect 232618 105482 232740 105718
rect 189173 94518 189493 94560
rect 189173 94282 189215 94518
rect 189451 94282 189493 94518
rect 189173 94240 189493 94282
rect 214173 94518 214493 94560
rect 214173 94282 214215 94518
rect 214451 94282 214493 94518
rect 214173 94240 214493 94282
rect 186507 83318 186827 83360
rect 186507 83082 186549 83318
rect 186785 83082 186827 83318
rect 186507 83040 186827 83082
rect 211507 83318 211827 83360
rect 211507 83082 211549 83318
rect 211785 83082 211827 83318
rect 211507 83040 211827 83082
rect 228740 83318 232740 105482
rect 228740 83082 228862 83318
rect 229098 83082 229182 83318
rect 229418 83082 229502 83318
rect 229738 83082 229822 83318
rect 230058 83082 230142 83318
rect 230378 83082 230462 83318
rect 230698 83082 230782 83318
rect 231018 83082 231102 83318
rect 231338 83082 231422 83318
rect 231658 83082 231742 83318
rect 231978 83082 232062 83318
rect 232298 83082 232382 83318
rect 232618 83082 232740 83318
rect 201499 69444 201565 69445
rect 201499 69380 201500 69444
rect 201564 69380 201565 69444
rect 201499 69379 201565 69380
rect 176843 69308 176909 69309
rect 176843 69244 176844 69308
rect 176908 69244 176909 69308
rect 176843 69243 176909 69244
rect 201502 65634 201562 69379
rect 201502 65574 201746 65634
rect 145840 60918 146160 60960
rect 145840 60682 145882 60918
rect 146118 60682 146160 60918
rect 145840 60640 146160 60682
rect 182507 60918 182827 60960
rect 182507 60682 182549 60918
rect 182785 60682 182827 60918
rect 182507 60640 182827 60682
rect 150840 49718 151160 49760
rect 150840 49482 150882 49718
rect 151118 49482 151160 49718
rect 150840 49440 151160 49482
rect 187173 49718 187493 49760
rect 187173 49482 187215 49718
rect 187451 49482 187493 49718
rect 187173 49440 187493 49482
rect 201686 41834 201746 65574
rect 201502 41774 201746 41834
rect 228740 60918 232740 83082
rect 228740 60682 228862 60918
rect 229098 60682 229182 60918
rect 229418 60682 229502 60918
rect 229738 60682 229822 60918
rect 230058 60682 230142 60918
rect 230378 60682 230462 60918
rect 230698 60682 230782 60918
rect 231018 60682 231102 60918
rect 231338 60682 231422 60918
rect 231658 60682 231742 60918
rect 231978 60682 232062 60918
rect 232298 60682 232382 60918
rect 232618 60682 232740 60918
rect 66259 40476 66325 40477
rect 66259 40412 66260 40476
rect 66324 40412 66325 40476
rect 66259 40411 66325 40412
rect 108914 40414 109598 40474
rect 109686 40069 109746 40326
rect 109683 40068 109749 40069
rect 109683 40004 109684 40068
rect 109748 40004 109749 40068
rect 109683 40003 109749 40004
rect 136918 39797 136978 40326
rect 181446 40069 181506 40326
rect 181443 40068 181509 40069
rect 181443 40004 181444 40068
rect 181508 40004 181509 40068
rect 181443 40003 181509 40004
rect 136915 39796 136981 39797
rect 136915 39732 136916 39796
rect 136980 39732 136981 39796
rect 136915 39731 136981 39732
rect 201502 39202 201562 41774
rect 5000 38282 5122 38518
rect 5358 38282 5442 38518
rect 5678 38282 5762 38518
rect 5998 38282 6082 38518
rect 6318 38282 6402 38518
rect 6638 38282 6722 38518
rect 6958 38282 7042 38518
rect 7278 38282 7362 38518
rect 7598 38282 7682 38518
rect 7918 38282 8002 38518
rect 8238 38282 8322 38518
rect 8558 38282 8642 38518
rect 8878 38282 9000 38518
rect 5000 16118 9000 38282
rect 228740 38518 232740 60682
rect 228740 38282 228862 38518
rect 229098 38282 229182 38518
rect 229418 38282 229502 38518
rect 229738 38282 229822 38518
rect 230058 38282 230142 38518
rect 230378 38282 230462 38518
rect 230698 38282 230782 38518
rect 231018 38282 231102 38518
rect 231338 38282 231422 38518
rect 231658 38282 231742 38518
rect 231978 38282 232062 38518
rect 232298 38282 232382 38518
rect 232618 38282 232740 38518
rect 78840 27318 79160 27360
rect 78840 27082 78882 27318
rect 79118 27082 79160 27318
rect 78840 27040 79160 27082
rect 150840 27318 151160 27360
rect 150840 27082 150882 27318
rect 151118 27082 151160 27318
rect 150840 27040 151160 27082
rect 5000 15882 5122 16118
rect 5358 15882 5442 16118
rect 5678 15882 5762 16118
rect 5998 15882 6082 16118
rect 6318 15882 6402 16118
rect 6638 15882 6722 16118
rect 6958 15882 7042 16118
rect 7278 15882 7362 16118
rect 7598 15882 7682 16118
rect 7918 15882 8002 16118
rect 8238 15882 8322 16118
rect 8558 15882 8642 16118
rect 8878 15882 9000 16118
rect 5000 8878 9000 15882
rect 73840 16118 74160 16160
rect 73840 15882 73882 16118
rect 74118 15882 74160 16118
rect 73840 15840 74160 15882
rect 145840 16118 146160 16160
rect 145840 15882 145882 16118
rect 146118 15882 146160 16118
rect 145840 15840 146160 15882
rect 228740 16118 232740 38282
rect 228740 15882 228862 16118
rect 229098 15882 229182 16118
rect 229418 15882 229502 16118
rect 229738 15882 229822 16118
rect 230058 15882 230142 16118
rect 230378 15882 230462 16118
rect 230698 15882 230782 16118
rect 231018 15882 231102 16118
rect 231338 15882 231422 16118
rect 231658 15882 231742 16118
rect 231978 15882 232062 16118
rect 232298 15882 232382 16118
rect 232618 15882 232740 16118
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 9000 8878
rect 5000 8558 9000 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 9000 8558
rect 5000 8238 9000 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 9000 8238
rect 5000 7918 9000 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 9000 7918
rect 5000 7598 9000 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 9000 7598
rect 5000 7278 9000 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 9000 7278
rect 5000 6958 9000 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 9000 6958
rect 5000 6638 9000 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 9000 6638
rect 5000 6318 9000 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 9000 6318
rect 5000 5998 9000 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 9000 5998
rect 5000 5678 9000 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 9000 5678
rect 5000 5358 9000 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 9000 5358
rect 5000 5000 9000 5122
rect 228740 8878 232740 15882
rect 228740 8642 228862 8878
rect 229098 8642 229182 8878
rect 229418 8642 229502 8878
rect 229738 8642 229822 8878
rect 230058 8642 230142 8878
rect 230378 8642 230462 8878
rect 230698 8642 230782 8878
rect 231018 8642 231102 8878
rect 231338 8642 231422 8878
rect 231658 8642 231742 8878
rect 231978 8642 232062 8878
rect 232298 8642 232382 8878
rect 232618 8642 232740 8878
rect 228740 8558 232740 8642
rect 228740 8322 228862 8558
rect 229098 8322 229182 8558
rect 229418 8322 229502 8558
rect 229738 8322 229822 8558
rect 230058 8322 230142 8558
rect 230378 8322 230462 8558
rect 230698 8322 230782 8558
rect 231018 8322 231102 8558
rect 231338 8322 231422 8558
rect 231658 8322 231742 8558
rect 231978 8322 232062 8558
rect 232298 8322 232382 8558
rect 232618 8322 232740 8558
rect 228740 8238 232740 8322
rect 228740 8002 228862 8238
rect 229098 8002 229182 8238
rect 229418 8002 229502 8238
rect 229738 8002 229822 8238
rect 230058 8002 230142 8238
rect 230378 8002 230462 8238
rect 230698 8002 230782 8238
rect 231018 8002 231102 8238
rect 231338 8002 231422 8238
rect 231658 8002 231742 8238
rect 231978 8002 232062 8238
rect 232298 8002 232382 8238
rect 232618 8002 232740 8238
rect 228740 7918 232740 8002
rect 228740 7682 228862 7918
rect 229098 7682 229182 7918
rect 229418 7682 229502 7918
rect 229738 7682 229822 7918
rect 230058 7682 230142 7918
rect 230378 7682 230462 7918
rect 230698 7682 230782 7918
rect 231018 7682 231102 7918
rect 231338 7682 231422 7918
rect 231658 7682 231742 7918
rect 231978 7682 232062 7918
rect 232298 7682 232382 7918
rect 232618 7682 232740 7918
rect 228740 7598 232740 7682
rect 228740 7362 228862 7598
rect 229098 7362 229182 7598
rect 229418 7362 229502 7598
rect 229738 7362 229822 7598
rect 230058 7362 230142 7598
rect 230378 7362 230462 7598
rect 230698 7362 230782 7598
rect 231018 7362 231102 7598
rect 231338 7362 231422 7598
rect 231658 7362 231742 7598
rect 231978 7362 232062 7598
rect 232298 7362 232382 7598
rect 232618 7362 232740 7598
rect 228740 7278 232740 7362
rect 228740 7042 228862 7278
rect 229098 7042 229182 7278
rect 229418 7042 229502 7278
rect 229738 7042 229822 7278
rect 230058 7042 230142 7278
rect 230378 7042 230462 7278
rect 230698 7042 230782 7278
rect 231018 7042 231102 7278
rect 231338 7042 231422 7278
rect 231658 7042 231742 7278
rect 231978 7042 232062 7278
rect 232298 7042 232382 7278
rect 232618 7042 232740 7278
rect 228740 6958 232740 7042
rect 228740 6722 228862 6958
rect 229098 6722 229182 6958
rect 229418 6722 229502 6958
rect 229738 6722 229822 6958
rect 230058 6722 230142 6958
rect 230378 6722 230462 6958
rect 230698 6722 230782 6958
rect 231018 6722 231102 6958
rect 231338 6722 231422 6958
rect 231658 6722 231742 6958
rect 231978 6722 232062 6958
rect 232298 6722 232382 6958
rect 232618 6722 232740 6958
rect 228740 6638 232740 6722
rect 228740 6402 228862 6638
rect 229098 6402 229182 6638
rect 229418 6402 229502 6638
rect 229738 6402 229822 6638
rect 230058 6402 230142 6638
rect 230378 6402 230462 6638
rect 230698 6402 230782 6638
rect 231018 6402 231102 6638
rect 231338 6402 231422 6638
rect 231658 6402 231742 6638
rect 231978 6402 232062 6638
rect 232298 6402 232382 6638
rect 232618 6402 232740 6638
rect 228740 6318 232740 6402
rect 228740 6082 228862 6318
rect 229098 6082 229182 6318
rect 229418 6082 229502 6318
rect 229738 6082 229822 6318
rect 230058 6082 230142 6318
rect 230378 6082 230462 6318
rect 230698 6082 230782 6318
rect 231018 6082 231102 6318
rect 231338 6082 231422 6318
rect 231658 6082 231742 6318
rect 231978 6082 232062 6318
rect 232298 6082 232382 6318
rect 232618 6082 232740 6318
rect 228740 5998 232740 6082
rect 228740 5762 228862 5998
rect 229098 5762 229182 5998
rect 229418 5762 229502 5998
rect 229738 5762 229822 5998
rect 230058 5762 230142 5998
rect 230378 5762 230462 5998
rect 230698 5762 230782 5998
rect 231018 5762 231102 5998
rect 231338 5762 231422 5998
rect 231658 5762 231742 5998
rect 231978 5762 232062 5998
rect 232298 5762 232382 5998
rect 232618 5762 232740 5998
rect 228740 5678 232740 5762
rect 228740 5442 228862 5678
rect 229098 5442 229182 5678
rect 229418 5442 229502 5678
rect 229738 5442 229822 5678
rect 230058 5442 230142 5678
rect 230378 5442 230462 5678
rect 230698 5442 230782 5678
rect 231018 5442 231102 5678
rect 231338 5442 231422 5678
rect 231658 5442 231742 5678
rect 231978 5442 232062 5678
rect 232298 5442 232382 5678
rect 232618 5442 232740 5678
rect 228740 5358 232740 5442
rect 228740 5122 228862 5358
rect 229098 5122 229182 5358
rect 229418 5122 229502 5358
rect 229738 5122 229822 5358
rect 230058 5122 230142 5358
rect 230378 5122 230462 5358
rect 230698 5122 230782 5358
rect 231018 5122 231102 5358
rect 231338 5122 231422 5358
rect 231658 5122 231742 5358
rect 231978 5122 232062 5358
rect 232298 5122 232382 5358
rect 232618 5122 232740 5358
rect 228740 5000 232740 5122
rect 233740 228918 237740 251498
rect 233740 228682 233862 228918
rect 234098 228682 234182 228918
rect 234418 228682 234502 228918
rect 234738 228682 234822 228918
rect 235058 228682 235142 228918
rect 235378 228682 235462 228918
rect 235698 228682 235782 228918
rect 236018 228682 236102 228918
rect 236338 228682 236422 228918
rect 236658 228682 236742 228918
rect 236978 228682 237062 228918
rect 237298 228682 237382 228918
rect 237618 228682 237740 228918
rect 233740 206518 237740 228682
rect 233740 206282 233862 206518
rect 234098 206282 234182 206518
rect 234418 206282 234502 206518
rect 234738 206282 234822 206518
rect 235058 206282 235142 206518
rect 235378 206282 235462 206518
rect 235698 206282 235782 206518
rect 236018 206282 236102 206518
rect 236338 206282 236422 206518
rect 236658 206282 236742 206518
rect 236978 206282 237062 206518
rect 237298 206282 237382 206518
rect 237618 206282 237740 206518
rect 233740 184118 237740 206282
rect 233740 183882 233862 184118
rect 234098 183882 234182 184118
rect 234418 183882 234502 184118
rect 234738 183882 234822 184118
rect 235058 183882 235142 184118
rect 235378 183882 235462 184118
rect 235698 183882 235782 184118
rect 236018 183882 236102 184118
rect 236338 183882 236422 184118
rect 236658 183882 236742 184118
rect 236978 183882 237062 184118
rect 237298 183882 237382 184118
rect 237618 183882 237740 184118
rect 233740 161718 237740 183882
rect 233740 161482 233862 161718
rect 234098 161482 234182 161718
rect 234418 161482 234502 161718
rect 234738 161482 234822 161718
rect 235058 161482 235142 161718
rect 235378 161482 235462 161718
rect 235698 161482 235782 161718
rect 236018 161482 236102 161718
rect 236338 161482 236422 161718
rect 236658 161482 236742 161718
rect 236978 161482 237062 161718
rect 237298 161482 237382 161718
rect 237618 161482 237740 161718
rect 233740 139318 237740 161482
rect 233740 139082 233862 139318
rect 234098 139082 234182 139318
rect 234418 139082 234502 139318
rect 234738 139082 234822 139318
rect 235058 139082 235142 139318
rect 235378 139082 235462 139318
rect 235698 139082 235782 139318
rect 236018 139082 236102 139318
rect 236338 139082 236422 139318
rect 236658 139082 236742 139318
rect 236978 139082 237062 139318
rect 237298 139082 237382 139318
rect 237618 139082 237740 139318
rect 233740 116918 237740 139082
rect 233740 116682 233862 116918
rect 234098 116682 234182 116918
rect 234418 116682 234502 116918
rect 234738 116682 234822 116918
rect 235058 116682 235142 116918
rect 235378 116682 235462 116918
rect 235698 116682 235782 116918
rect 236018 116682 236102 116918
rect 236338 116682 236422 116918
rect 236658 116682 236742 116918
rect 236978 116682 237062 116918
rect 237298 116682 237382 116918
rect 237618 116682 237740 116918
rect 233740 94518 237740 116682
rect 233740 94282 233862 94518
rect 234098 94282 234182 94518
rect 234418 94282 234502 94518
rect 234738 94282 234822 94518
rect 235058 94282 235142 94518
rect 235378 94282 235462 94518
rect 235698 94282 235782 94518
rect 236018 94282 236102 94518
rect 236338 94282 236422 94518
rect 236658 94282 236742 94518
rect 236978 94282 237062 94518
rect 237298 94282 237382 94518
rect 237618 94282 237740 94518
rect 233740 72118 237740 94282
rect 233740 71882 233862 72118
rect 234098 71882 234182 72118
rect 234418 71882 234502 72118
rect 234738 71882 234822 72118
rect 235058 71882 235142 72118
rect 235378 71882 235462 72118
rect 235698 71882 235782 72118
rect 236018 71882 236102 72118
rect 236338 71882 236422 72118
rect 236658 71882 236742 72118
rect 236978 71882 237062 72118
rect 237298 71882 237382 72118
rect 237618 71882 237740 72118
rect 233740 49718 237740 71882
rect 233740 49482 233862 49718
rect 234098 49482 234182 49718
rect 234418 49482 234502 49718
rect 234738 49482 234822 49718
rect 235058 49482 235142 49718
rect 235378 49482 235462 49718
rect 235698 49482 235782 49718
rect 236018 49482 236102 49718
rect 236338 49482 236422 49718
rect 236658 49482 236742 49718
rect 236978 49482 237062 49718
rect 237298 49482 237382 49718
rect 237618 49482 237740 49718
rect 233740 27318 237740 49482
rect 233740 27082 233862 27318
rect 234098 27082 234182 27318
rect 234418 27082 234502 27318
rect 234738 27082 234822 27318
rect 235058 27082 235142 27318
rect 235378 27082 235462 27318
rect 235698 27082 235782 27318
rect 236018 27082 236102 27318
rect 236338 27082 236422 27318
rect 236658 27082 236742 27318
rect 236978 27082 237062 27318
rect 237298 27082 237382 27318
rect 237618 27082 237740 27318
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 4000 3878
rect 0 3558 4000 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 4000 3558
rect 0 3238 4000 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 4000 3238
rect 0 2918 4000 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 4000 2918
rect 0 2598 4000 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 4000 2598
rect 0 2278 4000 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 4000 2278
rect 0 1958 4000 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 4000 1958
rect 0 1638 4000 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 4000 1638
rect 0 1318 4000 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 4000 1318
rect 0 998 4000 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 4000 998
rect 0 678 4000 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 4000 678
rect 0 358 4000 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 4000 358
rect 0 0 4000 122
rect 233740 3878 237740 27082
rect 233740 3642 233862 3878
rect 234098 3642 234182 3878
rect 234418 3642 234502 3878
rect 234738 3642 234822 3878
rect 235058 3642 235142 3878
rect 235378 3642 235462 3878
rect 235698 3642 235782 3878
rect 236018 3642 236102 3878
rect 236338 3642 236422 3878
rect 236658 3642 236742 3878
rect 236978 3642 237062 3878
rect 237298 3642 237382 3878
rect 237618 3642 237740 3878
rect 233740 3558 237740 3642
rect 233740 3322 233862 3558
rect 234098 3322 234182 3558
rect 234418 3322 234502 3558
rect 234738 3322 234822 3558
rect 235058 3322 235142 3558
rect 235378 3322 235462 3558
rect 235698 3322 235782 3558
rect 236018 3322 236102 3558
rect 236338 3322 236422 3558
rect 236658 3322 236742 3558
rect 236978 3322 237062 3558
rect 237298 3322 237382 3558
rect 237618 3322 237740 3558
rect 233740 3238 237740 3322
rect 233740 3002 233862 3238
rect 234098 3002 234182 3238
rect 234418 3002 234502 3238
rect 234738 3002 234822 3238
rect 235058 3002 235142 3238
rect 235378 3002 235462 3238
rect 235698 3002 235782 3238
rect 236018 3002 236102 3238
rect 236338 3002 236422 3238
rect 236658 3002 236742 3238
rect 236978 3002 237062 3238
rect 237298 3002 237382 3238
rect 237618 3002 237740 3238
rect 233740 2918 237740 3002
rect 233740 2682 233862 2918
rect 234098 2682 234182 2918
rect 234418 2682 234502 2918
rect 234738 2682 234822 2918
rect 235058 2682 235142 2918
rect 235378 2682 235462 2918
rect 235698 2682 235782 2918
rect 236018 2682 236102 2918
rect 236338 2682 236422 2918
rect 236658 2682 236742 2918
rect 236978 2682 237062 2918
rect 237298 2682 237382 2918
rect 237618 2682 237740 2918
rect 233740 2598 237740 2682
rect 233740 2362 233862 2598
rect 234098 2362 234182 2598
rect 234418 2362 234502 2598
rect 234738 2362 234822 2598
rect 235058 2362 235142 2598
rect 235378 2362 235462 2598
rect 235698 2362 235782 2598
rect 236018 2362 236102 2598
rect 236338 2362 236422 2598
rect 236658 2362 236742 2598
rect 236978 2362 237062 2598
rect 237298 2362 237382 2598
rect 237618 2362 237740 2598
rect 233740 2278 237740 2362
rect 233740 2042 233862 2278
rect 234098 2042 234182 2278
rect 234418 2042 234502 2278
rect 234738 2042 234822 2278
rect 235058 2042 235142 2278
rect 235378 2042 235462 2278
rect 235698 2042 235782 2278
rect 236018 2042 236102 2278
rect 236338 2042 236422 2278
rect 236658 2042 236742 2278
rect 236978 2042 237062 2278
rect 237298 2042 237382 2278
rect 237618 2042 237740 2278
rect 233740 1958 237740 2042
rect 233740 1722 233862 1958
rect 234098 1722 234182 1958
rect 234418 1722 234502 1958
rect 234738 1722 234822 1958
rect 235058 1722 235142 1958
rect 235378 1722 235462 1958
rect 235698 1722 235782 1958
rect 236018 1722 236102 1958
rect 236338 1722 236422 1958
rect 236658 1722 236742 1958
rect 236978 1722 237062 1958
rect 237298 1722 237382 1958
rect 237618 1722 237740 1958
rect 233740 1638 237740 1722
rect 233740 1402 233862 1638
rect 234098 1402 234182 1638
rect 234418 1402 234502 1638
rect 234738 1402 234822 1638
rect 235058 1402 235142 1638
rect 235378 1402 235462 1638
rect 235698 1402 235782 1638
rect 236018 1402 236102 1638
rect 236338 1402 236422 1638
rect 236658 1402 236742 1638
rect 236978 1402 237062 1638
rect 237298 1402 237382 1638
rect 237618 1402 237740 1638
rect 233740 1318 237740 1402
rect 233740 1082 233862 1318
rect 234098 1082 234182 1318
rect 234418 1082 234502 1318
rect 234738 1082 234822 1318
rect 235058 1082 235142 1318
rect 235378 1082 235462 1318
rect 235698 1082 235782 1318
rect 236018 1082 236102 1318
rect 236338 1082 236422 1318
rect 236658 1082 236742 1318
rect 236978 1082 237062 1318
rect 237298 1082 237382 1318
rect 237618 1082 237740 1318
rect 233740 998 237740 1082
rect 233740 762 233862 998
rect 234098 762 234182 998
rect 234418 762 234502 998
rect 234738 762 234822 998
rect 235058 762 235142 998
rect 235378 762 235462 998
rect 235698 762 235782 998
rect 236018 762 236102 998
rect 236338 762 236422 998
rect 236658 762 236742 998
rect 236978 762 237062 998
rect 237298 762 237382 998
rect 237618 762 237740 998
rect 233740 678 237740 762
rect 233740 442 233862 678
rect 234098 442 234182 678
rect 234418 442 234502 678
rect 234738 442 234822 678
rect 235058 442 235142 678
rect 235378 442 235462 678
rect 235698 442 235782 678
rect 236018 442 236102 678
rect 236338 442 236422 678
rect 236658 442 236742 678
rect 236978 442 237062 678
rect 237298 442 237382 678
rect 237618 442 237740 678
rect 233740 358 237740 442
rect 233740 122 233862 358
rect 234098 122 234182 358
rect 234418 122 234502 358
rect 234738 122 234822 358
rect 235058 122 235142 358
rect 235378 122 235462 358
rect 235698 122 235782 358
rect 236018 122 236102 358
rect 236338 122 236422 358
rect 236658 122 236742 358
rect 236978 122 237062 358
rect 237298 122 237382 358
rect 237618 122 237740 358
rect 233740 0 237740 122
<< via4 >>
rect 122 255018 358 255254
rect 442 255018 678 255254
rect 762 255018 998 255254
rect 1082 255018 1318 255254
rect 1402 255018 1638 255254
rect 1722 255018 1958 255254
rect 2042 255018 2278 255254
rect 2362 255018 2598 255254
rect 2682 255018 2918 255254
rect 3002 255018 3238 255254
rect 3322 255018 3558 255254
rect 3642 255018 3878 255254
rect 122 254698 358 254934
rect 442 254698 678 254934
rect 762 254698 998 254934
rect 1082 254698 1318 254934
rect 1402 254698 1638 254934
rect 1722 254698 1958 254934
rect 2042 254698 2278 254934
rect 2362 254698 2598 254934
rect 2682 254698 2918 254934
rect 3002 254698 3238 254934
rect 3322 254698 3558 254934
rect 3642 254698 3878 254934
rect 122 254378 358 254614
rect 442 254378 678 254614
rect 762 254378 998 254614
rect 1082 254378 1318 254614
rect 1402 254378 1638 254614
rect 1722 254378 1958 254614
rect 2042 254378 2278 254614
rect 2362 254378 2598 254614
rect 2682 254378 2918 254614
rect 3002 254378 3238 254614
rect 3322 254378 3558 254614
rect 3642 254378 3878 254614
rect 122 254058 358 254294
rect 442 254058 678 254294
rect 762 254058 998 254294
rect 1082 254058 1318 254294
rect 1402 254058 1638 254294
rect 1722 254058 1958 254294
rect 2042 254058 2278 254294
rect 2362 254058 2598 254294
rect 2682 254058 2918 254294
rect 3002 254058 3238 254294
rect 3322 254058 3558 254294
rect 3642 254058 3878 254294
rect 122 253738 358 253974
rect 442 253738 678 253974
rect 762 253738 998 253974
rect 1082 253738 1318 253974
rect 1402 253738 1638 253974
rect 1722 253738 1958 253974
rect 2042 253738 2278 253974
rect 2362 253738 2598 253974
rect 2682 253738 2918 253974
rect 3002 253738 3238 253974
rect 3322 253738 3558 253974
rect 3642 253738 3878 253974
rect 122 253418 358 253654
rect 442 253418 678 253654
rect 762 253418 998 253654
rect 1082 253418 1318 253654
rect 1402 253418 1638 253654
rect 1722 253418 1958 253654
rect 2042 253418 2278 253654
rect 2362 253418 2598 253654
rect 2682 253418 2918 253654
rect 3002 253418 3238 253654
rect 3322 253418 3558 253654
rect 3642 253418 3878 253654
rect 122 253098 358 253334
rect 442 253098 678 253334
rect 762 253098 998 253334
rect 1082 253098 1318 253334
rect 1402 253098 1638 253334
rect 1722 253098 1958 253334
rect 2042 253098 2278 253334
rect 2362 253098 2598 253334
rect 2682 253098 2918 253334
rect 3002 253098 3238 253334
rect 3322 253098 3558 253334
rect 3642 253098 3878 253334
rect 122 252778 358 253014
rect 442 252778 678 253014
rect 762 252778 998 253014
rect 1082 252778 1318 253014
rect 1402 252778 1638 253014
rect 1722 252778 1958 253014
rect 2042 252778 2278 253014
rect 2362 252778 2598 253014
rect 2682 252778 2918 253014
rect 3002 252778 3238 253014
rect 3322 252778 3558 253014
rect 3642 252778 3878 253014
rect 122 252458 358 252694
rect 442 252458 678 252694
rect 762 252458 998 252694
rect 1082 252458 1318 252694
rect 1402 252458 1638 252694
rect 1722 252458 1958 252694
rect 2042 252458 2278 252694
rect 2362 252458 2598 252694
rect 2682 252458 2918 252694
rect 3002 252458 3238 252694
rect 3322 252458 3558 252694
rect 3642 252458 3878 252694
rect 122 252138 358 252374
rect 442 252138 678 252374
rect 762 252138 998 252374
rect 1082 252138 1318 252374
rect 1402 252138 1638 252374
rect 1722 252138 1958 252374
rect 2042 252138 2278 252374
rect 2362 252138 2598 252374
rect 2682 252138 2918 252374
rect 3002 252138 3238 252374
rect 3322 252138 3558 252374
rect 3642 252138 3878 252374
rect 122 251818 358 252054
rect 442 251818 678 252054
rect 762 251818 998 252054
rect 1082 251818 1318 252054
rect 1402 251818 1638 252054
rect 1722 251818 1958 252054
rect 2042 251818 2278 252054
rect 2362 251818 2598 252054
rect 2682 251818 2918 252054
rect 3002 251818 3238 252054
rect 3322 251818 3558 252054
rect 3642 251818 3878 252054
rect 122 251498 358 251734
rect 442 251498 678 251734
rect 762 251498 998 251734
rect 1082 251498 1318 251734
rect 1402 251498 1638 251734
rect 1722 251498 1958 251734
rect 2042 251498 2278 251734
rect 2362 251498 2598 251734
rect 2682 251498 2918 251734
rect 3002 251498 3238 251734
rect 3322 251498 3558 251734
rect 3642 251498 3878 251734
rect 233862 255018 234098 255254
rect 234182 255018 234418 255254
rect 234502 255018 234738 255254
rect 234822 255018 235058 255254
rect 235142 255018 235378 255254
rect 235462 255018 235698 255254
rect 235782 255018 236018 255254
rect 236102 255018 236338 255254
rect 236422 255018 236658 255254
rect 236742 255018 236978 255254
rect 237062 255018 237298 255254
rect 237382 255018 237618 255254
rect 233862 254698 234098 254934
rect 234182 254698 234418 254934
rect 234502 254698 234738 254934
rect 234822 254698 235058 254934
rect 235142 254698 235378 254934
rect 235462 254698 235698 254934
rect 235782 254698 236018 254934
rect 236102 254698 236338 254934
rect 236422 254698 236658 254934
rect 236742 254698 236978 254934
rect 237062 254698 237298 254934
rect 237382 254698 237618 254934
rect 233862 254378 234098 254614
rect 234182 254378 234418 254614
rect 234502 254378 234738 254614
rect 234822 254378 235058 254614
rect 235142 254378 235378 254614
rect 235462 254378 235698 254614
rect 235782 254378 236018 254614
rect 236102 254378 236338 254614
rect 236422 254378 236658 254614
rect 236742 254378 236978 254614
rect 237062 254378 237298 254614
rect 237382 254378 237618 254614
rect 233862 254058 234098 254294
rect 234182 254058 234418 254294
rect 234502 254058 234738 254294
rect 234822 254058 235058 254294
rect 235142 254058 235378 254294
rect 235462 254058 235698 254294
rect 235782 254058 236018 254294
rect 236102 254058 236338 254294
rect 236422 254058 236658 254294
rect 236742 254058 236978 254294
rect 237062 254058 237298 254294
rect 237382 254058 237618 254294
rect 233862 253738 234098 253974
rect 234182 253738 234418 253974
rect 234502 253738 234738 253974
rect 234822 253738 235058 253974
rect 235142 253738 235378 253974
rect 235462 253738 235698 253974
rect 235782 253738 236018 253974
rect 236102 253738 236338 253974
rect 236422 253738 236658 253974
rect 236742 253738 236978 253974
rect 237062 253738 237298 253974
rect 237382 253738 237618 253974
rect 233862 253418 234098 253654
rect 234182 253418 234418 253654
rect 234502 253418 234738 253654
rect 234822 253418 235058 253654
rect 235142 253418 235378 253654
rect 235462 253418 235698 253654
rect 235782 253418 236018 253654
rect 236102 253418 236338 253654
rect 236422 253418 236658 253654
rect 236742 253418 236978 253654
rect 237062 253418 237298 253654
rect 237382 253418 237618 253654
rect 233862 253098 234098 253334
rect 234182 253098 234418 253334
rect 234502 253098 234738 253334
rect 234822 253098 235058 253334
rect 235142 253098 235378 253334
rect 235462 253098 235698 253334
rect 235782 253098 236018 253334
rect 236102 253098 236338 253334
rect 236422 253098 236658 253334
rect 236742 253098 236978 253334
rect 237062 253098 237298 253334
rect 237382 253098 237618 253334
rect 233862 252778 234098 253014
rect 234182 252778 234418 253014
rect 234502 252778 234738 253014
rect 234822 252778 235058 253014
rect 235142 252778 235378 253014
rect 235462 252778 235698 253014
rect 235782 252778 236018 253014
rect 236102 252778 236338 253014
rect 236422 252778 236658 253014
rect 236742 252778 236978 253014
rect 237062 252778 237298 253014
rect 237382 252778 237618 253014
rect 233862 252458 234098 252694
rect 234182 252458 234418 252694
rect 234502 252458 234738 252694
rect 234822 252458 235058 252694
rect 235142 252458 235378 252694
rect 235462 252458 235698 252694
rect 235782 252458 236018 252694
rect 236102 252458 236338 252694
rect 236422 252458 236658 252694
rect 236742 252458 236978 252694
rect 237062 252458 237298 252694
rect 237382 252458 237618 252694
rect 233862 252138 234098 252374
rect 234182 252138 234418 252374
rect 234502 252138 234738 252374
rect 234822 252138 235058 252374
rect 235142 252138 235378 252374
rect 235462 252138 235698 252374
rect 235782 252138 236018 252374
rect 236102 252138 236338 252374
rect 236422 252138 236658 252374
rect 236742 252138 236978 252374
rect 237062 252138 237298 252374
rect 237382 252138 237618 252374
rect 233862 251818 234098 252054
rect 234182 251818 234418 252054
rect 234502 251818 234738 252054
rect 234822 251818 235058 252054
rect 235142 251818 235378 252054
rect 235462 251818 235698 252054
rect 235782 251818 236018 252054
rect 236102 251818 236338 252054
rect 236422 251818 236658 252054
rect 236742 251818 236978 252054
rect 237062 251818 237298 252054
rect 237382 251818 237618 252054
rect 233862 251498 234098 251734
rect 234182 251498 234418 251734
rect 234502 251498 234738 251734
rect 234822 251498 235058 251734
rect 235142 251498 235378 251734
rect 235462 251498 235698 251734
rect 235782 251498 236018 251734
rect 236102 251498 236338 251734
rect 236422 251498 236658 251734
rect 236742 251498 236978 251734
rect 237062 251498 237298 251734
rect 237382 251498 237618 251734
rect 122 228682 358 228918
rect 442 228682 678 228918
rect 762 228682 998 228918
rect 1082 228682 1318 228918
rect 1402 228682 1638 228918
rect 1722 228682 1958 228918
rect 2042 228682 2278 228918
rect 2362 228682 2598 228918
rect 2682 228682 2918 228918
rect 3002 228682 3238 228918
rect 3322 228682 3558 228918
rect 3642 228682 3878 228918
rect 122 206282 358 206518
rect 442 206282 678 206518
rect 762 206282 998 206518
rect 1082 206282 1318 206518
rect 1402 206282 1638 206518
rect 1722 206282 1958 206518
rect 2042 206282 2278 206518
rect 2362 206282 2598 206518
rect 2682 206282 2918 206518
rect 3002 206282 3238 206518
rect 3322 206282 3558 206518
rect 3642 206282 3878 206518
rect 122 183882 358 184118
rect 442 183882 678 184118
rect 762 183882 998 184118
rect 1082 183882 1318 184118
rect 1402 183882 1638 184118
rect 1722 183882 1958 184118
rect 2042 183882 2278 184118
rect 2362 183882 2598 184118
rect 2682 183882 2918 184118
rect 3002 183882 3238 184118
rect 3322 183882 3558 184118
rect 3642 183882 3878 184118
rect 122 161482 358 161718
rect 442 161482 678 161718
rect 762 161482 998 161718
rect 1082 161482 1318 161718
rect 1402 161482 1638 161718
rect 1722 161482 1958 161718
rect 2042 161482 2278 161718
rect 2362 161482 2598 161718
rect 2682 161482 2918 161718
rect 3002 161482 3238 161718
rect 3322 161482 3558 161718
rect 3642 161482 3878 161718
rect 122 139082 358 139318
rect 442 139082 678 139318
rect 762 139082 998 139318
rect 1082 139082 1318 139318
rect 1402 139082 1638 139318
rect 1722 139082 1958 139318
rect 2042 139082 2278 139318
rect 2362 139082 2598 139318
rect 2682 139082 2918 139318
rect 3002 139082 3238 139318
rect 3322 139082 3558 139318
rect 3642 139082 3878 139318
rect 122 116682 358 116918
rect 442 116682 678 116918
rect 762 116682 998 116918
rect 1082 116682 1318 116918
rect 1402 116682 1638 116918
rect 1722 116682 1958 116918
rect 2042 116682 2278 116918
rect 2362 116682 2598 116918
rect 2682 116682 2918 116918
rect 3002 116682 3238 116918
rect 3322 116682 3558 116918
rect 3642 116682 3878 116918
rect 122 94282 358 94518
rect 442 94282 678 94518
rect 762 94282 998 94518
rect 1082 94282 1318 94518
rect 1402 94282 1638 94518
rect 1722 94282 1958 94518
rect 2042 94282 2278 94518
rect 2362 94282 2598 94518
rect 2682 94282 2918 94518
rect 3002 94282 3238 94518
rect 3322 94282 3558 94518
rect 3642 94282 3878 94518
rect 122 71882 358 72118
rect 442 71882 678 72118
rect 762 71882 998 72118
rect 1082 71882 1318 72118
rect 1402 71882 1638 72118
rect 1722 71882 1958 72118
rect 2042 71882 2278 72118
rect 2362 71882 2598 72118
rect 2682 71882 2918 72118
rect 3002 71882 3238 72118
rect 3322 71882 3558 72118
rect 3642 71882 3878 72118
rect 122 49482 358 49718
rect 442 49482 678 49718
rect 762 49482 998 49718
rect 1082 49482 1318 49718
rect 1402 49482 1638 49718
rect 1722 49482 1958 49718
rect 2042 49482 2278 49718
rect 2362 49482 2598 49718
rect 2682 49482 2918 49718
rect 3002 49482 3238 49718
rect 3322 49482 3558 49718
rect 3642 49482 3878 49718
rect 122 27082 358 27318
rect 442 27082 678 27318
rect 762 27082 998 27318
rect 1082 27082 1318 27318
rect 1402 27082 1638 27318
rect 1722 27082 1958 27318
rect 2042 27082 2278 27318
rect 2362 27082 2598 27318
rect 2682 27082 2918 27318
rect 3002 27082 3238 27318
rect 3322 27082 3558 27318
rect 3642 27082 3878 27318
rect 5122 250018 5358 250254
rect 5442 250018 5678 250254
rect 5762 250018 5998 250254
rect 6082 250018 6318 250254
rect 6402 250018 6638 250254
rect 6722 250018 6958 250254
rect 7042 250018 7278 250254
rect 7362 250018 7598 250254
rect 7682 250018 7918 250254
rect 8002 250018 8238 250254
rect 8322 250018 8558 250254
rect 8642 250018 8878 250254
rect 5122 249698 5358 249934
rect 5442 249698 5678 249934
rect 5762 249698 5998 249934
rect 6082 249698 6318 249934
rect 6402 249698 6638 249934
rect 6722 249698 6958 249934
rect 7042 249698 7278 249934
rect 7362 249698 7598 249934
rect 7682 249698 7918 249934
rect 8002 249698 8238 249934
rect 8322 249698 8558 249934
rect 8642 249698 8878 249934
rect 5122 249378 5358 249614
rect 5442 249378 5678 249614
rect 5762 249378 5998 249614
rect 6082 249378 6318 249614
rect 6402 249378 6638 249614
rect 6722 249378 6958 249614
rect 7042 249378 7278 249614
rect 7362 249378 7598 249614
rect 7682 249378 7918 249614
rect 8002 249378 8238 249614
rect 8322 249378 8558 249614
rect 8642 249378 8878 249614
rect 5122 249058 5358 249294
rect 5442 249058 5678 249294
rect 5762 249058 5998 249294
rect 6082 249058 6318 249294
rect 6402 249058 6638 249294
rect 6722 249058 6958 249294
rect 7042 249058 7278 249294
rect 7362 249058 7598 249294
rect 7682 249058 7918 249294
rect 8002 249058 8238 249294
rect 8322 249058 8558 249294
rect 8642 249058 8878 249294
rect 5122 248738 5358 248974
rect 5442 248738 5678 248974
rect 5762 248738 5998 248974
rect 6082 248738 6318 248974
rect 6402 248738 6638 248974
rect 6722 248738 6958 248974
rect 7042 248738 7278 248974
rect 7362 248738 7598 248974
rect 7682 248738 7918 248974
rect 8002 248738 8238 248974
rect 8322 248738 8558 248974
rect 8642 248738 8878 248974
rect 5122 248418 5358 248654
rect 5442 248418 5678 248654
rect 5762 248418 5998 248654
rect 6082 248418 6318 248654
rect 6402 248418 6638 248654
rect 6722 248418 6958 248654
rect 7042 248418 7278 248654
rect 7362 248418 7598 248654
rect 7682 248418 7918 248654
rect 8002 248418 8238 248654
rect 8322 248418 8558 248654
rect 8642 248418 8878 248654
rect 5122 248098 5358 248334
rect 5442 248098 5678 248334
rect 5762 248098 5998 248334
rect 6082 248098 6318 248334
rect 6402 248098 6638 248334
rect 6722 248098 6958 248334
rect 7042 248098 7278 248334
rect 7362 248098 7598 248334
rect 7682 248098 7918 248334
rect 8002 248098 8238 248334
rect 8322 248098 8558 248334
rect 8642 248098 8878 248334
rect 5122 247778 5358 248014
rect 5442 247778 5678 248014
rect 5762 247778 5998 248014
rect 6082 247778 6318 248014
rect 6402 247778 6638 248014
rect 6722 247778 6958 248014
rect 7042 247778 7278 248014
rect 7362 247778 7598 248014
rect 7682 247778 7918 248014
rect 8002 247778 8238 248014
rect 8322 247778 8558 248014
rect 8642 247778 8878 248014
rect 5122 247458 5358 247694
rect 5442 247458 5678 247694
rect 5762 247458 5998 247694
rect 6082 247458 6318 247694
rect 6402 247458 6638 247694
rect 6722 247458 6958 247694
rect 7042 247458 7278 247694
rect 7362 247458 7598 247694
rect 7682 247458 7918 247694
rect 8002 247458 8238 247694
rect 8322 247458 8558 247694
rect 8642 247458 8878 247694
rect 5122 247138 5358 247374
rect 5442 247138 5678 247374
rect 5762 247138 5998 247374
rect 6082 247138 6318 247374
rect 6402 247138 6638 247374
rect 6722 247138 6958 247374
rect 7042 247138 7278 247374
rect 7362 247138 7598 247374
rect 7682 247138 7918 247374
rect 8002 247138 8238 247374
rect 8322 247138 8558 247374
rect 8642 247138 8878 247374
rect 5122 246818 5358 247054
rect 5442 246818 5678 247054
rect 5762 246818 5998 247054
rect 6082 246818 6318 247054
rect 6402 246818 6638 247054
rect 6722 246818 6958 247054
rect 7042 246818 7278 247054
rect 7362 246818 7598 247054
rect 7682 246818 7918 247054
rect 8002 246818 8238 247054
rect 8322 246818 8558 247054
rect 8642 246818 8878 247054
rect 5122 246498 5358 246734
rect 5442 246498 5678 246734
rect 5762 246498 5998 246734
rect 6082 246498 6318 246734
rect 6402 246498 6638 246734
rect 6722 246498 6958 246734
rect 7042 246498 7278 246734
rect 7362 246498 7598 246734
rect 7682 246498 7918 246734
rect 8002 246498 8238 246734
rect 8322 246498 8558 246734
rect 8642 246498 8878 246734
rect 228862 250018 229098 250254
rect 229182 250018 229418 250254
rect 229502 250018 229738 250254
rect 229822 250018 230058 250254
rect 230142 250018 230378 250254
rect 230462 250018 230698 250254
rect 230782 250018 231018 250254
rect 231102 250018 231338 250254
rect 231422 250018 231658 250254
rect 231742 250018 231978 250254
rect 232062 250018 232298 250254
rect 232382 250018 232618 250254
rect 228862 249698 229098 249934
rect 229182 249698 229418 249934
rect 229502 249698 229738 249934
rect 229822 249698 230058 249934
rect 230142 249698 230378 249934
rect 230462 249698 230698 249934
rect 230782 249698 231018 249934
rect 231102 249698 231338 249934
rect 231422 249698 231658 249934
rect 231742 249698 231978 249934
rect 232062 249698 232298 249934
rect 232382 249698 232618 249934
rect 228862 249378 229098 249614
rect 229182 249378 229418 249614
rect 229502 249378 229738 249614
rect 229822 249378 230058 249614
rect 230142 249378 230378 249614
rect 230462 249378 230698 249614
rect 230782 249378 231018 249614
rect 231102 249378 231338 249614
rect 231422 249378 231658 249614
rect 231742 249378 231978 249614
rect 232062 249378 232298 249614
rect 232382 249378 232618 249614
rect 228862 249058 229098 249294
rect 229182 249058 229418 249294
rect 229502 249058 229738 249294
rect 229822 249058 230058 249294
rect 230142 249058 230378 249294
rect 230462 249058 230698 249294
rect 230782 249058 231018 249294
rect 231102 249058 231338 249294
rect 231422 249058 231658 249294
rect 231742 249058 231978 249294
rect 232062 249058 232298 249294
rect 232382 249058 232618 249294
rect 228862 248738 229098 248974
rect 229182 248738 229418 248974
rect 229502 248738 229738 248974
rect 229822 248738 230058 248974
rect 230142 248738 230378 248974
rect 230462 248738 230698 248974
rect 230782 248738 231018 248974
rect 231102 248738 231338 248974
rect 231422 248738 231658 248974
rect 231742 248738 231978 248974
rect 232062 248738 232298 248974
rect 232382 248738 232618 248974
rect 228862 248418 229098 248654
rect 229182 248418 229418 248654
rect 229502 248418 229738 248654
rect 229822 248418 230058 248654
rect 230142 248418 230378 248654
rect 230462 248418 230698 248654
rect 230782 248418 231018 248654
rect 231102 248418 231338 248654
rect 231422 248418 231658 248654
rect 231742 248418 231978 248654
rect 232062 248418 232298 248654
rect 232382 248418 232618 248654
rect 228862 248098 229098 248334
rect 229182 248098 229418 248334
rect 229502 248098 229738 248334
rect 229822 248098 230058 248334
rect 230142 248098 230378 248334
rect 230462 248098 230698 248334
rect 230782 248098 231018 248334
rect 231102 248098 231338 248334
rect 231422 248098 231658 248334
rect 231742 248098 231978 248334
rect 232062 248098 232298 248334
rect 232382 248098 232618 248334
rect 228862 247778 229098 248014
rect 229182 247778 229418 248014
rect 229502 247778 229738 248014
rect 229822 247778 230058 248014
rect 230142 247778 230378 248014
rect 230462 247778 230698 248014
rect 230782 247778 231018 248014
rect 231102 247778 231338 248014
rect 231422 247778 231658 248014
rect 231742 247778 231978 248014
rect 232062 247778 232298 248014
rect 232382 247778 232618 248014
rect 228862 247458 229098 247694
rect 229182 247458 229418 247694
rect 229502 247458 229738 247694
rect 229822 247458 230058 247694
rect 230142 247458 230378 247694
rect 230462 247458 230698 247694
rect 230782 247458 231018 247694
rect 231102 247458 231338 247694
rect 231422 247458 231658 247694
rect 231742 247458 231978 247694
rect 232062 247458 232298 247694
rect 232382 247458 232618 247694
rect 228862 247138 229098 247374
rect 229182 247138 229418 247374
rect 229502 247138 229738 247374
rect 229822 247138 230058 247374
rect 230142 247138 230378 247374
rect 230462 247138 230698 247374
rect 230782 247138 231018 247374
rect 231102 247138 231338 247374
rect 231422 247138 231658 247374
rect 231742 247138 231978 247374
rect 232062 247138 232298 247374
rect 232382 247138 232618 247374
rect 228862 246818 229098 247054
rect 229182 246818 229418 247054
rect 229502 246818 229738 247054
rect 229822 246818 230058 247054
rect 230142 246818 230378 247054
rect 230462 246818 230698 247054
rect 230782 246818 231018 247054
rect 231102 246818 231338 247054
rect 231422 246818 231658 247054
rect 231742 246818 231978 247054
rect 232062 246818 232298 247054
rect 232382 246818 232618 247054
rect 228862 246498 229098 246734
rect 229182 246498 229418 246734
rect 229502 246498 229738 246734
rect 229822 246498 230058 246734
rect 230142 246498 230378 246734
rect 230462 246498 230698 246734
rect 230782 246498 231018 246734
rect 231102 246498 231338 246734
rect 231422 246498 231658 246734
rect 231742 246498 231978 246734
rect 232062 246498 232298 246734
rect 232382 246498 232618 246734
rect 5122 239882 5358 240118
rect 5442 239882 5678 240118
rect 5762 239882 5998 240118
rect 6082 239882 6318 240118
rect 6402 239882 6638 240118
rect 6722 239882 6958 240118
rect 7042 239882 7278 240118
rect 7362 239882 7598 240118
rect 7682 239882 7918 240118
rect 8002 239882 8238 240118
rect 8322 239882 8558 240118
rect 8642 239882 8878 240118
rect 72816 239882 73052 240118
rect 144816 239882 145052 240118
rect 228862 239882 229098 240118
rect 229182 239882 229418 240118
rect 229502 239882 229738 240118
rect 229822 239882 230058 240118
rect 230142 239882 230378 240118
rect 230462 239882 230698 240118
rect 230782 239882 231018 240118
rect 231102 239882 231338 240118
rect 231422 239882 231658 240118
rect 231742 239882 231978 240118
rect 232062 239882 232298 240118
rect 232382 239882 232618 240118
rect 5122 217482 5358 217718
rect 5442 217482 5678 217718
rect 5762 217482 5998 217718
rect 6082 217482 6318 217718
rect 6402 217482 6638 217718
rect 6722 217482 6958 217718
rect 7042 217482 7278 217718
rect 7362 217482 7598 217718
rect 7682 217482 7918 217718
rect 8002 217482 8238 217718
rect 8322 217482 8558 217718
rect 8642 217482 8878 217718
rect 5122 195082 5358 195318
rect 5442 195082 5678 195318
rect 5762 195082 5998 195318
rect 6082 195082 6318 195318
rect 6402 195082 6638 195318
rect 6722 195082 6958 195318
rect 7042 195082 7278 195318
rect 7362 195082 7598 195318
rect 7682 195082 7918 195318
rect 8002 195082 8238 195318
rect 8322 195082 8558 195318
rect 8642 195082 8878 195318
rect 77816 228682 78052 228918
rect 149816 228682 150052 228918
rect 228862 217482 229098 217718
rect 229182 217482 229418 217718
rect 229502 217482 229738 217718
rect 229822 217482 230058 217718
rect 230142 217482 230378 217718
rect 230462 217482 230698 217718
rect 230782 217482 231018 217718
rect 231102 217482 231338 217718
rect 231422 217482 231658 217718
rect 231742 217482 231978 217718
rect 232062 217482 232298 217718
rect 232382 217482 232618 217718
rect 19990 183126 20226 183362
rect 17046 175646 17282 175882
rect 16310 173606 16546 173842
rect 5122 172682 5358 172918
rect 5442 172682 5678 172918
rect 5762 172682 5998 172918
rect 6082 172682 6318 172918
rect 6402 172682 6638 172918
rect 6722 172682 6958 172918
rect 7042 172682 7278 172918
rect 7362 172682 7598 172918
rect 7682 172682 7918 172918
rect 8002 172682 8238 172918
rect 8322 172682 8558 172918
rect 8642 172682 8878 172918
rect 28638 173606 28874 173842
rect 17549 172682 17785 172918
rect 17046 166126 17282 166362
rect 28638 162726 28874 162962
rect 20215 161482 20451 161718
rect 17046 153886 17282 154122
rect 28638 153886 28874 154122
rect 16494 151846 16730 152082
rect 5122 150282 5358 150518
rect 5442 150282 5678 150518
rect 5762 150282 5998 150518
rect 6082 150282 6318 150518
rect 6402 150282 6638 150518
rect 6722 150282 6958 150518
rect 7042 150282 7278 150518
rect 7362 150282 7598 150518
rect 7682 150282 7918 150518
rect 8002 150282 8238 150518
rect 8322 150282 8558 150518
rect 8642 150282 8878 150518
rect 28638 153206 28874 153442
rect 17549 150282 17785 150518
rect 42927 206282 43163 206518
rect 78882 206282 79118 206518
rect 150882 206282 151118 206518
rect 187215 206282 187451 206518
rect 38261 195082 38497 195318
rect 73882 195082 74118 195318
rect 145882 195082 146118 195318
rect 182549 195082 182785 195318
rect 228862 195082 229098 195318
rect 229182 195082 229418 195318
rect 229502 195082 229738 195318
rect 229822 195082 230058 195318
rect 230142 195082 230378 195318
rect 230462 195082 230698 195318
rect 230782 195082 231018 195318
rect 231102 195082 231338 195318
rect 231422 195082 231658 195318
rect 231742 195082 231978 195318
rect 232062 195082 232298 195318
rect 232382 195082 232618 195318
rect 42549 172682 42785 172918
rect 67146 172682 67382 172918
rect 114549 172682 114785 172918
rect 139146 172682 139382 172918
rect 186549 172682 186785 172918
rect 211549 172682 211785 172918
rect 228862 172682 229098 172918
rect 229182 172682 229418 172918
rect 229502 172682 229738 172918
rect 229822 172682 230058 172918
rect 230142 172682 230378 172918
rect 230462 172682 230698 172918
rect 230782 172682 231018 172918
rect 231102 172682 231338 172918
rect 231422 172682 231658 172918
rect 231742 172682 231978 172918
rect 232062 172682 232298 172918
rect 232382 172682 232618 172918
rect 45215 161482 45451 161718
rect 82506 161482 82742 161718
rect 117215 161482 117451 161718
rect 154506 161482 154742 161718
rect 189215 161482 189451 161718
rect 214215 161482 214451 161718
rect 42549 150282 42785 150518
rect 67146 150282 67382 150518
rect 114549 150282 114785 150518
rect 139146 150282 139382 150518
rect 186549 150282 186785 150518
rect 211549 150282 211785 150518
rect 228862 150282 229098 150518
rect 229182 150282 229418 150518
rect 229502 150282 229738 150518
rect 229822 150282 230058 150518
rect 230142 150282 230378 150518
rect 230462 150282 230698 150518
rect 230782 150282 231018 150518
rect 231102 150282 231338 150518
rect 231422 150282 231658 150518
rect 231742 150282 231978 150518
rect 232062 150282 232298 150518
rect 232382 150282 232618 150518
rect 5122 127882 5358 128118
rect 5442 127882 5678 128118
rect 5762 127882 5998 128118
rect 6082 127882 6318 128118
rect 6402 127882 6638 128118
rect 6722 127882 6958 128118
rect 7042 127882 7278 128118
rect 7362 127882 7598 128118
rect 7682 127882 7918 128118
rect 8002 127882 8238 128118
rect 8322 127882 8558 128118
rect 8642 127882 8878 128118
rect 43215 139082 43451 139318
rect 38549 127882 38785 128118
rect 73882 127882 74118 128118
rect 43215 116682 43451 116918
rect 31766 113766 32002 114002
rect 56790 113766 57026 114002
rect 71878 113236 72114 113322
rect 71878 113172 71964 113236
rect 71964 113172 72028 113236
rect 72028 113172 72114 113236
rect 71878 113086 72114 113172
rect 5122 105482 5358 105718
rect 5442 105482 5678 105718
rect 5762 105482 5998 105718
rect 6082 105482 6318 105718
rect 6402 105482 6638 105718
rect 6722 105482 6958 105718
rect 7042 105482 7278 105718
rect 7362 105482 7598 105718
rect 7682 105482 7918 105718
rect 8002 105482 8238 105718
rect 8322 105482 8558 105718
rect 8642 105482 8878 105718
rect 17549 105482 17785 105718
rect 42549 105482 42785 105718
rect 67146 105482 67382 105718
rect 20215 94282 20451 94518
rect 45215 94282 45451 94518
rect 82506 94282 82742 94518
rect 5122 83082 5358 83318
rect 5442 83082 5678 83318
rect 5762 83082 5998 83318
rect 6082 83082 6318 83318
rect 6402 83082 6638 83318
rect 6722 83082 6958 83318
rect 7042 83082 7278 83318
rect 7362 83082 7598 83318
rect 7682 83082 7918 83318
rect 8002 83082 8238 83318
rect 8322 83082 8558 83318
rect 8642 83082 8878 83318
rect 17549 83082 17785 83318
rect 42549 83082 42785 83318
rect 67146 83082 67382 83318
rect 115215 139082 115451 139318
rect 110549 127882 110785 128118
rect 145882 127882 146118 128118
rect 115215 116682 115451 116918
rect 114549 105482 114785 105718
rect 139146 105482 139382 105718
rect 117215 94282 117451 94518
rect 154506 94282 154742 94518
rect 114549 83082 114785 83318
rect 139146 83082 139382 83318
rect 5122 60682 5358 60918
rect 5442 60682 5678 60918
rect 5762 60682 5998 60918
rect 6082 60682 6318 60918
rect 6402 60682 6638 60918
rect 6722 60682 6958 60918
rect 7042 60682 7278 60918
rect 7362 60682 7598 60918
rect 7682 60682 7918 60918
rect 8002 60682 8238 60918
rect 8322 60682 8558 60918
rect 8642 60682 8878 60918
rect 38549 60682 38785 60918
rect 73882 60682 74118 60918
rect 110549 60682 110785 60918
rect 43215 49482 43451 49718
rect 78882 49482 79118 49718
rect 115215 49482 115451 49718
rect 31766 41006 32002 41242
rect 66174 41006 66410 41242
rect 187215 139082 187451 139318
rect 182549 127882 182785 128118
rect 228862 127882 229098 128118
rect 229182 127882 229418 128118
rect 229502 127882 229738 128118
rect 229822 127882 230058 128118
rect 230142 127882 230378 128118
rect 230462 127882 230698 128118
rect 230782 127882 231018 128118
rect 231102 127882 231338 128118
rect 231422 127882 231658 128118
rect 231742 127882 231978 128118
rect 232062 127882 232298 128118
rect 232382 127882 232618 128118
rect 187215 116682 187451 116918
rect 186549 105482 186785 105718
rect 211549 105482 211785 105718
rect 228862 105482 229098 105718
rect 229182 105482 229418 105718
rect 229502 105482 229738 105718
rect 229822 105482 230058 105718
rect 230142 105482 230378 105718
rect 230462 105482 230698 105718
rect 230782 105482 231018 105718
rect 231102 105482 231338 105718
rect 231422 105482 231658 105718
rect 231742 105482 231978 105718
rect 232062 105482 232298 105718
rect 232382 105482 232618 105718
rect 189215 94282 189451 94518
rect 214215 94282 214451 94518
rect 186549 83082 186785 83318
rect 211549 83082 211785 83318
rect 228862 83082 229098 83318
rect 229182 83082 229418 83318
rect 229502 83082 229738 83318
rect 229822 83082 230058 83318
rect 230142 83082 230378 83318
rect 230462 83082 230698 83318
rect 230782 83082 231018 83318
rect 231102 83082 231338 83318
rect 231422 83082 231658 83318
rect 231742 83082 231978 83318
rect 232062 83082 232298 83318
rect 232382 83082 232618 83318
rect 145882 60682 146118 60918
rect 182549 60682 182785 60918
rect 150882 49482 151118 49718
rect 187215 49482 187451 49718
rect 228862 60682 229098 60918
rect 229182 60682 229418 60918
rect 229502 60682 229738 60918
rect 229822 60682 230058 60918
rect 230142 60682 230378 60918
rect 230462 60682 230698 60918
rect 230782 60682 231018 60918
rect 231102 60682 231338 60918
rect 231422 60682 231658 60918
rect 231742 60682 231978 60918
rect 232062 60682 232298 60918
rect 232382 60682 232618 60918
rect 93774 40476 94010 40562
rect 93774 40412 93860 40476
rect 93860 40412 93924 40476
rect 93924 40412 94010 40476
rect 93774 40326 94010 40412
rect 108678 40326 108914 40562
rect 109598 40326 109834 40562
rect 129654 40326 129890 40562
rect 136830 40326 137066 40562
rect 181358 40326 181594 40562
rect 166086 39796 166322 39882
rect 166086 39732 166172 39796
rect 166172 39732 166236 39796
rect 166236 39732 166322 39796
rect 166086 39646 166322 39732
rect 201414 38966 201650 39202
rect 5122 38282 5358 38518
rect 5442 38282 5678 38518
rect 5762 38282 5998 38518
rect 6082 38282 6318 38518
rect 6402 38282 6638 38518
rect 6722 38282 6958 38518
rect 7042 38282 7278 38518
rect 7362 38282 7598 38518
rect 7682 38282 7918 38518
rect 8002 38282 8238 38518
rect 8322 38282 8558 38518
rect 8642 38282 8878 38518
rect 228862 38282 229098 38518
rect 229182 38282 229418 38518
rect 229502 38282 229738 38518
rect 229822 38282 230058 38518
rect 230142 38282 230378 38518
rect 230462 38282 230698 38518
rect 230782 38282 231018 38518
rect 231102 38282 231338 38518
rect 231422 38282 231658 38518
rect 231742 38282 231978 38518
rect 232062 38282 232298 38518
rect 232382 38282 232618 38518
rect 78882 27082 79118 27318
rect 150882 27082 151118 27318
rect 5122 15882 5358 16118
rect 5442 15882 5678 16118
rect 5762 15882 5998 16118
rect 6082 15882 6318 16118
rect 6402 15882 6638 16118
rect 6722 15882 6958 16118
rect 7042 15882 7278 16118
rect 7362 15882 7598 16118
rect 7682 15882 7918 16118
rect 8002 15882 8238 16118
rect 8322 15882 8558 16118
rect 8642 15882 8878 16118
rect 73882 15882 74118 16118
rect 145882 15882 146118 16118
rect 228862 15882 229098 16118
rect 229182 15882 229418 16118
rect 229502 15882 229738 16118
rect 229822 15882 230058 16118
rect 230142 15882 230378 16118
rect 230462 15882 230698 16118
rect 230782 15882 231018 16118
rect 231102 15882 231338 16118
rect 231422 15882 231658 16118
rect 231742 15882 231978 16118
rect 232062 15882 232298 16118
rect 232382 15882 232618 16118
rect 5122 8642 5358 8878
rect 5442 8642 5678 8878
rect 5762 8642 5998 8878
rect 6082 8642 6318 8878
rect 6402 8642 6638 8878
rect 6722 8642 6958 8878
rect 7042 8642 7278 8878
rect 7362 8642 7598 8878
rect 7682 8642 7918 8878
rect 8002 8642 8238 8878
rect 8322 8642 8558 8878
rect 8642 8642 8878 8878
rect 5122 8322 5358 8558
rect 5442 8322 5678 8558
rect 5762 8322 5998 8558
rect 6082 8322 6318 8558
rect 6402 8322 6638 8558
rect 6722 8322 6958 8558
rect 7042 8322 7278 8558
rect 7362 8322 7598 8558
rect 7682 8322 7918 8558
rect 8002 8322 8238 8558
rect 8322 8322 8558 8558
rect 8642 8322 8878 8558
rect 5122 8002 5358 8238
rect 5442 8002 5678 8238
rect 5762 8002 5998 8238
rect 6082 8002 6318 8238
rect 6402 8002 6638 8238
rect 6722 8002 6958 8238
rect 7042 8002 7278 8238
rect 7362 8002 7598 8238
rect 7682 8002 7918 8238
rect 8002 8002 8238 8238
rect 8322 8002 8558 8238
rect 8642 8002 8878 8238
rect 5122 7682 5358 7918
rect 5442 7682 5678 7918
rect 5762 7682 5998 7918
rect 6082 7682 6318 7918
rect 6402 7682 6638 7918
rect 6722 7682 6958 7918
rect 7042 7682 7278 7918
rect 7362 7682 7598 7918
rect 7682 7682 7918 7918
rect 8002 7682 8238 7918
rect 8322 7682 8558 7918
rect 8642 7682 8878 7918
rect 5122 7362 5358 7598
rect 5442 7362 5678 7598
rect 5762 7362 5998 7598
rect 6082 7362 6318 7598
rect 6402 7362 6638 7598
rect 6722 7362 6958 7598
rect 7042 7362 7278 7598
rect 7362 7362 7598 7598
rect 7682 7362 7918 7598
rect 8002 7362 8238 7598
rect 8322 7362 8558 7598
rect 8642 7362 8878 7598
rect 5122 7042 5358 7278
rect 5442 7042 5678 7278
rect 5762 7042 5998 7278
rect 6082 7042 6318 7278
rect 6402 7042 6638 7278
rect 6722 7042 6958 7278
rect 7042 7042 7278 7278
rect 7362 7042 7598 7278
rect 7682 7042 7918 7278
rect 8002 7042 8238 7278
rect 8322 7042 8558 7278
rect 8642 7042 8878 7278
rect 5122 6722 5358 6958
rect 5442 6722 5678 6958
rect 5762 6722 5998 6958
rect 6082 6722 6318 6958
rect 6402 6722 6638 6958
rect 6722 6722 6958 6958
rect 7042 6722 7278 6958
rect 7362 6722 7598 6958
rect 7682 6722 7918 6958
rect 8002 6722 8238 6958
rect 8322 6722 8558 6958
rect 8642 6722 8878 6958
rect 5122 6402 5358 6638
rect 5442 6402 5678 6638
rect 5762 6402 5998 6638
rect 6082 6402 6318 6638
rect 6402 6402 6638 6638
rect 6722 6402 6958 6638
rect 7042 6402 7278 6638
rect 7362 6402 7598 6638
rect 7682 6402 7918 6638
rect 8002 6402 8238 6638
rect 8322 6402 8558 6638
rect 8642 6402 8878 6638
rect 5122 6082 5358 6318
rect 5442 6082 5678 6318
rect 5762 6082 5998 6318
rect 6082 6082 6318 6318
rect 6402 6082 6638 6318
rect 6722 6082 6958 6318
rect 7042 6082 7278 6318
rect 7362 6082 7598 6318
rect 7682 6082 7918 6318
rect 8002 6082 8238 6318
rect 8322 6082 8558 6318
rect 8642 6082 8878 6318
rect 5122 5762 5358 5998
rect 5442 5762 5678 5998
rect 5762 5762 5998 5998
rect 6082 5762 6318 5998
rect 6402 5762 6638 5998
rect 6722 5762 6958 5998
rect 7042 5762 7278 5998
rect 7362 5762 7598 5998
rect 7682 5762 7918 5998
rect 8002 5762 8238 5998
rect 8322 5762 8558 5998
rect 8642 5762 8878 5998
rect 5122 5442 5358 5678
rect 5442 5442 5678 5678
rect 5762 5442 5998 5678
rect 6082 5442 6318 5678
rect 6402 5442 6638 5678
rect 6722 5442 6958 5678
rect 7042 5442 7278 5678
rect 7362 5442 7598 5678
rect 7682 5442 7918 5678
rect 8002 5442 8238 5678
rect 8322 5442 8558 5678
rect 8642 5442 8878 5678
rect 5122 5122 5358 5358
rect 5442 5122 5678 5358
rect 5762 5122 5998 5358
rect 6082 5122 6318 5358
rect 6402 5122 6638 5358
rect 6722 5122 6958 5358
rect 7042 5122 7278 5358
rect 7362 5122 7598 5358
rect 7682 5122 7918 5358
rect 8002 5122 8238 5358
rect 8322 5122 8558 5358
rect 8642 5122 8878 5358
rect 228862 8642 229098 8878
rect 229182 8642 229418 8878
rect 229502 8642 229738 8878
rect 229822 8642 230058 8878
rect 230142 8642 230378 8878
rect 230462 8642 230698 8878
rect 230782 8642 231018 8878
rect 231102 8642 231338 8878
rect 231422 8642 231658 8878
rect 231742 8642 231978 8878
rect 232062 8642 232298 8878
rect 232382 8642 232618 8878
rect 228862 8322 229098 8558
rect 229182 8322 229418 8558
rect 229502 8322 229738 8558
rect 229822 8322 230058 8558
rect 230142 8322 230378 8558
rect 230462 8322 230698 8558
rect 230782 8322 231018 8558
rect 231102 8322 231338 8558
rect 231422 8322 231658 8558
rect 231742 8322 231978 8558
rect 232062 8322 232298 8558
rect 232382 8322 232618 8558
rect 228862 8002 229098 8238
rect 229182 8002 229418 8238
rect 229502 8002 229738 8238
rect 229822 8002 230058 8238
rect 230142 8002 230378 8238
rect 230462 8002 230698 8238
rect 230782 8002 231018 8238
rect 231102 8002 231338 8238
rect 231422 8002 231658 8238
rect 231742 8002 231978 8238
rect 232062 8002 232298 8238
rect 232382 8002 232618 8238
rect 228862 7682 229098 7918
rect 229182 7682 229418 7918
rect 229502 7682 229738 7918
rect 229822 7682 230058 7918
rect 230142 7682 230378 7918
rect 230462 7682 230698 7918
rect 230782 7682 231018 7918
rect 231102 7682 231338 7918
rect 231422 7682 231658 7918
rect 231742 7682 231978 7918
rect 232062 7682 232298 7918
rect 232382 7682 232618 7918
rect 228862 7362 229098 7598
rect 229182 7362 229418 7598
rect 229502 7362 229738 7598
rect 229822 7362 230058 7598
rect 230142 7362 230378 7598
rect 230462 7362 230698 7598
rect 230782 7362 231018 7598
rect 231102 7362 231338 7598
rect 231422 7362 231658 7598
rect 231742 7362 231978 7598
rect 232062 7362 232298 7598
rect 232382 7362 232618 7598
rect 228862 7042 229098 7278
rect 229182 7042 229418 7278
rect 229502 7042 229738 7278
rect 229822 7042 230058 7278
rect 230142 7042 230378 7278
rect 230462 7042 230698 7278
rect 230782 7042 231018 7278
rect 231102 7042 231338 7278
rect 231422 7042 231658 7278
rect 231742 7042 231978 7278
rect 232062 7042 232298 7278
rect 232382 7042 232618 7278
rect 228862 6722 229098 6958
rect 229182 6722 229418 6958
rect 229502 6722 229738 6958
rect 229822 6722 230058 6958
rect 230142 6722 230378 6958
rect 230462 6722 230698 6958
rect 230782 6722 231018 6958
rect 231102 6722 231338 6958
rect 231422 6722 231658 6958
rect 231742 6722 231978 6958
rect 232062 6722 232298 6958
rect 232382 6722 232618 6958
rect 228862 6402 229098 6638
rect 229182 6402 229418 6638
rect 229502 6402 229738 6638
rect 229822 6402 230058 6638
rect 230142 6402 230378 6638
rect 230462 6402 230698 6638
rect 230782 6402 231018 6638
rect 231102 6402 231338 6638
rect 231422 6402 231658 6638
rect 231742 6402 231978 6638
rect 232062 6402 232298 6638
rect 232382 6402 232618 6638
rect 228862 6082 229098 6318
rect 229182 6082 229418 6318
rect 229502 6082 229738 6318
rect 229822 6082 230058 6318
rect 230142 6082 230378 6318
rect 230462 6082 230698 6318
rect 230782 6082 231018 6318
rect 231102 6082 231338 6318
rect 231422 6082 231658 6318
rect 231742 6082 231978 6318
rect 232062 6082 232298 6318
rect 232382 6082 232618 6318
rect 228862 5762 229098 5998
rect 229182 5762 229418 5998
rect 229502 5762 229738 5998
rect 229822 5762 230058 5998
rect 230142 5762 230378 5998
rect 230462 5762 230698 5998
rect 230782 5762 231018 5998
rect 231102 5762 231338 5998
rect 231422 5762 231658 5998
rect 231742 5762 231978 5998
rect 232062 5762 232298 5998
rect 232382 5762 232618 5998
rect 228862 5442 229098 5678
rect 229182 5442 229418 5678
rect 229502 5442 229738 5678
rect 229822 5442 230058 5678
rect 230142 5442 230378 5678
rect 230462 5442 230698 5678
rect 230782 5442 231018 5678
rect 231102 5442 231338 5678
rect 231422 5442 231658 5678
rect 231742 5442 231978 5678
rect 232062 5442 232298 5678
rect 232382 5442 232618 5678
rect 228862 5122 229098 5358
rect 229182 5122 229418 5358
rect 229502 5122 229738 5358
rect 229822 5122 230058 5358
rect 230142 5122 230378 5358
rect 230462 5122 230698 5358
rect 230782 5122 231018 5358
rect 231102 5122 231338 5358
rect 231422 5122 231658 5358
rect 231742 5122 231978 5358
rect 232062 5122 232298 5358
rect 232382 5122 232618 5358
rect 233862 228682 234098 228918
rect 234182 228682 234418 228918
rect 234502 228682 234738 228918
rect 234822 228682 235058 228918
rect 235142 228682 235378 228918
rect 235462 228682 235698 228918
rect 235782 228682 236018 228918
rect 236102 228682 236338 228918
rect 236422 228682 236658 228918
rect 236742 228682 236978 228918
rect 237062 228682 237298 228918
rect 237382 228682 237618 228918
rect 233862 206282 234098 206518
rect 234182 206282 234418 206518
rect 234502 206282 234738 206518
rect 234822 206282 235058 206518
rect 235142 206282 235378 206518
rect 235462 206282 235698 206518
rect 235782 206282 236018 206518
rect 236102 206282 236338 206518
rect 236422 206282 236658 206518
rect 236742 206282 236978 206518
rect 237062 206282 237298 206518
rect 237382 206282 237618 206518
rect 233862 183882 234098 184118
rect 234182 183882 234418 184118
rect 234502 183882 234738 184118
rect 234822 183882 235058 184118
rect 235142 183882 235378 184118
rect 235462 183882 235698 184118
rect 235782 183882 236018 184118
rect 236102 183882 236338 184118
rect 236422 183882 236658 184118
rect 236742 183882 236978 184118
rect 237062 183882 237298 184118
rect 237382 183882 237618 184118
rect 233862 161482 234098 161718
rect 234182 161482 234418 161718
rect 234502 161482 234738 161718
rect 234822 161482 235058 161718
rect 235142 161482 235378 161718
rect 235462 161482 235698 161718
rect 235782 161482 236018 161718
rect 236102 161482 236338 161718
rect 236422 161482 236658 161718
rect 236742 161482 236978 161718
rect 237062 161482 237298 161718
rect 237382 161482 237618 161718
rect 233862 139082 234098 139318
rect 234182 139082 234418 139318
rect 234502 139082 234738 139318
rect 234822 139082 235058 139318
rect 235142 139082 235378 139318
rect 235462 139082 235698 139318
rect 235782 139082 236018 139318
rect 236102 139082 236338 139318
rect 236422 139082 236658 139318
rect 236742 139082 236978 139318
rect 237062 139082 237298 139318
rect 237382 139082 237618 139318
rect 233862 116682 234098 116918
rect 234182 116682 234418 116918
rect 234502 116682 234738 116918
rect 234822 116682 235058 116918
rect 235142 116682 235378 116918
rect 235462 116682 235698 116918
rect 235782 116682 236018 116918
rect 236102 116682 236338 116918
rect 236422 116682 236658 116918
rect 236742 116682 236978 116918
rect 237062 116682 237298 116918
rect 237382 116682 237618 116918
rect 233862 94282 234098 94518
rect 234182 94282 234418 94518
rect 234502 94282 234738 94518
rect 234822 94282 235058 94518
rect 235142 94282 235378 94518
rect 235462 94282 235698 94518
rect 235782 94282 236018 94518
rect 236102 94282 236338 94518
rect 236422 94282 236658 94518
rect 236742 94282 236978 94518
rect 237062 94282 237298 94518
rect 237382 94282 237618 94518
rect 233862 71882 234098 72118
rect 234182 71882 234418 72118
rect 234502 71882 234738 72118
rect 234822 71882 235058 72118
rect 235142 71882 235378 72118
rect 235462 71882 235698 72118
rect 235782 71882 236018 72118
rect 236102 71882 236338 72118
rect 236422 71882 236658 72118
rect 236742 71882 236978 72118
rect 237062 71882 237298 72118
rect 237382 71882 237618 72118
rect 233862 49482 234098 49718
rect 234182 49482 234418 49718
rect 234502 49482 234738 49718
rect 234822 49482 235058 49718
rect 235142 49482 235378 49718
rect 235462 49482 235698 49718
rect 235782 49482 236018 49718
rect 236102 49482 236338 49718
rect 236422 49482 236658 49718
rect 236742 49482 236978 49718
rect 237062 49482 237298 49718
rect 237382 49482 237618 49718
rect 233862 27082 234098 27318
rect 234182 27082 234418 27318
rect 234502 27082 234738 27318
rect 234822 27082 235058 27318
rect 235142 27082 235378 27318
rect 235462 27082 235698 27318
rect 235782 27082 236018 27318
rect 236102 27082 236338 27318
rect 236422 27082 236658 27318
rect 236742 27082 236978 27318
rect 237062 27082 237298 27318
rect 237382 27082 237618 27318
rect 122 3642 358 3878
rect 442 3642 678 3878
rect 762 3642 998 3878
rect 1082 3642 1318 3878
rect 1402 3642 1638 3878
rect 1722 3642 1958 3878
rect 2042 3642 2278 3878
rect 2362 3642 2598 3878
rect 2682 3642 2918 3878
rect 3002 3642 3238 3878
rect 3322 3642 3558 3878
rect 3642 3642 3878 3878
rect 122 3322 358 3558
rect 442 3322 678 3558
rect 762 3322 998 3558
rect 1082 3322 1318 3558
rect 1402 3322 1638 3558
rect 1722 3322 1958 3558
rect 2042 3322 2278 3558
rect 2362 3322 2598 3558
rect 2682 3322 2918 3558
rect 3002 3322 3238 3558
rect 3322 3322 3558 3558
rect 3642 3322 3878 3558
rect 122 3002 358 3238
rect 442 3002 678 3238
rect 762 3002 998 3238
rect 1082 3002 1318 3238
rect 1402 3002 1638 3238
rect 1722 3002 1958 3238
rect 2042 3002 2278 3238
rect 2362 3002 2598 3238
rect 2682 3002 2918 3238
rect 3002 3002 3238 3238
rect 3322 3002 3558 3238
rect 3642 3002 3878 3238
rect 122 2682 358 2918
rect 442 2682 678 2918
rect 762 2682 998 2918
rect 1082 2682 1318 2918
rect 1402 2682 1638 2918
rect 1722 2682 1958 2918
rect 2042 2682 2278 2918
rect 2362 2682 2598 2918
rect 2682 2682 2918 2918
rect 3002 2682 3238 2918
rect 3322 2682 3558 2918
rect 3642 2682 3878 2918
rect 122 2362 358 2598
rect 442 2362 678 2598
rect 762 2362 998 2598
rect 1082 2362 1318 2598
rect 1402 2362 1638 2598
rect 1722 2362 1958 2598
rect 2042 2362 2278 2598
rect 2362 2362 2598 2598
rect 2682 2362 2918 2598
rect 3002 2362 3238 2598
rect 3322 2362 3558 2598
rect 3642 2362 3878 2598
rect 122 2042 358 2278
rect 442 2042 678 2278
rect 762 2042 998 2278
rect 1082 2042 1318 2278
rect 1402 2042 1638 2278
rect 1722 2042 1958 2278
rect 2042 2042 2278 2278
rect 2362 2042 2598 2278
rect 2682 2042 2918 2278
rect 3002 2042 3238 2278
rect 3322 2042 3558 2278
rect 3642 2042 3878 2278
rect 122 1722 358 1958
rect 442 1722 678 1958
rect 762 1722 998 1958
rect 1082 1722 1318 1958
rect 1402 1722 1638 1958
rect 1722 1722 1958 1958
rect 2042 1722 2278 1958
rect 2362 1722 2598 1958
rect 2682 1722 2918 1958
rect 3002 1722 3238 1958
rect 3322 1722 3558 1958
rect 3642 1722 3878 1958
rect 122 1402 358 1638
rect 442 1402 678 1638
rect 762 1402 998 1638
rect 1082 1402 1318 1638
rect 1402 1402 1638 1638
rect 1722 1402 1958 1638
rect 2042 1402 2278 1638
rect 2362 1402 2598 1638
rect 2682 1402 2918 1638
rect 3002 1402 3238 1638
rect 3322 1402 3558 1638
rect 3642 1402 3878 1638
rect 122 1082 358 1318
rect 442 1082 678 1318
rect 762 1082 998 1318
rect 1082 1082 1318 1318
rect 1402 1082 1638 1318
rect 1722 1082 1958 1318
rect 2042 1082 2278 1318
rect 2362 1082 2598 1318
rect 2682 1082 2918 1318
rect 3002 1082 3238 1318
rect 3322 1082 3558 1318
rect 3642 1082 3878 1318
rect 122 762 358 998
rect 442 762 678 998
rect 762 762 998 998
rect 1082 762 1318 998
rect 1402 762 1638 998
rect 1722 762 1958 998
rect 2042 762 2278 998
rect 2362 762 2598 998
rect 2682 762 2918 998
rect 3002 762 3238 998
rect 3322 762 3558 998
rect 3642 762 3878 998
rect 122 442 358 678
rect 442 442 678 678
rect 762 442 998 678
rect 1082 442 1318 678
rect 1402 442 1638 678
rect 1722 442 1958 678
rect 2042 442 2278 678
rect 2362 442 2598 678
rect 2682 442 2918 678
rect 3002 442 3238 678
rect 3322 442 3558 678
rect 3642 442 3878 678
rect 122 122 358 358
rect 442 122 678 358
rect 762 122 998 358
rect 1082 122 1318 358
rect 1402 122 1638 358
rect 1722 122 1958 358
rect 2042 122 2278 358
rect 2362 122 2598 358
rect 2682 122 2918 358
rect 3002 122 3238 358
rect 3322 122 3558 358
rect 3642 122 3878 358
rect 233862 3642 234098 3878
rect 234182 3642 234418 3878
rect 234502 3642 234738 3878
rect 234822 3642 235058 3878
rect 235142 3642 235378 3878
rect 235462 3642 235698 3878
rect 235782 3642 236018 3878
rect 236102 3642 236338 3878
rect 236422 3642 236658 3878
rect 236742 3642 236978 3878
rect 237062 3642 237298 3878
rect 237382 3642 237618 3878
rect 233862 3322 234098 3558
rect 234182 3322 234418 3558
rect 234502 3322 234738 3558
rect 234822 3322 235058 3558
rect 235142 3322 235378 3558
rect 235462 3322 235698 3558
rect 235782 3322 236018 3558
rect 236102 3322 236338 3558
rect 236422 3322 236658 3558
rect 236742 3322 236978 3558
rect 237062 3322 237298 3558
rect 237382 3322 237618 3558
rect 233862 3002 234098 3238
rect 234182 3002 234418 3238
rect 234502 3002 234738 3238
rect 234822 3002 235058 3238
rect 235142 3002 235378 3238
rect 235462 3002 235698 3238
rect 235782 3002 236018 3238
rect 236102 3002 236338 3238
rect 236422 3002 236658 3238
rect 236742 3002 236978 3238
rect 237062 3002 237298 3238
rect 237382 3002 237618 3238
rect 233862 2682 234098 2918
rect 234182 2682 234418 2918
rect 234502 2682 234738 2918
rect 234822 2682 235058 2918
rect 235142 2682 235378 2918
rect 235462 2682 235698 2918
rect 235782 2682 236018 2918
rect 236102 2682 236338 2918
rect 236422 2682 236658 2918
rect 236742 2682 236978 2918
rect 237062 2682 237298 2918
rect 237382 2682 237618 2918
rect 233862 2362 234098 2598
rect 234182 2362 234418 2598
rect 234502 2362 234738 2598
rect 234822 2362 235058 2598
rect 235142 2362 235378 2598
rect 235462 2362 235698 2598
rect 235782 2362 236018 2598
rect 236102 2362 236338 2598
rect 236422 2362 236658 2598
rect 236742 2362 236978 2598
rect 237062 2362 237298 2598
rect 237382 2362 237618 2598
rect 233862 2042 234098 2278
rect 234182 2042 234418 2278
rect 234502 2042 234738 2278
rect 234822 2042 235058 2278
rect 235142 2042 235378 2278
rect 235462 2042 235698 2278
rect 235782 2042 236018 2278
rect 236102 2042 236338 2278
rect 236422 2042 236658 2278
rect 236742 2042 236978 2278
rect 237062 2042 237298 2278
rect 237382 2042 237618 2278
rect 233862 1722 234098 1958
rect 234182 1722 234418 1958
rect 234502 1722 234738 1958
rect 234822 1722 235058 1958
rect 235142 1722 235378 1958
rect 235462 1722 235698 1958
rect 235782 1722 236018 1958
rect 236102 1722 236338 1958
rect 236422 1722 236658 1958
rect 236742 1722 236978 1958
rect 237062 1722 237298 1958
rect 237382 1722 237618 1958
rect 233862 1402 234098 1638
rect 234182 1402 234418 1638
rect 234502 1402 234738 1638
rect 234822 1402 235058 1638
rect 235142 1402 235378 1638
rect 235462 1402 235698 1638
rect 235782 1402 236018 1638
rect 236102 1402 236338 1638
rect 236422 1402 236658 1638
rect 236742 1402 236978 1638
rect 237062 1402 237298 1638
rect 237382 1402 237618 1638
rect 233862 1082 234098 1318
rect 234182 1082 234418 1318
rect 234502 1082 234738 1318
rect 234822 1082 235058 1318
rect 235142 1082 235378 1318
rect 235462 1082 235698 1318
rect 235782 1082 236018 1318
rect 236102 1082 236338 1318
rect 236422 1082 236658 1318
rect 236742 1082 236978 1318
rect 237062 1082 237298 1318
rect 237382 1082 237618 1318
rect 233862 762 234098 998
rect 234182 762 234418 998
rect 234502 762 234738 998
rect 234822 762 235058 998
rect 235142 762 235378 998
rect 235462 762 235698 998
rect 235782 762 236018 998
rect 236102 762 236338 998
rect 236422 762 236658 998
rect 236742 762 236978 998
rect 237062 762 237298 998
rect 237382 762 237618 998
rect 233862 442 234098 678
rect 234182 442 234418 678
rect 234502 442 234738 678
rect 234822 442 235058 678
rect 235142 442 235378 678
rect 235462 442 235698 678
rect 235782 442 236018 678
rect 236102 442 236338 678
rect 236422 442 236658 678
rect 236742 442 236978 678
rect 237062 442 237298 678
rect 237382 442 237618 678
rect 233862 122 234098 358
rect 234182 122 234418 358
rect 234502 122 234738 358
rect 234822 122 235058 358
rect 235142 122 235378 358
rect 235462 122 235698 358
rect 235782 122 236018 358
rect 236102 122 236338 358
rect 236422 122 236658 358
rect 236742 122 236978 358
rect 237062 122 237298 358
rect 237382 122 237618 358
<< metal5 >>
rect 0 255254 237740 255376
rect 0 255018 122 255254
rect 358 255018 442 255254
rect 678 255018 762 255254
rect 998 255018 1082 255254
rect 1318 255018 1402 255254
rect 1638 255018 1722 255254
rect 1958 255018 2042 255254
rect 2278 255018 2362 255254
rect 2598 255018 2682 255254
rect 2918 255018 3002 255254
rect 3238 255018 3322 255254
rect 3558 255018 3642 255254
rect 3878 255018 233862 255254
rect 234098 255018 234182 255254
rect 234418 255018 234502 255254
rect 234738 255018 234822 255254
rect 235058 255018 235142 255254
rect 235378 255018 235462 255254
rect 235698 255018 235782 255254
rect 236018 255018 236102 255254
rect 236338 255018 236422 255254
rect 236658 255018 236742 255254
rect 236978 255018 237062 255254
rect 237298 255018 237382 255254
rect 237618 255018 237740 255254
rect 0 254934 237740 255018
rect 0 254698 122 254934
rect 358 254698 442 254934
rect 678 254698 762 254934
rect 998 254698 1082 254934
rect 1318 254698 1402 254934
rect 1638 254698 1722 254934
rect 1958 254698 2042 254934
rect 2278 254698 2362 254934
rect 2598 254698 2682 254934
rect 2918 254698 3002 254934
rect 3238 254698 3322 254934
rect 3558 254698 3642 254934
rect 3878 254698 233862 254934
rect 234098 254698 234182 254934
rect 234418 254698 234502 254934
rect 234738 254698 234822 254934
rect 235058 254698 235142 254934
rect 235378 254698 235462 254934
rect 235698 254698 235782 254934
rect 236018 254698 236102 254934
rect 236338 254698 236422 254934
rect 236658 254698 236742 254934
rect 236978 254698 237062 254934
rect 237298 254698 237382 254934
rect 237618 254698 237740 254934
rect 0 254614 237740 254698
rect 0 254378 122 254614
rect 358 254378 442 254614
rect 678 254378 762 254614
rect 998 254378 1082 254614
rect 1318 254378 1402 254614
rect 1638 254378 1722 254614
rect 1958 254378 2042 254614
rect 2278 254378 2362 254614
rect 2598 254378 2682 254614
rect 2918 254378 3002 254614
rect 3238 254378 3322 254614
rect 3558 254378 3642 254614
rect 3878 254378 233862 254614
rect 234098 254378 234182 254614
rect 234418 254378 234502 254614
rect 234738 254378 234822 254614
rect 235058 254378 235142 254614
rect 235378 254378 235462 254614
rect 235698 254378 235782 254614
rect 236018 254378 236102 254614
rect 236338 254378 236422 254614
rect 236658 254378 236742 254614
rect 236978 254378 237062 254614
rect 237298 254378 237382 254614
rect 237618 254378 237740 254614
rect 0 254294 237740 254378
rect 0 254058 122 254294
rect 358 254058 442 254294
rect 678 254058 762 254294
rect 998 254058 1082 254294
rect 1318 254058 1402 254294
rect 1638 254058 1722 254294
rect 1958 254058 2042 254294
rect 2278 254058 2362 254294
rect 2598 254058 2682 254294
rect 2918 254058 3002 254294
rect 3238 254058 3322 254294
rect 3558 254058 3642 254294
rect 3878 254058 233862 254294
rect 234098 254058 234182 254294
rect 234418 254058 234502 254294
rect 234738 254058 234822 254294
rect 235058 254058 235142 254294
rect 235378 254058 235462 254294
rect 235698 254058 235782 254294
rect 236018 254058 236102 254294
rect 236338 254058 236422 254294
rect 236658 254058 236742 254294
rect 236978 254058 237062 254294
rect 237298 254058 237382 254294
rect 237618 254058 237740 254294
rect 0 253974 237740 254058
rect 0 253738 122 253974
rect 358 253738 442 253974
rect 678 253738 762 253974
rect 998 253738 1082 253974
rect 1318 253738 1402 253974
rect 1638 253738 1722 253974
rect 1958 253738 2042 253974
rect 2278 253738 2362 253974
rect 2598 253738 2682 253974
rect 2918 253738 3002 253974
rect 3238 253738 3322 253974
rect 3558 253738 3642 253974
rect 3878 253738 233862 253974
rect 234098 253738 234182 253974
rect 234418 253738 234502 253974
rect 234738 253738 234822 253974
rect 235058 253738 235142 253974
rect 235378 253738 235462 253974
rect 235698 253738 235782 253974
rect 236018 253738 236102 253974
rect 236338 253738 236422 253974
rect 236658 253738 236742 253974
rect 236978 253738 237062 253974
rect 237298 253738 237382 253974
rect 237618 253738 237740 253974
rect 0 253654 237740 253738
rect 0 253418 122 253654
rect 358 253418 442 253654
rect 678 253418 762 253654
rect 998 253418 1082 253654
rect 1318 253418 1402 253654
rect 1638 253418 1722 253654
rect 1958 253418 2042 253654
rect 2278 253418 2362 253654
rect 2598 253418 2682 253654
rect 2918 253418 3002 253654
rect 3238 253418 3322 253654
rect 3558 253418 3642 253654
rect 3878 253418 233862 253654
rect 234098 253418 234182 253654
rect 234418 253418 234502 253654
rect 234738 253418 234822 253654
rect 235058 253418 235142 253654
rect 235378 253418 235462 253654
rect 235698 253418 235782 253654
rect 236018 253418 236102 253654
rect 236338 253418 236422 253654
rect 236658 253418 236742 253654
rect 236978 253418 237062 253654
rect 237298 253418 237382 253654
rect 237618 253418 237740 253654
rect 0 253334 237740 253418
rect 0 253098 122 253334
rect 358 253098 442 253334
rect 678 253098 762 253334
rect 998 253098 1082 253334
rect 1318 253098 1402 253334
rect 1638 253098 1722 253334
rect 1958 253098 2042 253334
rect 2278 253098 2362 253334
rect 2598 253098 2682 253334
rect 2918 253098 3002 253334
rect 3238 253098 3322 253334
rect 3558 253098 3642 253334
rect 3878 253098 233862 253334
rect 234098 253098 234182 253334
rect 234418 253098 234502 253334
rect 234738 253098 234822 253334
rect 235058 253098 235142 253334
rect 235378 253098 235462 253334
rect 235698 253098 235782 253334
rect 236018 253098 236102 253334
rect 236338 253098 236422 253334
rect 236658 253098 236742 253334
rect 236978 253098 237062 253334
rect 237298 253098 237382 253334
rect 237618 253098 237740 253334
rect 0 253014 237740 253098
rect 0 252778 122 253014
rect 358 252778 442 253014
rect 678 252778 762 253014
rect 998 252778 1082 253014
rect 1318 252778 1402 253014
rect 1638 252778 1722 253014
rect 1958 252778 2042 253014
rect 2278 252778 2362 253014
rect 2598 252778 2682 253014
rect 2918 252778 3002 253014
rect 3238 252778 3322 253014
rect 3558 252778 3642 253014
rect 3878 252778 233862 253014
rect 234098 252778 234182 253014
rect 234418 252778 234502 253014
rect 234738 252778 234822 253014
rect 235058 252778 235142 253014
rect 235378 252778 235462 253014
rect 235698 252778 235782 253014
rect 236018 252778 236102 253014
rect 236338 252778 236422 253014
rect 236658 252778 236742 253014
rect 236978 252778 237062 253014
rect 237298 252778 237382 253014
rect 237618 252778 237740 253014
rect 0 252694 237740 252778
rect 0 252458 122 252694
rect 358 252458 442 252694
rect 678 252458 762 252694
rect 998 252458 1082 252694
rect 1318 252458 1402 252694
rect 1638 252458 1722 252694
rect 1958 252458 2042 252694
rect 2278 252458 2362 252694
rect 2598 252458 2682 252694
rect 2918 252458 3002 252694
rect 3238 252458 3322 252694
rect 3558 252458 3642 252694
rect 3878 252458 233862 252694
rect 234098 252458 234182 252694
rect 234418 252458 234502 252694
rect 234738 252458 234822 252694
rect 235058 252458 235142 252694
rect 235378 252458 235462 252694
rect 235698 252458 235782 252694
rect 236018 252458 236102 252694
rect 236338 252458 236422 252694
rect 236658 252458 236742 252694
rect 236978 252458 237062 252694
rect 237298 252458 237382 252694
rect 237618 252458 237740 252694
rect 0 252374 237740 252458
rect 0 252138 122 252374
rect 358 252138 442 252374
rect 678 252138 762 252374
rect 998 252138 1082 252374
rect 1318 252138 1402 252374
rect 1638 252138 1722 252374
rect 1958 252138 2042 252374
rect 2278 252138 2362 252374
rect 2598 252138 2682 252374
rect 2918 252138 3002 252374
rect 3238 252138 3322 252374
rect 3558 252138 3642 252374
rect 3878 252138 233862 252374
rect 234098 252138 234182 252374
rect 234418 252138 234502 252374
rect 234738 252138 234822 252374
rect 235058 252138 235142 252374
rect 235378 252138 235462 252374
rect 235698 252138 235782 252374
rect 236018 252138 236102 252374
rect 236338 252138 236422 252374
rect 236658 252138 236742 252374
rect 236978 252138 237062 252374
rect 237298 252138 237382 252374
rect 237618 252138 237740 252374
rect 0 252054 237740 252138
rect 0 251818 122 252054
rect 358 251818 442 252054
rect 678 251818 762 252054
rect 998 251818 1082 252054
rect 1318 251818 1402 252054
rect 1638 251818 1722 252054
rect 1958 251818 2042 252054
rect 2278 251818 2362 252054
rect 2598 251818 2682 252054
rect 2918 251818 3002 252054
rect 3238 251818 3322 252054
rect 3558 251818 3642 252054
rect 3878 251818 233862 252054
rect 234098 251818 234182 252054
rect 234418 251818 234502 252054
rect 234738 251818 234822 252054
rect 235058 251818 235142 252054
rect 235378 251818 235462 252054
rect 235698 251818 235782 252054
rect 236018 251818 236102 252054
rect 236338 251818 236422 252054
rect 236658 251818 236742 252054
rect 236978 251818 237062 252054
rect 237298 251818 237382 252054
rect 237618 251818 237740 252054
rect 0 251734 237740 251818
rect 0 251498 122 251734
rect 358 251498 442 251734
rect 678 251498 762 251734
rect 998 251498 1082 251734
rect 1318 251498 1402 251734
rect 1638 251498 1722 251734
rect 1958 251498 2042 251734
rect 2278 251498 2362 251734
rect 2598 251498 2682 251734
rect 2918 251498 3002 251734
rect 3238 251498 3322 251734
rect 3558 251498 3642 251734
rect 3878 251498 233862 251734
rect 234098 251498 234182 251734
rect 234418 251498 234502 251734
rect 234738 251498 234822 251734
rect 235058 251498 235142 251734
rect 235378 251498 235462 251734
rect 235698 251498 235782 251734
rect 236018 251498 236102 251734
rect 236338 251498 236422 251734
rect 236658 251498 236742 251734
rect 236978 251498 237062 251734
rect 237298 251498 237382 251734
rect 237618 251498 237740 251734
rect 0 251376 237740 251498
rect 5000 250254 232740 250376
rect 5000 250018 5122 250254
rect 5358 250018 5442 250254
rect 5678 250018 5762 250254
rect 5998 250018 6082 250254
rect 6318 250018 6402 250254
rect 6638 250018 6722 250254
rect 6958 250018 7042 250254
rect 7278 250018 7362 250254
rect 7598 250018 7682 250254
rect 7918 250018 8002 250254
rect 8238 250018 8322 250254
rect 8558 250018 8642 250254
rect 8878 250018 228862 250254
rect 229098 250018 229182 250254
rect 229418 250018 229502 250254
rect 229738 250018 229822 250254
rect 230058 250018 230142 250254
rect 230378 250018 230462 250254
rect 230698 250018 230782 250254
rect 231018 250018 231102 250254
rect 231338 250018 231422 250254
rect 231658 250018 231742 250254
rect 231978 250018 232062 250254
rect 232298 250018 232382 250254
rect 232618 250018 232740 250254
rect 5000 249934 232740 250018
rect 5000 249698 5122 249934
rect 5358 249698 5442 249934
rect 5678 249698 5762 249934
rect 5998 249698 6082 249934
rect 6318 249698 6402 249934
rect 6638 249698 6722 249934
rect 6958 249698 7042 249934
rect 7278 249698 7362 249934
rect 7598 249698 7682 249934
rect 7918 249698 8002 249934
rect 8238 249698 8322 249934
rect 8558 249698 8642 249934
rect 8878 249698 228862 249934
rect 229098 249698 229182 249934
rect 229418 249698 229502 249934
rect 229738 249698 229822 249934
rect 230058 249698 230142 249934
rect 230378 249698 230462 249934
rect 230698 249698 230782 249934
rect 231018 249698 231102 249934
rect 231338 249698 231422 249934
rect 231658 249698 231742 249934
rect 231978 249698 232062 249934
rect 232298 249698 232382 249934
rect 232618 249698 232740 249934
rect 5000 249614 232740 249698
rect 5000 249378 5122 249614
rect 5358 249378 5442 249614
rect 5678 249378 5762 249614
rect 5998 249378 6082 249614
rect 6318 249378 6402 249614
rect 6638 249378 6722 249614
rect 6958 249378 7042 249614
rect 7278 249378 7362 249614
rect 7598 249378 7682 249614
rect 7918 249378 8002 249614
rect 8238 249378 8322 249614
rect 8558 249378 8642 249614
rect 8878 249378 228862 249614
rect 229098 249378 229182 249614
rect 229418 249378 229502 249614
rect 229738 249378 229822 249614
rect 230058 249378 230142 249614
rect 230378 249378 230462 249614
rect 230698 249378 230782 249614
rect 231018 249378 231102 249614
rect 231338 249378 231422 249614
rect 231658 249378 231742 249614
rect 231978 249378 232062 249614
rect 232298 249378 232382 249614
rect 232618 249378 232740 249614
rect 5000 249294 232740 249378
rect 5000 249058 5122 249294
rect 5358 249058 5442 249294
rect 5678 249058 5762 249294
rect 5998 249058 6082 249294
rect 6318 249058 6402 249294
rect 6638 249058 6722 249294
rect 6958 249058 7042 249294
rect 7278 249058 7362 249294
rect 7598 249058 7682 249294
rect 7918 249058 8002 249294
rect 8238 249058 8322 249294
rect 8558 249058 8642 249294
rect 8878 249058 228862 249294
rect 229098 249058 229182 249294
rect 229418 249058 229502 249294
rect 229738 249058 229822 249294
rect 230058 249058 230142 249294
rect 230378 249058 230462 249294
rect 230698 249058 230782 249294
rect 231018 249058 231102 249294
rect 231338 249058 231422 249294
rect 231658 249058 231742 249294
rect 231978 249058 232062 249294
rect 232298 249058 232382 249294
rect 232618 249058 232740 249294
rect 5000 248974 232740 249058
rect 5000 248738 5122 248974
rect 5358 248738 5442 248974
rect 5678 248738 5762 248974
rect 5998 248738 6082 248974
rect 6318 248738 6402 248974
rect 6638 248738 6722 248974
rect 6958 248738 7042 248974
rect 7278 248738 7362 248974
rect 7598 248738 7682 248974
rect 7918 248738 8002 248974
rect 8238 248738 8322 248974
rect 8558 248738 8642 248974
rect 8878 248738 228862 248974
rect 229098 248738 229182 248974
rect 229418 248738 229502 248974
rect 229738 248738 229822 248974
rect 230058 248738 230142 248974
rect 230378 248738 230462 248974
rect 230698 248738 230782 248974
rect 231018 248738 231102 248974
rect 231338 248738 231422 248974
rect 231658 248738 231742 248974
rect 231978 248738 232062 248974
rect 232298 248738 232382 248974
rect 232618 248738 232740 248974
rect 5000 248654 232740 248738
rect 5000 248418 5122 248654
rect 5358 248418 5442 248654
rect 5678 248418 5762 248654
rect 5998 248418 6082 248654
rect 6318 248418 6402 248654
rect 6638 248418 6722 248654
rect 6958 248418 7042 248654
rect 7278 248418 7362 248654
rect 7598 248418 7682 248654
rect 7918 248418 8002 248654
rect 8238 248418 8322 248654
rect 8558 248418 8642 248654
rect 8878 248418 228862 248654
rect 229098 248418 229182 248654
rect 229418 248418 229502 248654
rect 229738 248418 229822 248654
rect 230058 248418 230142 248654
rect 230378 248418 230462 248654
rect 230698 248418 230782 248654
rect 231018 248418 231102 248654
rect 231338 248418 231422 248654
rect 231658 248418 231742 248654
rect 231978 248418 232062 248654
rect 232298 248418 232382 248654
rect 232618 248418 232740 248654
rect 5000 248334 232740 248418
rect 5000 248098 5122 248334
rect 5358 248098 5442 248334
rect 5678 248098 5762 248334
rect 5998 248098 6082 248334
rect 6318 248098 6402 248334
rect 6638 248098 6722 248334
rect 6958 248098 7042 248334
rect 7278 248098 7362 248334
rect 7598 248098 7682 248334
rect 7918 248098 8002 248334
rect 8238 248098 8322 248334
rect 8558 248098 8642 248334
rect 8878 248098 228862 248334
rect 229098 248098 229182 248334
rect 229418 248098 229502 248334
rect 229738 248098 229822 248334
rect 230058 248098 230142 248334
rect 230378 248098 230462 248334
rect 230698 248098 230782 248334
rect 231018 248098 231102 248334
rect 231338 248098 231422 248334
rect 231658 248098 231742 248334
rect 231978 248098 232062 248334
rect 232298 248098 232382 248334
rect 232618 248098 232740 248334
rect 5000 248014 232740 248098
rect 5000 247778 5122 248014
rect 5358 247778 5442 248014
rect 5678 247778 5762 248014
rect 5998 247778 6082 248014
rect 6318 247778 6402 248014
rect 6638 247778 6722 248014
rect 6958 247778 7042 248014
rect 7278 247778 7362 248014
rect 7598 247778 7682 248014
rect 7918 247778 8002 248014
rect 8238 247778 8322 248014
rect 8558 247778 8642 248014
rect 8878 247778 228862 248014
rect 229098 247778 229182 248014
rect 229418 247778 229502 248014
rect 229738 247778 229822 248014
rect 230058 247778 230142 248014
rect 230378 247778 230462 248014
rect 230698 247778 230782 248014
rect 231018 247778 231102 248014
rect 231338 247778 231422 248014
rect 231658 247778 231742 248014
rect 231978 247778 232062 248014
rect 232298 247778 232382 248014
rect 232618 247778 232740 248014
rect 5000 247694 232740 247778
rect 5000 247458 5122 247694
rect 5358 247458 5442 247694
rect 5678 247458 5762 247694
rect 5998 247458 6082 247694
rect 6318 247458 6402 247694
rect 6638 247458 6722 247694
rect 6958 247458 7042 247694
rect 7278 247458 7362 247694
rect 7598 247458 7682 247694
rect 7918 247458 8002 247694
rect 8238 247458 8322 247694
rect 8558 247458 8642 247694
rect 8878 247458 228862 247694
rect 229098 247458 229182 247694
rect 229418 247458 229502 247694
rect 229738 247458 229822 247694
rect 230058 247458 230142 247694
rect 230378 247458 230462 247694
rect 230698 247458 230782 247694
rect 231018 247458 231102 247694
rect 231338 247458 231422 247694
rect 231658 247458 231742 247694
rect 231978 247458 232062 247694
rect 232298 247458 232382 247694
rect 232618 247458 232740 247694
rect 5000 247374 232740 247458
rect 5000 247138 5122 247374
rect 5358 247138 5442 247374
rect 5678 247138 5762 247374
rect 5998 247138 6082 247374
rect 6318 247138 6402 247374
rect 6638 247138 6722 247374
rect 6958 247138 7042 247374
rect 7278 247138 7362 247374
rect 7598 247138 7682 247374
rect 7918 247138 8002 247374
rect 8238 247138 8322 247374
rect 8558 247138 8642 247374
rect 8878 247138 228862 247374
rect 229098 247138 229182 247374
rect 229418 247138 229502 247374
rect 229738 247138 229822 247374
rect 230058 247138 230142 247374
rect 230378 247138 230462 247374
rect 230698 247138 230782 247374
rect 231018 247138 231102 247374
rect 231338 247138 231422 247374
rect 231658 247138 231742 247374
rect 231978 247138 232062 247374
rect 232298 247138 232382 247374
rect 232618 247138 232740 247374
rect 5000 247054 232740 247138
rect 5000 246818 5122 247054
rect 5358 246818 5442 247054
rect 5678 246818 5762 247054
rect 5998 246818 6082 247054
rect 6318 246818 6402 247054
rect 6638 246818 6722 247054
rect 6958 246818 7042 247054
rect 7278 246818 7362 247054
rect 7598 246818 7682 247054
rect 7918 246818 8002 247054
rect 8238 246818 8322 247054
rect 8558 246818 8642 247054
rect 8878 246818 228862 247054
rect 229098 246818 229182 247054
rect 229418 246818 229502 247054
rect 229738 246818 229822 247054
rect 230058 246818 230142 247054
rect 230378 246818 230462 247054
rect 230698 246818 230782 247054
rect 231018 246818 231102 247054
rect 231338 246818 231422 247054
rect 231658 246818 231742 247054
rect 231978 246818 232062 247054
rect 232298 246818 232382 247054
rect 232618 246818 232740 247054
rect 5000 246734 232740 246818
rect 5000 246498 5122 246734
rect 5358 246498 5442 246734
rect 5678 246498 5762 246734
rect 5998 246498 6082 246734
rect 6318 246498 6402 246734
rect 6638 246498 6722 246734
rect 6958 246498 7042 246734
rect 7278 246498 7362 246734
rect 7598 246498 7682 246734
rect 7918 246498 8002 246734
rect 8238 246498 8322 246734
rect 8558 246498 8642 246734
rect 8878 246498 228862 246734
rect 229098 246498 229182 246734
rect 229418 246498 229502 246734
rect 229738 246498 229822 246734
rect 230058 246498 230142 246734
rect 230378 246498 230462 246734
rect 230698 246498 230782 246734
rect 231018 246498 231102 246734
rect 231338 246498 231422 246734
rect 231658 246498 231742 246734
rect 231978 246498 232062 246734
rect 232298 246498 232382 246734
rect 232618 246498 232740 246734
rect 5000 246376 232740 246498
rect 0 240118 237740 240160
rect 0 239882 5122 240118
rect 5358 239882 5442 240118
rect 5678 239882 5762 240118
rect 5998 239882 6082 240118
rect 6318 239882 6402 240118
rect 6638 239882 6722 240118
rect 6958 239882 7042 240118
rect 7278 239882 7362 240118
rect 7598 239882 7682 240118
rect 7918 239882 8002 240118
rect 8238 239882 8322 240118
rect 8558 239882 8642 240118
rect 8878 239882 72816 240118
rect 73052 239882 144816 240118
rect 145052 239882 228862 240118
rect 229098 239882 229182 240118
rect 229418 239882 229502 240118
rect 229738 239882 229822 240118
rect 230058 239882 230142 240118
rect 230378 239882 230462 240118
rect 230698 239882 230782 240118
rect 231018 239882 231102 240118
rect 231338 239882 231422 240118
rect 231658 239882 231742 240118
rect 231978 239882 232062 240118
rect 232298 239882 232382 240118
rect 232618 239882 237740 240118
rect 0 239840 237740 239882
rect 0 228918 237740 228960
rect 0 228682 122 228918
rect 358 228682 442 228918
rect 678 228682 762 228918
rect 998 228682 1082 228918
rect 1318 228682 1402 228918
rect 1638 228682 1722 228918
rect 1958 228682 2042 228918
rect 2278 228682 2362 228918
rect 2598 228682 2682 228918
rect 2918 228682 3002 228918
rect 3238 228682 3322 228918
rect 3558 228682 3642 228918
rect 3878 228682 77816 228918
rect 78052 228682 149816 228918
rect 150052 228682 233862 228918
rect 234098 228682 234182 228918
rect 234418 228682 234502 228918
rect 234738 228682 234822 228918
rect 235058 228682 235142 228918
rect 235378 228682 235462 228918
rect 235698 228682 235782 228918
rect 236018 228682 236102 228918
rect 236338 228682 236422 228918
rect 236658 228682 236742 228918
rect 236978 228682 237062 228918
rect 237298 228682 237382 228918
rect 237618 228682 237740 228918
rect 0 228640 237740 228682
rect 0 217718 237740 217760
rect 0 217482 5122 217718
rect 5358 217482 5442 217718
rect 5678 217482 5762 217718
rect 5998 217482 6082 217718
rect 6318 217482 6402 217718
rect 6638 217482 6722 217718
rect 6958 217482 7042 217718
rect 7278 217482 7362 217718
rect 7598 217482 7682 217718
rect 7918 217482 8002 217718
rect 8238 217482 8322 217718
rect 8558 217482 8642 217718
rect 8878 217482 228862 217718
rect 229098 217482 229182 217718
rect 229418 217482 229502 217718
rect 229738 217482 229822 217718
rect 230058 217482 230142 217718
rect 230378 217482 230462 217718
rect 230698 217482 230782 217718
rect 231018 217482 231102 217718
rect 231338 217482 231422 217718
rect 231658 217482 231742 217718
rect 231978 217482 232062 217718
rect 232298 217482 232382 217718
rect 232618 217482 237740 217718
rect 0 217440 237740 217482
rect 0 206518 237740 206560
rect 0 206282 122 206518
rect 358 206282 442 206518
rect 678 206282 762 206518
rect 998 206282 1082 206518
rect 1318 206282 1402 206518
rect 1638 206282 1722 206518
rect 1958 206282 2042 206518
rect 2278 206282 2362 206518
rect 2598 206282 2682 206518
rect 2918 206282 3002 206518
rect 3238 206282 3322 206518
rect 3558 206282 3642 206518
rect 3878 206282 42927 206518
rect 43163 206282 78882 206518
rect 79118 206282 150882 206518
rect 151118 206282 187215 206518
rect 187451 206282 233862 206518
rect 234098 206282 234182 206518
rect 234418 206282 234502 206518
rect 234738 206282 234822 206518
rect 235058 206282 235142 206518
rect 235378 206282 235462 206518
rect 235698 206282 235782 206518
rect 236018 206282 236102 206518
rect 236338 206282 236422 206518
rect 236658 206282 236742 206518
rect 236978 206282 237062 206518
rect 237298 206282 237382 206518
rect 237618 206282 237740 206518
rect 0 206240 237740 206282
rect 0 195318 237740 195360
rect 0 195082 5122 195318
rect 5358 195082 5442 195318
rect 5678 195082 5762 195318
rect 5998 195082 6082 195318
rect 6318 195082 6402 195318
rect 6638 195082 6722 195318
rect 6958 195082 7042 195318
rect 7278 195082 7362 195318
rect 7598 195082 7682 195318
rect 7918 195082 8002 195318
rect 8238 195082 8322 195318
rect 8558 195082 8642 195318
rect 8878 195082 38261 195318
rect 38497 195082 73882 195318
rect 74118 195082 145882 195318
rect 146118 195082 182549 195318
rect 182785 195082 228862 195318
rect 229098 195082 229182 195318
rect 229418 195082 229502 195318
rect 229738 195082 229822 195318
rect 230058 195082 230142 195318
rect 230378 195082 230462 195318
rect 230698 195082 230782 195318
rect 231018 195082 231102 195318
rect 231338 195082 231422 195318
rect 231658 195082 231742 195318
rect 231978 195082 232062 195318
rect 232298 195082 232382 195318
rect 232618 195082 237740 195318
rect 0 195040 237740 195082
rect 0 184118 237740 184160
rect 0 183882 122 184118
rect 358 183882 442 184118
rect 678 183882 762 184118
rect 998 183882 1082 184118
rect 1318 183882 1402 184118
rect 1638 183882 1722 184118
rect 1958 183882 2042 184118
rect 2278 183882 2362 184118
rect 2598 183882 2682 184118
rect 2918 183882 3002 184118
rect 3238 183882 3322 184118
rect 3558 183882 3642 184118
rect 3878 183882 233862 184118
rect 234098 183882 234182 184118
rect 234418 183882 234502 184118
rect 234738 183882 234822 184118
rect 235058 183882 235142 184118
rect 235378 183882 235462 184118
rect 235698 183882 235782 184118
rect 236018 183882 236102 184118
rect 236338 183882 236422 184118
rect 236658 183882 236742 184118
rect 236978 183882 237062 184118
rect 237298 183882 237382 184118
rect 237618 183882 237740 184118
rect 0 183840 237740 183882
rect 19948 183362 20636 183404
rect 19948 183126 19990 183362
rect 20226 183126 20636 183362
rect 19948 183084 20636 183126
rect 20316 175924 20636 183084
rect 17004 175882 20636 175924
rect 17004 175646 17046 175882
rect 17282 175646 20636 175882
rect 17004 175604 20636 175646
rect 16268 173842 28916 173884
rect 16268 173606 16310 173842
rect 16546 173606 28638 173842
rect 28874 173606 28916 173842
rect 16268 173564 28916 173606
rect 0 172918 237740 172960
rect 0 172682 5122 172918
rect 5358 172682 5442 172918
rect 5678 172682 5762 172918
rect 5998 172682 6082 172918
rect 6318 172682 6402 172918
rect 6638 172682 6722 172918
rect 6958 172682 7042 172918
rect 7278 172682 7362 172918
rect 7598 172682 7682 172918
rect 7918 172682 8002 172918
rect 8238 172682 8322 172918
rect 8558 172682 8642 172918
rect 8878 172682 17549 172918
rect 17785 172682 42549 172918
rect 42785 172682 67146 172918
rect 67382 172682 114549 172918
rect 114785 172682 139146 172918
rect 139382 172682 186549 172918
rect 186785 172682 211549 172918
rect 211785 172682 228862 172918
rect 229098 172682 229182 172918
rect 229418 172682 229502 172918
rect 229738 172682 229822 172918
rect 230058 172682 230142 172918
rect 230378 172682 230462 172918
rect 230698 172682 230782 172918
rect 231018 172682 231102 172918
rect 231338 172682 231422 172918
rect 231658 172682 231742 172918
rect 231978 172682 232062 172918
rect 232298 172682 232382 172918
rect 232618 172682 237740 172918
rect 0 172640 237740 172682
rect 17004 166362 19716 166404
rect 17004 166126 17046 166362
rect 17282 166126 19716 166362
rect 17004 166084 19716 166126
rect 19396 164364 19716 166084
rect 19396 164044 20636 164364
rect 20316 163004 20636 164044
rect 20316 162962 28916 163004
rect 20316 162726 28638 162962
rect 28874 162726 28916 162962
rect 20316 162684 28916 162726
rect 0 161718 237740 161760
rect 0 161482 122 161718
rect 358 161482 442 161718
rect 678 161482 762 161718
rect 998 161482 1082 161718
rect 1318 161482 1402 161718
rect 1638 161482 1722 161718
rect 1958 161482 2042 161718
rect 2278 161482 2362 161718
rect 2598 161482 2682 161718
rect 2918 161482 3002 161718
rect 3238 161482 3322 161718
rect 3558 161482 3642 161718
rect 3878 161482 20215 161718
rect 20451 161482 45215 161718
rect 45451 161482 82506 161718
rect 82742 161482 117215 161718
rect 117451 161482 154506 161718
rect 154742 161482 189215 161718
rect 189451 161482 214215 161718
rect 214451 161482 233862 161718
rect 234098 161482 234182 161718
rect 234418 161482 234502 161718
rect 234738 161482 234822 161718
rect 235058 161482 235142 161718
rect 235378 161482 235462 161718
rect 235698 161482 235782 161718
rect 236018 161482 236102 161718
rect 236338 161482 236422 161718
rect 236658 161482 236742 161718
rect 236978 161482 237062 161718
rect 237298 161482 237382 161718
rect 237618 161482 237740 161718
rect 0 161440 237740 161482
rect 17004 154122 28916 154164
rect 17004 153886 17046 154122
rect 17282 153886 28638 154122
rect 28874 153886 28916 154122
rect 17004 153844 28916 153886
rect 17556 153442 28916 153484
rect 17556 153206 28638 153442
rect 28874 153206 28916 153442
rect 17556 153164 28916 153206
rect 17556 152124 17876 153164
rect 16452 152082 17876 152124
rect 16452 151846 16494 152082
rect 16730 151846 17876 152082
rect 16452 151804 17876 151846
rect 0 150518 237740 150560
rect 0 150282 5122 150518
rect 5358 150282 5442 150518
rect 5678 150282 5762 150518
rect 5998 150282 6082 150518
rect 6318 150282 6402 150518
rect 6638 150282 6722 150518
rect 6958 150282 7042 150518
rect 7278 150282 7362 150518
rect 7598 150282 7682 150518
rect 7918 150282 8002 150518
rect 8238 150282 8322 150518
rect 8558 150282 8642 150518
rect 8878 150282 17549 150518
rect 17785 150282 42549 150518
rect 42785 150282 67146 150518
rect 67382 150282 114549 150518
rect 114785 150282 139146 150518
rect 139382 150282 186549 150518
rect 186785 150282 211549 150518
rect 211785 150282 228862 150518
rect 229098 150282 229182 150518
rect 229418 150282 229502 150518
rect 229738 150282 229822 150518
rect 230058 150282 230142 150518
rect 230378 150282 230462 150518
rect 230698 150282 230782 150518
rect 231018 150282 231102 150518
rect 231338 150282 231422 150518
rect 231658 150282 231742 150518
rect 231978 150282 232062 150518
rect 232298 150282 232382 150518
rect 232618 150282 237740 150518
rect 0 150240 237740 150282
rect 0 139318 237740 139360
rect 0 139082 122 139318
rect 358 139082 442 139318
rect 678 139082 762 139318
rect 998 139082 1082 139318
rect 1318 139082 1402 139318
rect 1638 139082 1722 139318
rect 1958 139082 2042 139318
rect 2278 139082 2362 139318
rect 2598 139082 2682 139318
rect 2918 139082 3002 139318
rect 3238 139082 3322 139318
rect 3558 139082 3642 139318
rect 3878 139082 43215 139318
rect 43451 139082 115215 139318
rect 115451 139082 187215 139318
rect 187451 139082 233862 139318
rect 234098 139082 234182 139318
rect 234418 139082 234502 139318
rect 234738 139082 234822 139318
rect 235058 139082 235142 139318
rect 235378 139082 235462 139318
rect 235698 139082 235782 139318
rect 236018 139082 236102 139318
rect 236338 139082 236422 139318
rect 236658 139082 236742 139318
rect 236978 139082 237062 139318
rect 237298 139082 237382 139318
rect 237618 139082 237740 139318
rect 0 139040 237740 139082
rect 0 128118 237740 128160
rect 0 127882 5122 128118
rect 5358 127882 5442 128118
rect 5678 127882 5762 128118
rect 5998 127882 6082 128118
rect 6318 127882 6402 128118
rect 6638 127882 6722 128118
rect 6958 127882 7042 128118
rect 7278 127882 7362 128118
rect 7598 127882 7682 128118
rect 7918 127882 8002 128118
rect 8238 127882 8322 128118
rect 8558 127882 8642 128118
rect 8878 127882 38549 128118
rect 38785 127882 73882 128118
rect 74118 127882 110549 128118
rect 110785 127882 145882 128118
rect 146118 127882 182549 128118
rect 182785 127882 228862 128118
rect 229098 127882 229182 128118
rect 229418 127882 229502 128118
rect 229738 127882 229822 128118
rect 230058 127882 230142 128118
rect 230378 127882 230462 128118
rect 230698 127882 230782 128118
rect 231018 127882 231102 128118
rect 231338 127882 231422 128118
rect 231658 127882 231742 128118
rect 231978 127882 232062 128118
rect 232298 127882 232382 128118
rect 232618 127882 237740 128118
rect 0 127840 237740 127882
rect 0 116918 237740 116960
rect 0 116682 122 116918
rect 358 116682 442 116918
rect 678 116682 762 116918
rect 998 116682 1082 116918
rect 1318 116682 1402 116918
rect 1638 116682 1722 116918
rect 1958 116682 2042 116918
rect 2278 116682 2362 116918
rect 2598 116682 2682 116918
rect 2918 116682 3002 116918
rect 3238 116682 3322 116918
rect 3558 116682 3642 116918
rect 3878 116682 43215 116918
rect 43451 116682 115215 116918
rect 115451 116682 187215 116918
rect 187451 116682 233862 116918
rect 234098 116682 234182 116918
rect 234418 116682 234502 116918
rect 234738 116682 234822 116918
rect 235058 116682 235142 116918
rect 235378 116682 235462 116918
rect 235698 116682 235782 116918
rect 236018 116682 236102 116918
rect 236338 116682 236422 116918
rect 236658 116682 236742 116918
rect 236978 116682 237062 116918
rect 237298 116682 237382 116918
rect 237618 116682 237740 116918
rect 0 116640 237740 116682
rect 31724 114002 58172 114044
rect 31724 113766 31766 114002
rect 32002 113766 56790 114002
rect 57026 113766 58172 114002
rect 31724 113724 58172 113766
rect 57852 113364 58172 113724
rect 57852 113322 72156 113364
rect 57852 113086 71878 113322
rect 72114 113086 72156 113322
rect 57852 113044 72156 113086
rect 0 105718 237740 105760
rect 0 105482 5122 105718
rect 5358 105482 5442 105718
rect 5678 105482 5762 105718
rect 5998 105482 6082 105718
rect 6318 105482 6402 105718
rect 6638 105482 6722 105718
rect 6958 105482 7042 105718
rect 7278 105482 7362 105718
rect 7598 105482 7682 105718
rect 7918 105482 8002 105718
rect 8238 105482 8322 105718
rect 8558 105482 8642 105718
rect 8878 105482 17549 105718
rect 17785 105482 42549 105718
rect 42785 105482 67146 105718
rect 67382 105482 114549 105718
rect 114785 105482 139146 105718
rect 139382 105482 186549 105718
rect 186785 105482 211549 105718
rect 211785 105482 228862 105718
rect 229098 105482 229182 105718
rect 229418 105482 229502 105718
rect 229738 105482 229822 105718
rect 230058 105482 230142 105718
rect 230378 105482 230462 105718
rect 230698 105482 230782 105718
rect 231018 105482 231102 105718
rect 231338 105482 231422 105718
rect 231658 105482 231742 105718
rect 231978 105482 232062 105718
rect 232298 105482 232382 105718
rect 232618 105482 237740 105718
rect 0 105440 237740 105482
rect 0 94518 237740 94560
rect 0 94282 122 94518
rect 358 94282 442 94518
rect 678 94282 762 94518
rect 998 94282 1082 94518
rect 1318 94282 1402 94518
rect 1638 94282 1722 94518
rect 1958 94282 2042 94518
rect 2278 94282 2362 94518
rect 2598 94282 2682 94518
rect 2918 94282 3002 94518
rect 3238 94282 3322 94518
rect 3558 94282 3642 94518
rect 3878 94282 20215 94518
rect 20451 94282 45215 94518
rect 45451 94282 82506 94518
rect 82742 94282 117215 94518
rect 117451 94282 154506 94518
rect 154742 94282 189215 94518
rect 189451 94282 214215 94518
rect 214451 94282 233862 94518
rect 234098 94282 234182 94518
rect 234418 94282 234502 94518
rect 234738 94282 234822 94518
rect 235058 94282 235142 94518
rect 235378 94282 235462 94518
rect 235698 94282 235782 94518
rect 236018 94282 236102 94518
rect 236338 94282 236422 94518
rect 236658 94282 236742 94518
rect 236978 94282 237062 94518
rect 237298 94282 237382 94518
rect 237618 94282 237740 94518
rect 0 94240 237740 94282
rect 0 83318 237740 83360
rect 0 83082 5122 83318
rect 5358 83082 5442 83318
rect 5678 83082 5762 83318
rect 5998 83082 6082 83318
rect 6318 83082 6402 83318
rect 6638 83082 6722 83318
rect 6958 83082 7042 83318
rect 7278 83082 7362 83318
rect 7598 83082 7682 83318
rect 7918 83082 8002 83318
rect 8238 83082 8322 83318
rect 8558 83082 8642 83318
rect 8878 83082 17549 83318
rect 17785 83082 42549 83318
rect 42785 83082 67146 83318
rect 67382 83082 114549 83318
rect 114785 83082 139146 83318
rect 139382 83082 186549 83318
rect 186785 83082 211549 83318
rect 211785 83082 228862 83318
rect 229098 83082 229182 83318
rect 229418 83082 229502 83318
rect 229738 83082 229822 83318
rect 230058 83082 230142 83318
rect 230378 83082 230462 83318
rect 230698 83082 230782 83318
rect 231018 83082 231102 83318
rect 231338 83082 231422 83318
rect 231658 83082 231742 83318
rect 231978 83082 232062 83318
rect 232298 83082 232382 83318
rect 232618 83082 237740 83318
rect 0 83040 237740 83082
rect 0 72118 237740 72160
rect 0 71882 122 72118
rect 358 71882 442 72118
rect 678 71882 762 72118
rect 998 71882 1082 72118
rect 1318 71882 1402 72118
rect 1638 71882 1722 72118
rect 1958 71882 2042 72118
rect 2278 71882 2362 72118
rect 2598 71882 2682 72118
rect 2918 71882 3002 72118
rect 3238 71882 3322 72118
rect 3558 71882 3642 72118
rect 3878 71882 233862 72118
rect 234098 71882 234182 72118
rect 234418 71882 234502 72118
rect 234738 71882 234822 72118
rect 235058 71882 235142 72118
rect 235378 71882 235462 72118
rect 235698 71882 235782 72118
rect 236018 71882 236102 72118
rect 236338 71882 236422 72118
rect 236658 71882 236742 72118
rect 236978 71882 237062 72118
rect 237298 71882 237382 72118
rect 237618 71882 237740 72118
rect 0 71840 237740 71882
rect 0 60918 237740 60960
rect 0 60682 5122 60918
rect 5358 60682 5442 60918
rect 5678 60682 5762 60918
rect 5998 60682 6082 60918
rect 6318 60682 6402 60918
rect 6638 60682 6722 60918
rect 6958 60682 7042 60918
rect 7278 60682 7362 60918
rect 7598 60682 7682 60918
rect 7918 60682 8002 60918
rect 8238 60682 8322 60918
rect 8558 60682 8642 60918
rect 8878 60682 38549 60918
rect 38785 60682 73882 60918
rect 74118 60682 110549 60918
rect 110785 60682 145882 60918
rect 146118 60682 182549 60918
rect 182785 60682 228862 60918
rect 229098 60682 229182 60918
rect 229418 60682 229502 60918
rect 229738 60682 229822 60918
rect 230058 60682 230142 60918
rect 230378 60682 230462 60918
rect 230698 60682 230782 60918
rect 231018 60682 231102 60918
rect 231338 60682 231422 60918
rect 231658 60682 231742 60918
rect 231978 60682 232062 60918
rect 232298 60682 232382 60918
rect 232618 60682 237740 60918
rect 0 60640 237740 60682
rect 0 49718 237740 49760
rect 0 49482 122 49718
rect 358 49482 442 49718
rect 678 49482 762 49718
rect 998 49482 1082 49718
rect 1318 49482 1402 49718
rect 1638 49482 1722 49718
rect 1958 49482 2042 49718
rect 2278 49482 2362 49718
rect 2598 49482 2682 49718
rect 2918 49482 3002 49718
rect 3238 49482 3322 49718
rect 3558 49482 3642 49718
rect 3878 49482 43215 49718
rect 43451 49482 78882 49718
rect 79118 49482 115215 49718
rect 115451 49482 150882 49718
rect 151118 49482 187215 49718
rect 187451 49482 233862 49718
rect 234098 49482 234182 49718
rect 234418 49482 234502 49718
rect 234738 49482 234822 49718
rect 235058 49482 235142 49718
rect 235378 49482 235462 49718
rect 235698 49482 235782 49718
rect 236018 49482 236102 49718
rect 236338 49482 236422 49718
rect 236658 49482 236742 49718
rect 236978 49482 237062 49718
rect 237298 49482 237382 49718
rect 237618 49482 237740 49718
rect 0 49440 237740 49482
rect 31724 41242 66452 41284
rect 31724 41006 31766 41242
rect 32002 41006 66174 41242
rect 66410 41006 66452 41242
rect 31724 40964 66452 41006
rect 93732 40562 108956 40604
rect 93732 40326 93774 40562
rect 94010 40326 108678 40562
rect 108914 40326 108956 40562
rect 93732 40284 108956 40326
rect 109556 40562 118708 40604
rect 109556 40326 109598 40562
rect 109834 40326 118708 40562
rect 109556 40284 118708 40326
rect 99252 38924 99756 40284
rect 118388 39244 118708 40284
rect 128508 40562 137108 40604
rect 128508 40326 129654 40562
rect 129890 40326 136830 40562
rect 137066 40326 137108 40562
rect 128508 40284 137108 40326
rect 171380 40562 190652 40604
rect 171380 40326 181358 40562
rect 181594 40326 190652 40562
rect 171380 40284 190652 40326
rect 128508 39244 128828 40284
rect 171380 39924 171700 40284
rect 166044 39882 171700 39924
rect 166044 39646 166086 39882
rect 166322 39646 171700 39882
rect 166044 39604 171700 39646
rect 118388 38924 128828 39244
rect 190332 39244 190652 40284
rect 190332 39202 201692 39244
rect 190332 38966 201414 39202
rect 201650 38966 201692 39202
rect 190332 38924 201692 38966
rect 0 38518 237740 38560
rect 0 38282 5122 38518
rect 5358 38282 5442 38518
rect 5678 38282 5762 38518
rect 5998 38282 6082 38518
rect 6318 38282 6402 38518
rect 6638 38282 6722 38518
rect 6958 38282 7042 38518
rect 7278 38282 7362 38518
rect 7598 38282 7682 38518
rect 7918 38282 8002 38518
rect 8238 38282 8322 38518
rect 8558 38282 8642 38518
rect 8878 38282 228862 38518
rect 229098 38282 229182 38518
rect 229418 38282 229502 38518
rect 229738 38282 229822 38518
rect 230058 38282 230142 38518
rect 230378 38282 230462 38518
rect 230698 38282 230782 38518
rect 231018 38282 231102 38518
rect 231338 38282 231422 38518
rect 231658 38282 231742 38518
rect 231978 38282 232062 38518
rect 232298 38282 232382 38518
rect 232618 38282 237740 38518
rect 0 38240 237740 38282
rect 0 27318 237740 27360
rect 0 27082 122 27318
rect 358 27082 442 27318
rect 678 27082 762 27318
rect 998 27082 1082 27318
rect 1318 27082 1402 27318
rect 1638 27082 1722 27318
rect 1958 27082 2042 27318
rect 2278 27082 2362 27318
rect 2598 27082 2682 27318
rect 2918 27082 3002 27318
rect 3238 27082 3322 27318
rect 3558 27082 3642 27318
rect 3878 27082 78882 27318
rect 79118 27082 150882 27318
rect 151118 27082 233862 27318
rect 234098 27082 234182 27318
rect 234418 27082 234502 27318
rect 234738 27082 234822 27318
rect 235058 27082 235142 27318
rect 235378 27082 235462 27318
rect 235698 27082 235782 27318
rect 236018 27082 236102 27318
rect 236338 27082 236422 27318
rect 236658 27082 236742 27318
rect 236978 27082 237062 27318
rect 237298 27082 237382 27318
rect 237618 27082 237740 27318
rect 0 27040 237740 27082
rect 0 16118 237740 16160
rect 0 15882 5122 16118
rect 5358 15882 5442 16118
rect 5678 15882 5762 16118
rect 5998 15882 6082 16118
rect 6318 15882 6402 16118
rect 6638 15882 6722 16118
rect 6958 15882 7042 16118
rect 7278 15882 7362 16118
rect 7598 15882 7682 16118
rect 7918 15882 8002 16118
rect 8238 15882 8322 16118
rect 8558 15882 8642 16118
rect 8878 15882 73882 16118
rect 74118 15882 145882 16118
rect 146118 15882 228862 16118
rect 229098 15882 229182 16118
rect 229418 15882 229502 16118
rect 229738 15882 229822 16118
rect 230058 15882 230142 16118
rect 230378 15882 230462 16118
rect 230698 15882 230782 16118
rect 231018 15882 231102 16118
rect 231338 15882 231422 16118
rect 231658 15882 231742 16118
rect 231978 15882 232062 16118
rect 232298 15882 232382 16118
rect 232618 15882 237740 16118
rect 0 15840 237740 15882
rect 5000 8878 232740 9000
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 228862 8878
rect 229098 8642 229182 8878
rect 229418 8642 229502 8878
rect 229738 8642 229822 8878
rect 230058 8642 230142 8878
rect 230378 8642 230462 8878
rect 230698 8642 230782 8878
rect 231018 8642 231102 8878
rect 231338 8642 231422 8878
rect 231658 8642 231742 8878
rect 231978 8642 232062 8878
rect 232298 8642 232382 8878
rect 232618 8642 232740 8878
rect 5000 8558 232740 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 228862 8558
rect 229098 8322 229182 8558
rect 229418 8322 229502 8558
rect 229738 8322 229822 8558
rect 230058 8322 230142 8558
rect 230378 8322 230462 8558
rect 230698 8322 230782 8558
rect 231018 8322 231102 8558
rect 231338 8322 231422 8558
rect 231658 8322 231742 8558
rect 231978 8322 232062 8558
rect 232298 8322 232382 8558
rect 232618 8322 232740 8558
rect 5000 8238 232740 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 228862 8238
rect 229098 8002 229182 8238
rect 229418 8002 229502 8238
rect 229738 8002 229822 8238
rect 230058 8002 230142 8238
rect 230378 8002 230462 8238
rect 230698 8002 230782 8238
rect 231018 8002 231102 8238
rect 231338 8002 231422 8238
rect 231658 8002 231742 8238
rect 231978 8002 232062 8238
rect 232298 8002 232382 8238
rect 232618 8002 232740 8238
rect 5000 7918 232740 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 228862 7918
rect 229098 7682 229182 7918
rect 229418 7682 229502 7918
rect 229738 7682 229822 7918
rect 230058 7682 230142 7918
rect 230378 7682 230462 7918
rect 230698 7682 230782 7918
rect 231018 7682 231102 7918
rect 231338 7682 231422 7918
rect 231658 7682 231742 7918
rect 231978 7682 232062 7918
rect 232298 7682 232382 7918
rect 232618 7682 232740 7918
rect 5000 7598 232740 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 228862 7598
rect 229098 7362 229182 7598
rect 229418 7362 229502 7598
rect 229738 7362 229822 7598
rect 230058 7362 230142 7598
rect 230378 7362 230462 7598
rect 230698 7362 230782 7598
rect 231018 7362 231102 7598
rect 231338 7362 231422 7598
rect 231658 7362 231742 7598
rect 231978 7362 232062 7598
rect 232298 7362 232382 7598
rect 232618 7362 232740 7598
rect 5000 7278 232740 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 228862 7278
rect 229098 7042 229182 7278
rect 229418 7042 229502 7278
rect 229738 7042 229822 7278
rect 230058 7042 230142 7278
rect 230378 7042 230462 7278
rect 230698 7042 230782 7278
rect 231018 7042 231102 7278
rect 231338 7042 231422 7278
rect 231658 7042 231742 7278
rect 231978 7042 232062 7278
rect 232298 7042 232382 7278
rect 232618 7042 232740 7278
rect 5000 6958 232740 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 228862 6958
rect 229098 6722 229182 6958
rect 229418 6722 229502 6958
rect 229738 6722 229822 6958
rect 230058 6722 230142 6958
rect 230378 6722 230462 6958
rect 230698 6722 230782 6958
rect 231018 6722 231102 6958
rect 231338 6722 231422 6958
rect 231658 6722 231742 6958
rect 231978 6722 232062 6958
rect 232298 6722 232382 6958
rect 232618 6722 232740 6958
rect 5000 6638 232740 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 228862 6638
rect 229098 6402 229182 6638
rect 229418 6402 229502 6638
rect 229738 6402 229822 6638
rect 230058 6402 230142 6638
rect 230378 6402 230462 6638
rect 230698 6402 230782 6638
rect 231018 6402 231102 6638
rect 231338 6402 231422 6638
rect 231658 6402 231742 6638
rect 231978 6402 232062 6638
rect 232298 6402 232382 6638
rect 232618 6402 232740 6638
rect 5000 6318 232740 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 228862 6318
rect 229098 6082 229182 6318
rect 229418 6082 229502 6318
rect 229738 6082 229822 6318
rect 230058 6082 230142 6318
rect 230378 6082 230462 6318
rect 230698 6082 230782 6318
rect 231018 6082 231102 6318
rect 231338 6082 231422 6318
rect 231658 6082 231742 6318
rect 231978 6082 232062 6318
rect 232298 6082 232382 6318
rect 232618 6082 232740 6318
rect 5000 5998 232740 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 228862 5998
rect 229098 5762 229182 5998
rect 229418 5762 229502 5998
rect 229738 5762 229822 5998
rect 230058 5762 230142 5998
rect 230378 5762 230462 5998
rect 230698 5762 230782 5998
rect 231018 5762 231102 5998
rect 231338 5762 231422 5998
rect 231658 5762 231742 5998
rect 231978 5762 232062 5998
rect 232298 5762 232382 5998
rect 232618 5762 232740 5998
rect 5000 5678 232740 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 228862 5678
rect 229098 5442 229182 5678
rect 229418 5442 229502 5678
rect 229738 5442 229822 5678
rect 230058 5442 230142 5678
rect 230378 5442 230462 5678
rect 230698 5442 230782 5678
rect 231018 5442 231102 5678
rect 231338 5442 231422 5678
rect 231658 5442 231742 5678
rect 231978 5442 232062 5678
rect 232298 5442 232382 5678
rect 232618 5442 232740 5678
rect 5000 5358 232740 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 228862 5358
rect 229098 5122 229182 5358
rect 229418 5122 229502 5358
rect 229738 5122 229822 5358
rect 230058 5122 230142 5358
rect 230378 5122 230462 5358
rect 230698 5122 230782 5358
rect 231018 5122 231102 5358
rect 231338 5122 231422 5358
rect 231658 5122 231742 5358
rect 231978 5122 232062 5358
rect 232298 5122 232382 5358
rect 232618 5122 232740 5358
rect 5000 5000 232740 5122
rect 0 3878 237740 4000
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 233862 3878
rect 234098 3642 234182 3878
rect 234418 3642 234502 3878
rect 234738 3642 234822 3878
rect 235058 3642 235142 3878
rect 235378 3642 235462 3878
rect 235698 3642 235782 3878
rect 236018 3642 236102 3878
rect 236338 3642 236422 3878
rect 236658 3642 236742 3878
rect 236978 3642 237062 3878
rect 237298 3642 237382 3878
rect 237618 3642 237740 3878
rect 0 3558 237740 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 233862 3558
rect 234098 3322 234182 3558
rect 234418 3322 234502 3558
rect 234738 3322 234822 3558
rect 235058 3322 235142 3558
rect 235378 3322 235462 3558
rect 235698 3322 235782 3558
rect 236018 3322 236102 3558
rect 236338 3322 236422 3558
rect 236658 3322 236742 3558
rect 236978 3322 237062 3558
rect 237298 3322 237382 3558
rect 237618 3322 237740 3558
rect 0 3238 237740 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 233862 3238
rect 234098 3002 234182 3238
rect 234418 3002 234502 3238
rect 234738 3002 234822 3238
rect 235058 3002 235142 3238
rect 235378 3002 235462 3238
rect 235698 3002 235782 3238
rect 236018 3002 236102 3238
rect 236338 3002 236422 3238
rect 236658 3002 236742 3238
rect 236978 3002 237062 3238
rect 237298 3002 237382 3238
rect 237618 3002 237740 3238
rect 0 2918 237740 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 233862 2918
rect 234098 2682 234182 2918
rect 234418 2682 234502 2918
rect 234738 2682 234822 2918
rect 235058 2682 235142 2918
rect 235378 2682 235462 2918
rect 235698 2682 235782 2918
rect 236018 2682 236102 2918
rect 236338 2682 236422 2918
rect 236658 2682 236742 2918
rect 236978 2682 237062 2918
rect 237298 2682 237382 2918
rect 237618 2682 237740 2918
rect 0 2598 237740 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 233862 2598
rect 234098 2362 234182 2598
rect 234418 2362 234502 2598
rect 234738 2362 234822 2598
rect 235058 2362 235142 2598
rect 235378 2362 235462 2598
rect 235698 2362 235782 2598
rect 236018 2362 236102 2598
rect 236338 2362 236422 2598
rect 236658 2362 236742 2598
rect 236978 2362 237062 2598
rect 237298 2362 237382 2598
rect 237618 2362 237740 2598
rect 0 2278 237740 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 233862 2278
rect 234098 2042 234182 2278
rect 234418 2042 234502 2278
rect 234738 2042 234822 2278
rect 235058 2042 235142 2278
rect 235378 2042 235462 2278
rect 235698 2042 235782 2278
rect 236018 2042 236102 2278
rect 236338 2042 236422 2278
rect 236658 2042 236742 2278
rect 236978 2042 237062 2278
rect 237298 2042 237382 2278
rect 237618 2042 237740 2278
rect 0 1958 237740 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 233862 1958
rect 234098 1722 234182 1958
rect 234418 1722 234502 1958
rect 234738 1722 234822 1958
rect 235058 1722 235142 1958
rect 235378 1722 235462 1958
rect 235698 1722 235782 1958
rect 236018 1722 236102 1958
rect 236338 1722 236422 1958
rect 236658 1722 236742 1958
rect 236978 1722 237062 1958
rect 237298 1722 237382 1958
rect 237618 1722 237740 1958
rect 0 1638 237740 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 233862 1638
rect 234098 1402 234182 1638
rect 234418 1402 234502 1638
rect 234738 1402 234822 1638
rect 235058 1402 235142 1638
rect 235378 1402 235462 1638
rect 235698 1402 235782 1638
rect 236018 1402 236102 1638
rect 236338 1402 236422 1638
rect 236658 1402 236742 1638
rect 236978 1402 237062 1638
rect 237298 1402 237382 1638
rect 237618 1402 237740 1638
rect 0 1318 237740 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 233862 1318
rect 234098 1082 234182 1318
rect 234418 1082 234502 1318
rect 234738 1082 234822 1318
rect 235058 1082 235142 1318
rect 235378 1082 235462 1318
rect 235698 1082 235782 1318
rect 236018 1082 236102 1318
rect 236338 1082 236422 1318
rect 236658 1082 236742 1318
rect 236978 1082 237062 1318
rect 237298 1082 237382 1318
rect 237618 1082 237740 1318
rect 0 998 237740 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 233862 998
rect 234098 762 234182 998
rect 234418 762 234502 998
rect 234738 762 234822 998
rect 235058 762 235142 998
rect 235378 762 235462 998
rect 235698 762 235782 998
rect 236018 762 236102 998
rect 236338 762 236422 998
rect 236658 762 236742 998
rect 236978 762 237062 998
rect 237298 762 237382 998
rect 237618 762 237740 998
rect 0 678 237740 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 233862 678
rect 234098 442 234182 678
rect 234418 442 234502 678
rect 234738 442 234822 678
rect 235058 442 235142 678
rect 235378 442 235462 678
rect 235698 442 235782 678
rect 236018 442 236102 678
rect 236338 442 236422 678
rect 236658 442 236742 678
rect 236978 442 237062 678
rect 237298 442 237382 678
rect 237618 442 237740 678
rect 0 358 237740 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 233862 358
rect 234098 122 234182 358
rect 234418 122 234502 358
rect 234738 122 234822 358
rect 235058 122 235142 358
rect 235378 122 235462 358
rect 235698 122 235782 358
rect 236018 122 236102 358
rect 236338 122 236422 358
rect 236658 122 236742 358
rect 236978 122 237062 358
rect 237298 122 237382 358
rect 237618 122 237740 358
rect 0 0 237740 122
use sb_0__0_  sb_0__0_
timestamp 1604441278
transform 1 0 32896 0 1 39824
box 0 0 28000 27720
use grid_io_bottom  grid_io_bottom_1__0_
timestamp 1604441278
transform 1 0 67896 0 1 12824
box 0 0 28926 24000
use cbx_1__0_  cbx_1__0_
timestamp 1604441278
transform 1 0 67896 0 1 41824
box 0 0 30000 24000
use sb_1__0_  sb_1__0_
timestamp 1604441278
transform 1 0 104896 0 1 39824
box 0 0 28000 28000
use grid_io_bottom  grid_io_bottom_2__0_
timestamp 1604441278
transform 1 0 139896 0 1 12824
box 0 0 28926 24000
use cbx_1__0_  cbx_2__0_
timestamp 1604441278
transform 1 0 139896 0 1 41824
box 0 0 30000 24000
use sb_2__0_  sb_2__0_
timestamp 1604441278
transform 1 0 176896 0 1 39824
box 0 0 27678 28000
use grid_io_left  grid_io_left_0__1_
timestamp 1604441278
transform 1 0 13896 0 1 70824
box 0 0 16000 37584
use cby_0__1_  cby_0__1_
timestamp 1604441278
transform 1 0 38896 0 1 70824
box 0 0 16000 40000
use grid_clb  grid_clb_1__1_
timestamp 1604441278
transform 1 0 62896 0 1 70824
box 0 0 40000 39432
use cby_1__1_  cby_1__1_
timestamp 1604441278
transform 1 0 110896 0 1 70824
box 0 0 16000 40000
use grid_clb  grid_clb_2__1_
timestamp 1604441278
transform 1 0 134896 0 1 70824
box 0 0 40000 39432
use grid_io_right  grid_io_right_3__1_
timestamp 1604441278
transform 1 0 207896 0 1 70824
box 0 0 16000 37584
use cby_1__1_  cby_2__1_
timestamp 1604441278
transform 1 0 182896 0 1 70824
box 0 0 16000 40000
use grid_io_left  grid_io_left_0__2_
timestamp 1604441278
transform 1 0 13896 0 1 144824
box 0 0 16000 37584
use sb_0__1_  sb_0__1_
timestamp 1604441278
transform 1 0 32896 0 1 113824
box 0 0 28000 28000
use cby_0__1_  cby_0__2_
timestamp 1604441278
transform 1 0 38896 0 1 144824
box 0 0 16000 40000
use grid_clb  grid_clb_1__2_
timestamp 1604441278
transform 1 0 62896 0 1 144824
box 0 0 40000 39432
use cbx_1__1_  cbx_1__1_
timestamp 1604441278
transform 1 0 67896 0 1 115824
box 0 0 30000 24000
use sb_1__1_  sb_1__1_
timestamp 1604441278
transform 1 0 104896 0 1 113824
box 0 0 28000 28000
use cby_1__1_  cby_1__2_
timestamp 1604441278
transform 1 0 110896 0 1 144824
box 0 0 16000 40000
use grid_clb  grid_clb_2__2_
timestamp 1604441278
transform 1 0 134896 0 1 144824
box 0 0 40000 39432
use cbx_1__1_  cbx_2__1_
timestamp 1604441278
transform 1 0 139896 0 1 115824
box 0 0 30000 24000
use grid_io_right  grid_io_right_3__2_
timestamp 1604441278
transform 1 0 207896 0 1 144824
box 0 0 16000 37584
use sb_2__1_  sb_2__1_
timestamp 1604441278
transform 1 0 176896 0 1 113824
box 0 0 28000 28000
use cby_1__1_  cby_2__2_
timestamp 1604441278
transform 1 0 182896 0 1 144824
box 0 0 16000 40000
use sb_0__2_  sb_0__2_
timestamp 1604441278
transform 1 0 32895 0 1 187824
box 1 0 27712 28000
use cbx_1__2_  cbx_1__2_
timestamp 1604441278
transform 1 0 67896 0 1 189823
box 0 1 30000 23970
use sb_1__2_  sb_1__2_
timestamp 1604441278
transform 1 0 104896 0 1 187824
box 0 0 28000 28000
use cbx_1__2_  cbx_2__2_
timestamp 1604441278
transform 1 0 139896 0 1 189823
box 0 1 30000 23970
use sb_2__2_  sb_2__2_
timestamp 1604441278
transform 1 0 176896 0 1 187824
box 0 0 28000 27600
use grid_io_top  grid_io_top_1__3_
timestamp 1604441278
transform 1 0 67896 0 1 218824
box 0 0 28934 24000
use grid_io_top  grid_io_top_2__3_
timestamp 1604441278
transform 1 0 139896 0 1 218824
box 0 0 28934 24000
<< labels >>
rlabel metal3 s 9896 214192 10376 214312 6 Test_en
port 0 nsew default input
rlabel metal3 s 227416 211064 227896 211184 6 ccff_head
port 1 nsew default input
rlabel metal3 s 9896 19576 10376 19696 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 9896 235816 10376 235936 6 clk
port 3 nsew default input
rlabel metal2 s 23530 246344 23586 246824 6 gfpga_pad_GPIO_A[0]
port 4 nsew default tristate
rlabel metal2 s 50762 246344 50818 246824 6 gfpga_pad_GPIO_A[1]
port 5 nsew default tristate
rlabel metal3 s 227416 20664 227896 20784 6 gfpga_pad_GPIO_A[2]
port 6 nsew default tristate
rlabel metal3 s 227416 44464 227896 44584 6 gfpga_pad_GPIO_A[3]
port 7 nsew default tristate
rlabel metal2 s 23530 8824 23586 9304 6 gfpga_pad_GPIO_A[4]
port 8 nsew default tristate
rlabel metal2 s 50762 8824 50818 9304 6 gfpga_pad_GPIO_A[5]
port 9 nsew default tristate
rlabel metal3 s 9896 41200 10376 41320 6 gfpga_pad_GPIO_A[6]
port 10 nsew default tristate
rlabel metal3 s 9896 62824 10376 62944 6 gfpga_pad_GPIO_A[7]
port 11 nsew default tristate
rlabel metal2 s 77994 246344 78050 246824 6 gfpga_pad_GPIO_IE[0]
port 12 nsew default tristate
rlabel metal2 s 105226 246344 105282 246824 6 gfpga_pad_GPIO_IE[1]
port 13 nsew default tristate
rlabel metal3 s 227416 68264 227896 68384 6 gfpga_pad_GPIO_IE[2]
port 14 nsew default tristate
rlabel metal3 s 227416 92064 227896 92184 6 gfpga_pad_GPIO_IE[3]
port 15 nsew default tristate
rlabel metal2 s 77994 8824 78050 9304 6 gfpga_pad_GPIO_IE[4]
port 16 nsew default tristate
rlabel metal2 s 105226 8824 105282 9304 6 gfpga_pad_GPIO_IE[5]
port 17 nsew default tristate
rlabel metal3 s 9896 84448 10376 84568 6 gfpga_pad_GPIO_IE[6]
port 18 nsew default tristate
rlabel metal3 s 9896 106072 10376 106192 6 gfpga_pad_GPIO_IE[7]
port 19 nsew default tristate
rlabel metal2 s 132550 246344 132606 246824 6 gfpga_pad_GPIO_OE[0]
port 20 nsew default tristate
rlabel metal2 s 159782 246344 159838 246824 6 gfpga_pad_GPIO_OE[1]
port 21 nsew default tristate
rlabel metal3 s 227416 115864 227896 115984 6 gfpga_pad_GPIO_OE[2]
port 22 nsew default tristate
rlabel metal3 s 227416 139664 227896 139784 6 gfpga_pad_GPIO_OE[3]
port 23 nsew default tristate
rlabel metal2 s 132550 8824 132606 9304 6 gfpga_pad_GPIO_OE[4]
port 24 nsew default tristate
rlabel metal2 s 159782 8824 159838 9304 6 gfpga_pad_GPIO_OE[5]
port 25 nsew default tristate
rlabel metal3 s 9896 127696 10376 127816 6 gfpga_pad_GPIO_OE[6]
port 26 nsew default tristate
rlabel metal3 s 9896 149320 10376 149440 6 gfpga_pad_GPIO_OE[7]
port 27 nsew default tristate
rlabel metal2 s 187014 246344 187070 246824 6 gfpga_pad_GPIO_Y[0]
port 28 nsew default bidirectional
rlabel metal2 s 214246 246344 214302 246824 6 gfpga_pad_GPIO_Y[1]
port 29 nsew default bidirectional
rlabel metal3 s 227416 163464 227896 163584 6 gfpga_pad_GPIO_Y[2]
port 30 nsew default bidirectional
rlabel metal3 s 227416 187264 227896 187384 6 gfpga_pad_GPIO_Y[3]
port 31 nsew default bidirectional
rlabel metal2 s 187014 8824 187070 9304 6 gfpga_pad_GPIO_Y[4]
port 32 nsew default bidirectional
rlabel metal2 s 214246 8824 214302 9304 6 gfpga_pad_GPIO_Y[5]
port 33 nsew default bidirectional
rlabel metal3 s 9896 170944 10376 171064 6 gfpga_pad_GPIO_Y[6]
port 34 nsew default bidirectional
rlabel metal3 s 9896 192568 10376 192688 6 gfpga_pad_GPIO_Y[7]
port 35 nsew default bidirectional
rlabel metal3 s 227416 234864 227896 234984 6 prog_clk
port 36 nsew default input
rlabel metal5 s 5000 5000 232740 9000 8 vpwr
port 37 nsew default input
rlabel metal5 s 0 0 237740 4000 8 vgnd
port 38 nsew default input
<< properties >>
string FIXED_BBOX 0 0 237740 255376
<< end >>
