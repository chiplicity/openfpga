* NGSPICE file created from cby_0__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

.subckt cby_0__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_grid_pin_0_ left_grid_pin_10_ left_grid_pin_12_ left_grid_pin_14_ left_grid_pin_2_
+ left_grid_pin_4_ left_grid_pin_6_ left_grid_pin_8_ right_grid_pin_3_ right_grid_pin_7_
+ vpwr vgnd
XFILLER_26_41 vpwr vgnd scs8hd_fill_2
XANTENNA__113__B _116_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[5] mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_29 vgnd vpwr scs8hd_decap_4
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XFILLER_10_125 vgnd vpwr scs8hd_decap_12
XFILLER_37_40 vpwr vgnd scs8hd_fill_2
XFILLER_37_95 vgnd vpwr scs8hd_fill_1
XANTENNA__108__B _108_/B vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _124_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_2_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_062_ address[1] address[2] address[0] _062_/X vgnd vpwr scs8hd_or3_4
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_23_86 vpwr vgnd scs8hd_fill_2
X_131_ _139_/A _131_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_48_61 vpwr vgnd scs8hd_fill_2
XFILLER_2_143 vgnd vpwr scs8hd_decap_3
XANTENNA__110__C _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_88 vgnd vpwr scs8hd_decap_4
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
XFILLER_56_117 vgnd vpwr scs8hd_decap_12
XFILLER_18_64 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_0_.latch/Q mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_30 vgnd vpwr scs8hd_fill_1
XFILLER_34_85 vgnd vpwr scs8hd_decap_6
X_114_ _122_/A _116_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_59_82 vpwr vgnd scs8hd_fill_2
XFILLER_38_106 vgnd vpwr scs8hd_decap_4
XANTENNA__121__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_19 vpwr vgnd scs8hd_fill_2
XFILLER_44_109 vgnd vpwr scs8hd_decap_12
XFILLER_29_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_2.LATCH_1_.latch data_in mem_right_ipin_2.LATCH_1_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_10 vpwr vgnd scs8hd_fill_2
XFILLER_20_43 vpwr vgnd scs8hd_fill_2
XFILLER_29_30 vpwr vgnd scs8hd_fill_2
XFILLER_45_62 vpwr vgnd scs8hd_fill_2
XANTENNA__116__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XFILLER_6_78 vgnd vpwr scs8hd_fill_1
XFILLER_6_45 vgnd vpwr scs8hd_decap_8
XANTENNA__132__A _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_4.LATCH_4_.latch data_in mem_right_ipin_4.LATCH_4_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_109 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_31_42 vpwr vgnd scs8hd_fill_2
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_4.LATCH_4_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__127__A address[5] vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_134 vgnd vpwr scs8hd_decap_12
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_105 vgnd vpwr scs8hd_decap_4
XFILLER_13_112 vgnd vpwr scs8hd_decap_8
XFILLER_13_123 vpwr vgnd scs8hd_fill_2
XFILLER_13_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_64 vpwr vgnd scs8hd_fill_2
XFILLER_26_75 vpwr vgnd scs8hd_fill_2
XFILLER_26_86 vgnd vpwr scs8hd_decap_3
XFILLER_42_85 vgnd vpwr scs8hd_decap_6
XFILLER_42_41 vpwr vgnd scs8hd_fill_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XFILLER_10_137 vgnd vpwr scs8hd_decap_8
XFILLER_53_62 vgnd vpwr scs8hd_decap_12
XFILLER_53_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _175_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__124__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _140_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_32 vgnd vpwr scs8hd_fill_1
X_130_ _138_/A _131_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_65 vpwr vgnd scs8hd_fill_2
XFILLER_48_40 vgnd vpwr scs8hd_fill_1
XFILLER_64_94 vgnd vpwr scs8hd_decap_12
XFILLER_0_47 vpwr vgnd scs8hd_fill_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XFILLER_9_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.LATCH_5_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__135__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_43_3 vpwr vgnd scs8hd_fill_2
XFILLER_56_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _145_/A mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_21 vpwr vgnd scs8hd_fill_2
XFILLER_18_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_113_ _121_/A _116_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_64 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_5.LATCH_0_.latch data_in mem_right_ipin_5.LATCH_0_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_61_143 vgnd vpwr scs8hd_decap_3
XFILLER_61_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_77 vpwr vgnd scs8hd_fill_2
XFILLER_45_85 vpwr vgnd scs8hd_fill_2
XFILLER_43_143 vgnd vpwr scs8hd_decap_3
XFILLER_43_121 vgnd vpwr scs8hd_fill_1
XFILLER_61_62 vgnd vpwr scs8hd_decap_12
XFILLER_61_51 vgnd vpwr scs8hd_decap_8
Xmem_right_ipin_7.LATCH_3_.latch data_in mem_right_ipin_7.LATCH_3_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_57 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__132__B _131_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_102 vgnd vpwr scs8hd_decap_8
XFILLER_25_121 vgnd vpwr scs8hd_fill_1
XFILLER_31_21 vpwr vgnd scs8hd_fill_2
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_113 vpwr vgnd scs8hd_fill_2
XANTENNA__143__A _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_102 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_4
XFILLER_42_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_47 vpwr vgnd scs8hd_fill_2
XFILLER_3_14 vpwr vgnd scs8hd_fill_2
XANTENNA__138__A _138_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_0_.latch/Q mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_45 vgnd vpwr scs8hd_fill_1
XFILLER_37_75 vpwr vgnd scs8hd_fill_2
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
XFILLER_53_74 vgnd vpwr scs8hd_decap_12
XFILLER_38_6 vgnd vpwr scs8hd_decap_4
XANTENNA__140__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_11 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_101 vgnd vpwr scs8hd_decap_8
XFILLER_48_96 vgnd vpwr scs8hd_decap_3
X_189_ chany_bottom_in[8] chany_top_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__135__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA__151__A _137_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_108 vgnd vpwr scs8hd_decap_12
XFILLER_34_21 vpwr vgnd scs8hd_fill_2
XFILLER_34_43 vpwr vgnd scs8hd_fill_2
X_112_ _112_/A _116_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_59_73 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_0.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[2] mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__146__A _146_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_7_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_20_89 vgnd vpwr scs8hd_fill_1
XFILLER_28_130 vgnd vpwr scs8hd_decap_12
XFILLER_45_53 vpwr vgnd scs8hd_fill_2
XFILLER_61_74 vgnd vpwr scs8hd_decap_12
XFILLER_20_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.LATCH_5_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_130 vgnd vpwr scs8hd_decap_4
XFILLER_19_141 vgnd vpwr scs8hd_decap_4
XFILLER_40_114 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_45 vpwr vgnd scs8hd_fill_2
XFILLER_15_56 vgnd vpwr scs8hd_decap_3
XFILLER_31_88 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__127__C _154_/C vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _143_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_125 vpwr vgnd scs8hd_fill_2
XFILLER_26_22 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_0.LATCH_4_.latch data_in mem_right_ipin_0.LATCH_4_.latch/Q _072_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__138__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__154__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_8_140 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_ipin_0.LATCH_3_.latch/Q mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_10_106 vgnd vpwr scs8hd_decap_4
XFILLER_12_24 vgnd vpwr scs8hd_decap_3
XFILLER_12_68 vgnd vpwr scs8hd_fill_1
XANTENNA__064__A _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_53_86 vgnd vpwr scs8hd_decap_12
XFILLER_5_121 vgnd vpwr scs8hd_fill_1
XFILLER_5_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _176_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__149__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_59_139 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_135 vgnd vpwr scs8hd_decap_8
XFILLER_2_124 vgnd vpwr scs8hd_decap_8
XFILLER_2_113 vgnd vpwr scs8hd_decap_8
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_58 vgnd vpwr scs8hd_decap_3
XANTENNA__135__C _066_/C vgnd vpwr scs8hd_diode_2
X_188_ chany_top_in[0] chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_3
XFILLER_34_77 vpwr vgnd scs8hd_fill_2
XFILLER_50_32 vgnd vpwr scs8hd_decap_12
X_111_ _110_/X _116_/B vgnd vpwr scs8hd_buf_1
XFILLER_59_41 vpwr vgnd scs8hd_fill_2
XFILLER_61_123 vgnd vpwr scs8hd_decap_12
XANTENNA__162__A _161_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_120 vpwr vgnd scs8hd_fill_2
XFILLER_29_109 vpwr vgnd scs8hd_fill_2
XFILLER_52_145 vgnd vpwr scs8hd_fill_1
XANTENNA__072__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_11 vpwr vgnd scs8hd_fill_2
XFILLER_45_21 vpwr vgnd scs8hd_fill_2
XFILLER_43_123 vgnd vpwr scs8hd_decap_12
XFILLER_43_101 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_142 vgnd vpwr scs8hd_decap_4
XFILLER_29_88 vgnd vpwr scs8hd_decap_4
XFILLER_61_86 vgnd vpwr scs8hd_decap_12
XFILLER_45_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_0_.latch/Q mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__157__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_34_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_1.LATCH_0_.latch data_in mem_right_ipin_1.LATCH_0_.latch/Q _089_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_123 vpwr vgnd scs8hd_fill_2
XFILLER_40_126 vgnd vpwr scs8hd_decap_12
XANTENNA__067__A _066_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_24 vpwr vgnd scs8hd_fill_2
XFILLER_15_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_145 vgnd vpwr scs8hd_fill_1
XFILLER_16_145 vgnd vpwr scs8hd_fill_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_126 vpwr vgnd scs8hd_fill_2
XANTENNA__143__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_1_.latch/Q mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_ipin_3.LATCH_3_.latch data_in mem_right_ipin_3.LATCH_3_.latch/Q _106_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_45 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_11 vgnd vpwr scs8hd_fill_1
XFILLER_3_27 vpwr vgnd scs8hd_fill_2
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XANTENNA__154__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__064__B _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA__080__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_58 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_5.INVTX1_3_.scs8hd_inv_1 chany_top_in[6] mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_44 vgnd vpwr scs8hd_decap_3
XFILLER_37_22 vgnd vpwr scs8hd_decap_3
XFILLER_37_11 vgnd vpwr scs8hd_fill_1
XFILLER_37_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_81 vpwr vgnd scs8hd_fill_2
XFILLER_23_24 vpwr vgnd scs8hd_fill_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XANTENNA__075__A _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_32 vgnd vpwr scs8hd_decap_8
XFILLER_48_65 vpwr vgnd scs8hd_fill_2
XFILLER_64_75 vgnd vpwr scs8hd_decap_12
XFILLER_9_48 vgnd vpwr scs8hd_decap_4
XANTENNA__135__D _143_/B vgnd vpwr scs8hd_diode_2
X_187_ chany_top_in[1] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_0.LATCH_4_.latch data_in mem_left_ipin_0.LATCH_4_.latch/Q _159_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_143 vgnd vpwr scs8hd_decap_3
XFILLER_55_110 vgnd vpwr scs8hd_decap_12
X_110_ _110_/A address[3] _102_/A _110_/X vgnd vpwr scs8hd_or3_4
XFILLER_50_44 vgnd vpwr scs8hd_decap_8
XFILLER_59_97 vpwr vgnd scs8hd_fill_2
XFILLER_59_86 vgnd vpwr scs8hd_decap_6
XFILLER_61_135 vgnd vpwr scs8hd_decap_8
XFILLER_41_3 vgnd vpwr scs8hd_decap_3
XFILLER_37_143 vgnd vpwr scs8hd_decap_3
XFILLER_1_71 vpwr vgnd scs8hd_fill_2
XANTENNA__072__B _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_47 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_29_34 vpwr vgnd scs8hd_fill_2
XFILLER_45_66 vpwr vgnd scs8hd_fill_2
XFILLER_45_11 vgnd vpwr scs8hd_decap_3
XFILLER_43_135 vgnd vpwr scs8hd_decap_8
XFILLER_43_113 vgnd vpwr scs8hd_decap_8
XFILLER_61_98 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_7 vgnd vpwr scs8hd_fill_1
XANTENNA__157__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_102 vpwr vgnd scs8hd_fill_2
XFILLER_34_113 vgnd vpwr scs8hd_decap_12
XFILLER_25_102 vgnd vpwr scs8hd_decap_4
XFILLER_25_113 vpwr vgnd scs8hd_fill_2
XFILLER_40_138 vgnd vpwr scs8hd_decap_8
XANTENNA__083__A _082_/X vgnd vpwr scs8hd_diode_2
XFILLER_31_46 vpwr vgnd scs8hd_fill_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_6.LATCH_2_.latch data_in mem_right_ipin_6.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_32 vgnd vpwr scs8hd_decap_12
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_102 vgnd vpwr scs8hd_decap_8
XFILLER_16_113 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_105 vpwr vgnd scs8hd_fill_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _167_/X vgnd vpwr scs8hd_diode_2
XANTENNA__078__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_105 vgnd vpwr scs8hd_decap_4
XFILLER_13_127 vgnd vpwr scs8hd_decap_12
XFILLER_26_79 vgnd vpwr scs8hd_decap_4
XFILLER_42_45 vgnd vpwr scs8hd_decap_4
XFILLER_42_23 vpwr vgnd scs8hd_fill_2
XFILLER_9_109 vgnd vpwr scs8hd_fill_1
XANTENNA__154__C _154_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_48 vgnd vpwr scs8hd_fill_1
XANTENNA__080__B _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_1.LATCH_0_.latch data_in _146_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _177_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__149__C _161_/C vgnd vpwr scs8hd_diode_2
XANTENNA__181__A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_2.LATCH_2_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_23_69 vpwr vgnd scs8hd_fill_2
XFILLER_58_141 vgnd vpwr scs8hd_decap_4
XFILLER_48_44 vpwr vgnd scs8hd_fill_2
XFILLER_64_87 vgnd vpwr scs8hd_decap_6
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_0_.latch/Q mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_27 vpwr vgnd scs8hd_fill_2
X_186_ chany_top_in[2] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
Xmux_right_ipin_3.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_25 vgnd vpwr scs8hd_decap_4
XFILLER_18_47 vpwr vgnd scs8hd_fill_2
XANTENNA__086__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_50_89 vgnd vpwr scs8hd_decap_3
XFILLER_50_78 vgnd vpwr scs8hd_fill_1
XFILLER_1_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
X_169_ _169_/A _141_/A _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XFILLER_45_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_100 vpwr vgnd scs8hd_fill_2
XFILLER_19_111 vpwr vgnd scs8hd_fill_2
XANTENNA__157__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_125 vgnd vpwr scs8hd_decap_12
XFILLER_31_25 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB _074_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_69 vpwr vgnd scs8hd_fill_2
XFILLER_56_44 vgnd vpwr scs8hd_decap_12
XPHY_120 vgnd vpwr scs8hd_decap_3
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vgnd vpwr scs8hd_decap_12
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_117 vgnd vpwr scs8hd_decap_4
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__184__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_7_82 vpwr vgnd scs8hd_fill_2
XANTENNA__078__B _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_139 vgnd vpwr scs8hd_decap_6
XANTENNA__094__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_58 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _146_/A mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XANTENNA__089__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_135 vgnd vpwr scs8hd_decap_8
XFILLER_5_113 vgnd vpwr scs8hd_decap_8
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XANTENNA__091__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_48_78 vgnd vpwr scs8hd_decap_12
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
X_185_ chany_top_in[3] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_13_92 vgnd vpwr scs8hd_fill_1
XFILLER_64_145 vgnd vpwr scs8hd_fill_1
XFILLER_49_120 vpwr vgnd scs8hd_fill_2
XANTENNA__192__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_55_123 vgnd vpwr scs8hd_decap_12
XANTENNA__086__B _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_25 vgnd vpwr scs8hd_decap_3
XFILLER_34_47 vpwr vgnd scs8hd_fill_2
XFILLER_59_77 vgnd vpwr scs8hd_fill_1
XFILLER_59_66 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_145 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_ipin_7.LATCH_3_.latch/Q mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_40_90 vpwr vgnd scs8hd_fill_2
XFILLER_24_80 vpwr vgnd scs8hd_fill_2
XFILLER_24_91 vgnd vpwr scs8hd_fill_1
X_168_ _167_/X _141_/A vgnd vpwr scs8hd_buf_1
X_099_ _091_/A address[6] _066_/C _102_/A vgnd vpwr scs8hd_or3_4
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_37_112 vgnd vpwr scs8hd_decap_8
XANTENNA__187__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.INVTX1_3_.scs8hd_inv_1 chany_top_in[3] mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_2_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XFILLER_29_47 vpwr vgnd scs8hd_fill_2
XFILLER_29_69 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_57 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_145 vgnd vpwr scs8hd_fill_1
XFILLER_34_137 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_16 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_56_56 vgnd vpwr scs8hd_decap_12
XFILLER_16_137 vgnd vpwr scs8hd_decap_8
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_7_50 vpwr vgnd scs8hd_fill_2
XFILLER_26_26 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_0_.latch/Q mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_58 vgnd vpwr scs8hd_decap_4
XANTENNA__094__B _096_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_100 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_2.LATCH_2_.latch data_in mem_right_ipin_2.LATCH_2_.latch/Q _096_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__195__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__089__B _083_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_3_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_4.LATCH_5_.latch data_in mem_right_ipin_4.LATCH_5_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _178_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XFILLER_4_73 vpwr vgnd scs8hd_fill_2
XFILLER_4_40 vgnd vpwr scs8hd_fill_1
XANTENNA__091__C _154_/C vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_1_.latch/Q mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_56 vgnd vpwr scs8hd_decap_6
X_184_ chany_top_in[4] chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_135 vgnd vpwr scs8hd_decap_8
XFILLER_59_45 vgnd vpwr scs8hd_decap_12
XFILLER_46_113 vgnd vpwr scs8hd_decap_12
XFILLER_46_102 vgnd vpwr scs8hd_decap_8
X_098_ _125_/A _096_/B _098_/Y vgnd vpwr scs8hd_nor2_4
X_167_ address[1] address[2] _161_/C _167_/X vgnd vpwr scs8hd_or3_4
XFILLER_52_105 vgnd vpwr scs8hd_decap_12
XFILLER_37_135 vgnd vpwr scs8hd_decap_8
XFILLER_29_15 vpwr vgnd scs8hd_fill_2
XANTENNA__097__B _096_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_102 vpwr vgnd scs8hd_fill_2
XFILLER_6_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_4_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_0_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_28 vpwr vgnd scs8hd_fill_2
XFILLER_25_127 vgnd vpwr scs8hd_decap_12
XFILLER_31_38 vpwr vgnd scs8hd_fill_2
XFILLER_56_68 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_decap_3
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_93 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_22_119 vgnd vpwr scs8hd_decap_4
XFILLER_30_130 vgnd vpwr scs8hd_decap_12
XFILLER_7_95 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_5.LATCH_1_.latch data_in mem_right_ipin_5.LATCH_1_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_130 vpwr vgnd scs8hd_fill_2
XFILLER_21_141 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_70 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_7.LATCH_4_.latch data_in mem_right_ipin_7.LATCH_4_.latch/Q _138_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_29 vpwr vgnd scs8hd_fill_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_ipin_6.LATCH_3_.latch/Q mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_ipin_6.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_85 vgnd vpwr scs8hd_decap_4
XFILLER_4_52 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_5_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_28 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _171_/HI _145_/Y mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_183_ chany_top_in[5] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_49_100 vgnd vpwr scs8hd_decap_12
XFILLER_64_125 vgnd vpwr scs8hd_decap_12
XFILLER_38_91 vgnd vpwr scs8hd_fill_1
XFILLER_18_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_50_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_57 vpwr vgnd scs8hd_fill_2
XFILLER_59_35 vpwr vgnd scs8hd_fill_2
XFILLER_46_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
X_097_ _124_/A _096_/B _097_/Y vgnd vpwr scs8hd_nor2_4
X_166_ _169_/A _140_/A _166_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_0_.latch/Q mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_52_117 vgnd vpwr scs8hd_decap_12
XFILLER_1_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_84 vgnd vpwr scs8hd_decap_8
XFILLER_34_106 vgnd vpwr scs8hd_decap_4
XFILLER_35_92 vgnd vpwr scs8hd_fill_1
X_149_ address[1] _149_/B _161_/C _149_/X vgnd vpwr scs8hd_or3_4
XFILLER_25_117 vgnd vpwr scs8hd_decap_4
XFILLER_25_139 vgnd vpwr scs8hd_decap_6
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_109 vpwr vgnd scs8hd_fill_2
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_1_.latch/Q mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_109 vgnd vpwr scs8hd_fill_1
XFILLER_26_17 vgnd vpwr scs8hd_decap_3
XFILLER_42_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_61 vgnd vpwr scs8hd_fill_1
XFILLER_57_90 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_49 vgnd vpwr scs8hd_fill_1
XFILLER_37_27 vpwr vgnd scs8hd_fill_2
XFILLER_53_59 vpwr vgnd scs8hd_fill_2
XFILLER_53_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_105 vpwr vgnd scs8hd_fill_2
XFILLER_27_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _179_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_48_48 vpwr vgnd scs8hd_fill_2
XFILLER_48_15 vgnd vpwr scs8hd_decap_12
XFILLER_58_145 vgnd vpwr scs8hd_fill_1
X_182_ chany_top_in[6] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_13_40 vpwr vgnd scs8hd_fill_2
XFILLER_13_73 vpwr vgnd scs8hd_fill_2
XFILLER_13_95 vgnd vpwr scs8hd_fill_1
XFILLER_49_123 vgnd vpwr scs8hd_decap_12
XFILLER_49_112 vgnd vpwr scs8hd_decap_8
XFILLER_1_130 vpwr vgnd scs8hd_fill_2
XFILLER_1_141 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_137 vgnd vpwr scs8hd_decap_8
XFILLER_54_80 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_0.LATCH_5_.latch data_in mem_right_ipin_0.LATCH_5_.latch/Q _070_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_4.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_50_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_137 vgnd vpwr scs8hd_decap_8
X_165_ _164_/X _140_/A vgnd vpwr scs8hd_buf_1
XFILLER_41_8 vpwr vgnd scs8hd_fill_2
XFILLER_40_82 vgnd vpwr scs8hd_decap_8
X_096_ _123_/A _096_/B _096_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_7 vgnd vpwr scs8hd_decap_3
XFILLER_52_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_6.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_61_59 vpwr vgnd scs8hd_fill_2
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_52 vpwr vgnd scs8hd_fill_2
XFILLER_19_83 vpwr vgnd scs8hd_fill_2
XFILLER_19_104 vpwr vgnd scs8hd_fill_2
XFILLER_19_115 vpwr vgnd scs8hd_fill_2
XFILLER_19_126 vpwr vgnd scs8hd_fill_2
XFILLER_19_137 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_71 vpwr vgnd scs8hd_fill_2
XFILLER_51_70 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
X_148_ address[0] _161_/C vgnd vpwr scs8hd_inv_8
Xmux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_ipin_5.LATCH_3_.latch/Q mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
X_079_ _142_/A _125_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_15 vgnd vpwr scs8hd_decap_12
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_51 vpwr vgnd scs8hd_fill_2
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_80 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_ipin_0.LATCH_4_.latch/Q mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_16_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_53_27 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_1.LATCH_1_.latch data_in mem_right_ipin_1.LATCH_1_.latch/Q _088_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_0_.latch/Q mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_71 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XFILLER_4_10 vpwr vgnd scs8hd_fill_2
XFILLER_48_27 vgnd vpwr scs8hd_decap_4
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_3.LATCH_4_.latch data_in mem_right_ipin_3.LATCH_4_.latch/Q _105_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_181_ chany_top_in[7] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_49_135 vgnd vpwr scs8hd_decap_8
XFILLER_38_71 vgnd vpwr scs8hd_fill_1
XANTENNA__100__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_15 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_40_61 vgnd vpwr scs8hd_decap_4
X_095_ _122_/A _096_/B _095_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_84 vgnd vpwr scs8hd_decap_4
X_164_ _161_/A address[2] address[0] _164_/X vgnd vpwr scs8hd_or3_4
Xmux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_8_ vgnd vpwr scs8hd_inv_1
Xmux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_1_.latch/Q mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_105 vgnd vpwr scs8hd_decap_4
XFILLER_1_88 vgnd vpwr scs8hd_decap_6
XANTENNA__111__A _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_60_141 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_62 vgnd vpwr scs8hd_decap_4
XFILLER_51_82 vgnd vpwr scs8hd_decap_12
X_078_ _124_/A _069_/X _078_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A _122_/A vgnd vpwr scs8hd_diode_2
X_147_ address[2] _149_/B vgnd vpwr scs8hd_inv_8
XFILLER_18_3 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_2_.latch/Q mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_27 vgnd vpwr scs8hd_decap_4
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_ipin_0.LATCH_5_.latch data_in mem_left_ipin_0.LATCH_5_.latch/Q _156_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_130 vgnd vpwr scs8hd_decap_12
XFILLER_21_30 vpwr vgnd scs8hd_fill_2
XFILLER_21_74 vpwr vgnd scs8hd_fill_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_54 vgnd vpwr scs8hd_decap_4
XFILLER_8_104 vgnd vpwr scs8hd_decap_12
XFILLER_12_144 vpwr vgnd scs8hd_fill_2
XFILLER_32_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_5.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_4.LATCH_0_.latch data_in mem_right_ipin_4.LATCH_0_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_39 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_0_.latch/Q mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_50 vpwr vgnd scs8hd_fill_2
XFILLER_27_51 vpwr vgnd scs8hd_fill_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_3
XANTENNA__114__A _122_/A vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_6.LATCH_3_.latch data_in mem_right_ipin_6.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
X_180_ chany_top_in[8] chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_ipin_4.LATCH_3_.latch/Q mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_64_106 vgnd vpwr scs8hd_decap_12
XFILLER_38_83 vgnd vpwr scs8hd_decap_8
XFILLER_54_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_59_27 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_9 vpwr vgnd scs8hd_fill_2
XFILLER_24_41 vgnd vpwr scs8hd_decap_3
XFILLER_40_51 vgnd vpwr scs8hd_fill_1
X_163_ _169_/A _139_/A _163_/Y vgnd vpwr scs8hd_nor2_4
X_094_ _121_/A _096_/B _094_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_49_71 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_1.LATCH_1_.latch data_in _145_/A _143_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_ipin_3.LATCH_1_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_106 vgnd vpwr scs8hd_decap_4
XFILLER_61_39 vgnd vpwr scs8hd_decap_12
XFILLER_10_32 vpwr vgnd scs8hd_fill_2
XFILLER_10_65 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_95 vgnd vpwr scs8hd_fill_1
XFILLER_51_94 vgnd vpwr scs8hd_decap_12
X_146_ _146_/A _146_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__106__B _108_/B vgnd vpwr scs8hd_diode_2
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
X_077_ _141_/A _124_/A vgnd vpwr scs8hd_buf_1
XFILLER_32_6 vpwr vgnd scs8hd_fill_2
XFILLER_25_109 vpwr vgnd scs8hd_fill_2
XFILLER_33_120 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_0_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_126 vgnd vpwr scs8hd_decap_3
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_decap_3
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_62_93 vgnd vpwr scs8hd_decap_12
XANTENNA__117__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_66 vgnd vpwr scs8hd_fill_1
XFILLER_7_33 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_99 vgnd vpwr scs8hd_decap_4
X_129_ _137_/A _131_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_112 vpwr vgnd scs8hd_fill_2
XFILLER_21_145 vgnd vpwr scs8hd_fill_1
XFILLER_16_64 vpwr vgnd scs8hd_fill_2
XFILLER_8_116 vgnd vpwr scs8hd_decap_12
XFILLER_37_19 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_6.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_1_.latch/Q mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_2_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__114__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_89 vgnd vpwr scs8hd_fill_1
XFILLER_4_56 vpwr vgnd scs8hd_fill_2
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
XANTENNA__130__A _138_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_100 vpwr vgnd scs8hd_fill_2
XFILLER_64_118 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__109__B _108_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _125_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
X_162_ _161_/X _139_/A vgnd vpwr scs8hd_buf_1
XFILLER_24_64 vgnd vpwr scs8hd_decap_3
XFILLER_40_41 vgnd vpwr scs8hd_decap_8
X_093_ _112_/A _096_/B _093_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_24 vpwr vgnd scs8hd_fill_2
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
XFILLER_51_143 vgnd vpwr scs8hd_decap_3
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_51_62 vgnd vpwr scs8hd_decap_4
X_145_ _145_/A _145_/Y vgnd vpwr scs8hd_inv_8
X_076_ _123_/A _069_/X _076_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__122__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_0_.latch/Q mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_decap_3
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_43 vpwr vgnd scs8hd_fill_2
XFILLER_21_65 vpwr vgnd scs8hd_fill_2
XFILLER_46_84 vgnd vpwr scs8hd_decap_8
XFILLER_46_62 vgnd vpwr scs8hd_fill_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_143 vgnd vpwr scs8hd_decap_3
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XANTENNA__117__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_78 vpwr vgnd scs8hd_fill_2
XFILLER_7_12 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A _141_/A vgnd vpwr scs8hd_diode_2
X_128_ _128_/A _131_/B vgnd vpwr scs8hd_buf_1
XFILLER_23_3 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _146_/Y mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_ipin_3.LATCH_3_.latch/Q mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_12_102 vpwr vgnd scs8hd_fill_2
XFILLER_12_113 vgnd vpwr scs8hd_decap_8
XFILLER_12_124 vgnd vpwr scs8hd_decap_12
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XFILLER_16_43 vgnd vpwr scs8hd_decap_4
XFILLER_8_128 vgnd vpwr scs8hd_decap_12
XANTENNA__128__A _128_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_109 vpwr vgnd scs8hd_fill_2
XFILLER_27_31 vpwr vgnd scs8hd_fill_2
XFILLER_27_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_3_ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _131_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.LATCH_0_.latch data_in mem_right_ipin_0.LATCH_0_.latch/Q _080_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_4.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_88 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_ipin_7.LATCH_4_.latch/Q mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_38_41 vgnd vpwr scs8hd_decap_3
XFILLER_1_145 vgnd vpwr scs8hd_fill_1
XANTENNA__125__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _141_/A vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_2.LATCH_3_.latch data_in mem_right_ipin_2.LATCH_3_.latch/Q _095_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_54_141 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_5.INVTX1_5_.scs8hd_inv_1 chany_top_in[7] mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB _064_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_10 vpwr vgnd scs8hd_fill_2
XFILLER_24_76 vpwr vgnd scs8hd_fill_2
X_161_ _161_/A address[2] _161_/C _161_/X vgnd vpwr scs8hd_or3_4
X_092_ _092_/A _096_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mem_right_ipin_6.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XANTENNA__136__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_119 vgnd vpwr scs8hd_decap_8
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_19_32 vpwr vgnd scs8hd_fill_2
XFILLER_19_87 vpwr vgnd scs8hd_fill_2
XFILLER_19_119 vgnd vpwr scs8hd_decap_3
XFILLER_27_130 vpwr vgnd scs8hd_fill_2
XFILLER_27_141 vgnd vpwr scs8hd_decap_4
XFILLER_35_31 vpwr vgnd scs8hd_fill_2
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XFILLER_35_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_144_ _143_/A _143_/B address[0] _144_/Y vgnd vpwr scs8hd_nor3_4
X_075_ _140_/A _123_/A vgnd vpwr scs8hd_buf_1
Xmux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_1_.latch/Q mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XPHY_106 vgnd vpwr scs8hd_decap_3
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_55 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_8 vgnd vpwr scs8hd_decap_3
X_127_ address[5] _127_/B _154_/C _128_/A vgnd vpwr scs8hd_or3_4
XFILLER_7_46 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_136 vgnd vpwr scs8hd_decap_8
XFILLER_16_88 vpwr vgnd scs8hd_fill_2
XFILLER_32_10 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vpwr vgnd scs8hd_fill_2
XFILLER_32_65 vgnd vpwr scs8hd_decap_3
XFILLER_57_62 vgnd vpwr scs8hd_decap_12
XFILLER_57_51 vgnd vpwr scs8hd_decap_8
XANTENNA__144__A _143_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_3_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_2_.latch/Q mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_76 vpwr vgnd scs8hd_fill_2
XFILLER_43_75 vgnd vpwr scs8hd_decap_3
XFILLER_4_36 vpwr vgnd scs8hd_fill_2
XFILLER_4_69 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_117 vgnd vpwr scs8hd_decap_12
XFILLER_13_23 vpwr vgnd scs8hd_fill_2
XFILLER_1_113 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_5.LATCH_2_.latch data_in mem_right_ipin_5.LATCH_2_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_64 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_0_.latch/Q mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__141__B _142_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_7.LATCH_5_.latch data_in mem_right_ipin_7.LATCH_5_.latch/Q _137_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_21 vgnd vpwr scs8hd_decap_8
X_091_ _091_/A address[6] _154_/C _092_/A vgnd vpwr scs8hd_or3_4
XFILLER_24_88 vgnd vpwr scs8hd_fill_1
X_160_ address[1] _161_/A vgnd vpwr scs8hd_inv_8
XFILLER_40_65 vgnd vpwr scs8hd_fill_1
XFILLER_45_120 vpwr vgnd scs8hd_fill_2
XFILLER_37_109 vgnd vpwr scs8hd_fill_1
XFILLER_60_145 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__152__A enable vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_1_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_2.LATCH_3_.latch/Q mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_51_123 vgnd vpwr scs8hd_decap_12
XFILLER_36_131 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_2.LATCH_4_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__062__A address[1] vgnd vpwr scs8hd_diode_2
X_074_ _122_/A _069_/X _074_/Y vgnd vpwr scs8hd_nor2_4
X_143_ _143_/A _143_/B _161_/C _143_/Y vgnd vpwr scs8hd_nor3_4
Xmem_left_ipin_0.LATCH_0_.latch data_in mem_left_ipin_0.LATCH_0_.latch/Q _064_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.INVTX1_5_.scs8hd_inv_1 chany_top_in[5] mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_112 vgnd vpwr scs8hd_decap_8
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XANTENNA__147__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
XPHY_129 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XPHY_107 vgnd vpwr scs8hd_decap_3
XFILLER_21_89 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_101 vgnd vpwr scs8hd_decap_4
XFILLER_15_112 vpwr vgnd scs8hd_fill_2
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
X_126_ address[6] _127_/B vgnd vpwr scs8hd_inv_8
XFILLER_7_58 vgnd vpwr scs8hd_fill_1
XFILLER_30_6 vpwr vgnd scs8hd_fill_2
XFILLER_21_126 vpwr vgnd scs8hd_fill_2
XFILLER_21_137 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_ipin_6.LATCH_4_.latch/Q mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_88 vpwr vgnd scs8hd_fill_2
XFILLER_57_74 vpwr vgnd scs8hd_fill_2
XANTENNA__144__B _143_/B vgnd vpwr scs8hd_diode_2
XANTENNA__160__A address[1] vgnd vpwr scs8hd_diode_2
X_109_ _125_/A _108_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__070__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_43_10 vpwr vgnd scs8hd_fill_2
XFILLER_27_55 vgnd vpwr scs8hd_decap_4
XFILLER_43_54 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB _070_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _155_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _171_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__065__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_1_.latch/Q mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_143 vgnd vpwr scs8hd_decap_3
XFILLER_63_110 vgnd vpwr scs8hd_decap_12
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
X_090_ address[5] _091_/A vgnd vpwr scs8hd_inv_8
XFILLER_49_75 vpwr vgnd scs8hd_fill_2
XFILLER_49_53 vpwr vgnd scs8hd_fill_2
XFILLER_49_42 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_3
XFILLER_45_143 vgnd vpwr scs8hd_decap_3
XFILLER_39_3 vgnd vpwr scs8hd_decap_4
XFILLER_51_135 vgnd vpwr scs8hd_decap_8
XFILLER_36_143 vgnd vpwr scs8hd_decap_3
XFILLER_10_36 vgnd vpwr scs8hd_fill_1
XANTENNA__062__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_42_102 vgnd vpwr scs8hd_decap_12
XFILLER_51_10 vgnd vpwr scs8hd_decap_12
X_142_ _142_/A _142_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_35_88 vgnd vpwr scs8hd_decap_4
XFILLER_35_99 vgnd vpwr scs8hd_decap_4
X_073_ _139_/A _122_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_8
XANTENNA__163__A _169_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_2_.latch/Q mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_81 vpwr vgnd scs8hd_fill_2
XFILLER_24_102 vgnd vpwr scs8hd_decap_8
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
XFILLER_21_13 vgnd vpwr scs8hd_fill_1
XANTENNA__073__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_46_65 vgnd vpwr scs8hd_decap_3
XFILLER_46_54 vpwr vgnd scs8hd_fill_2
XFILLER_15_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_125_ _125_/A _123_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_116 vgnd vpwr scs8hd_decap_6
XANTENNA__158__A _157_/X vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.INVTX1_5_.scs8hd_inv_1 chany_top_in[7] mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_4_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__068__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_57 vgnd vpwr scs8hd_decap_4
XFILLER_16_68 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_0_.latch/Q mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_23 vpwr vgnd scs8hd_fill_2
XANTENNA__144__C address[0] vgnd vpwr scs8hd_diode_2
X_108_ _124_/A _108_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_3 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_0.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__070__B _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_12 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_7.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_ipin_1.LATCH_3_.latch/Q mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_4_145 vgnd vpwr scs8hd_fill_1
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_13_36 vpwr vgnd scs8hd_fill_2
XFILLER_13_69 vpwr vgnd scs8hd_fill_2
XFILLER_1_104 vgnd vpwr scs8hd_decap_3
XFILLER_1_126 vpwr vgnd scs8hd_fill_2
XFILLER_1_137 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_54_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_92 vpwr vgnd scs8hd_fill_2
XANTENNA__076__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_46 vgnd vpwr scs8hd_decap_4
XFILLER_40_78 vpwr vgnd scs8hd_fill_2
XFILLER_1_28 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_5.LATCH_5_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_1.LATCH_2_.latch data_in mem_right_ipin_1.LATCH_2_.latch/Q _087_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_90 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_ipin_5.LATCH_4_.latch/Q mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_36_100 vpwr vgnd scs8hd_fill_2
XANTENNA__062__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_10_48 vpwr vgnd scs8hd_fill_2
XFILLER_19_13 vpwr vgnd scs8hd_fill_2
XFILLER_42_114 vgnd vpwr scs8hd_decap_12
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XFILLER_19_68 vpwr vgnd scs8hd_fill_2
XFILLER_35_12 vpwr vgnd scs8hd_fill_2
XFILLER_51_66 vgnd vpwr scs8hd_fill_1
XFILLER_51_22 vgnd vpwr scs8hd_decap_12
X_141_ _141_/A _142_/B _141_/Y vgnd vpwr scs8hd_nor2_4
X_072_ _121_/A _069_/X _072_/Y vgnd vpwr scs8hd_nor2_4
Xmem_right_ipin_3.LATCH_5_.latch data_in mem_right_ipin_3.LATCH_5_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_144 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _139_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _170_/HI mem_left_ipin_0.LATCH_5_.latch/Q
+ mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_93 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_decap_3
XFILLER_21_47 vpwr vgnd scs8hd_fill_2
XFILLER_21_69 vgnd vpwr scs8hd_decap_3
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XFILLER_30_106 vgnd vpwr scs8hd_decap_4
X_124_ _124_/A _123_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_23_7 vpwr vgnd scs8hd_fill_2
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
XFILLER_21_106 vgnd vpwr scs8hd_decap_4
XANTENNA__068__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_12_106 vgnd vpwr scs8hd_decap_4
XFILLER_16_47 vgnd vpwr scs8hd_fill_1
XANTENNA__084__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_46 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_1_.latch/Q mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_143 vgnd vpwr scs8hd_decap_3
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
X_107_ _123_/A _108_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_3 vgnd vpwr scs8hd_decap_4
XANTENNA__169__A _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__079__A _142_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_35 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_89 vgnd vpwr scs8hd_decap_12
XFILLER_43_34 vgnd vpwr scs8hd_decap_3
XFILLER_4_113 vgnd vpwr scs8hd_decap_12
XFILLER_4_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XFILLER_38_23 vgnd vpwr scs8hd_decap_4
XFILLER_38_12 vpwr vgnd scs8hd_fill_2
XFILLER_54_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_2_.latch/Q mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_5.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[6] mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_63_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__166__B _140_/A vgnd vpwr scs8hd_diode_2
XANTENNA__182__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XFILLER_54_145 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_4.LATCH_1_.latch data_in mem_right_ipin_4.LATCH_1_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__076__B _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_49_88 vgnd vpwr scs8hd_decap_12
XFILLER_45_123 vgnd vpwr scs8hd_decap_12
XFILLER_45_112 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_0_.latch/Q mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_6.LATCH_4_.latch data_in mem_right_ipin_6.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_36 vgnd vpwr scs8hd_decap_4
XFILLER_42_126 vgnd vpwr scs8hd_decap_12
XANTENNA__087__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_112 vpwr vgnd scs8hd_fill_2
XFILLER_27_145 vgnd vpwr scs8hd_fill_1
XFILLER_35_35 vgnd vpwr scs8hd_decap_4
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
XFILLER_51_34 vgnd vpwr scs8hd_decap_12
X_140_ _140_/A _142_/B _140_/Y vgnd vpwr scs8hd_nor2_4
X_071_ _138_/A _121_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_104 vpwr vgnd scs8hd_fill_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_8
XFILLER_21_26 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_ipin_0.LATCH_3_.latch/Q mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XFILLER_46_23 vpwr vgnd scs8hd_fill_2
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
X_123_ _123_/A _123_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__190__A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__068__C _143_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_1_.latch/Q mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__084__B _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_36 vgnd vpwr scs8hd_fill_1
X_106_ _122_/A _108_/B _106_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__169__B _141_/A vgnd vpwr scs8hd_diode_2
XANTENNA__185__A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _146_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_46 vpwr vgnd scs8hd_fill_2
XANTENNA__095__A _122_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_4.LATCH_4_.latch/Q mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_4_125 vgnd vpwr scs8hd_decap_12
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_57_143 vgnd vpwr scs8hd_decap_3
XFILLER_38_68 vgnd vpwr scs8hd_fill_1
XFILLER_38_46 vgnd vpwr scs8hd_fill_1
XFILLER_1_117 vgnd vpwr scs8hd_decap_3
XFILLER_54_56 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_7.LATCH_0_.latch data_in mem_right_ipin_7.LATCH_0_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_135 vgnd vpwr scs8hd_decap_8
XFILLER_39_143 vgnd vpwr scs8hd_decap_3
XFILLER_24_59 vgnd vpwr scs8hd_decap_3
XFILLER_45_135 vgnd vpwr scs8hd_decap_8
XFILLER_45_102 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_60_105 vgnd vpwr scs8hd_decap_12
XANTENNA__193__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_1_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_3.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_138 vgnd vpwr scs8hd_decap_8
XANTENNA__087__B _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_51_46 vgnd vpwr scs8hd_decap_12
X_070_ _112_/A _069_/X _070_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_102 vgnd vpwr scs8hd_decap_8
XFILLER_18_113 vpwr vgnd scs8hd_fill_2
XFILLER_18_124 vgnd vpwr scs8hd_decap_12
XPHY_91 vgnd vpwr scs8hd_decap_3
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_51 vpwr vgnd scs8hd_fill_2
XANTENNA__188__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_16 vgnd vpwr scs8hd_fill_1
XFILLER_46_79 vgnd vpwr scs8hd_decap_3
XFILLER_46_35 vgnd vpwr scs8hd_decap_6
XFILLER_15_116 vgnd vpwr scs8hd_decap_6
XANTENNA__098__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_62_56 vgnd vpwr scs8hd_decap_12
XFILLER_30_119 vgnd vpwr scs8hd_decap_8
XFILLER_7_29 vpwr vgnd scs8hd_fill_2
XFILLER_11_71 vpwr vgnd scs8hd_fill_2
X_122_ _122_/A _123_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_57_78 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_2_.latch/Q mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_11_130 vgnd vpwr scs8hd_decap_12
XFILLER_22_70 vgnd vpwr scs8hd_decap_4
X_105_ _121_/A _108_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB _076_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_14 vpwr vgnd scs8hd_fill_2
XFILLER_43_58 vgnd vpwr scs8hd_fill_1
XANTENNA__095__B _096_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_137 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_92 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_0_.latch/Q mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__196__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_58 vgnd vpwr scs8hd_decap_4
XFILLER_54_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_111 vpwr vgnd scs8hd_fill_2
XFILLER_39_100 vpwr vgnd scs8hd_fill_2
XFILLER_24_27 vpwr vgnd scs8hd_fill_2
XFILLER_49_57 vpwr vgnd scs8hd_fill_2
XFILLER_49_46 vpwr vgnd scs8hd_fill_2
XFILLER_60_117 vgnd vpwr scs8hd_decap_12
XFILLER_39_7 vgnd vpwr scs8hd_fill_1
XFILLER_51_106 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_1_.latch/Q mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.LATCH_1_.latch data_in mem_right_ipin_0.LATCH_1_.latch/Q _078_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_136 vgnd vpwr scs8hd_decap_8
XPHY_92 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_51_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_85 vgnd vpwr scs8hd_decap_6
Xmux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_ipin_3.LATCH_4_.latch/Q mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_46_58 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_2.LATCH_4_.latch data_in mem_right_ipin_2.LATCH_4_.latch/Q _094_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__098__B _096_/B vgnd vpwr scs8hd_diode_2
XFILLER_62_68 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[3] mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_121_ _121_/A _123_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_91 vgnd vpwr scs8hd_fill_1
XFILLER_16_39 vpwr vgnd scs8hd_fill_2
XFILLER_20_131 vgnd vpwr scs8hd_decap_12
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_135 vgnd vpwr scs8hd_decap_8
XFILLER_11_142 vgnd vpwr scs8hd_decap_4
X_104_ _112_/A _108_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_27_16 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _179_/HI mem_right_ipin_7.LATCH_5_.latch/Q
+ mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_6
XFILLER_57_123 vgnd vpwr scs8hd_decap_12
XFILLER_38_37 vpwr vgnd scs8hd_fill_2
XFILLER_48_101 vgnd vpwr scs8hd_decap_12
XFILLER_48_145 vgnd vpwr scs8hd_fill_1
XFILLER_28_81 vgnd vpwr scs8hd_decap_3
XFILLER_44_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_5.LATCH_2_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_6_8 vpwr vgnd scs8hd_fill_2
XFILLER_60_129 vgnd vpwr scs8hd_decap_12
XFILLER_14_50 vpwr vgnd scs8hd_fill_2
XFILLER_14_72 vgnd vpwr scs8hd_decap_4
XFILLER_51_118 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_3.LATCH_0_.latch data_in mem_right_ipin_3.LATCH_0_.latch/Q _109_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_17 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_2_.latch/Q mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_104 vpwr vgnd scs8hd_fill_2
XFILLER_27_126 vpwr vgnd scs8hd_fill_2
XFILLER_27_137 vpwr vgnd scs8hd_fill_2
XFILLER_35_16 vpwr vgnd scs8hd_fill_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
X_197_ chany_bottom_in[0] chany_top_out[0] vgnd vpwr scs8hd_buf_2
XPHY_93 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_5.LATCH_3_.latch data_in mem_right_ipin_5.LATCH_3_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_15 vgnd vpwr scs8hd_decap_4
X_120_ _137_/A _123_/B _120_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_0_.latch/Q mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_80 vgnd vpwr scs8hd_decap_12
XFILLER_42_3 vgnd vpwr scs8hd_decap_8
XFILLER_20_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_3.LATCH_3_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_22_83 vgnd vpwr scs8hd_decap_3
X_103_ _103_/A _108_/B vgnd vpwr scs8hd_buf_1
XFILLER_47_91 vpwr vgnd scs8hd_fill_2
XFILLER_8_96 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_0.LATCH_1_.latch data_in mem_left_ipin_0.LATCH_1_.latch/Q _169_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_106 vgnd vpwr scs8hd_decap_4
XFILLER_17_50 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_1_.latch/Q mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_19 vpwr vgnd scs8hd_fill_2
XFILLER_57_102 vgnd vpwr scs8hd_decap_12
XFILLER_38_16 vgnd vpwr scs8hd_decap_4
XFILLER_57_135 vgnd vpwr scs8hd_decap_8
XFILLER_54_15 vgnd vpwr scs8hd_decap_12
XFILLER_48_113 vgnd vpwr scs8hd_decap_12
XFILLER_0_120 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_60 vgnd vpwr scs8hd_decap_8
XFILLER_60_91 vgnd vpwr scs8hd_fill_1
XFILLER_44_81 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_ipin_2.LATCH_4_.latch/Q mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_2_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_54_105 vgnd vpwr scs8hd_decap_12
XFILLER_39_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.INVTX1_3_.scs8hd_inv_1 chany_top_in[7] mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_49_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_1.LATCH_4_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_72 vgnd vpwr scs8hd_fill_1
XANTENNA__101__A _100_/X vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_116 vgnd vpwr scs8hd_decap_6
XFILLER_35_39 vgnd vpwr scs8hd_fill_1
XFILLER_50_141 vgnd vpwr scs8hd_decap_4
XFILLER_4_6 vpwr vgnd scs8hd_fill_2
XPHY_94 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_33_108 vpwr vgnd scs8hd_fill_2
XPHY_72 vgnd vpwr scs8hd_decap_3
X_196_ chany_bottom_in[1] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_41_71 vpwr vgnd scs8hd_fill_2
XFILLER_2_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _145_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_119 vgnd vpwr scs8hd_decap_8
XFILLER_32_130 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _178_/HI mem_right_ipin_6.LATCH_5_.latch/Q
+ mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_46_27 vgnd vpwr scs8hd_decap_4
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_108 vpwr vgnd scs8hd_fill_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_179_ _179_/HI _179_/LO vgnd vpwr scs8hd_conb_1
XFILLER_57_15 vgnd vpwr scs8hd_decap_12
XFILLER_57_59 vpwr vgnd scs8hd_fill_2
X_102_ _102_/A _143_/B _103_/A vgnd vpwr scs8hd_or2_4
XFILLER_21_9 vgnd vpwr scs8hd_decap_4
XFILLER_8_64 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_72 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_2_.latch/Q mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__104__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_80 vgnd vpwr scs8hd_decap_12
XFILLER_57_114 vgnd vpwr scs8hd_decap_8
XFILLER_54_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_125 vgnd vpwr scs8hd_decap_12
XFILLER_0_132 vgnd vpwr scs8hd_decap_12
XFILLER_44_93 vpwr vgnd scs8hd_fill_2
XFILLER_5_32 vpwr vgnd scs8hd_fill_2
XFILLER_54_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_0_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_27 vgnd vpwr scs8hd_decap_12
XFILLER_14_41 vgnd vpwr scs8hd_decap_3
XFILLER_30_84 vpwr vgnd scs8hd_fill_2
XFILLER_18_117 vgnd vpwr scs8hd_decap_4
XPHY_95 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_4.INVTX1_3_.scs8hd_inv_1 chany_top_in[5] mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
X_195_ chany_bottom_in[2] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_37_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_22 vpwr vgnd scs8hd_fill_2
XANTENNA__112__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_1_.latch/Q mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_42 vpwr vgnd scs8hd_fill_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_75 vpwr vgnd scs8hd_fill_2
XFILLER_36_83 vpwr vgnd scs8hd_fill_2
XFILLER_36_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_52_93 vgnd vpwr scs8hd_decap_12
XANTENNA__107__A _123_/A vgnd vpwr scs8hd_diode_2
X_178_ _178_/HI _178_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_right_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_3 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_1.LATCH_3_.latch data_in mem_right_ipin_1.LATCH_3_.latch/Q _086_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_57_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_ipin_1.LATCH_4_.latch/Q mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
X_101_ _100_/X _143_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_14_9 vpwr vgnd scs8hd_fill_2
XFILLER_8_54 vpwr vgnd scs8hd_fill_2
XFILLER_8_43 vpwr vgnd scs8hd_fill_2
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_43_29 vgnd vpwr scs8hd_decap_3
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_3
XFILLER_3_130 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _108_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _137_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_29 vpwr vgnd scs8hd_fill_2
XFILLER_0_144 vpwr vgnd scs8hd_fill_2
XFILLER_0_111 vgnd vpwr scs8hd_fill_1
XFILLER_48_137 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_60_93 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _177_/HI mem_right_ipin_5.LATCH_5_.latch/Q
+ mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__115__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_115 vpwr vgnd scs8hd_fill_2
XFILLER_39_104 vpwr vgnd scs8hd_fill_2
XFILLER_5_88 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_54_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_4.LATCH_5_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_83 vpwr vgnd scs8hd_fill_2
XFILLER_36_107 vgnd vpwr scs8hd_decap_12
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_143 vgnd vpwr scs8hd_decap_3
XFILLER_41_121 vgnd vpwr scs8hd_fill_1
XFILLER_41_40 vpwr vgnd scs8hd_fill_2
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_85 vpwr vgnd scs8hd_fill_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
X_194_ chany_bottom_in[3] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_41_51 vpwr vgnd scs8hd_fill_2
XANTENNA__112__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_2_.latch/Q mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_4.LATCH_2_.latch data_in mem_right_ipin_4.LATCH_2_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_177_ _177_/HI _177_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__107__B _108_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XFILLER_57_39 vgnd vpwr scs8hd_decap_12
XFILLER_7_106 vpwr vgnd scs8hd_fill_2
X_100_ address[4] _118_/B _100_/X vgnd vpwr scs8hd_or2_4
Xmem_right_ipin_6.LATCH_5_.latch data_in mem_right_ipin_6.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__118__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_88 vpwr vgnd scs8hd_fill_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_6
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_41 vgnd vpwr scs8hd_decap_6
XFILLER_3_142 vgnd vpwr scs8hd_decap_4
XFILLER_58_93 vgnd vpwr scs8hd_decap_12
XANTENNA__120__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_30 vgnd vpwr scs8hd_fill_1
XFILLER_44_62 vpwr vgnd scs8hd_fill_2
XANTENNA__115__B _116_/B vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_62_141 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_1_.latch/Q mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_54 vgnd vpwr scs8hd_decap_3
XFILLER_14_76 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _146_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_53 vpwr vgnd scs8hd_fill_2
XFILLER_30_64 vgnd vpwr scs8hd_decap_8
XFILLER_39_62 vgnd vpwr scs8hd_decap_4
XFILLER_39_40 vpwr vgnd scs8hd_fill_2
XFILLER_36_119 vgnd vpwr scs8hd_decap_12
XANTENNA__126__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_108 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_ipin_0.LATCH_4_.latch/Q mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_31 vpwr vgnd scs8hd_fill_2
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
X_193_ chany_bottom_in[4] chany_top_out[4] vgnd vpwr scs8hd_buf_2
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_75 vpwr vgnd scs8hd_fill_2
XFILLER_2_68 vpwr vgnd scs8hd_fill_2
XFILLER_17_130 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_7.LATCH_1_.latch data_in mem_right_ipin_7.LATCH_1_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_19 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_2_.latch/Q mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_144 vpwr vgnd scs8hd_fill_2
XFILLER_11_22 vpwr vgnd scs8hd_fill_2
XFILLER_11_88 vpwr vgnd scs8hd_fill_2
XFILLER_36_96 vpwr vgnd scs8hd_fill_2
XFILLER_14_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_3.LATCH_0_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
X_176_ _176_/HI _176_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__123__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_10 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _176_/HI mem_right_ipin_4.LATCH_5_.latch/Q
+ mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_95 vpwr vgnd scs8hd_fill_2
XFILLER_47_62 vgnd vpwr scs8hd_fill_1
XFILLER_47_40 vpwr vgnd scs8hd_fill_2
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_78 vgnd vpwr scs8hd_decap_8
X_159_ _169_/A _138_/A _159_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__A _142_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_12_ vgnd vpwr scs8hd_inv_1
XFILLER_33_3 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_0.INVTX1_3_.scs8hd_inv_1 chany_top_in[2] mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_54 vgnd vpwr scs8hd_decap_4
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__A _137_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_86 vgnd vpwr scs8hd_decap_6
Xmux_right_ipin_6.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA__131__B _131_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_2_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_0.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_22 vgnd vpwr scs8hd_decap_6
XFILLER_30_10 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_7.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_62 vgnd vpwr scs8hd_decap_12
XFILLER_55_51 vgnd vpwr scs8hd_decap_8
XANTENNA__142__A _142_/A vgnd vpwr scs8hd_diode_2
XFILLER_50_145 vgnd vpwr scs8hd_fill_1
XPHY_98 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_decap_3
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_25_10 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
X_192_ chany_bottom_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_41_75 vpwr vgnd scs8hd_fill_2
XFILLER_25_98 vpwr vgnd scs8hd_fill_2
XFILLER_2_47 vpwr vgnd scs8hd_fill_2
XFILLER_17_120 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A _137_/A vgnd vpwr scs8hd_diode_2
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_112 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_175_ _175_/HI _175_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_126 vpwr vgnd scs8hd_fill_2
XFILLER_22_66 vpwr vgnd scs8hd_fill_2
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
XFILLER_47_74 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_1_.latch/Q mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
XFILLER_8_35 vpwr vgnd scs8hd_fill_2
XANTENNA__118__C _102_/A vgnd vpwr scs8hd_diode_2
X_089_ _125_/A _083_/X _089_/Y vgnd vpwr scs8hd_nor2_4
Xmem_right_ipin_0.LATCH_2_.latch data_in mem_right_ipin_0.LATCH_2_.latch/Q _076_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_158_ _157_/X _138_/A vgnd vpwr scs8hd_buf_1
XANTENNA__134__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_3
XANTENNA__150__A _149_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_33 vpwr vgnd scs8hd_fill_2
XFILLER_17_88 vpwr vgnd scs8hd_fill_2
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_21 vgnd vpwr scs8hd_decap_4
XFILLER_33_87 vpwr vgnd scs8hd_fill_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_111 vpwr vgnd scs8hd_fill_2
XFILLER_3_100 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_2.LATCH_5_.latch data_in mem_right_ipin_2.LATCH_5_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__129__B _131_/B vgnd vpwr scs8hd_diode_2
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_103 vgnd vpwr scs8hd_decap_8
XFILLER_28_43 vpwr vgnd scs8hd_fill_2
XFILLER_44_97 vgnd vpwr scs8hd_decap_12
XFILLER_5_36 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_2_.latch/Q mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_53_143 vgnd vpwr scs8hd_decap_3
XFILLER_53_110 vgnd vpwr scs8hd_decap_12
XFILLER_30_88 vgnd vpwr scs8hd_decap_4
XFILLER_44_121 vgnd vpwr scs8hd_decap_12
XFILLER_39_53 vpwr vgnd scs8hd_fill_2
XFILLER_55_74 vgnd vpwr scs8hd_decap_12
XANTENNA__142__B _142_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_143 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _175_/HI mem_right_ipin_3.LATCH_5_.latch/Q
+ mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_99 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_decap_3
XFILLER_41_135 vgnd vpwr scs8hd_decap_8
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
X_191_ chany_bottom_in[6] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_41_21 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_26 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_102 vpwr vgnd scs8hd_fill_2
XANTENNA__137__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_5.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__153__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA__063__A _062_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_87 vgnd vpwr scs8hd_decap_4
XFILLER_36_76 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_14_102 vpwr vgnd scs8hd_fill_2
XFILLER_14_113 vgnd vpwr scs8hd_decap_8
XFILLER_36_10 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_fill_1
XFILLER_14_124 vgnd vpwr scs8hd_decap_12
X_174_ _174_/HI _174_/LO vgnd vpwr scs8hd_conb_1
XFILLER_28_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__148__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _170_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_105 vpwr vgnd scs8hd_fill_2
XFILLER_22_23 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_3.LATCH_1_.latch data_in mem_right_ipin_3.LATCH_1_.latch/Q _108_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_47_53 vpwr vgnd scs8hd_fill_2
XFILLER_63_74 vgnd vpwr scs8hd_decap_12
XFILLER_8_58 vgnd vpwr scs8hd_decap_4
X_157_ address[1] _149_/B address[0] _157_/X vgnd vpwr scs8hd_or3_4
X_088_ _124_/A _083_/X _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_5.LATCH_4_.latch data_in mem_right_ipin_5.LATCH_4_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_2_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__071__A _138_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_141 vgnd vpwr scs8hd_decap_4
XFILLER_28_22 vpwr vgnd scs8hd_fill_2
XFILLER_28_77 vpwr vgnd scs8hd_fill_2
XFILLER_60_75 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vpwr vgnd scs8hd_fill_2
XFILLER_39_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__156__A _112_/A vgnd vpwr scs8hd_diode_2
XANTENNA__066__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_14_46 vpwr vgnd scs8hd_fill_2
XFILLER_14_79 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_0.LATCH_2_.latch data_in mem_left_ipin_0.LATCH_2_.latch/Q _166_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_23 vgnd vpwr scs8hd_decap_6
XFILLER_30_45 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_55_86 vgnd vpwr scs8hd_decap_12
XFILLER_44_133 vgnd vpwr scs8hd_decap_12
XFILLER_39_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_130 vpwr vgnd scs8hd_fill_2
XFILLER_29_141 vgnd vpwr scs8hd_decap_4
XPHY_12 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_1_.latch/Q mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_144 vpwr vgnd scs8hd_fill_2
X_190_ chany_bottom_in[7] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XPHY_89 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XFILLER_41_88 vgnd vpwr scs8hd_decap_6
XFILLER_41_55 vgnd vpwr scs8hd_decap_4
XFILLER_41_44 vpwr vgnd scs8hd_fill_2
XANTENNA__153__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_23_136 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_2.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_36_55 vgnd vpwr scs8hd_decap_8
XFILLER_14_136 vgnd vpwr scs8hd_decap_8
XFILLER_52_32 vgnd vpwr scs8hd_decap_12
X_173_ _173_/HI _173_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_right_ipin_2.LATCH_3_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_6.LATCH_0_.latch data_in mem_right_ipin_6.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_106 vgnd vpwr scs8hd_decap_4
XANTENNA__164__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_117 vgnd vpwr scs8hd_decap_3
XANTENNA__074__A _122_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_47_21 vgnd vpwr scs8hd_fill_1
XFILLER_63_86 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_2_.latch/Q mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_087_ _123_/A _083_/X _087_/Y vgnd vpwr scs8hd_nor2_4
X_156_ _112_/A _169_/A _156_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__159__A _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _069_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _145_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _174_/HI mem_right_ipin_2.LATCH_5_.latch/Q
+ mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_139_ _139_/A _142_/B _139_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_31_3 vgnd vpwr scs8hd_decap_3
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_44_66 vpwr vgnd scs8hd_fill_2
XFILLER_44_11 vgnd vpwr scs8hd_fill_1
XFILLER_60_87 vgnd vpwr scs8hd_decap_4
XFILLER_60_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_49 vpwr vgnd scs8hd_fill_2
XFILLER_47_120 vpwr vgnd scs8hd_fill_2
XFILLER_10_8 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB _072_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_53_123 vgnd vpwr scs8hd_decap_12
XANTENNA__066__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__082__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_55_98 vgnd vpwr scs8hd_decap_12
XFILLER_44_145 vgnd vpwr scs8hd_fill_1
XANTENNA__167__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XFILLER_6_81 vgnd vpwr scs8hd_decap_4
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_25_35 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _141_/A vgnd vpwr scs8hd_diode_2
XPHY_79 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_25_79 vgnd vpwr scs8hd_decap_4
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XFILLER_17_112 vgnd vpwr scs8hd_decap_8
XFILLER_17_134 vgnd vpwr scs8hd_decap_12
XANTENNA__153__C _066_/C vgnd vpwr scs8hd_diode_2
XFILLER_11_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_23 vgnd vpwr scs8hd_decap_8
XFILLER_52_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_172_ _172_/HI _172_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__164__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XANTENNA__180__A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_3_71 vpwr vgnd scs8hd_fill_2
XANTENNA__074__B _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_36 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_63_98 vgnd vpwr scs8hd_decap_12
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_155_ _155_/A _169_/A vgnd vpwr scs8hd_buf_1
XFILLER_12_80 vpwr vgnd scs8hd_fill_2
X_086_ _122_/A _083_/X _086_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__159__B _138_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_14 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_58 vgnd vpwr scs8hd_fill_1
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XFILLER_33_68 vpwr vgnd scs8hd_fill_2
XFILLER_58_32 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_3_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_90 vpwr vgnd scs8hd_fill_2
X_138_ _138_/A _142_/B _138_/Y vgnd vpwr scs8hd_nor2_4
X_069_ _069_/A _069_/X vgnd vpwr scs8hd_buf_1
XANTENNA__161__C _161_/C vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_1_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XFILLER_9_92 vgnd vpwr scs8hd_fill_1
XFILLER_0_128 vpwr vgnd scs8hd_fill_2
XFILLER_44_23 vpwr vgnd scs8hd_fill_2
XFILLER_60_44 vgnd vpwr scs8hd_decap_12
XFILLER_44_45 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_1.LATCH_4_.latch data_in mem_right_ipin_1.LATCH_4_.latch/Q _085_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_47_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_53_135 vgnd vpwr scs8hd_decap_8
XANTENNA__066__C _066_/C vgnd vpwr scs8hd_diode_2
XANTENNA__082__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_135 vgnd vpwr scs8hd_decap_8
XFILLER_50_105 vgnd vpwr scs8hd_decap_12
XANTENNA__183__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__167__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_41_105 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_2_.latch/Q mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_25_14 vgnd vpwr scs8hd_decap_4
XFILLER_26_102 vgnd vpwr scs8hd_decap_8
XFILLER_26_113 vgnd vpwr scs8hd_decap_8
XFILLER_26_124 vgnd vpwr scs8hd_decap_12
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XANTENNA__093__A _112_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_105 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_5.LATCH_4_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__088__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_52_56 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _173_/HI mem_right_ipin_1.LATCH_5_.latch/Q
+ mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
X_171_ _171_/HI _171_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_120 vpwr vgnd scs8hd_fill_2
XFILLER_20_119 vgnd vpwr scs8hd_decap_12
XANTENNA__164__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_47_78 vpwr vgnd scs8hd_fill_2
XFILLER_8_39 vpwr vgnd scs8hd_fill_2
XFILLER_40_9 vgnd vpwr scs8hd_fill_1
X_154_ address[5] address[6] _154_/C _155_/A vgnd vpwr scs8hd_or3_4
X_085_ _121_/A _083_/X _085_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__191__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_2.LATCH_0_.latch data_in mem_right_ipin_2.LATCH_0_.latch/Q _098_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_37 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__B _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_33_25 vgnd vpwr scs8hd_fill_1
XFILLER_33_47 vgnd vpwr scs8hd_fill_1
XFILLER_3_126 vpwr vgnd scs8hd_fill_2
XFILLER_3_115 vpwr vgnd scs8hd_fill_2
XFILLER_3_104 vgnd vpwr scs8hd_decap_4
XFILLER_58_44 vgnd vpwr scs8hd_decap_12
X_137_ _137_/A _142_/B _137_/Y vgnd vpwr scs8hd_nor2_4
X_068_ _110_/A address[3] _143_/A _069_/A vgnd vpwr scs8hd_or3_4
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_4.LATCH_3_.latch data_in mem_right_ipin_4.LATCH_3_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__186__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_84 vpwr vgnd scs8hd_fill_2
XFILLER_9_71 vpwr vgnd scs8hd_fill_2
XFILLER_28_47 vpwr vgnd scs8hd_fill_2
XFILLER_44_57 vgnd vpwr scs8hd_decap_3
XFILLER_44_35 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_5_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_60_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__082__C _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_68 vpwr vgnd scs8hd_fill_2
XFILLER_39_57 vpwr vgnd scs8hd_fill_2
XFILLER_20_81 vpwr vgnd scs8hd_fill_2
XANTENNA__167__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_103 vgnd vpwr scs8hd_fill_1
XFILLER_50_117 vgnd vpwr scs8hd_decap_12
XFILLER_6_61 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_5.INVTX1_1_.scs8hd_inv_1 chany_top_in[2] mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_26_136 vgnd vpwr scs8hd_decap_8
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_41_25 vpwr vgnd scs8hd_fill_2
XANTENNA__093__B _096_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_106 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__194__A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_36 vgnd vpwr scs8hd_decap_6
XANTENNA__088__B _083_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_52_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_170_ _170_/HI _170_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_106 vgnd vpwr scs8hd_decap_4
XFILLER_26_91 vgnd vpwr scs8hd_fill_1
XFILLER_9_143 vgnd vpwr scs8hd_decap_3
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XANTENNA__189__A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_3_95 vgnd vpwr scs8hd_fill_1
XFILLER_3_51 vgnd vpwr scs8hd_decap_4
XFILLER_11_109 vgnd vpwr scs8hd_decap_8
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
XFILLER_22_49 vgnd vpwr scs8hd_decap_8
XANTENNA__099__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_57 vpwr vgnd scs8hd_fill_2
XFILLER_6_102 vgnd vpwr scs8hd_decap_12
X_153_ address[4] address[3] _066_/C _154_/C vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _172_/HI vgnd vpwr
+ scs8hd_diode_2
X_084_ _112_/A _083_/X _084_/Y vgnd vpwr scs8hd_nor2_4
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_37 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_7.LATCH_2_.latch data_in mem_right_ipin_7.LATCH_2_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_58_56 vgnd vpwr scs8hd_decap_12
X_136_ _136_/A _142_/B vgnd vpwr scs8hd_buf_1
X_067_ _066_/X _143_/A vgnd vpwr scs8hd_buf_1
Xmux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_2_.latch/Q mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_145 vgnd vpwr scs8hd_fill_1
XFILLER_28_26 vpwr vgnd scs8hd_fill_2
XANTENNA__096__B _096_/B vgnd vpwr scs8hd_diode_2
XFILLER_60_68 vgnd vpwr scs8hd_decap_3
XFILLER_5_19 vpwr vgnd scs8hd_fill_2
XFILLER_47_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_70 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_91 vgnd vpwr scs8hd_fill_1
X_119_ _119_/A _123_/B vgnd vpwr scs8hd_buf_1
XFILLER_38_145 vgnd vpwr scs8hd_fill_1
XANTENNA__197__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _172_/HI mem_right_ipin_0.LATCH_5_.latch/Q
+ mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_28 vgnd vpwr scs8hd_fill_1
XFILLER_39_36 vpwr vgnd scs8hd_fill_2
XFILLER_29_145 vgnd vpwr scs8hd_fill_1
XFILLER_20_60 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_25_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_17_126 vpwr vgnd scs8hd_fill_2
XFILLER_31_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_18 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_91 vgnd vpwr scs8hd_fill_1
XFILLER_47_36 vpwr vgnd scs8hd_fill_2
XFILLER_47_25 vpwr vgnd scs8hd_fill_2
XANTENNA__099__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_6_114 vgnd vpwr scs8hd_decap_12
X_152_ enable _066_/C vgnd vpwr scs8hd_inv_8
X_083_ _082_/X _083_/X vgnd vpwr scs8hd_buf_1
Xmux_right_ipin_4.INVTX1_5_.scs8hd_inv_1 chany_top_in[6] mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_59_121 vgnd vpwr scs8hd_fill_1
XFILLER_58_68 vgnd vpwr scs8hd_decap_8
X_066_ address[5] address[6] _066_/C _066_/X vgnd vpwr scs8hd_or3_4
X_135_ address[5] _127_/B _066_/C _143_/B _136_/A vgnd vpwr scs8hd_or4_4
XANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_6 vpwr vgnd scs8hd_fill_2
XFILLER_48_90 vpwr vgnd scs8hd_fill_2
XFILLER_9_95 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XFILLER_62_105 vgnd vpwr scs8hd_decap_12
XFILLER_47_135 vgnd vpwr scs8hd_decap_8
XFILLER_18_60 vpwr vgnd scs8hd_fill_2
XFILLER_34_81 vpwr vgnd scs8hd_fill_2
X_118_ _110_/A _118_/B _102_/A _119_/A vgnd vpwr scs8hd_or3_4
XFILLER_38_113 vgnd vpwr scs8hd_decap_12
XFILLER_38_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.LATCH_3_.latch data_in mem_right_ipin_0.LATCH_3_.latch/Q _074_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_92 vgnd vpwr scs8hd_fill_1
XFILLER_6_41 vpwr vgnd scs8hd_fill_2
XFILLER_6_85 vgnd vpwr scs8hd_fill_1
XFILLER_6_74 vgnd vpwr scs8hd_decap_4
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_17_105 vgnd vpwr scs8hd_decap_4
XFILLER_32_119 vgnd vpwr scs8hd_decap_8
XFILLER_15_83 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_130 vpwr vgnd scs8hd_fill_2
XFILLER_52_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_130 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_2_.latch/Q mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_112 vgnd vpwr scs8hd_decap_8
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_42_81 vpwr vgnd scs8hd_fill_2
XFILLER_3_75 vpwr vgnd scs8hd_fill_2
XFILLER_3_31 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_0_.latch/Q mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_15 vgnd vpwr scs8hd_decap_6
XANTENNA__099__C _066_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_126 vgnd vpwr scs8hd_decap_12
X_082_ _110_/A _118_/B _143_/A _082_/X vgnd vpwr scs8hd_or3_4
XFILLER_12_84 vgnd vpwr scs8hd_decap_6
X_151_ _137_/A _112_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _173_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_92 vgnd vpwr scs8hd_fill_1
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[2] mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_ipin_7.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_18 vpwr vgnd scs8hd_fill_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_065_ address[4] _110_/A vgnd vpwr scs8hd_inv_8
X_134_ _142_/A _131_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
XFILLER_31_8 vpwr vgnd scs8hd_fill_2
XFILLER_0_43 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_76 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
XFILLER_62_117 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_3.LATCH_2_.latch data_in mem_right_ipin_3.LATCH_2_.latch/Q _107_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_117_ _125_/A _116_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_60 vpwr vgnd scs8hd_fill_2
XFILLER_50_81 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_125 vgnd vpwr scs8hd_decap_12
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
XFILLER_55_59 vpwr vgnd scs8hd_fill_2
XFILLER_55_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_5.LATCH_5_.latch data_in mem_right_ipin_5.LATCH_5_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_106 vgnd vpwr scs8hd_decap_12
XFILLER_45_81 vpwr vgnd scs8hd_fill_2
XFILLER_6_64 vgnd vpwr scs8hd_fill_1
XFILLER_6_53 vgnd vpwr scs8hd_fill_1
XFILLER_41_109 vgnd vpwr scs8hd_decap_12
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_8 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_5.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_23_109 vgnd vpwr scs8hd_fill_1
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_142 vgnd vpwr scs8hd_decap_4
XFILLER_9_135 vgnd vpwr scs8hd_decap_8
XFILLER_13_120 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_0.LATCH_3_.latch data_in mem_left_ipin_0.LATCH_3_.latch/Q _163_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_83 vgnd vpwr scs8hd_fill_1
XFILLER_42_93 vgnd vpwr scs8hd_decap_3
XFILLER_3_10 vpwr vgnd scs8hd_fill_2
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
X_150_ _149_/X _137_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_138 vgnd vpwr scs8hd_decap_8
X_081_ address[3] _118_/B vgnd vpwr scs8hd_inv_8
XFILLER_10_145 vgnd vpwr scs8hd_fill_1
XFILLER_12_41 vgnd vpwr scs8hd_decap_4
XFILLER_37_71 vpwr vgnd scs8hd_fill_2
XFILLER_45_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_119 vgnd vpwr scs8hd_decap_3
XFILLER_59_145 vgnd vpwr scs8hd_fill_1
XFILLER_59_123 vgnd vpwr scs8hd_decap_8
XFILLER_59_101 vgnd vpwr scs8hd_decap_12
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_40 vpwr vgnd scs8hd_fill_2
XFILLER_23_73 vpwr vgnd scs8hd_fill_2
X_133_ _141_/A _131_/B _133_/Y vgnd vpwr scs8hd_nor2_4
X_064_ _169_/A _142_/A _064_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_2_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_88 vgnd vpwr scs8hd_decap_3
XFILLER_9_31 vgnd vpwr scs8hd_decap_4
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
XFILLER_28_18 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_6.LATCH_1_.latch data_in mem_right_ipin_6.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_44_39 vgnd vpwr scs8hd_decap_4
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_62_129 vgnd vpwr scs8hd_decap_12
XFILLER_18_84 vgnd vpwr scs8hd_decap_6
XFILLER_50_93 vgnd vpwr scs8hd_decap_12
X_116_ _124_/A _116_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_137 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_2_.latch/Q mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_126 vpwr vgnd scs8hd_fill_2
XFILLER_29_137 vpwr vgnd scs8hd_fill_2
XFILLER_55_27 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.INVTX1_5_.scs8hd_inv_1 chany_top_in[6] mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_85 vgnd vpwr scs8hd_decap_4
XFILLER_35_118 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_15_41 vpwr vgnd scs8hd_fill_2
XFILLER_15_52 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[7] mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_62 vpwr vgnd scs8hd_fill_2
XFILLER_31_73 vpwr vgnd scs8hd_fill_2
XANTENNA__102__B _143_/B vgnd vpwr scs8hd_diode_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_1.LATCH_3_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__113__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_88 vgnd vpwr scs8hd_decap_4
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
X_080_ _125_/A _069_/X _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_102 vpwr vgnd scs8hd_fill_2
XFILLER_10_113 vgnd vpwr scs8hd_decap_12
XFILLER_12_20 vpwr vgnd scs8hd_fill_2
XFILLER_5_3 vgnd vpwr scs8hd_decap_3
XFILLER_12_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _174_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__108__A _124_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_135 vpwr vgnd scs8hd_fill_2
XFILLER_59_113 vgnd vpwr scs8hd_decap_8
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
X_063_ _062_/X _142_/A vgnd vpwr scs8hd_buf_1
X_132_ _140_/A _131_/B _132_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_9_54 vpwr vgnd scs8hd_fill_2
XFILLER_56_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_72 vgnd vpwr scs8hd_decap_6
XFILLER_50_61 vgnd vpwr scs8hd_decap_8
X_115_ _123_/A _116_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__B _108_/B vgnd vpwr scs8hd_diode_2
XFILLER_59_92 vgnd vpwr scs8hd_fill_1
XFILLER_59_70 vgnd vpwr scs8hd_fill_1
XFILLER_22_6 vpwr vgnd scs8hd_fill_2
XANTENNA__121__A _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_39 vgnd vpwr scs8hd_decap_12
XFILLER_29_105 vpwr vgnd scs8hd_fill_2
XFILLER_52_141 vgnd vpwr scs8hd_decap_4
XFILLER_29_51 vgnd vpwr scs8hd_decap_4
XFILLER_29_62 vpwr vgnd scs8hd_fill_2
XFILLER_29_73 vpwr vgnd scs8hd_fill_2
XFILLER_29_95 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__116__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_88 vgnd vpwr scs8hd_decap_4
XFILLER_15_20 vpwr vgnd scs8hd_fill_2
XFILLER_15_75 vpwr vgnd scs8hd_fill_2
XFILLER_15_97 vpwr vgnd scs8hd_fill_2
XFILLER_56_93 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_1.LATCH_5_.latch data_in mem_right_ipin_1.LATCH_5_.latch/Q _084_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

