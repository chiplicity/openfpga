* NGSPICE file created from sb_1__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

.subckt sb_1__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_bottom_in[0]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] data_in enable left_bottom_grid_pin_12_
+ left_top_grid_pin_11_ left_top_grid_pin_13_ left_top_grid_pin_15_ left_top_grid_pin_1_
+ left_top_grid_pin_3_ left_top_grid_pin_5_ left_top_grid_pin_7_ left_top_grid_pin_9_
+ right_bottom_grid_pin_12_ right_top_grid_pin_11_ right_top_grid_pin_13_ right_top_grid_pin_15_
+ right_top_grid_pin_1_ right_top_grid_pin_3_ right_top_grid_pin_5_ right_top_grid_pin_7_
+ right_top_grid_pin_9_ vpwr vgnd
XFILLER_22_166 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_41 vgnd vpwr scs8hd_decap_3
XFILLER_9_115 vgnd vpwr scs8hd_fill_1
XFILLER_13_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__113__B _113_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_258 vgnd vpwr scs8hd_decap_12
XFILLER_27_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
XFILLER_33_206 vpwr vgnd scs8hd_fill_2
XANTENNA__108__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _110_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_32_250 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_131_ _110_/A _131_/B _131_/Y vgnd vpwr scs8hd_nor2_4
X_062_ address[3] _134_/A vgnd vpwr scs8hd_inv_8
XFILLER_23_75 vpwr vgnd scs8hd_fill_2
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XFILLER_17_9 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _112_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _190_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _066_/Y mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_264 vgnd vpwr scs8hd_decap_8
XFILLER_18_97 vpwr vgnd scs8hd_fill_2
X_114_ _086_/A _118_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XANTENNA__105__C _105_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__121__B _122_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_106 vpwr vgnd scs8hd_fill_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_29_30 vpwr vgnd scs8hd_fill_2
XFILLER_28_172 vgnd vpwr scs8hd_decap_6
XANTENNA__116__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_78 vgnd vpwr scs8hd_decap_12
XANTENNA__132__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_4
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _103_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_194 vpwr vgnd scs8hd_fill_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_15_10 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_42 vpwr vgnd scs8hd_fill_2
XFILLER_0_230 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _080_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_274 vgnd vpwr scs8hd_decap_3
XFILLER_31_156 vpwr vgnd scs8hd_fill_2
XFILLER_31_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_186 vgnd vpwr scs8hd_decap_4
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _113_/A vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_223 vpwr vgnd scs8hd_fill_2
XFILLER_39_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_64 vgnd vpwr scs8hd_decap_8
XFILLER_13_134 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XANTENNA__113__C _085_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_104 vgnd vpwr scs8hd_fill_1
XFILLER_10_137 vgnd vpwr scs8hd_decap_12
XFILLER_10_159 vpwr vgnd scs8hd_fill_2
XFILLER_12_77 vpwr vgnd scs8hd_fill_2
XFILLER_12_88 vgnd vpwr scs8hd_fill_1
XFILLER_37_85 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__124__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _066_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__140__A address[6] vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_262 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_15_207 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_130_ _090_/B _131_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_061_ address[5] _113_/B vgnd vpwr scs8hd_inv_8
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XANTENNA__119__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_23 vgnd vpwr scs8hd_fill_1
XFILLER_9_67 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _082_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_4
XFILLER_34_75 vgnd vpwr scs8hd_decap_6
X_113_ _113_/A _113_/B _085_/C _118_/B vgnd vpwr scs8hd_or3_4
XFILLER_11_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XFILLER_38_129 vgnd vpwr scs8hd_decap_6
XFILLER_15_7 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_7_ mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_118 vgnd vpwr scs8hd_fill_1
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_66 vpwr vgnd scs8hd_fill_2
XFILLER_29_53 vgnd vpwr scs8hd_decap_4
XFILLER_29_42 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_151 vpwr vgnd scs8hd_fill_2
XANTENNA__132__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_132 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vpwr vgnd scs8hd_fill_2
XFILLER_34_165 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_121 vgnd vpwr scs8hd_fill_1
XFILLER_31_76 vpwr vgnd scs8hd_fill_2
XFILLER_15_77 vgnd vpwr scs8hd_decap_4
XFILLER_31_98 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_5_ mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XFILLER_31_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _068_/A vgnd
+ vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_143 vgnd vpwr scs8hd_decap_8
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XFILLER_16_176 vgnd vpwr scs8hd_fill_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__127__B _113_/B vgnd vpwr scs8hd_diode_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_39_257 vgnd vpwr scs8hd_decap_12
XFILLER_26_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _186_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_8_150 vgnd vpwr scs8hd_decap_3
XFILLER_27_238 vgnd vpwr scs8hd_decap_6
XFILLER_10_116 vpwr vgnd scs8hd_fill_2
XFILLER_6_109 vgnd vpwr scs8hd_decap_12
XFILLER_10_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_219 vpwr vgnd scs8hd_fill_2
XANTENNA__140__B _113_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_274 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_219 vpwr vgnd scs8hd_fill_2
XFILLER_23_33 vgnd vpwr scs8hd_decap_4
XFILLER_23_252 vgnd vpwr scs8hd_decap_3
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
X_060_ address[6] _113_/A vgnd vpwr scs8hd_inv_8
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _066_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_48 vgnd vpwr scs8hd_decap_12
XFILLER_9_35 vpwr vgnd scs8hd_fill_2
X_189_ _189_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__135__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA__151__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_200 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__061__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_77 vpwr vgnd scs8hd_fill_2
X_112_ _112_/A _110_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_270 vgnd vpwr scs8hd_decap_4
XFILLER_37_196 vgnd vpwr scs8hd_decap_8
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_87 vgnd vpwr scs8hd_decap_4
XFILLER_28_163 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_251 vpwr vgnd scs8hd_fill_2
XFILLER_34_111 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_141 vpwr vgnd scs8hd_fill_2
XFILLER_19_163 vpwr vgnd scs8hd_fill_2
XFILLER_34_177 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_144 vpwr vgnd scs8hd_fill_2
XFILLER_15_23 vpwr vgnd scs8hd_fill_2
XFILLER_15_34 vpwr vgnd scs8hd_fill_2
XFILLER_15_45 vpwr vgnd scs8hd_fill_2
XFILLER_31_22 vgnd vpwr scs8hd_decap_3
XFILLER_31_11 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _165_/HI mem_right_track_0.LATCH_2_.latch/Q
+ mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_16_122 vpwr vgnd scs8hd_fill_2
XFILLER_31_169 vgnd vpwr scs8hd_decap_4
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _106_/C vgnd vpwr scs8hd_diode_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _113_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vpwr vgnd scs8hd_fill_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_88 vpwr vgnd scs8hd_fill_2
XFILLER_9_107 vpwr vgnd scs8hd_fill_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_169 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__138__B _113_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_217 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__064__A enable vgnd vpwr scs8hd_diode_2
XFILLER_12_57 vgnd vpwr scs8hd_decap_4
XFILLER_37_10 vgnd vpwr scs8hd_decap_12
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XANTENNA__140__C _120_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__149__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_250 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _081_/A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XANTENNA__059__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_23_12 vpwr vgnd scs8hd_fill_2
XFILLER_23_56 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_9_58 vgnd vpwr scs8hd_decap_3
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_188_ _188_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA__135__C _143_/C vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_6
XANTENNA__151__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_20_212 vpwr vgnd scs8hd_fill_2
XFILLER_18_56 vpwr vgnd scs8hd_fill_2
XFILLER_11_201 vgnd vpwr scs8hd_decap_12
X_111_ _118_/A _110_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__146__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_37_131 vpwr vgnd scs8hd_fill_2
XANTENNA__072__A _072_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_46 vgnd vpwr scs8hd_decap_3
XFILLER_28_131 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_37 vgnd vpwr scs8hd_decap_4
XFILLER_6_15 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_7 vgnd vpwr scs8hd_decap_3
XFILLER_34_189 vpwr vgnd scs8hd_fill_2
XFILLER_34_145 vgnd vpwr scs8hd_decap_8
XFILLER_34_101 vgnd vpwr scs8hd_fill_1
XFILLER_19_175 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_40_137 vgnd vpwr scs8hd_decap_12
XFILLER_25_178 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_0_244 vgnd vpwr scs8hd_decap_4
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__C _143_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_204 vgnd vpwr scs8hd_decap_12
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_104 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_270 vgnd vpwr scs8hd_decap_4
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_126 vpwr vgnd scs8hd_fill_2
XFILLER_13_148 vpwr vgnd scs8hd_fill_2
XFILLER_36_229 vgnd vpwr scs8hd_decap_12
XFILLER_36_218 vpwr vgnd scs8hd_fill_2
XANTENNA__138__C _085_/C vgnd vpwr scs8hd_diode_2
XANTENNA__170__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_229 vgnd vpwr scs8hd_decap_3
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _110_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__080__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_22 vgnd vpwr scs8hd_decap_12
XFILLER_18_218 vpwr vgnd scs8hd_fill_2
XFILLER_18_229 vgnd vpwr scs8hd_decap_8
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
XFILLER_26_240 vgnd vpwr scs8hd_decap_8
XANTENNA__140__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__149__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_243 vgnd vpwr scs8hd_fill_1
XANTENNA__075__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA__135__D _083_/C vgnd vpwr scs8hd_diode_2
XANTENNA__151__C _143_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_110_ _110_/A _110_/B _110_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_213 vgnd vpwr scs8hd_decap_12
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _079_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__146__C _085_/C vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_121 vgnd vpwr scs8hd_fill_1
XFILLER_20_58 vpwr vgnd scs8hd_fill_2
XFILLER_29_78 vpwr vgnd scs8hd_fill_2
XFILLER_29_34 vpwr vgnd scs8hd_fill_2
XFILLER_28_187 vpwr vgnd scs8hd_fill_2
XFILLER_28_110 vgnd vpwr scs8hd_fill_1
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_275 vpwr vgnd scs8hd_fill_2
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XFILLER_34_157 vpwr vgnd scs8hd_fill_2
XANTENNA__173__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_25_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_149 vgnd vpwr scs8hd_decap_4
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XANTENNA__083__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_138 vpwr vgnd scs8hd_fill_2
XFILLER_24_190 vgnd vpwr scs8hd_decap_4
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _065_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__D _083_/C vgnd vpwr scs8hd_diode_2
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_216 vgnd vpwr scs8hd_decap_3
XFILLER_39_227 vgnd vpwr scs8hd_decap_12
XANTENNA__168__A _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_149 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_26_46 vgnd vpwr scs8hd_decap_3
XFILLER_13_138 vgnd vpwr scs8hd_fill_1
XANTENNA__078__A _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__138__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_16_90 vpwr vgnd scs8hd_fill_2
XFILLER_12_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _081_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_9_ mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_89 vgnd vpwr scs8hd_decap_12
XFILLER_37_34 vgnd vpwr scs8hd_decap_12
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _094_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__149__C _106_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_263 vpwr vgnd scs8hd_fill_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_4_71 vgnd vpwr scs8hd_decap_12
XFILLER_23_222 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA__151__D _083_/C vgnd vpwr scs8hd_diode_2
X_186_ _186_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_36_6 vgnd vpwr scs8hd_decap_12
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_25 vpwr vgnd scs8hd_fill_2
XFILLER_18_36 vgnd vpwr scs8hd_fill_1
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_4
XFILLER_11_225 vgnd vpwr scs8hd_decap_12
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _067_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_251 vgnd vpwr scs8hd_decap_4
X_169_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA__146__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_166 vgnd vpwr scs8hd_decap_12
XFILLER_37_144 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_7.LATCH_0_.latch data_in _072_/A _142_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_13 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_114 vgnd vpwr scs8hd_decap_4
XFILLER_31_36 vgnd vpwr scs8hd_decap_4
XANTENNA__083__B _083_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_169 vgnd vpwr scs8hd_decap_4
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_239 vgnd vpwr scs8hd_decap_4
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__184__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_58 vgnd vpwr scs8hd_decap_4
XANTENNA__094__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_172 vgnd vpwr scs8hd_decap_4
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XFILLER_8_121 vgnd vpwr scs8hd_decap_3
XANTENNA__179__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_12_27 vgnd vpwr scs8hd_fill_1
XFILLER_12_49 vpwr vgnd scs8hd_fill_2
XFILLER_37_79 vgnd vpwr scs8hd_decap_3
XFILLER_37_46 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__089__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XFILLER_32_212 vpwr vgnd scs8hd_fill_2
XFILLER_32_201 vpwr vgnd scs8hd_fill_2
XANTENNA__149__D _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_4_83 vgnd vpwr scs8hd_decap_8
XFILLER_3_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XANTENNA__091__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_17 vgnd vpwr scs8hd_decap_6
XFILLER_14_212 vpwr vgnd scs8hd_fill_2
X_185_ _185_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_9_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_204 vpwr vgnd scs8hd_fill_2
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XANTENNA__086__B _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_237 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _079_/A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
X_168_ _168_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
X_099_ _086_/A _103_/B _099_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_178 vgnd vpwr scs8hd_decap_4
XFILLER_37_123 vgnd vpwr scs8hd_decap_8
XFILLER_37_101 vgnd vpwr scs8hd_decap_12
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
XFILLER_28_145 vgnd vpwr scs8hd_decap_4
XFILLER_28_123 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A _134_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_15.LATCH_0_.latch data_in _080_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_255 vgnd vpwr scs8hd_decap_12
XFILLER_10_82 vgnd vpwr scs8hd_decap_6
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_123 vgnd vpwr scs8hd_fill_1
XFILLER_19_145 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_4
XFILLER_33_170 vpwr vgnd scs8hd_fill_2
XFILLER_25_148 vgnd vpwr scs8hd_decap_4
XFILLER_25_126 vpwr vgnd scs8hd_fill_2
XFILLER_15_27 vgnd vpwr scs8hd_decap_4
XFILLER_15_49 vpwr vgnd scs8hd_fill_2
XANTENNA__083__C _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_236 vgnd vpwr scs8hd_fill_1
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XFILLER_24_170 vgnd vpwr scs8hd_decap_8
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_22_129 vgnd vpwr scs8hd_decap_3
XFILLER_30_195 vpwr vgnd scs8hd_fill_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XANTENNA__094__B _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_4
XFILLER_3_19 vgnd vpwr scs8hd_decap_12
XFILLER_32_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XFILLER_8_111 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__089__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_37_58 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _102_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_210 vpwr vgnd scs8hd_fill_2
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _192_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_232 vgnd vpwr scs8hd_decap_4
XFILLER_17_243 vgnd vpwr scs8hd_fill_1
XFILLER_17_254 vgnd vpwr scs8hd_fill_1
XFILLER_23_235 vpwr vgnd scs8hd_fill_2
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XANTENNA__091__C address[0] vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_224 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_11_ mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_184_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_13_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_249 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_91 vgnd vpwr scs8hd_fill_1
X_167_ _167_/HI _167_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_271 vgnd vpwr scs8hd_decap_4
X_098_ address[6] address[5] _120_/C _103_/B vgnd vpwr scs8hd_or3_4
XFILLER_37_113 vgnd vpwr scs8hd_decap_8
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_168 vpwr vgnd scs8hd_fill_2
XFILLER_28_113 vgnd vpwr scs8hd_fill_1
XANTENNA__097__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_267 vgnd vpwr scs8hd_decap_8
XFILLER_19_102 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_3.LATCH_0_.latch data_in _068_/A _138_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_93 vpwr vgnd scs8hd_fill_2
XFILLER_11_7 vpwr vgnd scs8hd_fill_2
XFILLER_30_130 vgnd vpwr scs8hd_decap_6
XPHY_2 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _082_/A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_22_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _082_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_62 vpwr vgnd scs8hd_fill_2
XFILLER_7_51 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_274 vgnd vpwr scs8hd_fill_1
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _163_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_274 vgnd vpwr scs8hd_decap_3
XFILLER_16_71 vpwr vgnd scs8hd_fill_2
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
XFILLER_35_233 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__089__C _083_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_15.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_81 vgnd vpwr scs8hd_decap_6
XFILLER_17_211 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _176_/A vgnd vpwr scs8hd_inv_1
XFILLER_23_39 vpwr vgnd scs8hd_fill_2
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _068_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_236 vgnd vpwr scs8hd_decap_8
XFILLER_14_247 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_50 vpwr vgnd scs8hd_fill_2
XFILLER_13_83 vgnd vpwr scs8hd_decap_4
X_183_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_49 vgnd vpwr scs8hd_decap_6
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _164_/HI vgnd vpwr
+ scs8hd_diode_2
X_166_ _166_/HI _166_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_097_ _134_/A address[4] _105_/C _120_/C vgnd vpwr scs8hd_or3_4
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_38 vpwr vgnd scs8hd_fill_2
XANTENNA__097__C _105_/C vgnd vpwr scs8hd_diode_2
XFILLER_19_60 vgnd vpwr scs8hd_fill_1
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_34_128 vpwr vgnd scs8hd_fill_2
X_149_ _113_/A address[5] _106_/C _083_/C _149_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _066_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _188_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_106 vpwr vgnd scs8hd_fill_2
XFILLER_16_117 vgnd vpwr scs8hd_decap_3
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_track_11.LATCH_0_.latch data_in _076_/A _146_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _070_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_142 vpwr vgnd scs8hd_fill_2
XFILLER_29_231 vpwr vgnd scs8hd_fill_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_6
XFILLER_12_186 vpwr vgnd scs8hd_fill_2
XFILLER_35_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_201 vgnd vpwr scs8hd_fill_1
XFILLER_17_245 vgnd vpwr scs8hd_decap_3
XFILLER_17_267 vgnd vpwr scs8hd_decap_8
XFILLER_32_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_42 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_204 vgnd vpwr scs8hd_decap_6
X_182_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_259 vgnd vpwr scs8hd_decap_12
XFILLER_29_9 vgnd vpwr scs8hd_fill_1
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _088_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.INVTX1_1_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _068_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_165_ _165_/HI _165_/LO vgnd vpwr scs8hd_conb_1
XFILLER_24_50 vpwr vgnd scs8hd_fill_2
XFILLER_10_251 vgnd vpwr scs8hd_decap_4
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ _088_/A _112_/A _096_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_148 vgnd vpwr scs8hd_decap_12
XFILLER_27_6 vpwr vgnd scs8hd_fill_2
XFILLER_1_98 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.INVTX1_0_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_17 vpwr vgnd scs8hd_fill_2
XFILLER_10_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_159 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _077_/A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_148_ _113_/A address[5] _120_/C address[0] _148_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_25_3 vpwr vgnd scs8hd_fill_2
X_079_ _079_/A _079_/Y vgnd vpwr scs8hd_inv_8
XFILLER_25_118 vgnd vpwr scs8hd_fill_1
XFILLER_33_184 vpwr vgnd scs8hd_fill_2
XFILLER_31_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_140 vpwr vgnd scs8hd_fill_2
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A right_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_40 vpwr vgnd scs8hd_fill_2
XFILLER_21_62 vpwr vgnd scs8hd_fill_2
XFILLER_21_73 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_3_ mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_154 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_162 vpwr vgnd scs8hd_fill_2
XFILLER_15_184 vgnd vpwr scs8hd_decap_4
XFILLER_7_86 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_110 vpwr vgnd scs8hd_fill_2
XFILLER_21_176 vgnd vpwr scs8hd_fill_1
XFILLER_29_254 vgnd vpwr scs8hd_decap_12
XFILLER_8_103 vpwr vgnd scs8hd_fill_2
XFILLER_12_110 vpwr vgnd scs8hd_fill_2
XFILLER_12_165 vgnd vpwr scs8hd_decap_8
XFILLER_16_84 vgnd vpwr scs8hd_decap_4
XFILLER_32_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _118_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_7_ mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _157_/HI _081_/Y mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_205 vgnd vpwr scs8hd_decap_4
XFILLER_4_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_205 vpwr vgnd scs8hd_fill_2
X_181_ _181_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__100__B _103_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_208 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_253 vpwr vgnd scs8hd_fill_2
XFILLER_18_19 vgnd vpwr scs8hd_decap_4
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _109_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_40 vgnd vpwr scs8hd_fill_1
XFILLER_40_61 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_164_ _164_/HI _164_/LO vgnd vpwr scs8hd_conb_1
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
XFILLER_24_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr
+ scs8hd_diode_2
X_095_ address[1] address[2] address[0] _112_/A vgnd vpwr scs8hd_or3_4
XANTENNA__111__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_28_127 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_11.INVTX1_1_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_160 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_40 vgnd vpwr scs8hd_decap_3
XFILLER_35_72 vpwr vgnd scs8hd_fill_2
XFILLER_27_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_147_ _113_/A address[5] _120_/C _083_/C _147_/Y vgnd vpwr scs8hd_nor4_4
X_078_ _078_/A _078_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__106__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_3
XFILLER_18_171 vgnd vpwr scs8hd_decap_3
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_196 vpwr vgnd scs8hd_fill_2
XFILLER_24_152 vgnd vpwr scs8hd_fill_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_111 vgnd vpwr scs8hd_decap_6
XFILLER_38_211 vgnd vpwr scs8hd_decap_3
XFILLER_21_155 vpwr vgnd scs8hd_fill_2
XFILLER_21_188 vgnd vpwr scs8hd_fill_1
XFILLER_29_266 vgnd vpwr scs8hd_decap_8
XFILLER_16_41 vpwr vgnd scs8hd_fill_2
XFILLER_32_62 vpwr vgnd scs8hd_fill_2
XFILLER_8_126 vgnd vpwr scs8hd_decap_12
XFILLER_12_199 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__103__B _103_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _080_/A mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_8
XFILLER_32_228 vgnd vpwr scs8hd_decap_8
XFILLER_27_73 vpwr vgnd scs8hd_fill_2
XFILLER_17_236 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__114__A _086_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_239 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_180_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__109__A _090_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_73 vgnd vpwr scs8hd_decap_12
X_163_ _163_/HI _163_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
X_094_ _088_/A _118_/A _094_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__111__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _081_/Y vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _092_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_106 vgnd vpwr scs8hd_decap_4
XFILLER_10_32 vpwr vgnd scs8hd_fill_2
XFILLER_10_65 vpwr vgnd scs8hd_fill_2
XFILLER_27_161 vpwr vgnd scs8hd_fill_2
XFILLER_19_52 vpwr vgnd scs8hd_fill_2
XFILLER_35_95 vpwr vgnd scs8hd_fill_2
XFILLER_35_62 vgnd vpwr scs8hd_fill_1
XANTENNA__122__A _088_/B vgnd vpwr scs8hd_diode_2
X_077_ _077_/A _077_/Y vgnd vpwr scs8hd_inv_8
X_146_ _113_/A address[5] _085_/C address[0] _146_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__106__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_33_175 vpwr vgnd scs8hd_fill_2
XFILLER_33_164 vgnd vpwr scs8hd_decap_4
XFILLER_18_183 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_97 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_189 vgnd vpwr scs8hd_decap_4
XFILLER_30_145 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_66 vgnd vpwr scs8hd_decap_12
XFILLER_7_55 vgnd vpwr scs8hd_decap_4
XFILLER_7_22 vgnd vpwr scs8hd_decap_3
XFILLER_30_3 vpwr vgnd scs8hd_fill_2
X_129_ _088_/B _131_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _067_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _073_/A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
XFILLER_21_134 vpwr vgnd scs8hd_fill_2
XFILLER_29_212 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_75 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_7.LATCH_1_.latch data_in _071_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_138 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_145 vgnd vpwr scs8hd_decap_8
XFILLER_35_204 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _167_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_171 vgnd vpwr scs8hd_decap_12
XFILLER_34_270 vgnd vpwr scs8hd_decap_4
XFILLER_26_215 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_30 vpwr vgnd scs8hd_fill_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_17_259 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _090_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_218 vpwr vgnd scs8hd_fill_2
XFILLER_31_273 vgnd vpwr scs8hd_decap_4
XFILLER_13_54 vgnd vpwr scs8hd_decap_4
XFILLER_22_273 vpwr vgnd scs8hd_fill_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__109__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_200 vgnd vpwr scs8hd_decap_12
XANTENNA__125__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_192 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_162_ _162_/HI _162_/LO vgnd vpwr scs8hd_conb_1
XFILLER_40_85 vgnd vpwr scs8hd_decap_6
XFILLER_6_258 vgnd vpwr scs8hd_decap_12
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ address[1] address[2] _083_/C _118_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _069_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_55 vgnd vpwr scs8hd_fill_1
XFILLER_10_88 vgnd vpwr scs8hd_fill_1
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_19_75 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__106__C _106_/C vgnd vpwr scs8hd_diode_2
X_145_ _113_/A address[5] _085_/C _083_/C _145_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_32_7 vgnd vpwr scs8hd_decap_12
X_076_ _076_/A _076_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__122__B _122_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _153_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_143 vpwr vgnd scs8hd_fill_2
XFILLER_30_168 vgnd vpwr scs8hd_decap_12
XANTENNA__117__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_89 vpwr vgnd scs8hd_fill_2
XFILLER_7_78 vgnd vpwr scs8hd_decap_8
XFILLER_7_34 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A _112_/A vgnd vpwr scs8hd_diode_2
X_128_ _086_/A _131_/B _128_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_3
X_059_ address[0] _083_/C vgnd vpwr scs8hd_inv_8
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _075_/A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_29_235 vpwr vgnd scs8hd_fill_2
XFILLER_12_124 vpwr vgnd scs8hd_fill_2
XFILLER_16_54 vgnd vpwr scs8hd_decap_6
XFILLER_35_249 vgnd vpwr scs8hd_decap_6
XFILLER_35_216 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_15.LATCH_1_.latch data_in _079_/A _149_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__128__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A left_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_271 vgnd vpwr scs8hd_decap_4
XFILLER_31_230 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _156_/HI _079_/Y mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_241 vgnd vpwr scs8hd_decap_12
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_212 vgnd vpwr scs8hd_decap_12
XFILLER_9_245 vgnd vpwr scs8hd_decap_8
XFILLER_13_230 vgnd vpwr scs8hd_decap_12
XFILLER_13_263 vgnd vpwr scs8hd_decap_12
XANTENNA__125__B _122_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A address[6] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_182 vgnd vpwr scs8hd_fill_1
XFILLER_24_54 vpwr vgnd scs8hd_fill_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_8
XFILLER_24_10 vpwr vgnd scs8hd_fill_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
X_161_ _161_/HI _161_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_092_ _088_/A _110_/A _092_/Y vgnd vpwr scs8hd_nor2_4
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _101_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__136__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_45 vpwr vgnd scs8hd_fill_2
XFILLER_19_98 vgnd vpwr scs8hd_decap_4
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XFILLER_35_31 vgnd vpwr scs8hd_decap_12
XFILLER_27_174 vgnd vpwr scs8hd_decap_3
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_075_ _075_/A _075_/Y vgnd vpwr scs8hd_inv_8
X_144_ address[6] _113_/B _143_/C address[0] _144_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_100 vpwr vgnd scs8hd_fill_2
XFILLER_18_130 vpwr vgnd scs8hd_fill_2
XFILLER_18_152 vgnd vpwr scs8hd_fill_1
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XFILLER_33_188 vgnd vpwr scs8hd_decap_3
XFILLER_24_166 vpwr vgnd scs8hd_fill_2
XFILLER_24_144 vgnd vpwr scs8hd_decap_8
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_77 vgnd vpwr scs8hd_decap_3
XFILLER_30_158 vgnd vpwr scs8hd_fill_1
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_166 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_058_ address[2] _083_/B vgnd vpwr scs8hd_inv_8
XANTENNA__133__B _131_/B vgnd vpwr scs8hd_diode_2
X_127_ _113_/A _113_/B _106_/C _131_/B vgnd vpwr scs8hd_or3_4
XFILLER_38_203 vgnd vpwr scs8hd_decap_8
XFILLER_16_3 vgnd vpwr scs8hd_decap_3
XFILLER_38_258 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _194_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_107 vgnd vpwr scs8hd_decap_4
XFILLER_12_114 vgnd vpwr scs8hd_decap_8
XFILLER_32_87 vgnd vpwr scs8hd_decap_4
XFILLER_32_43 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__144__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
XFILLER_26_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_209 vgnd vpwr scs8hd_fill_1
XFILLER_27_87 vgnd vpwr scs8hd_fill_1
XFILLER_27_10 vgnd vpwr scs8hd_decap_3
XFILLER_25_250 vgnd vpwr scs8hd_decap_12
XFILLER_17_228 vpwr vgnd scs8hd_fill_2
XFILLER_17_239 vgnd vpwr scs8hd_decap_4
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_4_47 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_3.LATCH_1_.latch data_in _067_/A _137_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__139__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_13_45 vgnd vpwr scs8hd_decap_3
XFILLER_22_253 vgnd vpwr scs8hd_decap_12
XFILLER_13_89 vpwr vgnd scs8hd_fill_2
XFILLER_38_64 vgnd vpwr scs8hd_decap_12
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _078_/A mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_13_242 vpwr vgnd scs8hd_fill_2
XFILLER_9_224 vgnd vpwr scs8hd_decap_12
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XFILLER_13_275 vpwr vgnd scs8hd_fill_2
XANTENNA__141__B _113_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_88 vpwr vgnd scs8hd_fill_2
X_091_ _091_/A address[2] address[0] _110_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
X_160_ _160_/HI _160_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XANTENNA__136__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_120 vgnd vpwr scs8hd_decap_3
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_13 vpwr vgnd scs8hd_fill_2
XFILLER_10_24 vgnd vpwr scs8hd_fill_1
XANTENNA__062__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_27_142 vpwr vgnd scs8hd_fill_2
XFILLER_27_120 vpwr vgnd scs8hd_fill_2
XFILLER_19_88 vgnd vpwr scs8hd_decap_8
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_76 vpwr vgnd scs8hd_fill_2
XFILLER_35_43 vgnd vpwr scs8hd_decap_4
XFILLER_27_197 vpwr vgnd scs8hd_fill_2
X_074_ _074_/A _074_/Y vgnd vpwr scs8hd_inv_8
X_143_ address[6] _113_/B _143_/C _083_/C _143_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XFILLER_33_145 vpwr vgnd scs8hd_fill_2
XFILLER_33_134 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _082_/Y mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__147__A _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_1_ mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_178 vgnd vpwr scs8hd_decap_3
XFILLER_24_123 vpwr vgnd scs8hd_fill_2
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__057__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_21_12 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_101 vpwr vgnd scs8hd_fill_2
XFILLER_15_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_126_ _112_/A _122_/B _126_/Y vgnd vpwr scs8hd_nor2_4
X_057_ address[1] _091_/A vgnd vpwr scs8hd_inv_8
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_21_159 vpwr vgnd scs8hd_fill_2
XFILLER_16_12 vpwr vgnd scs8hd_fill_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_16_45 vpwr vgnd scs8hd_fill_2
XFILLER_32_99 vgnd vpwr scs8hd_fill_1
XFILLER_32_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_229 vpwr vgnd scs8hd_fill_2
XANTENNA__144__B _113_/B vgnd vpwr scs8hd_diode_2
X_109_ _090_/B _110_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_196 vgnd vpwr scs8hd_decap_6
XFILLER_26_229 vgnd vpwr scs8hd_decap_8
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__070__A _070_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_77 vpwr vgnd scs8hd_fill_2
XFILLER_25_262 vgnd vpwr scs8hd_decap_12
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _071_/A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XFILLER_4_59 vgnd vpwr scs8hd_decap_12
XANTENNA__139__B _113_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_11.LATCH_1_.latch data_in _075_/A _145_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__065__A _065_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_24 vpwr vgnd scs8hd_fill_2
XFILLER_13_79 vpwr vgnd scs8hd_fill_2
XFILLER_22_265 vgnd vpwr scs8hd_decap_8
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_103 vpwr vgnd scs8hd_fill_2
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_76 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_236 vgnd vpwr scs8hd_decap_8
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _070_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__141__C _106_/C vgnd vpwr scs8hd_diode_2
XFILLER_24_67 vgnd vpwr scs8hd_decap_4
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
XFILLER_40_44 vpwr vgnd scs8hd_fill_2
X_090_ _088_/A _090_/B _090_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XANTENNA__136__C _143_/C vgnd vpwr scs8hd_diode_2
XANTENNA__152__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ _068_/A mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_69 vgnd vpwr scs8hd_decap_4
XFILLER_19_45 vpwr vgnd scs8hd_fill_2
XFILLER_19_56 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
X_142_ address[6] _113_/B _106_/C address[0] _142_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_073_ _073_/A _073_/Y vgnd vpwr scs8hd_inv_8
XFILLER_18_8 vpwr vgnd scs8hd_fill_2
XFILLER_33_179 vgnd vpwr scs8hd_decap_4
XANTENNA__147__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_18_110 vgnd vpwr scs8hd_decap_3
XFILLER_24_102 vgnd vpwr scs8hd_decap_3
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _068_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_149 vpwr vgnd scs8hd_fill_2
XFILLER_30_138 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_4
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_125_ _118_/A _122_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_7 vgnd vpwr scs8hd_decap_6
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_14_190 vpwr vgnd scs8hd_fill_2
XFILLER_21_138 vpwr vgnd scs8hd_fill_2
XFILLER_29_227 vpwr vgnd scs8hd_fill_2
XANTENNA__068__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_208 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _072_/A vgnd
+ vpwr scs8hd_diode_2
X_108_ _088_/B _110_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_193 vpwr vgnd scs8hd_fill_2
XANTENNA__144__C _143_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_230 vgnd vpwr scs8hd_decap_4
XFILLER_26_219 vgnd vpwr scs8hd_fill_1
XFILLER_34_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _076_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_34 vpwr vgnd scs8hd_fill_2
XFILLER_25_274 vgnd vpwr scs8hd_decap_3
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _128_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XANTENNA__139__C _120_/C vgnd vpwr scs8hd_diode_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__171__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_22_211 vgnd vpwr scs8hd_decap_3
XFILLER_13_58 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XANTENNA__081__A _081_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_88 vgnd vpwr scs8hd_decap_4
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _154_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__141__D _083_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__076__A _076_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _155_/HI _077_/Y mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__136__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__152__C _143_/C vgnd vpwr scs8hd_diode_2
XFILLER_36_144 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _074_/A mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_35_89 vgnd vpwr scs8hd_decap_4
X_141_ address[6] _113_/B _106_/C _083_/C _141_/Y vgnd vpwr scs8hd_nor4_4
X_072_ _072_/A _072_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_114 vpwr vgnd scs8hd_fill_2
XANTENNA__147__C _120_/C vgnd vpwr scs8hd_diode_2
XFILLER_18_188 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _158_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_36 vpwr vgnd scs8hd_fill_2
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_147 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
X_124_ _110_/A _122_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_38 vpwr vgnd scs8hd_fill_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _108_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__174__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_29_239 vgnd vpwr scs8hd_decap_3
XFILLER_32_79 vpwr vgnd scs8hd_fill_2
XANTENNA__084__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
X_107_ _086_/A _110_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_110 vpwr vgnd scs8hd_fill_2
XANTENNA__144__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__169__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_8_81 vgnd vpwr scs8hd_decap_8
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _079_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__D _083_/C vgnd vpwr scs8hd_diode_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_6
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_245 vpwr vgnd scs8hd_fill_2
XFILLER_0_160 vpwr vgnd scs8hd_fill_2
XANTENNA__182__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_8_271 vgnd vpwr scs8hd_decap_4
XFILLER_39_142 vgnd vpwr scs8hd_decap_12
XFILLER_39_131 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XFILLER_10_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_263 vgnd vpwr scs8hd_decap_12
XANTENNA__152__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_8
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _076_/A mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_189 vgnd vpwr scs8hd_decap_12
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_10_49 vgnd vpwr scs8hd_decap_6
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_123 vpwr vgnd scs8hd_fill_2
XFILLER_27_112 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A address[1] vgnd vpwr scs8hd_diode_2
X_071_ _071_/A _071_/Y vgnd vpwr scs8hd_inv_8
X_140_ address[6] _113_/B _120_/C address[0] _140_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_18_145 vgnd vpwr scs8hd_decap_4
XFILLER_18_167 vpwr vgnd scs8hd_fill_2
XFILLER_33_104 vgnd vpwr scs8hd_fill_1
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__147__D _083_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_123_ _090_/B _122_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_8 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _080_/Y mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_262 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _090_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_47 vpwr vgnd scs8hd_fill_2
XANTENNA__084__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_184 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
X_106_ address[6] address[5] _106_/C _110_/B vgnd vpwr scs8hd_or3_4
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_34_243 vgnd vpwr scs8hd_decap_12
XFILLER_19_251 vgnd vpwr scs8hd_decap_4
XFILLER_8_93 vgnd vpwr scs8hd_fill_1
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XFILLER_25_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_31_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_90 vgnd vpwr scs8hd_decap_4
XFILLER_22_224 vpwr vgnd scs8hd_fill_2
XFILLER_13_213 vpwr vgnd scs8hd_fill_2
XFILLER_28_90 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_3_ mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _069_/A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_39_154 vgnd vpwr scs8hd_decap_12
XANTENNA__092__B _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_205 vgnd vpwr scs8hd_decap_8
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_5_275 vpwr vgnd scs8hd_fill_2
XFILLER_36_168 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_19_15 vpwr vgnd scs8hd_fill_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XFILLER_27_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__087__B _083_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_070_ _070_/A _070_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_33_149 vpwr vgnd scs8hd_fill_2
XFILLER_33_138 vpwr vgnd scs8hd_fill_2
XFILLER_26_190 vgnd vpwr scs8hd_decap_4
XFILLER_25_80 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _161_/HI _073_/Y mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_182 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_16 vgnd vpwr scs8hd_decap_3
XANTENNA__098__A address[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ _066_/A mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_193 vpwr vgnd scs8hd_fill_2
X_122_ _088_/B _122_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_8 vpwr vgnd scs8hd_fill_2
XFILLER_14_160 vpwr vgnd scs8hd_fill_2
XFILLER_37_274 vgnd vpwr scs8hd_decap_3
XFILLER_29_208 vpwr vgnd scs8hd_fill_2
XANTENNA__084__C _105_/C vgnd vpwr scs8hd_diode_2
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_16_49 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_196 vpwr vgnd scs8hd_fill_2
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XFILLER_28_252 vgnd vpwr scs8hd_decap_8
XFILLER_28_241 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _069_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
X_105_ address[3] _063_/Y _105_/C _106_/C vgnd vpwr scs8hd_or3_4
XFILLER_22_70 vgnd vpwr scs8hd_decap_4
XFILLER_19_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_15 vpwr vgnd scs8hd_fill_2
XANTENNA__095__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_19 vgnd vpwr scs8hd_decap_12
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 left_top_grid_pin_15_ mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_107 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_203 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _159_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_184 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_251 vgnd vpwr scs8hd_decap_4
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_39_166 vgnd vpwr scs8hd_decap_12
XFILLER_39_188 vpwr vgnd scs8hd_fill_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XFILLER_14_82 vgnd vpwr scs8hd_decap_4
XFILLER_14_93 vpwr vgnd scs8hd_fill_2
XFILLER_36_147 vgnd vpwr scs8hd_decap_6
XFILLER_36_136 vgnd vpwr scs8hd_decap_8
XFILLER_36_125 vpwr vgnd scs8hd_fill_2
XFILLER_10_18 vgnd vpwr scs8hd_decap_6
XANTENNA__087__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _071_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_125 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _075_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _154_/HI _075_/Y mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__B address[5] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _072_/A mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_7_19 vgnd vpwr scs8hd_fill_1
X_121_ _086_/A _122_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_83 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_194 vpwr vgnd scs8hd_fill_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _100_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
X_104_ _112_/A _103_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XFILLER_7_102 vgnd vpwr scs8hd_decap_8
XFILLER_11_164 vpwr vgnd scs8hd_fill_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
XFILLER_11_197 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_60 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_231 vgnd vpwr scs8hd_fill_1
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XFILLER_21_7 vgnd vpwr scs8hd_decap_3
XFILLER_8_51 vgnd vpwr scs8hd_decap_8
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_27_38 vgnd vpwr scs8hd_decap_4
XFILLER_25_245 vgnd vpwr scs8hd_decap_3
XANTENNA__095__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_226 vpwr vgnd scs8hd_fill_2
XFILLER_31_204 vgnd vpwr scs8hd_decap_3
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XFILLER_17_82 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _164_/HI mem_left_track_9.LATCH_2_.latch/Q
+ mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_270 vgnd vpwr scs8hd_decap_4
XFILLER_13_18 vgnd vpwr scs8hd_decap_4
XFILLER_1_119 vgnd vpwr scs8hd_decap_3
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _155_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_270 vgnd vpwr scs8hd_decap_4
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_39_178 vgnd vpwr scs8hd_decap_4
XFILLER_39_123 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_49 vgnd vpwr scs8hd_decap_12
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_6
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_5_ mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_115 vgnd vpwr scs8hd_decap_4
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_107 vgnd vpwr scs8hd_decap_3
XANTENNA__098__C _120_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _113_/A _113_/B _120_/C _122_/B vgnd vpwr scs8hd_or3_4
XFILLER_23_162 vpwr vgnd scs8hd_fill_2
XFILLER_14_173 vgnd vpwr scs8hd_decap_8
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_143 vgnd vpwr scs8hd_decap_3
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_20_165 vpwr vgnd scs8hd_fill_2
XFILLER_20_176 vgnd vpwr scs8hd_decap_8
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
X_103_ _118_/A _103_/B _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_8_74 vgnd vpwr scs8hd_fill_1
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_235 vpwr vgnd scs8hd_fill_2
XFILLER_25_224 vpwr vgnd scs8hd_fill_2
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _078_/Y mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_16_202 vgnd vpwr scs8hd_decap_12
XFILLER_16_224 vgnd vpwr scs8hd_decap_8
XFILLER_16_235 vgnd vpwr scs8hd_decap_12
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_249 vgnd vpwr scs8hd_decap_12
XFILLER_31_238 vgnd vpwr scs8hd_decap_6
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_205 vgnd vpwr scs8hd_decap_4
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_249 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_153 vpwr vgnd scs8hd_fill_2
XFILLER_0_164 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vpwr vgnd scs8hd_fill_2
XFILLER_28_82 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_5_53 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_15.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _181_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_83 vgnd vpwr scs8hd_fill_1
XFILLER_30_72 vgnd vpwr scs8hd_decap_4
XFILLER_5_245 vgnd vpwr scs8hd_decap_8
XANTENNA__101__A _090_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_138 vpwr vgnd scs8hd_fill_2
XFILLER_27_116 vpwr vgnd scs8hd_fill_2
XFILLER_27_105 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _067_/A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_193 vpwr vgnd scs8hd_fill_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_149 vgnd vpwr scs8hd_fill_1
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_182 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _191_/A vgnd vpwr scs8hd_inv_1
XFILLER_37_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_119 vpwr vgnd scs8hd_fill_2
XFILLER_17_160 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_17_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_30 vpwr vgnd scs8hd_fill_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_179_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_35_3 vpwr vgnd scs8hd_fill_2
XFILLER_37_266 vgnd vpwr scs8hd_decap_8
XFILLER_32_29 vpwr vgnd scs8hd_fill_2
XFILLER_20_122 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _160_/HI _071_/Y mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_100 vpwr vgnd scs8hd_fill_2
XFILLER_11_111 vpwr vgnd scs8hd_fill_2
X_102_ _110_/A _103_/B _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_159 vgnd vpwr scs8hd_decap_12
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_211 vgnd vpwr scs8hd_fill_1
XFILLER_34_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_16_247 vgnd vpwr scs8hd_decap_12
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _112_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XFILLER_22_228 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_217 vpwr vgnd scs8hd_fill_2
XFILLER_28_50 vpwr vgnd scs8hd_fill_2
XFILLER_0_176 vgnd vpwr scs8hd_decap_8
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.LATCH_0_.latch data_in _074_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _158_/HI _068_/Y mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _072_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_191 vgnd vpwr scs8hd_decap_12
XFILLER_14_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _076_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__101__B _103_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_191 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_19 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.INVTX1_0_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_194 vgnd vpwr scs8hd_fill_1
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_84 vpwr vgnd scs8hd_fill_2
XFILLER_25_62 vgnd vpwr scs8hd_decap_3
XFILLER_25_40 vpwr vgnd scs8hd_fill_2
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XANTENNA__112__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
XFILLER_23_197 vgnd vpwr scs8hd_decap_8
XFILLER_11_20 vpwr vgnd scs8hd_fill_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_75 vgnd vpwr scs8hd_decap_6
XFILLER_14_120 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _086_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_178_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_37_212 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_19 vgnd vpwr scs8hd_decap_8
X_101_ _090_/B _103_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_123 vgnd vpwr scs8hd_decap_3
XFILLER_11_145 vpwr vgnd scs8hd_fill_2
XFILLER_22_74 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _070_/A mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_234 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_4
XFILLER_34_226 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vpwr vgnd scs8hd_fill_2
XFILLER_8_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _074_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _078_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_259 vgnd vpwr scs8hd_decap_12
XFILLER_17_41 vgnd vpwr scs8hd_fill_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_73 vpwr vgnd scs8hd_fill_2
XANTENNA__104__B _103_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
XANTENNA__120__A _113_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _107_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_1_ mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A right_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_240 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _187_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_111 vgnd vpwr scs8hd_decap_12
XFILLER_0_133 vgnd vpwr scs8hd_decap_12
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _160_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__115__A _088_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _074_/Y mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_0_.latch data_in _082_/A _152_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_162 vpwr vgnd scs8hd_fill_2
XFILLER_35_19 vgnd vpwr scs8hd_decap_12
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__112__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_165 vpwr vgnd scs8hd_fill_2
XFILLER_32_132 vpwr vgnd scs8hd_fill_2
XFILLER_23_143 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_11.INVTX1_0_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_154 vgnd vpwr scs8hd_decap_4
X_177_ _177_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__107__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_198 vgnd vpwr scs8hd_decap_3
XANTENNA__123__A _090_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_224 vgnd vpwr scs8hd_decap_12
XFILLER_28_224 vpwr vgnd scs8hd_fill_2
X_100_ _088_/B _103_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_168 vpwr vgnd scs8hd_fill_2
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
XFILLER_22_42 vpwr vgnd scs8hd_fill_2
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_77 vpwr vgnd scs8hd_fill_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 left_top_grid_pin_13_ mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XFILLER_33_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _113_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_252 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_123 vgnd vpwr scs8hd_fill_1
XFILLER_0_145 vgnd vpwr scs8hd_decap_8
XFILLER_28_41 vgnd vpwr scs8hd_decap_3
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _088_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_274 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _076_/Y mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__115__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _156_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_138 vpwr vgnd scs8hd_fill_2
XANTENNA__131__A _110_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_11_ mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_32 vgnd vpwr scs8hd_decap_4
XFILLER_14_65 vpwr vgnd scs8hd_fill_2
XFILLER_30_86 vgnd vpwr scs8hd_decap_6
XFILLER_5_259 vpwr vgnd scs8hd_fill_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_36_108 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_182 vgnd vpwr scs8hd_fill_1
XANTENNA__126__A _112_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_5.LATCH_0_.latch data_in _070_/A _140_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_97 vpwr vgnd scs8hd_fill_2
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ _193_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_1_262 vgnd vpwr scs8hd_decap_12
XFILLER_17_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_30 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _065_/A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_96 vgnd vpwr scs8hd_decap_12
X_176_ _176_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__123__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_258 vpwr vgnd scs8hd_fill_2
XFILLER_37_236 vgnd vpwr scs8hd_decap_8
XFILLER_20_169 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_247 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vgnd vpwr scs8hd_decap_4
XFILLER_22_10 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_206 vgnd vpwr scs8hd_decap_8
XFILLER_19_214 vpwr vgnd scs8hd_fill_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_23 vgnd vpwr scs8hd_decap_8
XFILLER_8_89 vgnd vpwr scs8hd_decap_3
XFILLER_10_180 vgnd vpwr scs8hd_decap_4
XANTENNA__134__A _134_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_159_ _159_/HI _159_/LO vgnd vpwr scs8hd_conb_1
XFILLER_25_239 vgnd vpwr scs8hd_decap_4
XFILLER_25_228 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _163_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XFILLER_33_31 vpwr vgnd scs8hd_fill_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_209 vpwr vgnd scs8hd_fill_2
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_87 vpwr vgnd scs8hd_fill_2
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XANTENNA__120__C _120_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _159_/HI _069_/Y mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__129__A _088_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_264 vgnd vpwr scs8hd_decap_12
XFILLER_0_102 vgnd vpwr scs8hd_fill_1
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XFILLER_12_231 vgnd vpwr scs8hd_decap_12
XANTENNA__131__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_35 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_88 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_8
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__126__B _122_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_35_142 vgnd vpwr scs8hd_fill_1
XFILLER_35_197 vgnd vpwr scs8hd_decap_4
XFILLER_35_175 vpwr vgnd scs8hd_fill_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_186 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_10 vpwr vgnd scs8hd_fill_2
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _153_/HI _066_/Y mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_1_274 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_13.LATCH_0_.latch data_in _078_/A _148_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_32_145 vgnd vpwr scs8hd_decap_6
XANTENNA__137__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_17_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _167_/HI mem_right_track_8.LATCH_2_.latch/Q
+ mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_45 vpwr vgnd scs8hd_fill_2
XFILLER_36_86 vgnd vpwr scs8hd_decap_6
XFILLER_14_145 vgnd vpwr scs8hd_decap_6
X_175_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_37_204 vgnd vpwr scs8hd_fill_1
XFILLER_35_7 vgnd vpwr scs8hd_decap_12
XFILLER_28_6 vpwr vgnd scs8hd_fill_2
XFILLER_20_126 vpwr vgnd scs8hd_fill_2
XFILLER_20_148 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_204 vpwr vgnd scs8hd_fill_2
XFILLER_36_270 vgnd vpwr scs8hd_decap_4
XFILLER_11_104 vpwr vgnd scs8hd_fill_2
XFILLER_11_115 vgnd vpwr scs8hd_decap_4
XFILLER_22_55 vgnd vpwr scs8hd_decap_3
XFILLER_22_66 vpwr vgnd scs8hd_fill_2
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_68 vgnd vpwr scs8hd_decap_6
X_158_ _158_/HI _158_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__134__B _063_/Y vgnd vpwr scs8hd_diode_2
X_089_ _091_/A address[2] _083_/C _090_/B vgnd vpwr scs8hd_or3_4
XANTENNA__150__A _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _071_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_262 vpwr vgnd scs8hd_fill_2
XFILLER_33_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__060__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_17_22 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _075_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _113_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _068_/A mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_221 vpwr vgnd scs8hd_fill_2
XFILLER_21_232 vpwr vgnd scs8hd_fill_2
XFILLER_21_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_65 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _099_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_10 vgnd vpwr scs8hd_decap_4
XFILLER_12_243 vgnd vpwr scs8hd_fill_1
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_162 vpwr vgnd scs8hd_fill_2
XFILLER_14_12 vpwr vgnd scs8hd_fill_2
XFILLER_30_99 vgnd vpwr scs8hd_fill_1
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_39_53 vpwr vgnd scs8hd_fill_2
XFILLER_29_162 vpwr vgnd scs8hd_fill_2
XFILLER_29_140 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _166_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__B _113_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_154 vgnd vpwr scs8hd_decap_6
XFILLER_35_132 vpwr vgnd scs8hd_fill_2
XFILLER_6_90 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _072_/Y mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_165 vpwr vgnd scs8hd_fill_2
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ _191_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A left_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_1_253 vpwr vgnd scs8hd_fill_2
XFILLER_32_113 vgnd vpwr scs8hd_decap_4
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XANTENNA__137__B _113_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _073_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_113 vpwr vgnd scs8hd_fill_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_24 vgnd vpwr scs8hd_decap_4
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA__063__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _077_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_65 vgnd vpwr scs8hd_decap_8
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_0_.latch data_in _066_/A _136_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_124 vpwr vgnd scs8hd_fill_2
XFILLER_22_190 vpwr vgnd scs8hd_fill_2
X_174_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__148__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_105 vpwr vgnd scs8hd_fill_2
XFILLER_11_149 vpwr vgnd scs8hd_fill_2
XFILLER_22_23 vpwr vgnd scs8hd_fill_2
XANTENNA__058__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_227 vgnd vpwr scs8hd_decap_4
XFILLER_19_238 vgnd vpwr scs8hd_decap_6
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XFILLER_8_36 vgnd vpwr scs8hd_decap_6
XFILLER_10_193 vgnd vpwr scs8hd_decap_12
X_157_ _157_/HI _157_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__134__C _105_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_088_ _088_/A _088_/B _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
XFILLER_33_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_230 vgnd vpwr scs8hd_decap_4
XFILLER_17_34 vgnd vpwr scs8hd_decap_4
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_33_77 vpwr vgnd scs8hd_fill_2
XFILLER_33_11 vgnd vpwr scs8hd_decap_12
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_230 vpwr vgnd scs8hd_fill_2
XANTENNA__145__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_81 vgnd vpwr scs8hd_fill_1
XANTENNA__071__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_259 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_7 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _161_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XANTENNA__066__A _066_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_24 vgnd vpwr scs8hd_decap_4
XFILLER_30_23 vgnd vpwr scs8hd_decap_4
XFILLER_14_46 vpwr vgnd scs8hd_fill_2
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
XANTENNA__142__C _106_/C vgnd vpwr scs8hd_diode_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_67 vpwr vgnd scs8hd_fill_2
XFILLER_25_34 vgnd vpwr scs8hd_decap_4
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_32_169 vpwr vgnd scs8hd_fill_2
XANTENNA__137__C _085_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 right_top_grid_pin_15_ mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_158 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
X_173_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_139 vpwr vgnd scs8hd_fill_2
XFILLER_9_173 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vpwr vgnd scs8hd_fill_2
XFILLER_28_228 vgnd vpwr scs8hd_decap_4
XANTENNA__074__A _074_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_8_15 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_087_ address[1] _083_/B address[0] _088_/B vgnd vpwr scs8hd_or3_4
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XFILLER_6_121 vgnd vpwr scs8hd_decap_12
X_156_ _156_/HI _156_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__150__C _106_/C vgnd vpwr scs8hd_diode_2
XFILLER_25_209 vpwr vgnd scs8hd_fill_2
XFILLER_33_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _069_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_23 vgnd vpwr scs8hd_decap_8
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__145__C _085_/C vgnd vpwr scs8hd_diode_2
X_139_ address[6] _113_/B _120_/C _083_/C _139_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XFILLER_0_60 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _162_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_49 vpwr vgnd scs8hd_fill_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _157_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _067_/Y mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _193_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_69 vpwr vgnd scs8hd_fill_2
XFILLER_30_79 vgnd vpwr scs8hd_decap_4
XFILLER_30_68 vpwr vgnd scs8hd_fill_2
XFILLER_30_13 vgnd vpwr scs8hd_fill_1
XANTENNA__082__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XFILLER_29_175 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_35_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_26_145 vpwr vgnd scs8hd_fill_2
XFILLER_26_112 vpwr vgnd scs8hd_fill_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _077_/A vgnd vpwr scs8hd_diode_2
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vgnd vpwr scs8hd_decap_4
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XFILLER_17_112 vgnd vpwr scs8hd_decap_4
XANTENNA__137__D _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_3
XFILLER_17_145 vpwr vgnd scs8hd_fill_2
XFILLER_17_156 vpwr vgnd scs8hd_fill_2
XFILLER_17_178 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_192 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_9.LATCH_1_.latch data_in _073_/A _143_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB _146_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_104 vpwr vgnd scs8hd_fill_2
XFILLER_14_115 vgnd vpwr scs8hd_decap_3
X_172_ _172_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_22_170 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__148__C _120_/C vgnd vpwr scs8hd_diode_2
XANTENNA__180__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_22_36 vgnd vpwr scs8hd_decap_4
XANTENNA__090__A _088_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _126_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_262 vpwr vgnd scs8hd_fill_2
XFILLER_27_251 vgnd vpwr scs8hd_decap_4
XFILLER_19_207 vgnd vpwr scs8hd_decap_4
X_086_ _086_/A _088_/A _086_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_6_133 vgnd vpwr scs8hd_decap_12
X_155_ _155_/HI _155_/LO vgnd vpwr scs8hd_conb_1
XFILLER_12_91 vgnd vpwr scs8hd_fill_1
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XFILLER_26_6 vpwr vgnd scs8hd_fill_2
XANTENNA__150__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_240 vgnd vpwr scs8hd_decap_8
XFILLER_18_251 vgnd vpwr scs8hd_decap_8
XFILLER_18_262 vgnd vpwr scs8hd_decap_12
XANTENNA__175__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_243 vgnd vpwr scs8hd_decap_12
XANTENNA__085__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XFILLER_30_246 vgnd vpwr scs8hd_decap_12
XANTENNA__145__D _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_23_90 vpwr vgnd scs8hd_fill_2
X_138_ address[6] _113_/B _085_/C address[0] _138_/Y vgnd vpwr scs8hd_nor4_4
X_069_ _069_/A _069_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_3 vgnd vpwr scs8hd_decap_4
XFILLER_0_94 vgnd vpwr scs8hd_decap_8
XFILLER_21_202 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_46 vpwr vgnd scs8hd_fill_2
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _066_/A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_45 vgnd vpwr scs8hd_fill_1
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
XFILLER_29_121 vgnd vpwr scs8hd_fill_1
XFILLER_29_110 vgnd vpwr scs8hd_fill_1
XFILLER_29_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _074_/Y vgnd
+ vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_179 vpwr vgnd scs8hd_fill_2
XANTENNA__183__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _078_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_25_14 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_8
XFILLER_25_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__178__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_16_190 vgnd vpwr scs8hd_fill_1
XFILLER_11_49 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A _088_/A vgnd vpwr scs8hd_diode_2
X_171_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _070_/Y mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_37_208 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_1_.latch data_in _081_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__148__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_13_193 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_208 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_274 vgnd vpwr scs8hd_fill_1
XFILLER_36_241 vpwr vgnd scs8hd_fill_2
XFILLER_11_119 vgnd vpwr scs8hd_fill_1
XANTENNA__090__B _090_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_154_ _154_/HI _154_/LO vgnd vpwr scs8hd_conb_1
X_085_ address[6] address[5] _085_/C _088_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
XFILLER_6_145 vgnd vpwr scs8hd_decap_8
XFILLER_10_163 vgnd vpwr scs8hd_decap_4
XFILLER_33_266 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _189_/A vgnd vpwr scs8hd_inv_1
XFILLER_24_211 vgnd vpwr scs8hd_decap_3
XFILLER_17_26 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_36 vgnd vpwr scs8hd_decap_6
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__085__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_258 vgnd vpwr scs8hd_decap_12
X_137_ address[6] _113_/B _085_/C _083_/C _137_/Y vgnd vpwr scs8hd_nor4_4
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_068_ _068_/A _068_/Y vgnd vpwr scs8hd_inv_8
XFILLER_0_40 vgnd vpwr scs8hd_fill_1
XFILLER_17_3 vgnd vpwr scs8hd_decap_4
XFILLER_9_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _080_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_225 vpwr vgnd scs8hd_fill_2
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _168_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_107 vpwr vgnd scs8hd_fill_2
XFILLER_0_129 vpwr vgnd scs8hd_fill_2
XFILLER_28_69 vpwr vgnd scs8hd_fill_2
XFILLER_12_203 vgnd vpwr scs8hd_fill_1
XANTENNA__096__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_247 vgnd vpwr scs8hd_decap_8
XFILLER_12_258 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_16 vpwr vgnd scs8hd_fill_2
XFILLER_14_38 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_57 vgnd vpwr scs8hd_decap_4
XFILLER_29_144 vgnd vpwr scs8hd_decap_3
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_20_70 vgnd vpwr scs8hd_decap_3
XFILLER_35_136 vgnd vpwr scs8hd_decap_6
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _172_/A vgnd vpwr scs8hd_inv_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_169 vgnd vpwr scs8hd_decap_4
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _066_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__093__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_128 vpwr vgnd scs8hd_fill_2
XFILLER_31_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _086_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_180 vgnd vpwr scs8hd_decap_4
XFILLER_23_117 vgnd vpwr scs8hd_decap_3
XFILLER_23_139 vpwr vgnd scs8hd_fill_2
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _088_/B vgnd vpwr scs8hd_diode_2
X_170_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_132 vgnd vpwr scs8hd_decap_12
XFILLER_20_109 vpwr vgnd scs8hd_fill_2
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_120 vpwr vgnd scs8hd_fill_2
X_153_ _153_/HI _153_/LO vgnd vpwr scs8hd_conb_1
Xmem_bottom_track_5.LATCH_1_.latch data_in _069_/A _139_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_084_ address[3] address[4] _105_/C _085_/C vgnd vpwr scs8hd_or3_4
XFILLER_33_245 vgnd vpwr scs8hd_decap_8
XFILLER_33_223 vpwr vgnd scs8hd_fill_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_201 vpwr vgnd scs8hd_fill_2
XFILLER_17_38 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _166_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__C _085_/C vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vpwr vgnd scs8hd_fill_2
XFILLER_15_201 vgnd vpwr scs8hd_decap_6
XFILLER_15_223 vpwr vgnd scs8hd_fill_2
XFILLER_15_234 vpwr vgnd scs8hd_fill_2
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_136_ address[6] address[5] _143_/C address[0] _136_/Y vgnd vpwr scs8hd_nor4_4
X_067_ _067_/A _067_/Y vgnd vpwr scs8hd_inv_8
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_94 vpwr vgnd scs8hd_fill_2
XFILLER_21_248 vpwr vgnd scs8hd_fill_2
XFILLER_12_215 vpwr vgnd scs8hd_fill_2
XANTENNA__096__B _112_/A vgnd vpwr scs8hd_diode_2
X_119_ _112_/A _118_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_167 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_49 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_20_82 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_104 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA__093__C _083_/C vgnd vpwr scs8hd_diode_2
XFILLER_1_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _065_/Y mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_31_151 vgnd vpwr scs8hd_decap_3
XFILLER_23_129 vgnd vpwr scs8hd_fill_1
XFILLER_31_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _165_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_111 vgnd vpwr scs8hd_decap_4
XFILLER_9_144 vgnd vpwr scs8hd_decap_12
XFILLER_9_177 vgnd vpwr scs8hd_decap_6
XFILLER_9_188 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_173 vgnd vpwr scs8hd_decap_4
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_36_254 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__099__B _103_/B vgnd vpwr scs8hd_diode_2
X_083_ address[1] _083_/B _083_/C _086_/A vgnd vpwr scs8hd_or3_4
XFILLER_8_19 vgnd vpwr scs8hd_fill_1
XFILLER_10_154 vpwr vgnd scs8hd_fill_2
XFILLER_10_176 vpwr vgnd scs8hd_fill_2
XFILLER_12_61 vgnd vpwr scs8hd_fill_1
X_152_ _113_/A address[5] _143_/C address[0] _152_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_202 vpwr vgnd scs8hd_fill_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_13.LATCH_1_.latch data_in _077_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_7.INVTX1_1_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
X_066_ _066_/A _066_/Y vgnd vpwr scs8hd_inv_8
X_135_ address[6] address[5] _143_/C _083_/C _135_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_23_60 vgnd vpwr scs8hd_fill_1
XFILLER_23_71 vpwr vgnd scs8hd_fill_2
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_0_75 vgnd vpwr scs8hd_decap_6
XFILLER_9_62 vpwr vgnd scs8hd_fill_2
XFILLER_9_84 vgnd vpwr scs8hd_decap_8
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_18_60 vpwr vgnd scs8hd_fill_2
XFILLER_18_93 vpwr vgnd scs8hd_fill_2
X_118_ _118_/A _118_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_253 vpwr vgnd scs8hd_fill_2
XFILLER_7_242 vpwr vgnd scs8hd_fill_2
XFILLER_38_179 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_179 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_9_ mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_35_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_41 vgnd vpwr scs8hd_fill_1
XFILLER_26_149 vpwr vgnd scs8hd_fill_2
XFILLER_26_116 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_19_190 vpwr vgnd scs8hd_fill_2
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_34_193 vpwr vgnd scs8hd_fill_2
XPHY_39 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 right_top_grid_pin_13_ mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_7 vgnd vpwr scs8hd_decap_8
XFILLER_25_182 vgnd vpwr scs8hd_fill_1
XFILLER_17_149 vpwr vgnd scs8hd_fill_2
XFILLER_15_83 vgnd vpwr scs8hd_decap_3
XFILLER_31_93 vgnd vpwr scs8hd_decap_3
XFILLER_14_108 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_130 vpwr vgnd scs8hd_fill_2
XFILLER_13_152 vpwr vgnd scs8hd_fill_2
XFILLER_9_156 vpwr vgnd scs8hd_fill_2
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
XFILLER_3_31 vgnd vpwr scs8hd_decap_12
XFILLER_36_222 vgnd vpwr scs8hd_decap_4
XFILLER_27_266 vgnd vpwr scs8hd_decap_8
XFILLER_10_100 vpwr vgnd scs8hd_fill_2
X_082_ _082_/A _082_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_133 vpwr vgnd scs8hd_fill_2
XFILLER_12_73 vpwr vgnd scs8hd_fill_2
XFILLER_12_84 vgnd vpwr scs8hd_decap_4
X_151_ _113_/A address[5] _143_/C _083_/C _151_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_33_236 vpwr vgnd scs8hd_fill_2
XFILLER_18_200 vpwr vgnd scs8hd_fill_2
XFILLER_18_222 vpwr vgnd scs8hd_fill_2
XFILLER_33_258 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _068_/Y mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _162_/HI mem_left_track_1.LATCH_2_.latch/Q
+ mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _073_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_206 vgnd vpwr scs8hd_decap_8
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_065_ _065_/A _065_/Y vgnd vpwr scs8hd_inv_8
X_134_ _134_/A _063_/Y _105_/C _143_/C vgnd vpwr scs8hd_or3_4
XFILLER_23_94 vpwr vgnd scs8hd_fill_2
XFILLER_24_7 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_1.LATCH_1_.latch data_in _065_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _077_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_52 vgnd vpwr scs8hd_decap_4
XFILLER_12_206 vgnd vpwr scs8hd_decap_8
XFILLER_20_272 vgnd vpwr scs8hd_decap_3
XFILLER_34_93 vgnd vpwr scs8hd_decap_8
X_117_ _110_/A _118_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_210 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.INVTX1_1_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_3 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_29 vpwr vgnd scs8hd_fill_2
XFILLER_39_49 vpwr vgnd scs8hd_fill_2
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_29_136 vpwr vgnd scs8hd_fill_2
XFILLER_29_114 vgnd vpwr scs8hd_decap_4
XFILLER_29_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XFILLER_20_62 vpwr vgnd scs8hd_fill_2
XFILLER_35_117 vgnd vpwr scs8hd_decap_3
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _111_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_97 vgnd vpwr scs8hd_decap_12
XFILLER_34_161 vgnd vpwr scs8hd_decap_4
XFILLER_26_128 vgnd vpwr scs8hd_decap_6
XFILLER_25_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_34_183 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_109 vpwr vgnd scs8hd_fill_2
XFILLER_25_161 vpwr vgnd scs8hd_fill_2
XFILLER_15_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_109 vpwr vgnd scs8hd_fill_2
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_186 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_72 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _079_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_201 vgnd vpwr scs8hd_decap_12
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_3_43 vgnd vpwr scs8hd_decap_12
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
XFILLER_27_245 vgnd vpwr scs8hd_decap_4
XFILLER_27_234 vpwr vgnd scs8hd_fill_2
XFILLER_27_212 vgnd vpwr scs8hd_decap_3
X_150_ _113_/A address[5] _106_/C address[0] _150_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_081_ _081_/A _081_/Y vgnd vpwr scs8hd_inv_8
XFILLER_12_30 vgnd vpwr scs8hd_fill_1
XFILLER_37_71 vgnd vpwr scs8hd_decap_8
XFILLER_18_212 vpwr vgnd scs8hd_fill_2
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XFILLER_24_226 vpwr vgnd scs8hd_fill_2
XFILLER_24_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_229 vgnd vpwr scs8hd_decap_8
X_133_ _112_/A _131_/B _133_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
X_064_ enable _105_/C vgnd vpwr scs8hd_inv_8
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_44 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _065_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_72 vgnd vpwr scs8hd_fill_1
XFILLER_18_73 vpwr vgnd scs8hd_fill_2
XFILLER_18_84 vgnd vpwr scs8hd_decap_8
X_116_ _090_/B _118_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_222 vgnd vpwr scs8hd_decap_12
XANTENNA__105__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_137 vgnd vpwr scs8hd_fill_1
XFILLER_39_39 vgnd vpwr scs8hd_decap_6
XFILLER_20_41 vgnd vpwr scs8hd_decap_3
XFILLER_29_83 vpwr vgnd scs8hd_fill_2
XFILLER_29_72 vgnd vpwr scs8hd_decap_4
XFILLER_6_54 vgnd vpwr scs8hd_decap_12
XFILLER_6_32 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.INVTX1_1_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_19_170 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _096_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_184 vgnd vpwr scs8hd_decap_4
XFILLER_31_62 vgnd vpwr scs8hd_decap_3
XANTENNA__102__B _103_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_151 vpwr vgnd scs8hd_fill_2
XFILLER_16_173 vgnd vpwr scs8hd_fill_1
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_36_18 vgnd vpwr scs8hd_decap_12
XFILLER_22_121 vpwr vgnd scs8hd_fill_2
XFILLER_22_143 vgnd vpwr scs8hd_decap_4
XFILLER_22_154 vgnd vpwr scs8hd_decap_3
XFILLER_22_176 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vpwr vgnd scs8hd_fill_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_169 vpwr vgnd scs8hd_fill_2
XFILLER_13_165 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_213 vgnd vpwr scs8hd_fill_1
XFILLER_3_55 vgnd vpwr scs8hd_decap_6
XFILLER_36_246 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
X_080_ _080_/A _080_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _185_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_12_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _088_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_205 vgnd vpwr scs8hd_decap_4
XFILLER_30_219 vgnd vpwr scs8hd_fill_1
XFILLER_15_238 vgnd vpwr scs8hd_decap_6
X_063_ address[4] _063_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_52 vpwr vgnd scs8hd_fill_2
X_132_ _118_/A _131_/B _132_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__110__B _110_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _177_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_89 vgnd vpwr scs8hd_decap_4
XFILLER_14_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_12_219 vgnd vpwr scs8hd_decap_12
XFILLER_20_241 vgnd vpwr scs8hd_decap_8
XFILLER_20_252 vgnd vpwr scs8hd_decap_12
XFILLER_34_84 vgnd vpwr scs8hd_decap_8
X_115_ _088_/B _118_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_245 vgnd vpwr scs8hd_decap_8
XFILLER_7_234 vgnd vpwr scs8hd_decap_8
XANTENNA__105__B _063_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__121__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_6 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_160 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_182 vgnd vpwr scs8hd_fill_1
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_62 vgnd vpwr scs8hd_fill_1
XFILLER_20_86 vgnd vpwr scs8hd_decap_4
XANTENNA__116__A _090_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_66 vgnd vpwr scs8hd_decap_12
XFILLER_6_44 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_3 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_130 vgnd vpwr scs8hd_decap_3
XFILLER_17_108 vpwr vgnd scs8hd_fill_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_174 vpwr vgnd scs8hd_fill_2
XFILLER_15_31 vgnd vpwr scs8hd_fill_1
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_97 vpwr vgnd scs8hd_fill_2
XFILLER_0_240 vpwr vgnd scs8hd_fill_2
XFILLER_0_262 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_188 vpwr vgnd scs8hd_fill_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

