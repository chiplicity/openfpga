magic
tech EFS8A
magscale 1 2
timestamp 1602269747
<< locali >>
rect 9631 18785 9758 18819
rect 11471 18785 11506 18819
rect 4445 18275 4479 18377
rect 11287 17697 11322 17731
rect 1955 16745 1961 16779
rect 10051 16745 10057 16779
rect 1955 16677 1989 16745
rect 10051 16677 10085 16745
rect 4169 16609 4330 16643
rect 4169 16575 4203 16609
rect 16899 15521 16934 15555
rect 2047 14807 2081 14875
rect 2047 14773 2053 14807
rect 8217 13719 8251 14025
rect 9631 13345 9758 13379
rect 9683 12631 9717 12699
rect 9683 12597 9689 12631
rect 1863 12393 1869 12427
rect 6647 12393 6653 12427
rect 1863 12325 1897 12393
rect 6647 12325 6681 12393
rect 11931 12257 11966 12291
rect 3059 11543 3093 11611
rect 3059 11509 3065 11543
rect 4169 10999 4203 11305
rect 5083 11305 5089 11339
rect 5083 11237 5117 11305
rect 4445 10591 4479 10761
rect 3111 8993 3249 9027
rect 6101 8415 6135 8585
rect 5911 8041 5917 8075
rect 5911 7973 5945 8041
rect 14841 7939 14875 8041
rect 11471 7905 11598 7939
rect 16037 7905 16129 7939
rect 3111 7701 3249 7735
rect 12725 7327 12759 7497
rect 5951 6885 5996 6919
rect 12811 6103 12845 6171
rect 12811 6069 12817 6103
rect 6503 5729 6538 5763
rect 18463 5729 18498 5763
rect 7251 5185 7389 5219
rect 15669 5015 15703 5117
rect 13915 3927 13949 3995
rect 13915 3893 13921 3927
rect 12081 2839 12115 2941
rect 15577 2839 15611 3009
rect 16681 2873 16807 2907
rect 16773 2839 16807 2873
rect 8493 2499 8527 2601
rect 9321 2295 9355 2465
<< viali >>
rect 2559 19465 2593 19499
rect 2456 19261 2490 19295
rect 2881 19261 2915 19295
rect 5273 19261 5307 19295
rect 5825 19261 5859 19295
rect 8008 19261 8042 19295
rect 8401 19261 8435 19295
rect 9848 19261 9882 19295
rect 10828 19261 10862 19295
rect 11253 19261 11287 19295
rect 1869 19193 1903 19227
rect 5181 19193 5215 19227
rect 6009 19193 6043 19227
rect 1409 19125 1443 19159
rect 4077 19125 4111 19159
rect 6929 19125 6963 19159
rect 8079 19125 8113 19159
rect 9919 19125 9953 19159
rect 10333 19125 10367 19159
rect 10931 19125 10965 19159
rect 2237 18921 2271 18955
rect 4859 18921 4893 18955
rect 5273 18921 5307 18955
rect 7389 18921 7423 18955
rect 11575 18921 11609 18955
rect 2237 18785 2271 18819
rect 2421 18785 2455 18819
rect 4788 18785 4822 18819
rect 6009 18785 6043 18819
rect 6285 18785 6319 18819
rect 7573 18785 7607 18819
rect 7849 18785 7883 18819
rect 9597 18785 9631 18819
rect 11437 18785 11471 18819
rect 6377 18717 6411 18751
rect 1685 18581 1719 18615
rect 3065 18581 3099 18615
rect 9827 18581 9861 18615
rect 4261 18377 4295 18411
rect 4445 18377 4479 18411
rect 7849 18377 7883 18411
rect 13277 18377 13311 18411
rect 15669 18377 15703 18411
rect 17049 18377 17083 18411
rect 4445 18241 4479 18275
rect 5273 18241 5307 18275
rect 5825 18241 5859 18275
rect 6653 18241 6687 18275
rect 1409 18173 1443 18207
rect 1961 18173 1995 18207
rect 3065 18173 3099 18207
rect 3525 18173 3559 18207
rect 4997 18173 5031 18207
rect 5181 18173 5215 18207
rect 6837 18173 6871 18207
rect 7389 18173 7423 18207
rect 9045 18173 9079 18207
rect 9505 18173 9539 18207
rect 13093 18173 13127 18207
rect 13645 18173 13679 18207
rect 15485 18173 15519 18207
rect 16865 18173 16899 18207
rect 17417 18173 17451 18207
rect 2513 18105 2547 18139
rect 2881 18105 2915 18139
rect 4629 18105 4663 18139
rect 6193 18105 6227 18139
rect 9781 18105 9815 18139
rect 1685 18037 1719 18071
rect 3065 18037 3099 18071
rect 6929 18037 6963 18071
rect 8861 18037 8895 18071
rect 10057 18037 10091 18071
rect 10609 18037 10643 18071
rect 11437 18037 11471 18071
rect 16037 18037 16071 18071
rect 2513 17833 2547 17867
rect 9781 17833 9815 17867
rect 10701 17833 10735 17867
rect 15531 17833 15565 17867
rect 9045 17765 9079 17799
rect 1593 17697 1627 17731
rect 1869 17697 1903 17731
rect 3040 17697 3074 17731
rect 4077 17697 4111 17731
rect 5733 17697 5767 17731
rect 6285 17697 6319 17731
rect 8125 17697 8159 17731
rect 8585 17697 8619 17731
rect 9965 17697 9999 17731
rect 10149 17697 10183 17731
rect 11253 17697 11287 17731
rect 12332 17697 12366 17731
rect 13344 17697 13378 17731
rect 15428 17697 15462 17731
rect 1961 17629 1995 17663
rect 4445 17629 4479 17663
rect 6469 17629 6503 17663
rect 8769 17629 8803 17663
rect 3111 17561 3145 17595
rect 4242 17561 4276 17595
rect 7297 17561 7331 17595
rect 12403 17561 12437 17595
rect 2789 17493 2823 17527
rect 3525 17493 3559 17527
rect 4353 17493 4387 17527
rect 4537 17493 4571 17527
rect 5089 17493 5123 17527
rect 6837 17493 6871 17527
rect 7665 17493 7699 17527
rect 11391 17493 11425 17527
rect 13415 17493 13449 17527
rect 1685 17289 1719 17323
rect 5871 17289 5905 17323
rect 6285 17289 6319 17323
rect 12265 17289 12299 17323
rect 13461 17289 13495 17323
rect 3709 17221 3743 17255
rect 5641 17221 5675 17255
rect 4813 17153 4847 17187
rect 6929 17153 6963 17187
rect 10241 17153 10275 17187
rect 14289 17153 14323 17187
rect 14473 17153 14507 17187
rect 15945 17153 15979 17187
rect 2973 17085 3007 17119
rect 3985 17085 4019 17119
rect 4353 17085 4387 17119
rect 5800 17085 5834 17119
rect 8493 17085 8527 17119
rect 8861 17085 8895 17119
rect 9045 17085 9079 17119
rect 12449 17085 12483 17119
rect 12909 17085 12943 17119
rect 2329 17017 2363 17051
rect 2421 17017 2455 17051
rect 3341 17017 3375 17051
rect 7021 17017 7055 17051
rect 7573 17017 7607 17051
rect 9321 17017 9355 17051
rect 10333 17017 10367 17051
rect 10885 17017 10919 17051
rect 13185 17017 13219 17051
rect 14565 17017 14599 17051
rect 15117 17017 15151 17051
rect 1961 16949 1995 16983
rect 3893 16949 3927 16983
rect 5273 16949 5307 16983
rect 6561 16949 6595 16983
rect 8125 16949 8159 16983
rect 9781 16949 9815 16983
rect 11345 16949 11379 16983
rect 11805 16949 11839 16983
rect 15393 16949 15427 16983
rect 1961 16745 1995 16779
rect 2513 16745 2547 16779
rect 2881 16745 2915 16779
rect 6193 16745 6227 16779
rect 6929 16745 6963 16779
rect 8401 16745 8435 16779
rect 10057 16745 10091 16779
rect 10609 16745 10643 16779
rect 10885 16745 10919 16779
rect 12633 16745 12667 16779
rect 14105 16745 14139 16779
rect 14473 16745 14507 16779
rect 19257 16745 19291 16779
rect 5635 16677 5669 16711
rect 7481 16677 7515 16711
rect 13506 16677 13540 16711
rect 1593 16609 1627 16643
rect 5273 16609 5307 16643
rect 9689 16609 9723 16643
rect 11805 16609 11839 16643
rect 12081 16609 12115 16643
rect 15368 16609 15402 16643
rect 19073 16609 19107 16643
rect 4169 16541 4203 16575
rect 7389 16541 7423 16575
rect 12357 16541 12391 16575
rect 13185 16541 13219 16575
rect 3801 16473 3835 16507
rect 4399 16473 4433 16507
rect 5089 16473 5123 16507
rect 7941 16473 7975 16507
rect 9505 16473 9539 16507
rect 15439 16473 15473 16507
rect 3157 16405 3191 16439
rect 4813 16405 4847 16439
rect 8677 16405 8711 16439
rect 1593 16201 1627 16235
rect 2329 16201 2363 16235
rect 4261 16201 4295 16235
rect 6285 16201 6319 16235
rect 7757 16201 7791 16235
rect 8033 16201 8067 16235
rect 8401 16201 8435 16235
rect 8769 16201 8803 16235
rect 11253 16201 11287 16235
rect 12081 16201 12115 16235
rect 16267 16133 16301 16167
rect 4721 16065 4755 16099
rect 6837 16065 6871 16099
rect 9689 16065 9723 16099
rect 10885 16065 10919 16099
rect 1409 15997 1443 16031
rect 3617 15997 3651 16031
rect 8585 15997 8619 16031
rect 13369 15997 13403 16031
rect 14565 15997 14599 16031
rect 15184 15997 15218 16031
rect 16164 15997 16198 16031
rect 16589 15997 16623 16031
rect 2973 15929 3007 15963
rect 3065 15929 3099 15963
rect 3985 15929 4019 15963
rect 4813 15929 4847 15963
rect 5365 15929 5399 15963
rect 7158 15929 7192 15963
rect 9229 15929 9263 15963
rect 10010 15929 10044 15963
rect 12817 15929 12851 15963
rect 13185 15929 13219 15963
rect 13690 15929 13724 15963
rect 2053 15861 2087 15895
rect 2789 15861 2823 15895
rect 5733 15861 5767 15895
rect 6653 15861 6687 15895
rect 9505 15861 9539 15895
rect 10609 15861 10643 15895
rect 11621 15861 11655 15895
rect 14289 15861 14323 15895
rect 15255 15861 15289 15895
rect 15669 15861 15703 15895
rect 16037 15861 16071 15895
rect 19073 15861 19107 15895
rect 1685 15657 1719 15691
rect 2145 15657 2179 15691
rect 3157 15657 3191 15691
rect 5273 15657 5307 15691
rect 6469 15657 6503 15691
rect 9873 15657 9907 15691
rect 10977 15657 11011 15691
rect 13185 15657 13219 15691
rect 14381 15657 14415 15691
rect 2558 15589 2592 15623
rect 4261 15589 4295 15623
rect 6882 15589 6916 15623
rect 10378 15589 10412 15623
rect 11989 15589 12023 15623
rect 13782 15589 13816 15623
rect 15485 15589 15519 15623
rect 2237 15521 2271 15555
rect 6561 15521 6595 15555
rect 8344 15521 8378 15555
rect 10057 15521 10091 15555
rect 13461 15521 13495 15555
rect 16865 15521 16899 15555
rect 4169 15453 4203 15487
rect 4445 15453 4479 15487
rect 8447 15453 8481 15487
rect 11897 15453 11931 15487
rect 12357 15453 12391 15487
rect 15393 15453 15427 15487
rect 15669 15453 15703 15487
rect 7849 15385 7883 15419
rect 7481 15317 7515 15351
rect 11345 15317 11379 15351
rect 17003 15317 17037 15351
rect 2605 15113 2639 15147
rect 5089 15113 5123 15147
rect 5457 15113 5491 15147
rect 8309 15113 8343 15147
rect 10057 15113 10091 15147
rect 10609 15113 10643 15147
rect 11805 15113 11839 15147
rect 13829 15113 13863 15147
rect 14289 15113 14323 15147
rect 15485 15113 15519 15147
rect 7941 15045 7975 15079
rect 11345 15045 11379 15079
rect 15853 15045 15887 15079
rect 16221 15045 16255 15079
rect 1685 14977 1719 15011
rect 3433 14977 3467 15011
rect 3893 14977 3927 15011
rect 6561 14977 6595 15011
rect 7389 14977 7423 15011
rect 8953 14977 8987 15011
rect 9229 14977 9263 15011
rect 10793 14977 10827 15011
rect 13185 14977 13219 15011
rect 14565 14977 14599 15011
rect 15209 14977 15243 15011
rect 5692 14909 5726 14943
rect 12449 14909 12483 14943
rect 13001 14909 13035 14943
rect 16037 14909 16071 14943
rect 18096 14909 18130 14943
rect 18521 14909 18555 14943
rect 4214 14841 4248 14875
rect 5779 14841 5813 14875
rect 7481 14841 7515 14875
rect 8769 14841 8803 14875
rect 9045 14841 9079 14875
rect 10885 14841 10919 14875
rect 13461 14841 13495 14875
rect 14657 14841 14691 14875
rect 16681 14841 16715 14875
rect 2053 14773 2087 14807
rect 2881 14773 2915 14807
rect 3709 14773 3743 14807
rect 4813 14773 4847 14807
rect 6193 14773 6227 14807
rect 7205 14773 7239 14807
rect 12265 14773 12299 14807
rect 16957 14773 16991 14807
rect 18199 14773 18233 14807
rect 1777 14569 1811 14603
rect 2237 14569 2271 14603
rect 7389 14569 7423 14603
rect 8953 14569 8987 14603
rect 10057 14569 10091 14603
rect 11805 14569 11839 14603
rect 12173 14569 12207 14603
rect 14105 14569 14139 14603
rect 2513 14501 2547 14535
rect 3065 14501 3099 14535
rect 3893 14501 3927 14535
rect 4353 14501 4387 14535
rect 4445 14501 4479 14535
rect 6790 14501 6824 14535
rect 10793 14501 10827 14535
rect 11345 14501 11379 14535
rect 13087 14501 13121 14535
rect 15485 14501 15519 14535
rect 16037 14501 16071 14535
rect 6469 14433 6503 14467
rect 8252 14433 8286 14467
rect 16932 14433 16966 14467
rect 17912 14433 17946 14467
rect 2421 14365 2455 14399
rect 3341 14365 3375 14399
rect 4997 14365 5031 14399
rect 10701 14365 10735 14399
rect 12725 14365 12759 14399
rect 15393 14365 15427 14399
rect 12449 14297 12483 14331
rect 7757 14229 7791 14263
rect 8355 14229 8389 14263
rect 13645 14229 13679 14263
rect 14565 14229 14599 14263
rect 15025 14229 15059 14263
rect 17003 14229 17037 14263
rect 18015 14229 18049 14263
rect 5181 14025 5215 14059
rect 7205 14025 7239 14059
rect 8217 14025 8251 14059
rect 11483 14025 11517 14059
rect 18199 14025 18233 14059
rect 1961 13957 1995 13991
rect 3065 13957 3099 13991
rect 4813 13957 4847 13991
rect 4261 13889 4295 13923
rect 5549 13889 5583 13923
rect 5871 13889 5905 13923
rect 7389 13889 7423 13923
rect 8033 13889 8067 13923
rect 1460 13821 1494 13855
rect 5768 13821 5802 13855
rect 1547 13753 1581 13787
rect 2513 13753 2547 13787
rect 2605 13753 2639 13787
rect 3433 13753 3467 13787
rect 4077 13753 4111 13787
rect 4353 13753 4387 13787
rect 6193 13753 6227 13787
rect 7481 13753 7515 13787
rect 11161 13957 11195 13991
rect 19211 13957 19245 13991
rect 9045 13889 9079 13923
rect 9505 13889 9539 13923
rect 10793 13889 10827 13923
rect 12541 13889 12575 13923
rect 12817 13889 12851 13923
rect 14105 13889 14139 13923
rect 18521 13889 18555 13923
rect 19533 13889 19567 13923
rect 10425 13821 10459 13855
rect 11380 13821 11414 13855
rect 11805 13821 11839 13855
rect 15485 13821 15519 13855
rect 15577 13821 15611 13855
rect 16129 13821 16163 13855
rect 18096 13821 18130 13855
rect 19108 13821 19142 13855
rect 9413 13753 9447 13787
rect 9826 13753 9860 13787
rect 12265 13753 12299 13787
rect 12633 13753 12667 13787
rect 13553 13753 13587 13787
rect 13921 13753 13955 13787
rect 14197 13753 14231 13787
rect 14749 13753 14783 13787
rect 17785 13753 17819 13787
rect 2329 13685 2363 13719
rect 6653 13685 6687 13719
rect 8217 13685 8251 13719
rect 8309 13685 8343 13719
rect 15025 13685 15059 13719
rect 15669 13685 15703 13719
rect 16957 13685 16991 13719
rect 3617 13481 3651 13515
rect 6561 13481 6595 13515
rect 12449 13481 12483 13515
rect 12725 13481 12759 13515
rect 16957 13481 16991 13515
rect 18567 13481 18601 13515
rect 2006 13413 2040 13447
rect 4813 13413 4847 13447
rect 5365 13413 5399 13447
rect 6837 13413 6871 13447
rect 7297 13413 7331 13447
rect 10885 13413 10919 13447
rect 13271 13413 13305 13447
rect 15117 13413 15151 13447
rect 15485 13413 15519 13447
rect 2605 13345 2639 13379
rect 9597 13345 9631 13379
rect 17141 13345 17175 13379
rect 17417 13345 17451 13379
rect 18496 13345 18530 13379
rect 19508 13345 19542 13379
rect 1685 13277 1719 13311
rect 3249 13277 3283 13311
rect 4721 13277 4755 13311
rect 7205 13277 7239 13311
rect 10793 13277 10827 13311
rect 11069 13277 11103 13311
rect 12909 13277 12943 13311
rect 15393 13277 15427 13311
rect 16037 13277 16071 13311
rect 2881 13209 2915 13243
rect 7757 13209 7791 13243
rect 4261 13141 4295 13175
rect 9827 13141 9861 13175
rect 13829 13141 13863 13175
rect 14197 13141 14231 13175
rect 19579 13141 19613 13175
rect 4813 12937 4847 12971
rect 5089 12937 5123 12971
rect 5779 12937 5813 12971
rect 7757 12937 7791 12971
rect 8125 12937 8159 12971
rect 10885 12937 10919 12971
rect 12265 12937 12299 12971
rect 13921 12937 13955 12971
rect 15117 12937 15151 12971
rect 19625 12937 19659 12971
rect 5549 12869 5583 12903
rect 10517 12869 10551 12903
rect 14657 12869 14691 12903
rect 16221 12869 16255 12903
rect 2145 12801 2179 12835
rect 3065 12801 3099 12835
rect 6837 12801 6871 12835
rect 12541 12801 12575 12835
rect 12817 12801 12851 12835
rect 14105 12801 14139 12835
rect 15669 12801 15703 12835
rect 16957 12801 16991 12835
rect 3893 12733 3927 12767
rect 5708 12733 5742 12767
rect 6101 12733 6135 12767
rect 9321 12733 9355 12767
rect 11380 12733 11414 12767
rect 11805 12733 11839 12767
rect 18096 12733 18130 12767
rect 19140 12733 19174 12767
rect 2237 12665 2271 12699
rect 2789 12665 2823 12699
rect 3801 12665 3835 12699
rect 4255 12665 4289 12699
rect 6653 12665 6687 12699
rect 7199 12665 7233 12699
rect 9229 12665 9263 12699
rect 12633 12665 12667 12699
rect 14197 12665 14231 12699
rect 15761 12665 15795 12699
rect 18521 12665 18555 12699
rect 1777 12597 1811 12631
rect 9689 12597 9723 12631
rect 10241 12597 10275 12631
rect 11483 12597 11517 12631
rect 13553 12597 13587 12631
rect 15485 12597 15519 12631
rect 17233 12597 17267 12631
rect 18199 12597 18233 12631
rect 18889 12597 18923 12631
rect 19211 12597 19245 12631
rect 19901 12597 19935 12631
rect 1869 12393 1903 12427
rect 2421 12393 2455 12427
rect 2789 12393 2823 12427
rect 4169 12393 4203 12427
rect 6653 12393 6687 12427
rect 7481 12393 7515 12427
rect 10701 12393 10735 12427
rect 12357 12393 12391 12427
rect 12817 12393 12851 12427
rect 18521 12393 18555 12427
rect 8217 12325 8251 12359
rect 8769 12325 8803 12359
rect 10102 12325 10136 12359
rect 11069 12325 11103 12359
rect 11437 12325 11471 12359
rect 13271 12325 13305 12359
rect 15485 12325 15519 12359
rect 16037 12325 16071 12359
rect 16405 12325 16439 12359
rect 4077 12257 4111 12291
rect 4537 12257 4571 12291
rect 6285 12257 6319 12291
rect 7205 12257 7239 12291
rect 11897 12257 11931 12291
rect 12909 12257 12943 12291
rect 13829 12257 13863 12291
rect 17141 12257 17175 12291
rect 17325 12257 17359 12291
rect 18429 12257 18463 12291
rect 18889 12257 18923 12291
rect 1501 12189 1535 12223
rect 8125 12189 8159 12223
rect 9781 12189 9815 12223
rect 14657 12189 14691 12223
rect 15393 12189 15427 12223
rect 17417 12189 17451 12223
rect 7941 12121 7975 12155
rect 12035 12121 12069 12155
rect 15025 12121 15059 12155
rect 3065 12053 3099 12087
rect 5089 12053 5123 12087
rect 9413 12053 9447 12087
rect 14105 12053 14139 12087
rect 4169 11849 4203 11883
rect 6009 11849 6043 11883
rect 6377 11849 6411 11883
rect 8125 11849 8159 11883
rect 8493 11849 8527 11883
rect 16221 11849 16255 11883
rect 16911 11849 16945 11883
rect 18613 11849 18647 11883
rect 19257 11849 19291 11883
rect 11253 11781 11287 11815
rect 4997 11713 5031 11747
rect 7205 11713 7239 11747
rect 7849 11713 7883 11747
rect 10241 11713 10275 11747
rect 10885 11713 10919 11747
rect 11897 11713 11931 11747
rect 18061 11713 18095 11747
rect 1409 11645 1443 11679
rect 1961 11645 1995 11679
rect 2697 11645 2731 11679
rect 8712 11645 8746 11679
rect 9137 11645 9171 11679
rect 12484 11645 12518 11679
rect 12909 11645 12943 11679
rect 13461 11645 13495 11679
rect 15117 11645 15151 11679
rect 15209 11645 15243 11679
rect 15669 11645 15703 11679
rect 16808 11645 16842 11679
rect 17601 11645 17635 11679
rect 19073 11645 19107 11679
rect 19625 11645 19659 11679
rect 4537 11577 4571 11611
rect 4629 11577 4663 11611
rect 7297 11577 7331 11611
rect 10333 11577 10367 11611
rect 12587 11577 12621 11611
rect 13782 11577 13816 11611
rect 16589 11577 16623 11611
rect 17325 11577 17359 11611
rect 1593 11509 1627 11543
rect 2421 11509 2455 11543
rect 3065 11509 3099 11543
rect 3617 11509 3651 11543
rect 5457 11509 5491 11543
rect 8815 11509 8849 11543
rect 9781 11509 9815 11543
rect 13277 11509 13311 11543
rect 14381 11509 14415 11543
rect 14657 11509 14691 11543
rect 15301 11509 15335 11543
rect 18889 11509 18923 11543
rect 4169 11305 4203 11339
rect 2415 11237 2449 11271
rect 2053 11101 2087 11135
rect 3617 11101 3651 11135
rect 3249 11033 3283 11067
rect 5089 11305 5123 11339
rect 7481 11305 7515 11339
rect 10241 11305 10275 11339
rect 13001 11305 13035 11339
rect 16957 11305 16991 11339
rect 6653 11237 6687 11271
rect 8217 11237 8251 11271
rect 8769 11237 8803 11271
rect 10425 11237 10459 11271
rect 10517 11237 10551 11271
rect 11069 11237 11103 11271
rect 12081 11237 12115 11271
rect 13782 11237 13816 11271
rect 15485 11237 15519 11271
rect 5641 11169 5675 11203
rect 16865 11169 16899 11203
rect 17325 11169 17359 11203
rect 19073 11169 19107 11203
rect 4721 11101 4755 11135
rect 6377 11101 6411 11135
rect 6561 11101 6595 11135
rect 6837 11101 6871 11135
rect 7941 11101 7975 11135
rect 8125 11101 8159 11135
rect 11989 11101 12023 11135
rect 13461 11101 13495 11135
rect 15393 11101 15427 11135
rect 16037 11101 16071 11135
rect 12541 11033 12575 11067
rect 1869 10965 1903 10999
rect 2973 10965 3007 10999
rect 4169 10965 4203 10999
rect 4353 10965 4387 10999
rect 5917 10965 5951 10999
rect 13369 10965 13403 10999
rect 14381 10965 14415 10999
rect 15117 10965 15151 10999
rect 19257 10965 19291 10999
rect 2421 10761 2455 10795
rect 4445 10761 4479 10795
rect 4721 10761 4755 10795
rect 6285 10761 6319 10795
rect 8217 10761 8251 10795
rect 10333 10761 10367 10795
rect 11897 10761 11931 10795
rect 15025 10761 15059 10795
rect 19165 10761 19199 10795
rect 2053 10693 2087 10727
rect 4307 10625 4341 10659
rect 12909 10693 12943 10727
rect 5273 10625 5307 10659
rect 7021 10625 7055 10659
rect 11069 10625 11103 10659
rect 13369 10625 13403 10659
rect 16589 10625 16623 10659
rect 1409 10557 1443 10591
rect 4077 10557 4111 10591
rect 4220 10557 4254 10591
rect 4445 10557 4479 10591
rect 8953 10557 8987 10591
rect 16748 10557 16782 10591
rect 17141 10557 17175 10591
rect 18061 10557 18095 10591
rect 18521 10557 18555 10591
rect 2697 10489 2731 10523
rect 2789 10489 2823 10523
rect 3341 10489 3375 10523
rect 5365 10489 5399 10523
rect 5917 10489 5951 10523
rect 6653 10489 6687 10523
rect 7383 10489 7417 10523
rect 8861 10489 8895 10523
rect 9315 10489 9349 10523
rect 10793 10489 10827 10523
rect 10885 10489 10919 10523
rect 13690 10489 13724 10523
rect 15209 10489 15243 10523
rect 15301 10489 15335 10523
rect 15853 10489 15887 10523
rect 1593 10421 1627 10455
rect 3617 10421 3651 10455
rect 5089 10421 5123 10455
rect 7941 10421 7975 10455
rect 9873 10421 9907 10455
rect 13277 10421 13311 10455
rect 14289 10421 14323 10455
rect 14565 10421 14599 10455
rect 16129 10421 16163 10455
rect 16819 10421 16853 10455
rect 17877 10421 17911 10455
rect 18153 10421 18187 10455
rect 19625 10421 19659 10455
rect 1547 10217 1581 10251
rect 1961 10217 1995 10251
rect 3433 10217 3467 10251
rect 5457 10217 5491 10251
rect 9505 10217 9539 10251
rect 10609 10217 10643 10251
rect 10885 10217 10919 10251
rect 12449 10217 12483 10251
rect 15025 10217 15059 10251
rect 16957 10217 16991 10251
rect 18521 10217 18555 10251
rect 2605 10149 2639 10183
rect 4261 10149 4295 10183
rect 4813 10149 4847 10183
rect 5825 10149 5859 10183
rect 7849 10149 7883 10183
rect 8401 10149 8435 10183
rect 10010 10149 10044 10183
rect 11253 10149 11287 10183
rect 11621 10149 11655 10183
rect 13829 10149 13863 10183
rect 15485 10149 15519 10183
rect 16037 10149 16071 10183
rect 1476 10081 1510 10115
rect 16865 10081 16899 10115
rect 17325 10081 17359 10115
rect 18429 10081 18463 10115
rect 18889 10081 18923 10115
rect 2513 10013 2547 10047
rect 3801 10013 3835 10047
rect 4169 10013 4203 10047
rect 5733 10013 5767 10047
rect 6009 10013 6043 10047
rect 6929 10013 6963 10047
rect 7757 10013 7791 10047
rect 9689 10013 9723 10047
rect 11529 10013 11563 10047
rect 11805 10013 11839 10047
rect 13737 10013 13771 10047
rect 14381 10013 14415 10047
rect 15393 10013 15427 10047
rect 18061 10013 18095 10047
rect 3065 9945 3099 9979
rect 2237 9877 2271 9911
rect 5181 9877 5215 9911
rect 7297 9877 7331 9911
rect 9045 9877 9079 9911
rect 13461 9877 13495 9911
rect 14749 9877 14783 9911
rect 2605 9673 2639 9707
rect 2881 9673 2915 9707
rect 3249 9673 3283 9707
rect 5549 9673 5583 9707
rect 5825 9673 5859 9707
rect 6285 9673 6319 9707
rect 11621 9673 11655 9707
rect 13829 9673 13863 9707
rect 14105 9673 14139 9707
rect 14473 9673 14507 9707
rect 17325 9673 17359 9707
rect 3617 9605 3651 9639
rect 9689 9605 9723 9639
rect 10885 9605 10919 9639
rect 15301 9605 15335 9639
rect 6653 9537 6687 9571
rect 7941 9537 7975 9571
rect 8493 9537 8527 9571
rect 11897 9537 11931 9571
rect 14749 9537 14783 9571
rect 19763 9537 19797 9571
rect 1685 9469 1719 9503
rect 3433 9469 3467 9503
rect 4629 9469 4663 9503
rect 6837 9469 6871 9503
rect 7389 9469 7423 9503
rect 9137 9469 9171 9503
rect 9965 9469 9999 9503
rect 12909 9469 12943 9503
rect 16221 9469 16255 9503
rect 16773 9469 16807 9503
rect 18061 9469 18095 9503
rect 18521 9469 18555 9503
rect 19660 9469 19694 9503
rect 20085 9469 20119 9503
rect 2047 9401 2081 9435
rect 4537 9401 4571 9435
rect 4991 9401 5025 9435
rect 8585 9401 8619 9435
rect 10286 9401 10320 9435
rect 11161 9401 11195 9435
rect 12725 9401 12759 9435
rect 13230 9401 13264 9435
rect 14841 9401 14875 9435
rect 16129 9401 16163 9435
rect 19073 9401 19107 9435
rect 4077 9333 4111 9367
rect 6929 9333 6963 9367
rect 8309 9333 8343 9367
rect 15669 9333 15703 9367
rect 16313 9333 16347 9367
rect 17785 9333 17819 9367
rect 18153 9333 18187 9367
rect 1685 9129 1719 9163
rect 3525 9129 3559 9163
rect 6837 9129 6871 9163
rect 7941 9129 7975 9163
rect 8493 9129 8527 9163
rect 12909 9129 12943 9163
rect 15393 9129 15427 9163
rect 16957 9129 16991 9163
rect 18889 9129 18923 9163
rect 5273 9061 5307 9095
rect 5457 9061 5491 9095
rect 5549 9061 5583 9095
rect 6101 9061 6135 9095
rect 7113 9061 7147 9095
rect 9873 9061 9907 9095
rect 10425 9061 10459 9095
rect 11345 9061 11379 9095
rect 11437 9061 11471 9095
rect 11989 9061 12023 9095
rect 13553 9061 13587 9095
rect 13829 9061 13863 9095
rect 14381 9061 14415 9095
rect 15117 9061 15151 9095
rect 18061 9061 18095 9095
rect 1409 8993 1443 9027
rect 1869 8993 1903 9027
rect 3008 8993 3042 9027
rect 3249 8993 3283 9027
rect 4388 8993 4422 9027
rect 8652 8993 8686 9027
rect 9505 8993 9539 9027
rect 15301 8993 15335 9027
rect 15853 8993 15887 9027
rect 16865 8993 16899 9027
rect 17325 8993 17359 9027
rect 18496 8993 18530 9027
rect 19476 8993 19510 9027
rect 2513 8925 2547 8959
rect 4491 8925 4525 8959
rect 7021 8925 7055 8959
rect 9781 8925 9815 8959
rect 10793 8925 10827 8959
rect 13737 8925 13771 8959
rect 16313 8925 16347 8959
rect 7573 8857 7607 8891
rect 9045 8857 9079 8891
rect 2881 8789 2915 8823
rect 3893 8789 3927 8823
rect 4813 8789 4847 8823
rect 6377 8789 6411 8823
rect 8723 8789 8757 8823
rect 11069 8789 11103 8823
rect 14749 8789 14783 8823
rect 16681 8789 16715 8823
rect 18567 8789 18601 8823
rect 19579 8789 19613 8823
rect 2789 8585 2823 8619
rect 5641 8585 5675 8619
rect 6101 8585 6135 8619
rect 8585 8585 8619 8619
rect 9597 8585 9631 8619
rect 9873 8585 9907 8619
rect 11713 8585 11747 8619
rect 12725 8585 12759 8619
rect 13737 8585 13771 8619
rect 14013 8585 14047 8619
rect 19763 8585 19797 8619
rect 4445 8517 4479 8551
rect 4077 8449 4111 8483
rect 7205 8449 7239 8483
rect 11069 8449 11103 8483
rect 12265 8449 12299 8483
rect 12817 8449 12851 8483
rect 14933 8449 14967 8483
rect 15669 8449 15703 8483
rect 16037 8449 16071 8483
rect 17785 8449 17819 8483
rect 1685 8381 1719 8415
rect 1961 8381 1995 8415
rect 3249 8381 3283 8415
rect 3525 8381 3559 8415
rect 4537 8381 4571 8415
rect 5089 8381 5123 8415
rect 6101 8381 6135 8415
rect 8217 8381 8251 8415
rect 8677 8381 8711 8415
rect 16129 8381 16163 8415
rect 16589 8381 16623 8415
rect 17141 8381 17175 8415
rect 18153 8381 18187 8415
rect 19692 8381 19726 8415
rect 20085 8381 20119 8415
rect 2145 8313 2179 8347
rect 6285 8313 6319 8347
rect 6929 8313 6963 8347
rect 7021 8313 7055 8347
rect 9039 8313 9073 8347
rect 10793 8313 10827 8347
rect 10885 8313 10919 8347
rect 13138 8313 13172 8347
rect 14657 8313 14691 8347
rect 14749 8313 14783 8347
rect 19441 8313 19475 8347
rect 2513 8245 2547 8279
rect 3065 8245 3099 8279
rect 4629 8245 4663 8279
rect 6653 8245 6687 8279
rect 10609 8245 10643 8279
rect 14381 8245 14415 8279
rect 16221 8245 16255 8279
rect 18521 8245 18555 8279
rect 19073 8245 19107 8279
rect 1501 8041 1535 8075
rect 2513 8041 2547 8075
rect 3433 8041 3467 8075
rect 4445 8041 4479 8075
rect 5917 8041 5951 8075
rect 11989 8041 12023 8075
rect 14565 8041 14599 8075
rect 14841 8041 14875 8075
rect 15025 8041 15059 8075
rect 19073 8041 19107 8075
rect 2789 7973 2823 8007
rect 5365 7973 5399 8007
rect 7481 7973 7515 8007
rect 9505 7973 9539 8007
rect 10102 7973 10136 8007
rect 11345 7973 11379 8007
rect 13046 7973 13080 8007
rect 14013 7973 14047 8007
rect 15485 7973 15519 8007
rect 16773 7973 16807 8007
rect 1593 7905 1627 7939
rect 1961 7905 1995 7939
rect 3040 7905 3074 7939
rect 4169 7905 4203 7939
rect 4353 7905 4387 7939
rect 6469 7905 6503 7939
rect 8769 7905 8803 7939
rect 11437 7905 11471 7939
rect 13645 7905 13679 7939
rect 14841 7905 14875 7939
rect 16129 7905 16163 7939
rect 16957 7905 16991 7939
rect 18429 7905 18463 7939
rect 5549 7837 5583 7871
rect 7389 7837 7423 7871
rect 7665 7837 7699 7871
rect 9781 7837 9815 7871
rect 12725 7837 12759 7871
rect 15393 7837 15427 7871
rect 16865 7837 16899 7871
rect 18797 7837 18831 7871
rect 6929 7769 6963 7803
rect 10701 7769 10735 7803
rect 3249 7701 3283 7735
rect 3893 7701 3927 7735
rect 5089 7701 5123 7735
rect 8401 7701 8435 7735
rect 9045 7701 9079 7735
rect 11667 7701 11701 7735
rect 16313 7701 16347 7735
rect 18567 7701 18601 7735
rect 18705 7701 18739 7735
rect 1685 7497 1719 7531
rect 9689 7497 9723 7531
rect 12725 7497 12759 7531
rect 12909 7497 12943 7531
rect 13277 7497 13311 7531
rect 16313 7497 16347 7531
rect 3065 7429 3099 7463
rect 3985 7429 4019 7463
rect 4215 7429 4249 7463
rect 4353 7429 4387 7463
rect 5089 7429 5123 7463
rect 5641 7429 5675 7463
rect 10977 7429 11011 7463
rect 3617 7361 3651 7395
rect 4445 7361 4479 7395
rect 4813 7361 4847 7395
rect 9965 7361 9999 7395
rect 13829 7361 13863 7395
rect 14473 7361 14507 7395
rect 15209 7361 15243 7395
rect 18061 7361 18095 7395
rect 2421 7293 2455 7327
rect 5784 7293 5818 7327
rect 6193 7293 6227 7327
rect 8309 7293 8343 7327
rect 8585 7293 8619 7327
rect 8953 7293 8987 7327
rect 12516 7293 12550 7327
rect 12725 7293 12759 7327
rect 15301 7293 15335 7327
rect 15853 7293 15887 7327
rect 16900 7293 16934 7327
rect 17325 7293 17359 7327
rect 17785 7293 17819 7327
rect 18153 7293 18187 7327
rect 19441 7293 19475 7327
rect 1777 7225 1811 7259
rect 4077 7225 4111 7259
rect 5871 7225 5905 7259
rect 6929 7225 6963 7259
rect 7021 7225 7055 7259
rect 7573 7225 7607 7259
rect 8401 7225 8435 7259
rect 10057 7225 10091 7259
rect 10609 7225 10643 7259
rect 11621 7225 11655 7259
rect 13921 7225 13955 7259
rect 19625 7225 19659 7259
rect 6561 7157 6595 7191
rect 7849 7157 7883 7191
rect 9321 7157 9355 7191
rect 12587 7157 12621 7191
rect 14749 7157 14783 7191
rect 15393 7157 15427 7191
rect 16681 7157 16715 7191
rect 17003 7157 17037 7191
rect 19073 7157 19107 7191
rect 2973 6953 3007 6987
rect 5181 6953 5215 6987
rect 9505 6953 9539 6987
rect 10701 6953 10735 6987
rect 12725 6953 12759 6987
rect 14657 6953 14691 6987
rect 18889 6953 18923 6987
rect 19257 6953 19291 6987
rect 1777 6885 1811 6919
rect 5917 6885 5951 6919
rect 9873 6885 9907 6919
rect 10425 6885 10459 6919
rect 11437 6885 11471 6919
rect 13737 6885 13771 6919
rect 15117 6885 15151 6919
rect 18567 6885 18601 6919
rect 4077 6817 4111 6851
rect 5457 6817 5491 6851
rect 5641 6817 5675 6851
rect 7481 6817 7515 6851
rect 7941 6817 7975 6851
rect 15301 6817 15335 6851
rect 15761 6817 15795 6851
rect 16865 6817 16899 6851
rect 17141 6817 17175 6851
rect 18480 6817 18514 6851
rect 19508 6817 19542 6851
rect 1685 6749 1719 6783
rect 4224 6749 4258 6783
rect 4445 6749 4479 6783
rect 8217 6749 8251 6783
rect 9781 6749 9815 6783
rect 11345 6749 11379 6783
rect 11621 6749 11655 6783
rect 13645 6749 13679 6783
rect 15853 6749 15887 6783
rect 16957 6749 16991 6783
rect 17325 6749 17359 6783
rect 2237 6681 2271 6715
rect 4537 6681 4571 6715
rect 11069 6681 11103 6715
rect 14197 6681 14231 6715
rect 19579 6681 19613 6715
rect 2697 6613 2731 6647
rect 3433 6613 3467 6647
rect 3893 6613 3927 6647
rect 4353 6613 4387 6647
rect 6561 6613 6595 6647
rect 6837 6613 6871 6647
rect 7297 6613 7331 6647
rect 8585 6613 8619 6647
rect 8861 6613 8895 6647
rect 1685 6409 1719 6443
rect 3709 6409 3743 6443
rect 5733 6409 5767 6443
rect 6009 6409 6043 6443
rect 8033 6409 8067 6443
rect 11345 6409 11379 6443
rect 12265 6409 12299 6443
rect 13369 6409 13403 6443
rect 13737 6409 13771 6443
rect 14013 6409 14047 6443
rect 15301 6409 15335 6443
rect 16865 6409 16899 6443
rect 17601 6409 17635 6443
rect 18613 6409 18647 6443
rect 19625 6409 19659 6443
rect 19901 6409 19935 6443
rect 3433 6341 3467 6375
rect 9137 6341 9171 6375
rect 19211 6341 19245 6375
rect 2053 6273 2087 6307
rect 2329 6273 2363 6307
rect 5365 6273 5399 6307
rect 7389 6273 7423 6307
rect 10333 6273 10367 6307
rect 14289 6273 14323 6307
rect 3525 6205 3559 6239
rect 4905 6205 4939 6239
rect 5457 6205 5491 6239
rect 6561 6205 6595 6239
rect 7021 6205 7055 6239
rect 8217 6205 8251 6239
rect 11897 6205 11931 6239
rect 12449 6205 12483 6239
rect 15761 6205 15795 6239
rect 16221 6205 16255 6239
rect 19140 6205 19174 6239
rect 2145 6137 2179 6171
rect 3065 6137 3099 6171
rect 4537 6137 4571 6171
rect 6837 6137 6871 6171
rect 7665 6137 7699 6171
rect 8538 6137 8572 6171
rect 10057 6137 10091 6171
rect 10149 6137 10183 6171
rect 14381 6137 14415 6171
rect 14933 6137 14967 6171
rect 17233 6137 17267 6171
rect 4077 6069 4111 6103
rect 9413 6069 9447 6103
rect 9781 6069 9815 6103
rect 12817 6069 12851 6103
rect 15577 6069 15611 6103
rect 16037 6069 16071 6103
rect 18061 6069 18095 6103
rect 2881 5865 2915 5899
rect 4261 5865 4295 5899
rect 5457 5865 5491 5899
rect 8769 5865 8803 5899
rect 9505 5865 9539 5899
rect 10701 5865 10735 5899
rect 11391 5865 11425 5899
rect 16957 5865 16991 5899
rect 2323 5797 2357 5831
rect 7481 5797 7515 5831
rect 8170 5797 8204 5831
rect 9045 5797 9079 5831
rect 9781 5797 9815 5831
rect 9873 5797 9907 5831
rect 12862 5797 12896 5831
rect 15485 5797 15519 5831
rect 16313 5797 16347 5831
rect 4813 5729 4847 5763
rect 5365 5729 5399 5763
rect 6469 5729 6503 5763
rect 11288 5729 11322 5763
rect 11713 5729 11747 5763
rect 13461 5729 13495 5763
rect 13829 5729 13863 5763
rect 14289 5729 14323 5763
rect 15117 5729 15151 5763
rect 16865 5729 16899 5763
rect 17325 5729 17359 5763
rect 18429 5729 18463 5763
rect 19476 5729 19510 5763
rect 1961 5661 1995 5695
rect 5273 5661 5307 5695
rect 7849 5661 7883 5695
rect 10149 5661 10183 5695
rect 12541 5661 12575 5695
rect 15393 5661 15427 5695
rect 15669 5661 15703 5695
rect 19579 5661 19613 5695
rect 3433 5593 3467 5627
rect 18567 5593 18601 5627
rect 1685 5525 1719 5559
rect 3801 5525 3835 5559
rect 6009 5525 6043 5559
rect 6377 5525 6411 5559
rect 6607 5525 6641 5559
rect 7021 5525 7055 5559
rect 11069 5525 11103 5559
rect 2513 5321 2547 5355
rect 4445 5321 4479 5355
rect 8033 5321 8067 5355
rect 9321 5321 9355 5355
rect 9781 5321 9815 5355
rect 11253 5321 11287 5355
rect 12265 5321 12299 5355
rect 15393 5321 15427 5355
rect 17325 5321 17359 5355
rect 19211 5321 19245 5355
rect 7573 5253 7607 5287
rect 10517 5253 10551 5287
rect 11621 5253 11655 5287
rect 12725 5253 12759 5287
rect 13921 5253 13955 5287
rect 19533 5253 19567 5287
rect 2053 5185 2087 5219
rect 5181 5185 5215 5219
rect 7389 5185 7423 5219
rect 9965 5185 9999 5219
rect 12909 5185 12943 5219
rect 13553 5185 13587 5219
rect 15945 5185 15979 5219
rect 19901 5185 19935 5219
rect 3249 5117 3283 5151
rect 3617 5117 3651 5151
rect 4123 5117 4157 5151
rect 4353 5117 4387 5151
rect 5273 5117 5307 5151
rect 5457 5117 5491 5151
rect 7180 5117 7214 5151
rect 8125 5117 8159 5151
rect 15669 5117 15703 5151
rect 16037 5117 16071 5151
rect 18128 5117 18162 5151
rect 18889 5117 18923 5151
rect 19140 5117 19174 5151
rect 1593 5049 1627 5083
rect 1685 5049 1719 5083
rect 6193 5049 6227 5083
rect 8446 5049 8480 5083
rect 10057 5049 10091 5083
rect 13001 5049 13035 5083
rect 14473 5049 14507 5083
rect 14565 5049 14599 5083
rect 15117 5049 15151 5083
rect 4813 4981 4847 5015
rect 5549 4981 5583 5015
rect 6469 4981 6503 5015
rect 9045 4981 9079 5015
rect 10885 4981 10919 5015
rect 14289 4981 14323 5015
rect 15669 4981 15703 5015
rect 15761 4981 15795 5015
rect 17049 4981 17083 5015
rect 18199 4981 18233 5015
rect 18521 4981 18555 5015
rect 2881 4777 2915 4811
rect 3433 4777 3467 4811
rect 4169 4777 4203 4811
rect 7021 4777 7055 4811
rect 7481 4777 7515 4811
rect 7849 4777 7883 4811
rect 8953 4777 8987 4811
rect 9321 4777 9355 4811
rect 10701 4777 10735 4811
rect 12173 4777 12207 4811
rect 14381 4777 14415 4811
rect 16957 4777 16991 4811
rect 1955 4709 1989 4743
rect 9873 4709 9907 4743
rect 11615 4709 11649 4743
rect 12909 4709 12943 4743
rect 13185 4709 13219 4743
rect 13737 4709 13771 4743
rect 1593 4641 1627 4675
rect 3893 4641 3927 4675
rect 4353 4641 4387 4675
rect 4905 4641 4939 4675
rect 5089 4641 5123 4675
rect 6009 4641 6043 4675
rect 6285 4641 6319 4675
rect 7941 4641 7975 4675
rect 8401 4641 8435 4675
rect 15025 4641 15059 4675
rect 15393 4641 15427 4675
rect 15761 4641 15795 4675
rect 16865 4641 16899 4675
rect 17325 4641 17359 4675
rect 18429 4641 18463 4675
rect 19568 4641 19602 4675
rect 6745 4573 6779 4607
rect 8677 4573 8711 4607
rect 9781 4573 9815 4607
rect 10149 4573 10183 4607
rect 11253 4573 11287 4607
rect 13093 4573 13127 4607
rect 15853 4573 15887 4607
rect 2513 4505 2547 4539
rect 5549 4505 5583 4539
rect 6101 4505 6135 4539
rect 11069 4505 11103 4539
rect 12449 4505 12483 4539
rect 19671 4505 19705 4539
rect 5917 4437 5951 4471
rect 14105 4437 14139 4471
rect 18613 4437 18647 4471
rect 2697 4233 2731 4267
rect 3525 4233 3559 4267
rect 6653 4233 6687 4267
rect 8217 4233 8251 4267
rect 9873 4233 9907 4267
rect 12587 4233 12621 4267
rect 13369 4233 13403 4267
rect 14473 4233 14507 4267
rect 14749 4233 14783 4267
rect 16681 4233 16715 4267
rect 19165 4233 19199 4267
rect 20085 4233 20119 4267
rect 5273 4165 5307 4199
rect 11345 4165 11379 4199
rect 11713 4165 11747 4199
rect 18337 4165 18371 4199
rect 1685 4097 1719 4131
rect 2053 4097 2087 4131
rect 4353 4097 4387 4131
rect 8309 4097 8343 4131
rect 10149 4097 10183 4131
rect 10425 4097 10459 4131
rect 12265 4097 12299 4131
rect 13553 4097 13587 4131
rect 3893 4029 3927 4063
rect 4077 4029 4111 4063
rect 5181 4029 5215 4063
rect 5457 4029 5491 4063
rect 6837 4029 6871 4063
rect 7021 4029 7055 4063
rect 7389 4029 7423 4063
rect 9229 4029 9263 4063
rect 12516 4029 12550 4063
rect 17785 4029 17819 4063
rect 18337 4029 18371 4063
rect 19660 4029 19694 4063
rect 20453 4029 20487 4063
rect 1777 3961 1811 3995
rect 7665 3961 7699 3995
rect 8650 3961 8684 3995
rect 10241 3961 10275 3995
rect 13001 3961 13035 3995
rect 15393 3961 15427 3995
rect 15485 3961 15519 3995
rect 16037 3961 16071 3995
rect 19763 3961 19797 3995
rect 3157 3893 3191 3927
rect 4721 3893 4755 3927
rect 5089 3893 5123 3927
rect 5641 3893 5675 3927
rect 6193 3893 6227 3927
rect 9505 3893 9539 3927
rect 13921 3893 13955 3927
rect 15117 3893 15151 3927
rect 16313 3893 16347 3927
rect 16865 3893 16899 3927
rect 17325 3893 17359 3927
rect 2145 3689 2179 3723
rect 3709 3689 3743 3723
rect 4629 3689 4663 3723
rect 7573 3689 7607 3723
rect 9413 3689 9447 3723
rect 10701 3689 10735 3723
rect 13093 3689 13127 3723
rect 14381 3689 14415 3723
rect 16313 3689 16347 3723
rect 16957 3689 16991 3723
rect 7205 3621 7239 3655
rect 8217 3621 8251 3655
rect 9873 3621 9907 3655
rect 12081 3621 12115 3655
rect 13823 3621 13857 3655
rect 2605 3553 2639 3587
rect 3065 3553 3099 3587
rect 4123 3553 4157 3587
rect 4905 3553 4939 3587
rect 5089 3553 5123 3587
rect 5365 3553 5399 3587
rect 6653 3553 6687 3587
rect 6837 3553 6871 3587
rect 12633 3553 12667 3587
rect 15025 3553 15059 3587
rect 15577 3553 15611 3587
rect 17141 3553 17175 3587
rect 17325 3553 17359 3587
rect 19073 3553 19107 3587
rect 5825 3485 5859 3519
rect 7849 3485 7883 3519
rect 8125 3485 8159 3519
rect 9137 3485 9171 3519
rect 9781 3485 9815 3519
rect 11989 3485 12023 3519
rect 13461 3485 13495 3519
rect 15301 3485 15335 3519
rect 18429 3485 18463 3519
rect 4215 3417 4249 3451
rect 5181 3417 5215 3451
rect 6561 3417 6595 3451
rect 8677 3417 8711 3451
rect 10333 3417 10367 3451
rect 11805 3417 11839 3451
rect 1685 3349 1719 3383
rect 2421 3349 2455 3383
rect 6193 3349 6227 3383
rect 11069 3349 11103 3383
rect 14657 3349 14691 3383
rect 1961 3145 1995 3179
rect 2191 3145 2225 3179
rect 6193 3145 6227 3179
rect 8677 3145 8711 3179
rect 9689 3145 9723 3179
rect 9965 3145 9999 3179
rect 13921 3145 13955 3179
rect 17325 3145 17359 3179
rect 2329 3077 2363 3111
rect 3525 3077 3559 3111
rect 7941 3077 7975 3111
rect 10333 3077 10367 3111
rect 14289 3077 14323 3111
rect 2421 3009 2455 3043
rect 2789 3009 2823 3043
rect 4261 3009 4295 3043
rect 7021 3009 7055 3043
rect 8769 3009 8803 3043
rect 10517 3009 10551 3043
rect 14473 3009 14507 3043
rect 15577 3009 15611 3043
rect 18061 3009 18095 3043
rect 2053 2941 2087 2975
rect 3617 2941 3651 2975
rect 3709 2941 3743 2975
rect 3893 2941 3927 2975
rect 5457 2941 5491 2975
rect 5641 2941 5675 2975
rect 5917 2941 5951 2975
rect 10609 2941 10643 2975
rect 12081 2941 12115 2975
rect 12449 2941 12483 2975
rect 12909 2941 12943 2975
rect 13553 2941 13587 2975
rect 15117 2941 15151 2975
rect 6561 2873 6595 2907
rect 7383 2873 7417 2907
rect 9090 2873 9124 2907
rect 12173 2873 12207 2907
rect 14565 2873 14599 2907
rect 16221 2941 16255 2975
rect 16405 2941 16439 2975
rect 16957 2941 16991 2975
rect 18153 2941 18187 2975
rect 15761 2873 15795 2907
rect 19625 2873 19659 2907
rect 3065 2805 3099 2839
rect 4721 2805 4755 2839
rect 5089 2805 5123 2839
rect 8309 2805 8343 2839
rect 11805 2805 11839 2839
rect 12081 2805 12115 2839
rect 12725 2805 12759 2839
rect 15393 2805 15427 2839
rect 15577 2805 15611 2839
rect 16773 2805 16807 2839
rect 17785 2805 17819 2839
rect 19073 2805 19107 2839
rect 3709 2601 3743 2635
rect 4353 2601 4387 2635
rect 8493 2601 8527 2635
rect 9873 2601 9907 2635
rect 10793 2601 10827 2635
rect 11161 2601 11195 2635
rect 12449 2601 12483 2635
rect 12817 2601 12851 2635
rect 13277 2601 13311 2635
rect 14289 2601 14323 2635
rect 16589 2601 16623 2635
rect 17601 2601 17635 2635
rect 18797 2601 18831 2635
rect 2973 2533 3007 2567
rect 4813 2533 4847 2567
rect 6653 2533 6687 2567
rect 9505 2533 9539 2567
rect 12081 2533 12115 2567
rect 13690 2533 13724 2567
rect 2237 2465 2271 2499
rect 2513 2465 2547 2499
rect 3341 2465 3375 2499
rect 4169 2465 4203 2499
rect 5273 2465 5307 2499
rect 5549 2465 5583 2499
rect 7205 2465 7239 2499
rect 7389 2465 7423 2499
rect 8309 2465 8343 2499
rect 8493 2465 8527 2499
rect 8585 2465 8619 2499
rect 9137 2465 9171 2499
rect 9321 2465 9355 2499
rect 9781 2465 9815 2499
rect 10241 2465 10275 2499
rect 11437 2465 11471 2499
rect 13369 2465 13403 2499
rect 15485 2465 15519 2499
rect 15577 2465 15611 2499
rect 15761 2465 15795 2499
rect 17049 2465 17083 2499
rect 18429 2465 18463 2499
rect 6009 2397 6043 2431
rect 6377 2397 6411 2431
rect 7481 2397 7515 2431
rect 2329 2329 2363 2363
rect 5365 2329 5399 2363
rect 8769 2329 8803 2363
rect 15945 2397 15979 2431
rect 11621 2329 11655 2363
rect 1685 2261 1719 2295
rect 2053 2261 2087 2295
rect 5089 2261 5123 2295
rect 8033 2261 8067 2295
rect 9321 2261 9355 2295
rect 14841 2261 14875 2295
rect 15209 2261 15243 2295
rect 17233 2261 17267 2295
rect 18061 2261 18095 2295
<< metal1 >>
rect 1104 19610 20884 19632
rect 1104 19558 4648 19610
rect 4700 19558 4712 19610
rect 4764 19558 4776 19610
rect 4828 19558 4840 19610
rect 4892 19558 11982 19610
rect 12034 19558 12046 19610
rect 12098 19558 12110 19610
rect 12162 19558 12174 19610
rect 12226 19558 19315 19610
rect 19367 19558 19379 19610
rect 19431 19558 19443 19610
rect 19495 19558 19507 19610
rect 19559 19558 20884 19610
rect 1104 19536 20884 19558
rect 2547 19499 2605 19505
rect 2547 19465 2559 19499
rect 2593 19496 2605 19499
rect 2866 19496 2872 19508
rect 2593 19468 2872 19496
rect 2593 19465 2605 19468
rect 2547 19459 2605 19465
rect 2866 19456 2872 19468
rect 2924 19456 2930 19508
rect 1118 19252 1124 19304
rect 1176 19292 1182 19304
rect 2444 19295 2502 19301
rect 2444 19292 2456 19295
rect 1176 19264 2456 19292
rect 1176 19252 1182 19264
rect 2444 19261 2456 19264
rect 2490 19292 2502 19295
rect 2869 19295 2927 19301
rect 2869 19292 2881 19295
rect 2490 19264 2881 19292
rect 2490 19261 2502 19264
rect 2444 19255 2502 19261
rect 2869 19261 2881 19264
rect 2915 19261 2927 19295
rect 5258 19292 5264 19304
rect 5219 19264 5264 19292
rect 2869 19255 2927 19261
rect 5258 19252 5264 19264
rect 5316 19252 5322 19304
rect 5813 19295 5871 19301
rect 5813 19261 5825 19295
rect 5859 19292 5871 19295
rect 6270 19292 6276 19304
rect 5859 19264 6276 19292
rect 5859 19261 5871 19264
rect 5813 19255 5871 19261
rect 1302 19184 1308 19236
rect 1360 19224 1366 19236
rect 1857 19227 1915 19233
rect 1857 19224 1869 19227
rect 1360 19196 1869 19224
rect 1360 19184 1366 19196
rect 1857 19193 1869 19196
rect 1903 19193 1915 19227
rect 1857 19187 1915 19193
rect 5169 19227 5227 19233
rect 5169 19193 5181 19227
rect 5215 19224 5227 19227
rect 5828 19224 5856 19255
rect 6270 19252 6276 19264
rect 6328 19252 6334 19304
rect 7996 19295 8054 19301
rect 7996 19292 8008 19295
rect 6380 19264 8008 19292
rect 5994 19224 6000 19236
rect 5215 19196 5856 19224
rect 5955 19196 6000 19224
rect 5215 19193 5227 19196
rect 5169 19187 5227 19193
rect 5994 19184 6000 19196
rect 6052 19184 6058 19236
rect 1397 19159 1455 19165
rect 1397 19125 1409 19159
rect 1443 19156 1455 19159
rect 1486 19156 1492 19168
rect 1443 19128 1492 19156
rect 1443 19125 1455 19128
rect 1397 19119 1455 19125
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 4062 19156 4068 19168
rect 4023 19128 4068 19156
rect 4062 19116 4068 19128
rect 4120 19116 4126 19168
rect 5626 19116 5632 19168
rect 5684 19156 5690 19168
rect 6380 19156 6408 19264
rect 7996 19261 8008 19264
rect 8042 19292 8054 19295
rect 8389 19295 8447 19301
rect 8389 19292 8401 19295
rect 8042 19264 8401 19292
rect 8042 19261 8054 19264
rect 7996 19255 8054 19261
rect 8389 19261 8401 19264
rect 8435 19261 8447 19295
rect 8389 19255 8447 19261
rect 9836 19295 9894 19301
rect 9836 19261 9848 19295
rect 9882 19292 9894 19295
rect 10816 19295 10874 19301
rect 10816 19292 10828 19295
rect 9882 19264 10828 19292
rect 9882 19261 9894 19264
rect 9836 19255 9894 19261
rect 10336 19168 10364 19264
rect 10816 19261 10828 19264
rect 10862 19292 10874 19295
rect 11241 19295 11299 19301
rect 11241 19292 11253 19295
rect 10862 19264 11253 19292
rect 10862 19261 10874 19264
rect 10816 19255 10874 19261
rect 11241 19261 11253 19264
rect 11287 19261 11299 19295
rect 11241 19255 11299 19261
rect 6914 19156 6920 19168
rect 5684 19128 6408 19156
rect 6875 19128 6920 19156
rect 5684 19116 5690 19128
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 8067 19159 8125 19165
rect 8067 19125 8079 19159
rect 8113 19156 8125 19159
rect 8202 19156 8208 19168
rect 8113 19128 8208 19156
rect 8113 19125 8125 19128
rect 8067 19119 8125 19125
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 9214 19116 9220 19168
rect 9272 19156 9278 19168
rect 9907 19159 9965 19165
rect 9907 19156 9919 19159
rect 9272 19128 9919 19156
rect 9272 19116 9278 19128
rect 9907 19125 9919 19128
rect 9953 19125 9965 19159
rect 10318 19156 10324 19168
rect 10279 19128 10324 19156
rect 9907 19119 9965 19125
rect 10318 19116 10324 19128
rect 10376 19116 10382 19168
rect 10919 19159 10977 19165
rect 10919 19125 10931 19159
rect 10965 19156 10977 19159
rect 11146 19156 11152 19168
rect 10965 19128 11152 19156
rect 10965 19125 10977 19128
rect 10919 19119 10977 19125
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 1104 19066 20884 19088
rect 1104 19014 8315 19066
rect 8367 19014 8379 19066
rect 8431 19014 8443 19066
rect 8495 19014 8507 19066
rect 8559 19014 15648 19066
rect 15700 19014 15712 19066
rect 15764 19014 15776 19066
rect 15828 19014 15840 19066
rect 15892 19014 20884 19066
rect 1104 18992 20884 19014
rect 2222 18952 2228 18964
rect 2183 18924 2228 18952
rect 2222 18912 2228 18924
rect 2280 18912 2286 18964
rect 4847 18955 4905 18961
rect 4847 18921 4859 18955
rect 4893 18952 4905 18955
rect 5074 18952 5080 18964
rect 4893 18924 5080 18952
rect 4893 18921 4905 18924
rect 4847 18915 4905 18921
rect 5074 18912 5080 18924
rect 5132 18912 5138 18964
rect 5258 18952 5264 18964
rect 5219 18924 5264 18952
rect 5258 18912 5264 18924
rect 5316 18912 5322 18964
rect 6546 18912 6552 18964
rect 6604 18952 6610 18964
rect 7377 18955 7435 18961
rect 7377 18952 7389 18955
rect 6604 18924 7389 18952
rect 6604 18912 6610 18924
rect 7377 18921 7389 18924
rect 7423 18921 7435 18955
rect 7377 18915 7435 18921
rect 11563 18955 11621 18961
rect 11563 18921 11575 18955
rect 11609 18952 11621 18955
rect 21542 18952 21548 18964
rect 11609 18924 21548 18952
rect 11609 18921 11621 18924
rect 11563 18915 11621 18921
rect 21542 18912 21548 18924
rect 21600 18912 21606 18964
rect 2225 18819 2283 18825
rect 2225 18785 2237 18819
rect 2271 18816 2283 18819
rect 2314 18816 2320 18828
rect 2271 18788 2320 18816
rect 2271 18785 2283 18788
rect 2225 18779 2283 18785
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 2409 18819 2467 18825
rect 2409 18785 2421 18819
rect 2455 18785 2467 18819
rect 2409 18779 2467 18785
rect 4776 18819 4834 18825
rect 4776 18785 4788 18819
rect 4822 18816 4834 18819
rect 5074 18816 5080 18828
rect 4822 18788 5080 18816
rect 4822 18785 4834 18788
rect 4776 18779 4834 18785
rect 2424 18748 2452 18779
rect 5074 18776 5080 18788
rect 5132 18776 5138 18828
rect 5997 18819 6055 18825
rect 5997 18785 6009 18819
rect 6043 18816 6055 18819
rect 6086 18816 6092 18828
rect 6043 18788 6092 18816
rect 6043 18785 6055 18788
rect 5997 18779 6055 18785
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 6270 18816 6276 18828
rect 6231 18788 6276 18816
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 7558 18816 7564 18828
rect 7519 18788 7564 18816
rect 7558 18776 7564 18788
rect 7616 18776 7622 18828
rect 7834 18816 7840 18828
rect 7795 18788 7840 18816
rect 7834 18776 7840 18788
rect 7892 18776 7898 18828
rect 9585 18819 9643 18825
rect 9585 18785 9597 18819
rect 9631 18816 9643 18819
rect 9674 18816 9680 18828
rect 9631 18788 9680 18816
rect 9631 18785 9643 18788
rect 9585 18779 9643 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 11422 18816 11428 18828
rect 11383 18788 11428 18816
rect 11422 18776 11428 18788
rect 11480 18776 11486 18828
rect 6362 18748 6368 18760
rect 1872 18720 2452 18748
rect 6323 18720 6368 18748
rect 1872 18624 1900 18720
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 2682 18640 2688 18692
rect 2740 18680 2746 18692
rect 5258 18680 5264 18692
rect 2740 18652 5264 18680
rect 2740 18640 2746 18652
rect 5258 18640 5264 18652
rect 5316 18640 5322 18692
rect 1673 18615 1731 18621
rect 1673 18581 1685 18615
rect 1719 18612 1731 18615
rect 1854 18612 1860 18624
rect 1719 18584 1860 18612
rect 1719 18581 1731 18584
rect 1673 18575 1731 18581
rect 1854 18572 1860 18584
rect 1912 18572 1918 18624
rect 3050 18612 3056 18624
rect 3011 18584 3056 18612
rect 3050 18572 3056 18584
rect 3108 18572 3114 18624
rect 8938 18572 8944 18624
rect 8996 18612 9002 18624
rect 9815 18615 9873 18621
rect 9815 18612 9827 18615
rect 8996 18584 9827 18612
rect 8996 18572 9002 18584
rect 9815 18581 9827 18584
rect 9861 18581 9873 18615
rect 9815 18575 9873 18581
rect 1104 18522 20884 18544
rect 1104 18470 4648 18522
rect 4700 18470 4712 18522
rect 4764 18470 4776 18522
rect 4828 18470 4840 18522
rect 4892 18470 11982 18522
rect 12034 18470 12046 18522
rect 12098 18470 12110 18522
rect 12162 18470 12174 18522
rect 12226 18470 19315 18522
rect 19367 18470 19379 18522
rect 19431 18470 19443 18522
rect 19495 18470 19507 18522
rect 19559 18470 20884 18522
rect 1104 18448 20884 18470
rect 4249 18411 4307 18417
rect 4249 18377 4261 18411
rect 4295 18408 4307 18411
rect 4433 18411 4491 18417
rect 4433 18408 4445 18411
rect 4295 18380 4445 18408
rect 4295 18377 4307 18380
rect 4249 18371 4307 18377
rect 4433 18377 4445 18380
rect 4479 18408 4491 18411
rect 7834 18408 7840 18420
rect 4479 18380 5028 18408
rect 7795 18380 7840 18408
rect 4479 18377 4491 18380
rect 4433 18371 4491 18377
rect 3510 18300 3516 18352
rect 3568 18340 3574 18352
rect 5000 18340 5028 18380
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 13265 18411 13323 18417
rect 13265 18377 13277 18411
rect 13311 18408 13323 18411
rect 14274 18408 14280 18420
rect 13311 18380 14280 18408
rect 13311 18377 13323 18380
rect 13265 18371 13323 18377
rect 14274 18368 14280 18380
rect 14332 18368 14338 18420
rect 15657 18411 15715 18417
rect 15657 18377 15669 18411
rect 15703 18408 15715 18411
rect 16022 18408 16028 18420
rect 15703 18380 16028 18408
rect 15703 18377 15715 18380
rect 15657 18371 15715 18377
rect 16022 18368 16028 18380
rect 16080 18368 16086 18420
rect 17037 18411 17095 18417
rect 17037 18377 17049 18411
rect 17083 18408 17095 18411
rect 18322 18408 18328 18420
rect 17083 18380 18328 18408
rect 17083 18377 17095 18380
rect 17037 18371 17095 18377
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 8110 18340 8116 18352
rect 3568 18312 4660 18340
rect 3568 18300 3574 18312
rect 4433 18275 4491 18281
rect 4433 18272 4445 18275
rect 3068 18244 4445 18272
rect 3068 18216 3096 18244
rect 4433 18241 4445 18244
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 1302 18164 1308 18216
rect 1360 18204 1366 18216
rect 1397 18207 1455 18213
rect 1397 18204 1409 18207
rect 1360 18176 1409 18204
rect 1360 18164 1366 18176
rect 1397 18173 1409 18176
rect 1443 18173 1455 18207
rect 1397 18167 1455 18173
rect 1949 18207 2007 18213
rect 1949 18173 1961 18207
rect 1995 18173 2007 18207
rect 3050 18204 3056 18216
rect 3011 18176 3056 18204
rect 1949 18167 2007 18173
rect 1854 18096 1860 18148
rect 1912 18136 1918 18148
rect 1964 18136 1992 18167
rect 3050 18164 3056 18176
rect 3108 18164 3114 18216
rect 3513 18207 3571 18213
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 4338 18204 4344 18216
rect 3559 18176 4344 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 2501 18139 2559 18145
rect 2501 18136 2513 18139
rect 1912 18108 2513 18136
rect 1912 18096 1918 18108
rect 2501 18105 2513 18108
rect 2547 18136 2559 18139
rect 2869 18139 2927 18145
rect 2869 18136 2881 18139
rect 2547 18108 2881 18136
rect 2547 18105 2559 18108
rect 2501 18099 2559 18105
rect 2869 18105 2881 18108
rect 2915 18136 2927 18139
rect 3528 18136 3556 18167
rect 4338 18164 4344 18176
rect 4396 18164 4402 18216
rect 4632 18145 4660 18312
rect 5000 18312 8116 18340
rect 5000 18213 5028 18312
rect 8110 18300 8116 18312
rect 8168 18300 8174 18352
rect 5258 18272 5264 18284
rect 5219 18244 5264 18272
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 5813 18275 5871 18281
rect 5813 18241 5825 18275
rect 5859 18272 5871 18275
rect 6270 18272 6276 18284
rect 5859 18244 6276 18272
rect 5859 18241 5871 18244
rect 5813 18235 5871 18241
rect 4985 18207 5043 18213
rect 4985 18173 4997 18207
rect 5031 18173 5043 18207
rect 4985 18167 5043 18173
rect 5169 18207 5227 18213
rect 5169 18173 5181 18207
rect 5215 18204 5227 18207
rect 5828 18204 5856 18235
rect 6270 18232 6276 18244
rect 6328 18272 6334 18284
rect 6641 18275 6699 18281
rect 6641 18272 6653 18275
rect 6328 18244 6653 18272
rect 6328 18232 6334 18244
rect 6641 18241 6653 18244
rect 6687 18272 6699 18275
rect 6687 18244 7420 18272
rect 6687 18241 6699 18244
rect 6641 18235 6699 18241
rect 6822 18204 6828 18216
rect 5215 18176 5856 18204
rect 6783 18176 6828 18204
rect 5215 18173 5227 18176
rect 5169 18167 5227 18173
rect 2915 18108 3556 18136
rect 4617 18139 4675 18145
rect 2915 18105 2927 18108
rect 2869 18099 2927 18105
rect 4617 18105 4629 18139
rect 4663 18136 4675 18139
rect 5184 18136 5212 18167
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 7392 18213 7420 18244
rect 7377 18207 7435 18213
rect 7377 18173 7389 18207
rect 7423 18204 7435 18207
rect 7834 18204 7840 18216
rect 7423 18176 7840 18204
rect 7423 18173 7435 18176
rect 7377 18167 7435 18173
rect 7834 18164 7840 18176
rect 7892 18164 7898 18216
rect 9033 18207 9091 18213
rect 9033 18204 9045 18207
rect 8864 18176 9045 18204
rect 4663 18108 5212 18136
rect 4663 18105 4675 18108
rect 4617 18099 4675 18105
rect 6086 18096 6092 18148
rect 6144 18136 6150 18148
rect 6181 18139 6239 18145
rect 6181 18136 6193 18139
rect 6144 18108 6193 18136
rect 6144 18096 6150 18108
rect 6181 18105 6193 18108
rect 6227 18136 6239 18139
rect 7650 18136 7656 18148
rect 6227 18108 7656 18136
rect 6227 18105 6239 18108
rect 6181 18099 6239 18105
rect 7650 18096 7656 18108
rect 7708 18096 7714 18148
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 3050 18068 3056 18080
rect 3011 18040 3056 18068
rect 3050 18028 3056 18040
rect 3108 18028 3114 18080
rect 3142 18028 3148 18080
rect 3200 18068 3206 18080
rect 6104 18068 6132 18096
rect 3200 18040 6132 18068
rect 3200 18028 3206 18040
rect 6730 18028 6736 18080
rect 6788 18068 6794 18080
rect 6917 18071 6975 18077
rect 6917 18068 6929 18071
rect 6788 18040 6929 18068
rect 6788 18028 6794 18040
rect 6917 18037 6929 18040
rect 6963 18037 6975 18071
rect 6917 18031 6975 18037
rect 8662 18028 8668 18080
rect 8720 18068 8726 18080
rect 8864 18077 8892 18176
rect 9033 18173 9045 18176
rect 9079 18173 9091 18207
rect 9033 18167 9091 18173
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 9493 18207 9551 18213
rect 9493 18204 9505 18207
rect 9456 18176 9505 18204
rect 9456 18164 9462 18176
rect 9493 18173 9505 18176
rect 9539 18173 9551 18207
rect 9493 18167 9551 18173
rect 10686 18164 10692 18216
rect 10744 18204 10750 18216
rect 13081 18207 13139 18213
rect 13081 18204 13093 18207
rect 10744 18176 13093 18204
rect 10744 18164 10750 18176
rect 13081 18173 13093 18176
rect 13127 18204 13139 18207
rect 13630 18204 13636 18216
rect 13127 18176 13636 18204
rect 13127 18173 13139 18176
rect 13081 18167 13139 18173
rect 13630 18164 13636 18176
rect 13688 18164 13694 18216
rect 15473 18207 15531 18213
rect 15473 18173 15485 18207
rect 15519 18204 15531 18207
rect 16850 18204 16856 18216
rect 15519 18176 15976 18204
rect 16811 18176 16856 18204
rect 15519 18173 15531 18176
rect 15473 18167 15531 18173
rect 9766 18136 9772 18148
rect 9727 18108 9772 18136
rect 9766 18096 9772 18108
rect 9824 18096 9830 18148
rect 15948 18080 15976 18176
rect 16850 18164 16856 18176
rect 16908 18204 16914 18216
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 16908 18176 17417 18204
rect 16908 18164 16914 18176
rect 17405 18173 17417 18176
rect 17451 18173 17463 18207
rect 17405 18167 17463 18173
rect 8849 18071 8907 18077
rect 8849 18068 8861 18071
rect 8720 18040 8861 18068
rect 8720 18028 8726 18040
rect 8849 18037 8861 18040
rect 8895 18037 8907 18071
rect 8849 18031 8907 18037
rect 9674 18028 9680 18080
rect 9732 18068 9738 18080
rect 10045 18071 10103 18077
rect 10045 18068 10057 18071
rect 9732 18040 10057 18068
rect 9732 18028 9738 18040
rect 10045 18037 10057 18040
rect 10091 18037 10103 18071
rect 10594 18068 10600 18080
rect 10555 18040 10600 18068
rect 10045 18031 10103 18037
rect 10594 18028 10600 18040
rect 10652 18028 10658 18080
rect 10870 18028 10876 18080
rect 10928 18068 10934 18080
rect 11422 18068 11428 18080
rect 10928 18040 11428 18068
rect 10928 18028 10934 18040
rect 11422 18028 11428 18040
rect 11480 18028 11486 18080
rect 15930 18028 15936 18080
rect 15988 18068 15994 18080
rect 16025 18071 16083 18077
rect 16025 18068 16037 18071
rect 15988 18040 16037 18068
rect 15988 18028 15994 18040
rect 16025 18037 16037 18040
rect 16071 18037 16083 18071
rect 16025 18031 16083 18037
rect 1104 17978 20884 18000
rect 1104 17926 8315 17978
rect 8367 17926 8379 17978
rect 8431 17926 8443 17978
rect 8495 17926 8507 17978
rect 8559 17926 15648 17978
rect 15700 17926 15712 17978
rect 15764 17926 15776 17978
rect 15828 17926 15840 17978
rect 15892 17926 20884 17978
rect 1104 17904 20884 17926
rect 2314 17824 2320 17876
rect 2372 17864 2378 17876
rect 2501 17867 2559 17873
rect 2501 17864 2513 17867
rect 2372 17836 2513 17864
rect 2372 17824 2378 17836
rect 2501 17833 2513 17836
rect 2547 17864 2559 17867
rect 3142 17864 3148 17876
rect 2547 17836 3148 17864
rect 2547 17833 2559 17836
rect 2501 17827 2559 17833
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 7558 17864 7564 17876
rect 4217 17836 7564 17864
rect 2682 17796 2688 17808
rect 1596 17768 2688 17796
rect 1596 17740 1624 17768
rect 2682 17756 2688 17768
rect 2740 17756 2746 17808
rect 3970 17756 3976 17808
rect 4028 17796 4034 17808
rect 4217 17796 4245 17836
rect 7558 17824 7564 17836
rect 7616 17824 7622 17876
rect 9490 17824 9496 17876
rect 9548 17864 9554 17876
rect 9769 17867 9827 17873
rect 9769 17864 9781 17867
rect 9548 17836 9781 17864
rect 9548 17824 9554 17836
rect 9769 17833 9781 17836
rect 9815 17833 9827 17867
rect 9769 17827 9827 17833
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 10689 17867 10747 17873
rect 10689 17864 10701 17867
rect 10652 17836 10701 17864
rect 10652 17824 10658 17836
rect 10689 17833 10701 17836
rect 10735 17833 10747 17867
rect 10689 17827 10747 17833
rect 15519 17867 15577 17873
rect 15519 17833 15531 17867
rect 15565 17864 15577 17867
rect 20438 17864 20444 17876
rect 15565 17836 20444 17864
rect 15565 17833 15577 17836
rect 15519 17827 15577 17833
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 9033 17799 9091 17805
rect 9033 17796 9045 17799
rect 4028 17768 4245 17796
rect 5736 17768 9045 17796
rect 4028 17756 4034 17768
rect 5736 17740 5764 17768
rect 9033 17765 9045 17768
rect 9079 17796 9091 17799
rect 9398 17796 9404 17808
rect 9079 17768 9404 17796
rect 9079 17765 9091 17768
rect 9033 17759 9091 17765
rect 9398 17756 9404 17768
rect 9456 17756 9462 17808
rect 16850 17796 16856 17808
rect 12360 17768 16856 17796
rect 12360 17740 12388 17768
rect 16850 17756 16856 17768
rect 16908 17756 16914 17808
rect 1578 17728 1584 17740
rect 1539 17700 1584 17728
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 1854 17728 1860 17740
rect 1815 17700 1860 17728
rect 1854 17688 1860 17700
rect 1912 17688 1918 17740
rect 3028 17731 3086 17737
rect 3028 17697 3040 17731
rect 3074 17728 3086 17731
rect 3074 17700 3556 17728
rect 3074 17697 3086 17700
rect 3028 17691 3086 17697
rect 1762 17620 1768 17672
rect 1820 17660 1826 17672
rect 1949 17663 2007 17669
rect 1949 17660 1961 17663
rect 1820 17632 1961 17660
rect 1820 17620 1826 17632
rect 1949 17629 1961 17632
rect 1995 17629 2007 17663
rect 1949 17623 2007 17629
rect 2958 17552 2964 17604
rect 3016 17592 3022 17604
rect 3099 17595 3157 17601
rect 3099 17592 3111 17595
rect 3016 17564 3111 17592
rect 3016 17552 3022 17564
rect 3099 17561 3111 17564
rect 3145 17561 3157 17595
rect 3099 17555 3157 17561
rect 2774 17524 2780 17536
rect 2735 17496 2780 17524
rect 2774 17484 2780 17496
rect 2832 17484 2838 17536
rect 3528 17533 3556 17700
rect 3878 17688 3884 17740
rect 3936 17728 3942 17740
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 3936 17700 4077 17728
rect 3936 17688 3942 17700
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 4065 17691 4123 17697
rect 4154 17688 4160 17740
rect 4212 17688 4218 17740
rect 5718 17728 5724 17740
rect 5679 17700 5724 17728
rect 5718 17688 5724 17700
rect 5776 17688 5782 17740
rect 6270 17728 6276 17740
rect 6231 17700 6276 17728
rect 6270 17688 6276 17700
rect 6328 17688 6334 17740
rect 8110 17728 8116 17740
rect 8071 17700 8116 17728
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 8570 17728 8576 17740
rect 8531 17700 8576 17728
rect 8570 17688 8576 17700
rect 8628 17688 8634 17740
rect 9950 17728 9956 17740
rect 9911 17700 9956 17728
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 10137 17731 10195 17737
rect 10137 17728 10149 17731
rect 10060 17700 10149 17728
rect 3513 17527 3571 17533
rect 3513 17493 3525 17527
rect 3559 17524 3571 17527
rect 3602 17524 3608 17536
rect 3559 17496 3608 17524
rect 3559 17493 3571 17496
rect 3513 17487 3571 17493
rect 3602 17484 3608 17496
rect 3660 17484 3666 17536
rect 4172 17524 4200 17688
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 4522 17660 4528 17672
rect 4479 17632 4528 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 4522 17620 4528 17632
rect 4580 17620 4586 17672
rect 6454 17660 6460 17672
rect 6415 17632 6460 17660
rect 6454 17620 6460 17632
rect 6512 17620 6518 17672
rect 8754 17660 8760 17672
rect 8715 17632 8760 17660
rect 8754 17620 8760 17632
rect 8812 17620 8818 17672
rect 10060 17604 10088 17700
rect 10137 17697 10149 17700
rect 10183 17697 10195 17731
rect 10137 17691 10195 17697
rect 11241 17731 11299 17737
rect 11241 17697 11253 17731
rect 11287 17728 11299 17731
rect 11330 17728 11336 17740
rect 11287 17700 11336 17728
rect 11287 17697 11299 17700
rect 11241 17691 11299 17697
rect 11330 17688 11336 17700
rect 11388 17688 11394 17740
rect 12342 17737 12348 17740
rect 12320 17731 12348 17737
rect 12320 17728 12332 17731
rect 12255 17700 12332 17728
rect 12320 17697 12332 17700
rect 12320 17691 12348 17697
rect 12342 17688 12348 17691
rect 12400 17688 12406 17740
rect 13332 17731 13390 17737
rect 13332 17697 13344 17731
rect 13378 17728 13390 17731
rect 13446 17728 13452 17740
rect 13378 17700 13452 17728
rect 13378 17697 13390 17700
rect 13332 17691 13390 17697
rect 13446 17688 13452 17700
rect 13504 17688 13510 17740
rect 15286 17688 15292 17740
rect 15344 17728 15350 17740
rect 15416 17731 15474 17737
rect 15416 17728 15428 17731
rect 15344 17700 15428 17728
rect 15344 17688 15350 17700
rect 15416 17697 15428 17700
rect 15462 17697 15474 17731
rect 15416 17691 15474 17697
rect 4230 17595 4288 17601
rect 4230 17561 4242 17595
rect 4276 17592 4288 17595
rect 5166 17592 5172 17604
rect 4276 17564 5172 17592
rect 4276 17561 4288 17564
rect 4230 17555 4288 17561
rect 5166 17552 5172 17564
rect 5224 17552 5230 17604
rect 7285 17595 7343 17601
rect 7285 17561 7297 17595
rect 7331 17592 7343 17595
rect 7558 17592 7564 17604
rect 7331 17564 7564 17592
rect 7331 17561 7343 17564
rect 7285 17555 7343 17561
rect 7558 17552 7564 17564
rect 7616 17592 7622 17604
rect 10042 17592 10048 17604
rect 7616 17564 10048 17592
rect 7616 17552 7622 17564
rect 10042 17552 10048 17564
rect 10100 17552 10106 17604
rect 10134 17552 10140 17604
rect 10192 17592 10198 17604
rect 12391 17595 12449 17601
rect 12391 17592 12403 17595
rect 10192 17564 12403 17592
rect 10192 17552 10198 17564
rect 12391 17561 12403 17564
rect 12437 17561 12449 17595
rect 12391 17555 12449 17561
rect 4341 17527 4399 17533
rect 4341 17524 4353 17527
rect 4172 17496 4353 17524
rect 4341 17493 4353 17496
rect 4387 17493 4399 17527
rect 4341 17487 4399 17493
rect 4430 17484 4436 17536
rect 4488 17524 4494 17536
rect 4525 17527 4583 17533
rect 4525 17524 4537 17527
rect 4488 17496 4537 17524
rect 4488 17484 4494 17496
rect 4525 17493 4537 17496
rect 4571 17493 4583 17527
rect 5074 17524 5080 17536
rect 4987 17496 5080 17524
rect 4525 17487 4583 17493
rect 5074 17484 5080 17496
rect 5132 17524 5138 17536
rect 6178 17524 6184 17536
rect 5132 17496 6184 17524
rect 5132 17484 5138 17496
rect 6178 17484 6184 17496
rect 6236 17484 6242 17536
rect 6822 17524 6828 17536
rect 6783 17496 6828 17524
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 7653 17527 7711 17533
rect 7653 17524 7665 17527
rect 7432 17496 7665 17524
rect 7432 17484 7438 17496
rect 7653 17493 7665 17496
rect 7699 17493 7711 17527
rect 7653 17487 7711 17493
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 11379 17527 11437 17533
rect 11379 17524 11391 17527
rect 11020 17496 11391 17524
rect 11020 17484 11026 17496
rect 11379 17493 11391 17496
rect 11425 17493 11437 17527
rect 11379 17487 11437 17493
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 13403 17527 13461 17533
rect 13403 17524 13415 17527
rect 12584 17496 13415 17524
rect 12584 17484 12590 17496
rect 13403 17493 13415 17496
rect 13449 17493 13461 17527
rect 13403 17487 13461 17493
rect 1104 17434 20884 17456
rect 1104 17382 4648 17434
rect 4700 17382 4712 17434
rect 4764 17382 4776 17434
rect 4828 17382 4840 17434
rect 4892 17382 11982 17434
rect 12034 17382 12046 17434
rect 12098 17382 12110 17434
rect 12162 17382 12174 17434
rect 12226 17382 19315 17434
rect 19367 17382 19379 17434
rect 19431 17382 19443 17434
rect 19495 17382 19507 17434
rect 19559 17382 20884 17434
rect 1104 17360 20884 17382
rect 1673 17323 1731 17329
rect 1673 17289 1685 17323
rect 1719 17320 1731 17323
rect 1854 17320 1860 17332
rect 1719 17292 1860 17320
rect 1719 17289 1731 17292
rect 1673 17283 1731 17289
rect 1854 17280 1860 17292
rect 1912 17280 1918 17332
rect 5859 17323 5917 17329
rect 5859 17320 5871 17323
rect 1958 17292 5871 17320
rect 14 17212 20 17264
rect 72 17252 78 17264
rect 1958 17252 1986 17292
rect 5859 17289 5871 17292
rect 5905 17289 5917 17323
rect 6270 17320 6276 17332
rect 6231 17292 6276 17320
rect 5859 17283 5917 17289
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 6638 17280 6644 17332
rect 6696 17320 6702 17332
rect 12253 17323 12311 17329
rect 12253 17320 12265 17323
rect 6696 17292 12265 17320
rect 6696 17280 6702 17292
rect 12253 17289 12265 17292
rect 12299 17320 12311 17323
rect 12342 17320 12348 17332
rect 12299 17292 12348 17320
rect 12299 17289 12311 17292
rect 12253 17283 12311 17289
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 13446 17320 13452 17332
rect 13407 17292 13452 17320
rect 13446 17280 13452 17292
rect 13504 17320 13510 17332
rect 15930 17320 15936 17332
rect 13504 17292 15936 17320
rect 13504 17280 13510 17292
rect 15930 17280 15936 17292
rect 15988 17280 15994 17332
rect 72 17224 1986 17252
rect 3697 17255 3755 17261
rect 72 17212 78 17224
rect 3697 17221 3709 17255
rect 3743 17252 3755 17255
rect 4338 17252 4344 17264
rect 3743 17224 4344 17252
rect 3743 17221 3755 17224
rect 3697 17215 3755 17221
rect 4338 17212 4344 17224
rect 4396 17212 4402 17264
rect 5629 17255 5687 17261
rect 5629 17221 5641 17255
rect 5675 17252 5687 17255
rect 5675 17224 7604 17252
rect 5675 17221 5687 17224
rect 5629 17215 5687 17221
rect 3878 17144 3884 17196
rect 3936 17184 3942 17196
rect 4801 17187 4859 17193
rect 4801 17184 4813 17187
rect 3936 17156 4813 17184
rect 3936 17144 3942 17156
rect 4801 17153 4813 17156
rect 4847 17153 4859 17187
rect 4801 17147 4859 17153
rect 2961 17119 3019 17125
rect 2961 17085 2973 17119
rect 3007 17116 3019 17119
rect 3602 17116 3608 17128
rect 3007 17088 3608 17116
rect 3007 17085 3019 17088
rect 2961 17079 3019 17085
rect 3602 17076 3608 17088
rect 3660 17076 3666 17128
rect 3970 17116 3976 17128
rect 3931 17088 3976 17116
rect 3970 17076 3976 17088
rect 4028 17076 4034 17128
rect 4338 17116 4344 17128
rect 4299 17088 4344 17116
rect 4338 17076 4344 17088
rect 4396 17076 4402 17128
rect 5803 17125 5831 17224
rect 6914 17184 6920 17196
rect 6875 17156 6920 17184
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 5788 17119 5846 17125
rect 5788 17085 5800 17119
rect 5834 17085 5846 17119
rect 5788 17079 5846 17085
rect 2317 17051 2375 17057
rect 2317 17017 2329 17051
rect 2363 17017 2375 17051
rect 2317 17011 2375 17017
rect 2409 17051 2467 17057
rect 2409 17017 2421 17051
rect 2455 17048 2467 17051
rect 2774 17048 2780 17060
rect 2455 17020 2780 17048
rect 2455 17017 2467 17020
rect 2409 17011 2467 17017
rect 1578 16940 1584 16992
rect 1636 16980 1642 16992
rect 1854 16980 1860 16992
rect 1636 16952 1860 16980
rect 1636 16940 1642 16952
rect 1854 16940 1860 16952
rect 1912 16980 1918 16992
rect 1949 16983 2007 16989
rect 1949 16980 1961 16983
rect 1912 16952 1961 16980
rect 1912 16940 1918 16952
rect 1949 16949 1961 16952
rect 1995 16949 2007 16983
rect 2332 16980 2360 17011
rect 2774 17008 2780 17020
rect 2832 17008 2838 17060
rect 3329 17051 3387 17057
rect 3329 17017 3341 17051
rect 3375 17048 3387 17051
rect 4430 17048 4436 17060
rect 3375 17020 4436 17048
rect 3375 17017 3387 17020
rect 3329 17011 3387 17017
rect 4430 17008 4436 17020
rect 4488 17008 4494 17060
rect 6270 17008 6276 17060
rect 6328 17048 6334 17060
rect 7009 17051 7067 17057
rect 7009 17048 7021 17051
rect 6328 17020 7021 17048
rect 6328 17008 6334 17020
rect 7009 17017 7021 17020
rect 7055 17048 7067 17051
rect 7374 17048 7380 17060
rect 7055 17020 7380 17048
rect 7055 17017 7067 17020
rect 7009 17011 7067 17017
rect 7374 17008 7380 17020
rect 7432 17008 7438 17060
rect 7576 17057 7604 17224
rect 9398 17212 9404 17264
rect 9456 17252 9462 17264
rect 9456 17224 10891 17252
rect 9456 17212 9462 17224
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 10229 17187 10287 17193
rect 7708 17156 9076 17184
rect 7708 17144 7714 17156
rect 9048 17128 9076 17156
rect 10229 17153 10241 17187
rect 10275 17184 10287 17187
rect 10594 17184 10600 17196
rect 10275 17156 10600 17184
rect 10275 17153 10287 17156
rect 10229 17147 10287 17153
rect 10594 17144 10600 17156
rect 10652 17144 10658 17196
rect 10863 17184 10891 17224
rect 14277 17187 14335 17193
rect 10863 17156 12480 17184
rect 8481 17119 8539 17125
rect 8481 17085 8493 17119
rect 8527 17116 8539 17119
rect 8570 17116 8576 17128
rect 8527 17088 8576 17116
rect 8527 17085 8539 17088
rect 8481 17079 8539 17085
rect 8570 17076 8576 17088
rect 8628 17116 8634 17128
rect 8849 17119 8907 17125
rect 8849 17116 8861 17119
rect 8628 17088 8861 17116
rect 8628 17076 8634 17088
rect 8849 17085 8861 17088
rect 8895 17085 8907 17119
rect 9030 17116 9036 17128
rect 8991 17088 9036 17116
rect 8849 17079 8907 17085
rect 7561 17051 7619 17057
rect 7561 17017 7573 17051
rect 7607 17048 7619 17051
rect 7926 17048 7932 17060
rect 7607 17020 7932 17048
rect 7607 17017 7619 17020
rect 7561 17011 7619 17017
rect 7926 17008 7932 17020
rect 7984 17008 7990 17060
rect 2866 16980 2872 16992
rect 2332 16952 2872 16980
rect 1949 16943 2007 16949
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 3878 16980 3884 16992
rect 3839 16952 3884 16980
rect 3878 16940 3884 16952
rect 3936 16940 3942 16992
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 5261 16983 5319 16989
rect 5261 16980 5273 16983
rect 4212 16952 5273 16980
rect 4212 16940 4218 16952
rect 5261 16949 5273 16952
rect 5307 16980 5319 16983
rect 5350 16980 5356 16992
rect 5307 16952 5356 16980
rect 5307 16949 5319 16952
rect 5261 16943 5319 16949
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 5718 16940 5724 16992
rect 5776 16980 5782 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 5776 16952 6561 16980
rect 5776 16940 5782 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 8110 16980 8116 16992
rect 8071 16952 8116 16980
rect 6549 16943 6607 16949
rect 8110 16940 8116 16952
rect 8168 16940 8174 16992
rect 8864 16980 8892 17079
rect 9030 17076 9036 17088
rect 9088 17076 9094 17128
rect 12452 17125 12480 17156
rect 14277 17153 14289 17187
rect 14323 17184 14335 17187
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14323 17156 14473 17184
rect 14323 17153 14335 17156
rect 14277 17147 14335 17153
rect 14461 17153 14473 17156
rect 14507 17184 14519 17187
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 14507 17156 15945 17184
rect 14507 17153 14519 17156
rect 14461 17147 14519 17153
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 12437 17119 12495 17125
rect 12437 17085 12449 17119
rect 12483 17116 12495 17119
rect 12618 17116 12624 17128
rect 12483 17088 12624 17116
rect 12483 17085 12495 17088
rect 12437 17079 12495 17085
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 12897 17119 12955 17125
rect 12897 17085 12909 17119
rect 12943 17085 12955 17119
rect 12897 17079 12955 17085
rect 9306 17048 9312 17060
rect 9267 17020 9312 17048
rect 9306 17008 9312 17020
rect 9364 17008 9370 17060
rect 10321 17051 10379 17057
rect 10321 17017 10333 17051
rect 10367 17048 10379 17051
rect 10594 17048 10600 17060
rect 10367 17020 10600 17048
rect 10367 17017 10379 17020
rect 10321 17011 10379 17017
rect 10594 17008 10600 17020
rect 10652 17008 10658 17060
rect 10870 17048 10876 17060
rect 10831 17020 10876 17048
rect 10870 17008 10876 17020
rect 10928 17008 10934 17060
rect 12912 17048 12940 17079
rect 11808 17020 12940 17048
rect 13173 17051 13231 17057
rect 9769 16983 9827 16989
rect 9769 16980 9781 16983
rect 8864 16952 9781 16980
rect 9769 16949 9781 16952
rect 9815 16980 9827 16983
rect 9950 16980 9956 16992
rect 9815 16952 9956 16980
rect 9815 16949 9827 16952
rect 9769 16943 9827 16949
rect 9950 16940 9956 16952
rect 10008 16980 10014 16992
rect 10502 16980 10508 16992
rect 10008 16952 10508 16980
rect 10008 16940 10014 16952
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 11330 16980 11336 16992
rect 11291 16952 11336 16980
rect 11330 16940 11336 16952
rect 11388 16940 11394 16992
rect 11514 16940 11520 16992
rect 11572 16980 11578 16992
rect 11808 16989 11836 17020
rect 13173 17017 13185 17051
rect 13219 17048 13231 17051
rect 13446 17048 13452 17060
rect 13219 17020 13452 17048
rect 13219 17017 13231 17020
rect 13173 17011 13231 17017
rect 13446 17008 13452 17020
rect 13504 17008 13510 17060
rect 14550 17008 14556 17060
rect 14608 17048 14614 17060
rect 15105 17051 15163 17057
rect 14608 17020 14653 17048
rect 14608 17008 14614 17020
rect 15105 17017 15117 17051
rect 15151 17017 15163 17051
rect 15105 17011 15163 17017
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 11572 16952 11805 16980
rect 11572 16940 11578 16952
rect 11793 16949 11805 16952
rect 11839 16949 11851 16983
rect 15120 16980 15148 17011
rect 15286 16980 15292 16992
rect 15120 16952 15292 16980
rect 11793 16943 11851 16949
rect 15286 16940 15292 16952
rect 15344 16980 15350 16992
rect 15381 16983 15439 16989
rect 15381 16980 15393 16983
rect 15344 16952 15393 16980
rect 15344 16940 15350 16952
rect 15381 16949 15393 16952
rect 15427 16949 15439 16983
rect 15381 16943 15439 16949
rect 1104 16890 20884 16912
rect 1104 16838 8315 16890
rect 8367 16838 8379 16890
rect 8431 16838 8443 16890
rect 8495 16838 8507 16890
rect 8559 16838 15648 16890
rect 15700 16838 15712 16890
rect 15764 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 20884 16890
rect 1104 16816 20884 16838
rect 1946 16776 1952 16788
rect 1907 16748 1952 16776
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 2501 16779 2559 16785
rect 2501 16745 2513 16779
rect 2547 16776 2559 16779
rect 2774 16776 2780 16788
rect 2547 16748 2780 16776
rect 2547 16745 2559 16748
rect 2501 16739 2559 16745
rect 2774 16736 2780 16748
rect 2832 16736 2838 16788
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 4062 16776 4068 16788
rect 2924 16748 4068 16776
rect 2924 16736 2930 16748
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 6181 16779 6239 16785
rect 6181 16745 6193 16779
rect 6227 16776 6239 16779
rect 6270 16776 6276 16788
rect 6227 16748 6276 16776
rect 6227 16745 6239 16748
rect 6181 16739 6239 16745
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 6914 16776 6920 16788
rect 6875 16748 6920 16776
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 8389 16779 8447 16785
rect 8389 16745 8401 16779
rect 8435 16776 8447 16779
rect 8662 16776 8668 16788
rect 8435 16748 8668 16776
rect 8435 16745 8447 16748
rect 8389 16739 8447 16745
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10045 16779 10103 16785
rect 10045 16776 10057 16779
rect 10008 16748 10057 16776
rect 10008 16736 10014 16748
rect 10045 16745 10057 16748
rect 10091 16745 10103 16779
rect 10594 16776 10600 16788
rect 10555 16748 10600 16776
rect 10045 16739 10103 16745
rect 10594 16736 10600 16748
rect 10652 16776 10658 16788
rect 10873 16779 10931 16785
rect 10873 16776 10885 16779
rect 10652 16748 10885 16776
rect 10652 16736 10658 16748
rect 10873 16745 10885 16748
rect 10919 16745 10931 16779
rect 12618 16776 12624 16788
rect 12579 16748 12624 16776
rect 10873 16739 10931 16745
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 14093 16779 14151 16785
rect 14093 16745 14105 16779
rect 14139 16776 14151 16779
rect 14461 16779 14519 16785
rect 14461 16776 14473 16779
rect 14139 16748 14473 16776
rect 14139 16745 14151 16748
rect 14093 16739 14151 16745
rect 14461 16745 14473 16748
rect 14507 16776 14519 16779
rect 14550 16776 14556 16788
rect 14507 16748 14556 16776
rect 14507 16745 14519 16748
rect 14461 16739 14519 16745
rect 14550 16736 14556 16748
rect 14608 16736 14614 16788
rect 19242 16776 19248 16788
rect 19203 16748 19248 16776
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 5623 16711 5681 16717
rect 5623 16677 5635 16711
rect 5669 16708 5681 16711
rect 5718 16708 5724 16720
rect 5669 16680 5724 16708
rect 5669 16677 5681 16680
rect 5623 16671 5681 16677
rect 5718 16668 5724 16680
rect 5776 16668 5782 16720
rect 7466 16708 7472 16720
rect 7427 16680 7472 16708
rect 7466 16668 7472 16680
rect 7524 16668 7530 16720
rect 7650 16668 7656 16720
rect 7708 16708 7714 16720
rect 8110 16708 8116 16720
rect 7708 16680 8116 16708
rect 7708 16668 7714 16680
rect 8110 16668 8116 16680
rect 8168 16708 8174 16720
rect 8168 16680 11836 16708
rect 8168 16668 8174 16680
rect 11808 16652 11836 16680
rect 13262 16668 13268 16720
rect 13320 16708 13326 16720
rect 13494 16711 13552 16717
rect 13494 16708 13506 16711
rect 13320 16680 13506 16708
rect 13320 16668 13326 16680
rect 13494 16677 13506 16680
rect 13540 16677 13552 16711
rect 13494 16671 13552 16677
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16640 1639 16643
rect 2130 16640 2136 16652
rect 1627 16612 2136 16640
rect 1627 16609 1639 16612
rect 1581 16603 1639 16609
rect 2130 16600 2136 16612
rect 2188 16640 2194 16652
rect 3050 16640 3056 16652
rect 2188 16612 3056 16640
rect 2188 16600 2194 16612
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 5258 16640 5264 16652
rect 5219 16612 5264 16640
rect 5258 16600 5264 16612
rect 5316 16600 5322 16652
rect 8754 16600 8760 16652
rect 8812 16640 8818 16652
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 8812 16612 9689 16640
rect 8812 16600 8818 16612
rect 9677 16609 9689 16612
rect 9723 16640 9735 16643
rect 11238 16640 11244 16652
rect 9723 16612 11244 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 11790 16640 11796 16652
rect 11751 16612 11796 16640
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16609 12127 16643
rect 14918 16640 14924 16652
rect 12069 16603 12127 16609
rect 12268 16612 14924 16640
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16572 4215 16575
rect 4246 16572 4252 16584
rect 4203 16544 4252 16572
rect 4203 16541 4215 16544
rect 4157 16535 4215 16541
rect 4246 16532 4252 16544
rect 4304 16572 4310 16584
rect 5442 16572 5448 16584
rect 4304 16544 5448 16572
rect 4304 16532 4310 16544
rect 5442 16532 5448 16544
rect 5500 16572 5506 16584
rect 6638 16572 6644 16584
rect 5500 16544 6644 16572
rect 5500 16532 5506 16544
rect 6638 16532 6644 16544
rect 6696 16532 6702 16584
rect 7377 16575 7435 16581
rect 7377 16541 7389 16575
rect 7423 16572 7435 16575
rect 8018 16572 8024 16584
rect 7423 16544 8024 16572
rect 7423 16541 7435 16544
rect 7377 16535 7435 16541
rect 8018 16532 8024 16544
rect 8076 16572 8082 16584
rect 8386 16572 8392 16584
rect 8076 16544 8392 16572
rect 8076 16532 8082 16544
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 11514 16532 11520 16584
rect 11572 16572 11578 16584
rect 12084 16572 12112 16603
rect 11572 16544 12112 16572
rect 11572 16532 11578 16544
rect 3050 16464 3056 16516
rect 3108 16504 3114 16516
rect 3789 16507 3847 16513
rect 3789 16504 3801 16507
rect 3108 16476 3801 16504
rect 3108 16464 3114 16476
rect 3789 16473 3801 16476
rect 3835 16504 3847 16507
rect 3970 16504 3976 16516
rect 3835 16476 3976 16504
rect 3835 16473 3847 16476
rect 3789 16467 3847 16473
rect 3970 16464 3976 16476
rect 4028 16464 4034 16516
rect 4387 16507 4445 16513
rect 4387 16473 4399 16507
rect 4433 16504 4445 16507
rect 4522 16504 4528 16516
rect 4433 16476 4528 16504
rect 4433 16473 4445 16476
rect 4387 16467 4445 16473
rect 4522 16464 4528 16476
rect 4580 16504 4586 16516
rect 5077 16507 5135 16513
rect 5077 16504 5089 16507
rect 4580 16476 5089 16504
rect 4580 16464 4586 16476
rect 5077 16473 5089 16476
rect 5123 16473 5135 16507
rect 7926 16504 7932 16516
rect 7887 16476 7932 16504
rect 5077 16467 5135 16473
rect 7926 16464 7932 16476
rect 7984 16464 7990 16516
rect 9493 16507 9551 16513
rect 9493 16473 9505 16507
rect 9539 16504 9551 16507
rect 10042 16504 10048 16516
rect 9539 16476 10048 16504
rect 9539 16473 9551 16476
rect 9493 16467 9551 16473
rect 10042 16464 10048 16476
rect 10100 16504 10106 16516
rect 12268 16504 12296 16612
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 15356 16643 15414 16649
rect 15356 16609 15368 16643
rect 15402 16640 15414 16643
rect 16114 16640 16120 16652
rect 15402 16612 16120 16640
rect 15402 16609 15414 16612
rect 15356 16603 15414 16609
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 19058 16640 19064 16652
rect 19019 16612 19064 16640
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16572 12403 16575
rect 13170 16572 13176 16584
rect 12391 16544 13176 16572
rect 12391 16541 12403 16544
rect 12345 16535 12403 16541
rect 13170 16532 13176 16544
rect 13228 16532 13234 16584
rect 10100 16476 12296 16504
rect 10100 16464 10106 16476
rect 12434 16464 12440 16516
rect 12492 16504 12498 16516
rect 15427 16507 15485 16513
rect 15427 16504 15439 16507
rect 12492 16476 15439 16504
rect 12492 16464 12498 16476
rect 15427 16473 15439 16476
rect 15473 16473 15485 16507
rect 15427 16467 15485 16473
rect 2958 16396 2964 16448
rect 3016 16436 3022 16448
rect 3145 16439 3203 16445
rect 3145 16436 3157 16439
rect 3016 16408 3157 16436
rect 3016 16396 3022 16408
rect 3145 16405 3157 16408
rect 3191 16405 3203 16439
rect 3145 16399 3203 16405
rect 4801 16439 4859 16445
rect 4801 16405 4813 16439
rect 4847 16436 4859 16439
rect 5166 16436 5172 16448
rect 4847 16408 5172 16436
rect 4847 16405 4859 16408
rect 4801 16399 4859 16405
rect 5166 16396 5172 16408
rect 5224 16396 5230 16448
rect 8662 16436 8668 16448
rect 8623 16408 8668 16436
rect 8662 16396 8668 16408
rect 8720 16436 8726 16448
rect 9030 16436 9036 16448
rect 8720 16408 9036 16436
rect 8720 16396 8726 16408
rect 9030 16396 9036 16408
rect 9088 16396 9094 16448
rect 12618 16396 12624 16448
rect 12676 16436 12682 16448
rect 16666 16436 16672 16448
rect 12676 16408 16672 16436
rect 12676 16396 12682 16408
rect 16666 16396 16672 16408
rect 16724 16396 16730 16448
rect 1104 16346 20884 16368
rect 1104 16294 4648 16346
rect 4700 16294 4712 16346
rect 4764 16294 4776 16346
rect 4828 16294 4840 16346
rect 4892 16294 11982 16346
rect 12034 16294 12046 16346
rect 12098 16294 12110 16346
rect 12162 16294 12174 16346
rect 12226 16294 19315 16346
rect 19367 16294 19379 16346
rect 19431 16294 19443 16346
rect 19495 16294 19507 16346
rect 19559 16294 20884 16346
rect 1104 16272 20884 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 1946 16192 1952 16244
rect 2004 16232 2010 16244
rect 2317 16235 2375 16241
rect 2317 16232 2329 16235
rect 2004 16204 2329 16232
rect 2004 16192 2010 16204
rect 2317 16201 2329 16204
rect 2363 16201 2375 16235
rect 4246 16232 4252 16244
rect 4207 16204 4252 16232
rect 2317 16195 2375 16201
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 6273 16235 6331 16241
rect 6273 16201 6285 16235
rect 6319 16232 6331 16235
rect 6362 16232 6368 16244
rect 6319 16204 6368 16232
rect 6319 16201 6331 16204
rect 6273 16195 6331 16201
rect 6362 16192 6368 16204
rect 6420 16192 6426 16244
rect 7466 16192 7472 16244
rect 7524 16232 7530 16244
rect 7745 16235 7803 16241
rect 7745 16232 7757 16235
rect 7524 16204 7757 16232
rect 7524 16192 7530 16204
rect 7745 16201 7757 16204
rect 7791 16232 7803 16235
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 7791 16204 8033 16232
rect 7791 16201 7803 16204
rect 7745 16195 7803 16201
rect 8021 16201 8033 16204
rect 8067 16201 8079 16235
rect 8386 16232 8392 16244
rect 8347 16204 8392 16232
rect 8021 16195 8079 16201
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 8757 16235 8815 16241
rect 8757 16201 8769 16235
rect 8803 16232 8815 16235
rect 9858 16232 9864 16244
rect 8803 16204 9864 16232
rect 8803 16201 8815 16204
rect 8757 16195 8815 16201
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 11238 16232 11244 16244
rect 11199 16204 11244 16232
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 11790 16192 11796 16244
rect 11848 16232 11854 16244
rect 12069 16235 12127 16241
rect 12069 16232 12081 16235
rect 11848 16204 12081 16232
rect 11848 16192 11854 16204
rect 12069 16201 12081 16204
rect 12115 16232 12127 16235
rect 16482 16232 16488 16244
rect 12115 16204 16488 16232
rect 12115 16201 12127 16204
rect 12069 16195 12127 16201
rect 16482 16192 16488 16204
rect 16540 16192 16546 16244
rect 4430 16124 4436 16176
rect 4488 16164 4494 16176
rect 4614 16164 4620 16176
rect 4488 16136 4620 16164
rect 4488 16124 4494 16136
rect 4614 16124 4620 16136
rect 4672 16124 4678 16176
rect 4522 16056 4528 16108
rect 4580 16096 4586 16108
rect 4709 16099 4767 16105
rect 4709 16096 4721 16099
rect 4580 16068 4721 16096
rect 4580 16056 4586 16068
rect 4709 16065 4721 16068
rect 4755 16065 4767 16099
rect 6380 16096 6408 16192
rect 10410 16124 10416 16176
rect 10468 16164 10474 16176
rect 16255 16167 16313 16173
rect 16255 16164 16267 16167
rect 10468 16136 16267 16164
rect 10468 16124 10474 16136
rect 16255 16133 16267 16136
rect 16301 16133 16313 16167
rect 16255 16127 16313 16133
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 6380 16068 6837 16096
rect 4709 16059 4767 16065
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 9677 16099 9735 16105
rect 9677 16065 9689 16099
rect 9723 16096 9735 16099
rect 9766 16096 9772 16108
rect 9723 16068 9772 16096
rect 9723 16065 9735 16068
rect 9677 16059 9735 16065
rect 9766 16056 9772 16068
rect 9824 16096 9830 16108
rect 10873 16099 10931 16105
rect 10873 16096 10885 16099
rect 9824 16068 10885 16096
rect 9824 16056 9830 16068
rect 10873 16065 10885 16068
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 13630 16056 13636 16108
rect 13688 16096 13694 16108
rect 13688 16068 16195 16096
rect 13688 16056 13694 16068
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1443 16000 2084 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 2056 15904 2084 16000
rect 3602 15988 3608 16040
rect 3660 16028 3666 16040
rect 4430 16028 4436 16040
rect 3660 16000 4436 16028
rect 3660 15988 3666 16000
rect 4430 15988 4436 16000
rect 4488 15988 4494 16040
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 13354 16028 13360 16040
rect 8619 16000 9260 16028
rect 13315 16000 13360 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 2958 15960 2964 15972
rect 2919 15932 2964 15960
rect 2958 15920 2964 15932
rect 3016 15920 3022 15972
rect 3053 15963 3111 15969
rect 3053 15929 3065 15963
rect 3099 15929 3111 15963
rect 3053 15923 3111 15929
rect 3973 15963 4031 15969
rect 3973 15929 3985 15963
rect 4019 15960 4031 15963
rect 4801 15963 4859 15969
rect 4801 15960 4813 15963
rect 4019 15932 4813 15960
rect 4019 15929 4031 15932
rect 3973 15923 4031 15929
rect 4801 15929 4813 15932
rect 4847 15960 4859 15963
rect 5074 15960 5080 15972
rect 4847 15932 5080 15960
rect 4847 15929 4859 15932
rect 4801 15923 4859 15929
rect 2038 15892 2044 15904
rect 1999 15864 2044 15892
rect 2038 15852 2044 15864
rect 2096 15852 2102 15904
rect 2777 15895 2835 15901
rect 2777 15861 2789 15895
rect 2823 15892 2835 15895
rect 3068 15892 3096 15923
rect 5074 15920 5080 15932
rect 5132 15920 5138 15972
rect 5350 15960 5356 15972
rect 5311 15932 5356 15960
rect 5350 15920 5356 15932
rect 5408 15920 5414 15972
rect 9232 15969 9260 16000
rect 13354 15988 13360 16000
rect 13412 16028 13418 16040
rect 16167 16037 16195 16068
rect 14553 16031 14611 16037
rect 14553 16028 14565 16031
rect 13412 16000 14565 16028
rect 13412 15988 13418 16000
rect 14553 15997 14565 16000
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 15172 16031 15230 16037
rect 15172 15997 15184 16031
rect 15218 16028 15230 16031
rect 16152 16031 16210 16037
rect 15218 16000 15700 16028
rect 15218 15997 15230 16000
rect 15172 15991 15230 15997
rect 7146 15963 7204 15969
rect 7146 15960 7158 15963
rect 6656 15932 7158 15960
rect 6656 15904 6684 15932
rect 7146 15929 7158 15932
rect 7192 15960 7204 15963
rect 9217 15963 9275 15969
rect 7192 15932 9168 15960
rect 7192 15929 7204 15932
rect 7146 15923 7204 15929
rect 3142 15892 3148 15904
rect 2823 15864 3148 15892
rect 2823 15861 2835 15864
rect 2777 15855 2835 15861
rect 3142 15852 3148 15864
rect 3200 15852 3206 15904
rect 5718 15892 5724 15904
rect 5631 15864 5724 15892
rect 5718 15852 5724 15864
rect 5776 15892 5782 15904
rect 6638 15892 6644 15904
rect 5776 15864 6644 15892
rect 5776 15852 5782 15864
rect 6638 15852 6644 15864
rect 6696 15852 6702 15904
rect 9140 15892 9168 15932
rect 9217 15929 9229 15963
rect 9263 15960 9275 15963
rect 9582 15960 9588 15972
rect 9263 15932 9588 15960
rect 9263 15929 9275 15932
rect 9217 15923 9275 15929
rect 9582 15920 9588 15932
rect 9640 15920 9646 15972
rect 9998 15963 10056 15969
rect 9998 15960 10010 15963
rect 9876 15932 10010 15960
rect 9876 15904 9904 15932
rect 9998 15929 10010 15932
rect 10044 15960 10056 15963
rect 12805 15963 12863 15969
rect 12805 15960 12817 15963
rect 10044 15932 12817 15960
rect 10044 15929 10056 15932
rect 9998 15923 10056 15929
rect 12805 15929 12817 15932
rect 12851 15960 12863 15963
rect 13173 15963 13231 15969
rect 13173 15960 13185 15963
rect 12851 15932 13185 15960
rect 12851 15929 12863 15932
rect 12805 15923 12863 15929
rect 13173 15929 13185 15932
rect 13219 15960 13231 15963
rect 13262 15960 13268 15972
rect 13219 15932 13268 15960
rect 13219 15929 13231 15932
rect 13173 15923 13231 15929
rect 13262 15920 13268 15932
rect 13320 15960 13326 15972
rect 13678 15963 13736 15969
rect 13678 15960 13690 15963
rect 13320 15932 13690 15960
rect 13320 15920 13326 15932
rect 13678 15929 13690 15932
rect 13724 15929 13736 15963
rect 13678 15923 13736 15929
rect 9493 15895 9551 15901
rect 9493 15892 9505 15895
rect 9140 15864 9505 15892
rect 9493 15861 9505 15864
rect 9539 15892 9551 15895
rect 9858 15892 9864 15904
rect 9539 15864 9864 15892
rect 9539 15861 9551 15864
rect 9493 15855 9551 15861
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 10594 15892 10600 15904
rect 10555 15864 10600 15892
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 11609 15895 11667 15901
rect 11609 15892 11621 15895
rect 11572 15864 11621 15892
rect 11572 15852 11578 15864
rect 11609 15861 11621 15864
rect 11655 15861 11667 15895
rect 14274 15892 14280 15904
rect 14235 15864 14280 15892
rect 11609 15855 11667 15861
rect 14274 15852 14280 15864
rect 14332 15852 14338 15904
rect 14458 15852 14464 15904
rect 14516 15892 14522 15904
rect 15672 15901 15700 16000
rect 16152 15997 16164 16031
rect 16198 16028 16210 16031
rect 16577 16031 16635 16037
rect 16577 16028 16589 16031
rect 16198 16000 16589 16028
rect 16198 15997 16210 16000
rect 16152 15991 16210 15997
rect 16577 15997 16589 16000
rect 16623 15997 16635 16031
rect 16577 15991 16635 15997
rect 15243 15895 15301 15901
rect 15243 15892 15255 15895
rect 14516 15864 15255 15892
rect 14516 15852 14522 15864
rect 15243 15861 15255 15864
rect 15289 15861 15301 15895
rect 15243 15855 15301 15861
rect 15657 15895 15715 15901
rect 15657 15861 15669 15895
rect 15703 15892 15715 15895
rect 15930 15892 15936 15904
rect 15703 15864 15936 15892
rect 15703 15861 15715 15864
rect 15657 15855 15715 15861
rect 15930 15852 15936 15864
rect 15988 15852 15994 15904
rect 16025 15895 16083 15901
rect 16025 15861 16037 15895
rect 16071 15892 16083 15895
rect 16114 15892 16120 15904
rect 16071 15864 16120 15892
rect 16071 15861 16083 15864
rect 16025 15855 16083 15861
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 19058 15892 19064 15904
rect 19019 15864 19064 15892
rect 19058 15852 19064 15864
rect 19116 15852 19122 15904
rect 1104 15802 20884 15824
rect 1104 15750 8315 15802
rect 8367 15750 8379 15802
rect 8431 15750 8443 15802
rect 8495 15750 8507 15802
rect 8559 15750 15648 15802
rect 15700 15750 15712 15802
rect 15764 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 20884 15802
rect 1104 15728 20884 15750
rect 1670 15688 1676 15700
rect 1631 15660 1676 15688
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 2130 15688 2136 15700
rect 2091 15660 2136 15688
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 3142 15688 3148 15700
rect 3103 15660 3148 15688
rect 3142 15648 3148 15660
rect 3200 15648 3206 15700
rect 5258 15688 5264 15700
rect 5219 15660 5264 15688
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 6454 15688 6460 15700
rect 6415 15660 6460 15688
rect 6454 15648 6460 15660
rect 6512 15688 6518 15700
rect 9858 15688 9864 15700
rect 6512 15660 6592 15688
rect 9819 15660 9864 15688
rect 6512 15648 6518 15660
rect 1946 15580 1952 15632
rect 2004 15620 2010 15632
rect 2546 15623 2604 15629
rect 2546 15620 2558 15623
rect 2004 15592 2558 15620
rect 2004 15580 2010 15592
rect 2546 15589 2558 15592
rect 2592 15589 2604 15623
rect 4246 15620 4252 15632
rect 4207 15592 4252 15620
rect 2546 15583 2604 15589
rect 4246 15580 4252 15592
rect 4304 15580 4310 15632
rect 2222 15552 2228 15564
rect 2183 15524 2228 15552
rect 2222 15512 2228 15524
rect 2280 15512 2286 15564
rect 6564 15561 6592 15660
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 10965 15691 11023 15697
rect 10965 15657 10977 15691
rect 11011 15688 11023 15691
rect 11790 15688 11796 15700
rect 11011 15660 11796 15688
rect 11011 15657 11023 15660
rect 10965 15651 11023 15657
rect 11790 15648 11796 15660
rect 11848 15688 11854 15700
rect 13170 15688 13176 15700
rect 11848 15660 12020 15688
rect 13131 15660 13176 15688
rect 11848 15648 11854 15660
rect 6638 15580 6644 15632
rect 6696 15620 6702 15632
rect 6870 15623 6928 15629
rect 6870 15620 6882 15623
rect 6696 15592 6882 15620
rect 6696 15580 6702 15592
rect 6870 15589 6882 15592
rect 6916 15589 6928 15623
rect 9876 15620 9904 15648
rect 11992 15629 12020 15660
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 14369 15691 14427 15697
rect 14369 15657 14381 15691
rect 14415 15688 14427 15691
rect 14415 15660 15516 15688
rect 14415 15657 14427 15660
rect 14369 15651 14427 15657
rect 15488 15632 15516 15660
rect 10366 15623 10424 15629
rect 10366 15620 10378 15623
rect 9876 15592 10378 15620
rect 6870 15583 6928 15589
rect 10366 15589 10378 15592
rect 10412 15589 10424 15623
rect 10366 15583 10424 15589
rect 11977 15623 12035 15629
rect 11977 15589 11989 15623
rect 12023 15589 12035 15623
rect 11977 15583 12035 15589
rect 13262 15580 13268 15632
rect 13320 15620 13326 15632
rect 13770 15623 13828 15629
rect 13770 15620 13782 15623
rect 13320 15592 13782 15620
rect 13320 15580 13326 15592
rect 13770 15589 13782 15592
rect 13816 15589 13828 15623
rect 15470 15620 15476 15632
rect 15383 15592 15476 15620
rect 13770 15583 13828 15589
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 6549 15555 6607 15561
rect 6549 15521 6561 15555
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 7742 15512 7748 15564
rect 7800 15552 7806 15564
rect 8294 15552 8300 15564
rect 8352 15561 8358 15564
rect 8352 15555 8390 15561
rect 7800 15524 8300 15552
rect 7800 15512 7806 15524
rect 8294 15512 8300 15524
rect 8378 15521 8390 15555
rect 8352 15515 8390 15521
rect 8352 15512 8358 15515
rect 9306 15512 9312 15564
rect 9364 15552 9370 15564
rect 10042 15552 10048 15564
rect 9364 15524 10048 15552
rect 9364 15512 9370 15524
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 13446 15552 13452 15564
rect 13407 15524 13452 15552
rect 13446 15512 13452 15524
rect 13504 15512 13510 15564
rect 16853 15555 16911 15561
rect 16853 15521 16865 15555
rect 16899 15552 16911 15555
rect 16942 15552 16948 15564
rect 16899 15524 16948 15552
rect 16899 15521 16911 15524
rect 16853 15515 16911 15521
rect 16942 15512 16948 15524
rect 17000 15512 17006 15564
rect 3786 15444 3792 15496
rect 3844 15484 3850 15496
rect 4157 15487 4215 15493
rect 4157 15484 4169 15487
rect 3844 15456 4169 15484
rect 3844 15444 3850 15456
rect 4157 15453 4169 15456
rect 4203 15453 4215 15487
rect 4430 15484 4436 15496
rect 4391 15456 4436 15484
rect 4157 15447 4215 15453
rect 4430 15444 4436 15456
rect 4488 15444 4494 15496
rect 5534 15444 5540 15496
rect 5592 15484 5598 15496
rect 8435 15487 8493 15493
rect 8435 15484 8447 15487
rect 5592 15456 8447 15484
rect 5592 15444 5598 15456
rect 8435 15453 8447 15456
rect 8481 15453 8493 15487
rect 11882 15484 11888 15496
rect 11843 15456 11888 15484
rect 8435 15447 8493 15453
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 12342 15484 12348 15496
rect 12303 15456 12348 15484
rect 12342 15444 12348 15456
rect 12400 15444 12406 15496
rect 15378 15484 15384 15496
rect 15339 15456 15384 15484
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 15654 15484 15660 15496
rect 15615 15456 15660 15484
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 7374 15376 7380 15428
rect 7432 15416 7438 15428
rect 7834 15416 7840 15428
rect 7432 15388 7840 15416
rect 7432 15376 7438 15388
rect 7834 15376 7840 15388
rect 7892 15416 7898 15428
rect 9030 15416 9036 15428
rect 7892 15388 9036 15416
rect 7892 15376 7898 15388
rect 9030 15376 9036 15388
rect 9088 15376 9094 15428
rect 7466 15348 7472 15360
rect 7427 15320 7472 15348
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 11333 15351 11391 15357
rect 11333 15317 11345 15351
rect 11379 15348 11391 15351
rect 11606 15348 11612 15360
rect 11379 15320 11612 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 11606 15308 11612 15320
rect 11664 15308 11670 15360
rect 14090 15308 14096 15360
rect 14148 15348 14154 15360
rect 16991 15351 17049 15357
rect 16991 15348 17003 15351
rect 14148 15320 17003 15348
rect 14148 15308 14154 15320
rect 16991 15317 17003 15320
rect 17037 15317 17049 15351
rect 16991 15311 17049 15317
rect 1104 15258 20884 15280
rect 1104 15206 4648 15258
rect 4700 15206 4712 15258
rect 4764 15206 4776 15258
rect 4828 15206 4840 15258
rect 4892 15206 11982 15258
rect 12034 15206 12046 15258
rect 12098 15206 12110 15258
rect 12162 15206 12174 15258
rect 12226 15206 19315 15258
rect 19367 15206 19379 15258
rect 19431 15206 19443 15258
rect 19495 15206 19507 15258
rect 19559 15206 20884 15258
rect 1104 15184 20884 15206
rect 2593 15147 2651 15153
rect 2593 15113 2605 15147
rect 2639 15144 2651 15147
rect 4246 15144 4252 15156
rect 2639 15116 4252 15144
rect 2639 15113 2651 15116
rect 2593 15107 2651 15113
rect 4246 15104 4252 15116
rect 4304 15144 4310 15156
rect 5077 15147 5135 15153
rect 5077 15144 5089 15147
rect 4304 15116 5089 15144
rect 4304 15104 4310 15116
rect 5077 15113 5089 15116
rect 5123 15113 5135 15147
rect 5077 15107 5135 15113
rect 5350 15104 5356 15156
rect 5408 15144 5414 15156
rect 5445 15147 5503 15153
rect 5445 15144 5457 15147
rect 5408 15116 5457 15144
rect 5408 15104 5414 15116
rect 5445 15113 5457 15116
rect 5491 15113 5503 15147
rect 8294 15144 8300 15156
rect 8255 15116 8300 15144
rect 5445 15107 5503 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 9858 15104 9864 15156
rect 9916 15144 9922 15156
rect 10045 15147 10103 15153
rect 10045 15144 10057 15147
rect 9916 15116 10057 15144
rect 9916 15104 9922 15116
rect 10045 15113 10057 15116
rect 10091 15113 10103 15147
rect 10594 15144 10600 15156
rect 10555 15116 10600 15144
rect 10045 15107 10103 15113
rect 10594 15104 10600 15116
rect 10652 15104 10658 15156
rect 11790 15144 11796 15156
rect 11751 15116 11796 15144
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 13446 15104 13452 15156
rect 13504 15144 13510 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 13504 15116 13829 15144
rect 13504 15104 13510 15116
rect 13817 15113 13829 15116
rect 13863 15113 13875 15147
rect 14274 15144 14280 15156
rect 14235 15116 14280 15144
rect 13817 15107 13875 15113
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 15470 15144 15476 15156
rect 15431 15116 15476 15144
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 4706 15036 4712 15088
rect 4764 15076 4770 15088
rect 5368 15076 5396 15104
rect 7926 15076 7932 15088
rect 4764 15048 5396 15076
rect 7887 15048 7932 15076
rect 4764 15036 4770 15048
rect 7926 15036 7932 15048
rect 7984 15036 7990 15088
rect 8312 15076 8340 15104
rect 10686 15076 10692 15088
rect 8312 15048 10692 15076
rect 10686 15036 10692 15048
rect 10744 15036 10750 15088
rect 10870 15036 10876 15088
rect 10928 15076 10934 15088
rect 11333 15079 11391 15085
rect 11333 15076 11345 15079
rect 10928 15048 11345 15076
rect 10928 15036 10934 15048
rect 11333 15045 11345 15048
rect 11379 15076 11391 15079
rect 12342 15076 12348 15088
rect 11379 15048 12348 15076
rect 11379 15045 11391 15048
rect 11333 15039 11391 15045
rect 12342 15036 12348 15048
rect 12400 15036 12406 15088
rect 15378 15036 15384 15088
rect 15436 15076 15442 15088
rect 15841 15079 15899 15085
rect 15841 15076 15853 15079
rect 15436 15048 15853 15076
rect 15436 15036 15442 15048
rect 15841 15045 15853 15048
rect 15887 15076 15899 15079
rect 16022 15076 16028 15088
rect 15887 15048 16028 15076
rect 15887 15045 15899 15048
rect 15841 15039 15899 15045
rect 16022 15036 16028 15048
rect 16080 15036 16086 15088
rect 16209 15079 16267 15085
rect 16209 15045 16221 15079
rect 16255 15076 16267 15079
rect 21542 15076 21548 15088
rect 16255 15048 21548 15076
rect 16255 15045 16267 15048
rect 16209 15039 16267 15045
rect 21542 15036 21548 15048
rect 21600 15036 21606 15088
rect 1670 15008 1676 15020
rect 1631 14980 1676 15008
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 3878 15008 3884 15020
rect 3467 14980 3884 15008
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 4217 14980 6561 15008
rect 4217 14881 4245 14980
rect 6549 14977 6561 14980
rect 6595 15008 6607 15011
rect 6638 15008 6644 15020
rect 6595 14980 6644 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 7374 15008 7380 15020
rect 7335 14980 7380 15008
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 8938 15008 8944 15020
rect 8899 14980 8944 15008
rect 8938 14968 8944 14980
rect 8996 14968 9002 15020
rect 9030 14968 9036 15020
rect 9088 15008 9094 15020
rect 9217 15011 9275 15017
rect 9217 15008 9229 15011
rect 9088 14980 9229 15008
rect 9088 14968 9094 14980
rect 9217 14977 9229 14980
rect 9263 14977 9275 15011
rect 9217 14971 9275 14977
rect 10781 15011 10839 15017
rect 10781 14977 10793 15011
rect 10827 15008 10839 15011
rect 11606 15008 11612 15020
rect 10827 14980 11612 15008
rect 10827 14977 10839 14980
rect 10781 14971 10839 14977
rect 11606 14968 11612 14980
rect 11664 14968 11670 15020
rect 13173 15011 13231 15017
rect 13173 14977 13185 15011
rect 13219 15008 13231 15011
rect 13354 15008 13360 15020
rect 13219 14980 13360 15008
rect 13219 14977 13231 14980
rect 13173 14971 13231 14977
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 15008 14611 15011
rect 14734 15008 14740 15020
rect 14599 14980 14740 15008
rect 14599 14977 14611 14980
rect 14553 14971 14611 14977
rect 14734 14968 14740 14980
rect 14792 14968 14798 15020
rect 15197 15011 15255 15017
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 15286 15008 15292 15020
rect 15243 14980 15292 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 15286 14968 15292 14980
rect 15344 15008 15350 15020
rect 15654 15008 15660 15020
rect 15344 14980 15660 15008
rect 15344 14968 15350 14980
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 5680 14943 5738 14949
rect 5680 14909 5692 14943
rect 5726 14940 5738 14943
rect 5726 14912 6224 14940
rect 5726 14909 5738 14912
rect 5680 14903 5738 14909
rect 4202 14875 4260 14881
rect 4202 14872 4214 14875
rect 3712 14844 4214 14872
rect 1946 14764 1952 14816
rect 2004 14804 2010 14816
rect 3712 14813 3740 14844
rect 4202 14841 4214 14844
rect 4248 14841 4260 14875
rect 4202 14835 4260 14841
rect 4338 14832 4344 14884
rect 4396 14872 4402 14884
rect 5767 14875 5825 14881
rect 5767 14872 5779 14875
rect 4396 14844 5779 14872
rect 4396 14832 4402 14844
rect 5767 14841 5779 14844
rect 5813 14841 5825 14875
rect 5767 14835 5825 14841
rect 2041 14807 2099 14813
rect 2041 14804 2053 14807
rect 2004 14776 2053 14804
rect 2004 14764 2010 14776
rect 2041 14773 2053 14776
rect 2087 14804 2099 14807
rect 2869 14807 2927 14813
rect 2869 14804 2881 14807
rect 2087 14776 2881 14804
rect 2087 14773 2099 14776
rect 2041 14767 2099 14773
rect 2869 14773 2881 14776
rect 2915 14804 2927 14807
rect 3697 14807 3755 14813
rect 3697 14804 3709 14807
rect 2915 14776 3709 14804
rect 2915 14773 2927 14776
rect 2869 14767 2927 14773
rect 3697 14773 3709 14776
rect 3743 14773 3755 14807
rect 3697 14767 3755 14773
rect 3786 14764 3792 14816
rect 3844 14804 3850 14816
rect 4706 14804 4712 14816
rect 3844 14776 4712 14804
rect 3844 14764 3850 14776
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 4801 14807 4859 14813
rect 4801 14773 4813 14807
rect 4847 14804 4859 14807
rect 5074 14804 5080 14816
rect 4847 14776 5080 14804
rect 4847 14773 4859 14776
rect 4801 14767 4859 14773
rect 5074 14764 5080 14776
rect 5132 14764 5138 14816
rect 6196 14813 6224 14912
rect 12342 14900 12348 14952
rect 12400 14940 12406 14952
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12400 14912 12449 14940
rect 12400 14900 12406 14912
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12989 14943 13047 14949
rect 12989 14909 13001 14943
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 16025 14943 16083 14949
rect 16025 14909 16037 14943
rect 16071 14940 16083 14943
rect 16071 14912 16712 14940
rect 16071 14909 16083 14912
rect 16025 14903 16083 14909
rect 7466 14832 7472 14884
rect 7524 14872 7530 14884
rect 8754 14872 8760 14884
rect 7524 14844 7569 14872
rect 8667 14844 8760 14872
rect 7524 14832 7530 14844
rect 8754 14832 8760 14844
rect 8812 14872 8818 14884
rect 9033 14875 9091 14881
rect 9033 14872 9045 14875
rect 8812 14844 9045 14872
rect 8812 14832 8818 14844
rect 9033 14841 9045 14844
rect 9079 14841 9091 14875
rect 9033 14835 9091 14841
rect 10873 14875 10931 14881
rect 10873 14841 10885 14875
rect 10919 14841 10931 14875
rect 10873 14835 10931 14841
rect 6181 14807 6239 14813
rect 6181 14773 6193 14807
rect 6227 14804 6239 14807
rect 6454 14804 6460 14816
rect 6227 14776 6460 14804
rect 6227 14773 6239 14776
rect 6181 14767 6239 14773
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 7193 14807 7251 14813
rect 7193 14773 7205 14807
rect 7239 14804 7251 14807
rect 7484 14804 7512 14832
rect 7239 14776 7512 14804
rect 7239 14773 7251 14776
rect 7193 14767 7251 14773
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 10888 14804 10916 14835
rect 10652 14776 10916 14804
rect 10652 14764 10658 14776
rect 11514 14764 11520 14816
rect 11572 14804 11578 14816
rect 12253 14807 12311 14813
rect 12253 14804 12265 14807
rect 11572 14776 12265 14804
rect 11572 14764 11578 14776
rect 12253 14773 12265 14776
rect 12299 14804 12311 14807
rect 13004 14804 13032 14903
rect 13262 14832 13268 14884
rect 13320 14872 13326 14884
rect 13449 14875 13507 14881
rect 13449 14872 13461 14875
rect 13320 14844 13461 14872
rect 13320 14832 13326 14844
rect 13449 14841 13461 14844
rect 13495 14841 13507 14875
rect 13449 14835 13507 14841
rect 14274 14832 14280 14884
rect 14332 14872 14338 14884
rect 16684 14881 16712 14912
rect 16850 14900 16856 14952
rect 16908 14940 16914 14952
rect 18084 14943 18142 14949
rect 18084 14940 18096 14943
rect 16908 14912 18096 14940
rect 16908 14900 16914 14912
rect 18084 14909 18096 14912
rect 18130 14940 18142 14943
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18130 14912 18521 14940
rect 18130 14909 18142 14912
rect 18084 14903 18142 14909
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 14645 14875 14703 14881
rect 14645 14872 14657 14875
rect 14332 14844 14657 14872
rect 14332 14832 14338 14844
rect 14645 14841 14657 14844
rect 14691 14841 14703 14875
rect 14645 14835 14703 14841
rect 16669 14875 16727 14881
rect 16669 14841 16681 14875
rect 16715 14872 16727 14875
rect 18966 14872 18972 14884
rect 16715 14844 18972 14872
rect 16715 14841 16727 14844
rect 16669 14835 16727 14841
rect 18966 14832 18972 14844
rect 19024 14832 19030 14884
rect 15470 14804 15476 14816
rect 12299 14776 15476 14804
rect 12299 14773 12311 14776
rect 12253 14767 12311 14773
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 16942 14804 16948 14816
rect 16903 14776 16948 14804
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 17034 14764 17040 14816
rect 17092 14804 17098 14816
rect 18187 14807 18245 14813
rect 18187 14804 18199 14807
rect 17092 14776 18199 14804
rect 17092 14764 17098 14776
rect 18187 14773 18199 14776
rect 18233 14773 18245 14807
rect 18187 14767 18245 14773
rect 1104 14714 20884 14736
rect 1104 14662 8315 14714
rect 8367 14662 8379 14714
rect 8431 14662 8443 14714
rect 8495 14662 8507 14714
rect 8559 14662 15648 14714
rect 15700 14662 15712 14714
rect 15764 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 20884 14714
rect 1104 14640 20884 14662
rect 1765 14603 1823 14609
rect 1765 14569 1777 14603
rect 1811 14600 1823 14603
rect 1946 14600 1952 14612
rect 1811 14572 1952 14600
rect 1811 14569 1823 14572
rect 1765 14563 1823 14569
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 7190 14560 7196 14612
rect 7248 14600 7254 14612
rect 7377 14603 7435 14609
rect 7377 14600 7389 14603
rect 7248 14572 7389 14600
rect 7248 14560 7254 14572
rect 7377 14569 7389 14572
rect 7423 14600 7435 14603
rect 8754 14600 8760 14612
rect 7423 14572 8760 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 8754 14560 8760 14572
rect 8812 14560 8818 14612
rect 8938 14600 8944 14612
rect 8899 14572 8944 14600
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 10042 14600 10048 14612
rect 10003 14572 10048 14600
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 11348 14572 11805 14600
rect 2501 14535 2559 14541
rect 2501 14501 2513 14535
rect 2547 14532 2559 14535
rect 2590 14532 2596 14544
rect 2547 14504 2596 14532
rect 2547 14501 2559 14504
rect 2501 14495 2559 14501
rect 2590 14492 2596 14504
rect 2648 14492 2654 14544
rect 3053 14535 3111 14541
rect 3053 14501 3065 14535
rect 3099 14532 3111 14535
rect 3786 14532 3792 14544
rect 3099 14504 3792 14532
rect 3099 14501 3111 14504
rect 3053 14495 3111 14501
rect 3786 14492 3792 14504
rect 3844 14492 3850 14544
rect 3881 14535 3939 14541
rect 3881 14501 3893 14535
rect 3927 14532 3939 14535
rect 4338 14532 4344 14544
rect 3927 14504 4344 14532
rect 3927 14501 3939 14504
rect 3881 14495 3939 14501
rect 4338 14492 4344 14504
rect 4396 14492 4402 14544
rect 4433 14535 4491 14541
rect 4433 14501 4445 14535
rect 4479 14532 4491 14535
rect 5074 14532 5080 14544
rect 4479 14504 5080 14532
rect 4479 14501 4491 14504
rect 4433 14495 4491 14501
rect 5074 14492 5080 14504
rect 5132 14492 5138 14544
rect 6638 14492 6644 14544
rect 6696 14532 6702 14544
rect 6778 14535 6836 14541
rect 6778 14532 6790 14535
rect 6696 14504 6790 14532
rect 6696 14492 6702 14504
rect 6778 14501 6790 14504
rect 6824 14501 6836 14535
rect 10778 14532 10784 14544
rect 10739 14504 10784 14532
rect 6778 14495 6836 14501
rect 10778 14492 10784 14504
rect 10836 14492 10842 14544
rect 11054 14492 11060 14544
rect 11112 14532 11118 14544
rect 11348 14541 11376 14572
rect 11793 14569 11805 14572
rect 11839 14600 11851 14603
rect 11882 14600 11888 14612
rect 11839 14572 11888 14600
rect 11839 14569 11851 14572
rect 11793 14563 11851 14569
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 12161 14603 12219 14609
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 12526 14600 12532 14612
rect 12207 14572 12532 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 14090 14600 14096 14612
rect 14051 14572 14096 14600
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 11333 14535 11391 14541
rect 11333 14532 11345 14535
rect 11112 14504 11345 14532
rect 11112 14492 11118 14504
rect 11333 14501 11345 14504
rect 11379 14501 11391 14535
rect 11333 14495 11391 14501
rect 13075 14535 13133 14541
rect 13075 14501 13087 14535
rect 13121 14532 13133 14535
rect 13262 14532 13268 14544
rect 13121 14504 13268 14532
rect 13121 14501 13133 14504
rect 13075 14495 13133 14501
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 15102 14492 15108 14544
rect 15160 14532 15166 14544
rect 15473 14535 15531 14541
rect 15473 14532 15485 14535
rect 15160 14504 15485 14532
rect 15160 14492 15166 14504
rect 15473 14501 15485 14504
rect 15519 14501 15531 14535
rect 16022 14532 16028 14544
rect 15983 14504 16028 14532
rect 15473 14495 15531 14501
rect 16022 14492 16028 14504
rect 16080 14492 16086 14544
rect 6457 14467 6515 14473
rect 6457 14433 6469 14467
rect 6503 14464 6515 14467
rect 6546 14464 6552 14476
rect 6503 14436 6552 14464
rect 6503 14433 6515 14436
rect 6457 14427 6515 14433
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 8110 14424 8116 14476
rect 8168 14464 8174 14476
rect 8240 14467 8298 14473
rect 8240 14464 8252 14467
rect 8168 14436 8252 14464
rect 8168 14424 8174 14436
rect 8240 14433 8252 14436
rect 8286 14433 8298 14467
rect 14550 14464 14556 14476
rect 8240 14427 8298 14433
rect 12452 14436 14556 14464
rect 2409 14399 2467 14405
rect 2409 14365 2421 14399
rect 2455 14396 2467 14399
rect 3329 14399 3387 14405
rect 3329 14396 3341 14399
rect 2455 14368 3341 14396
rect 2455 14365 2467 14368
rect 2409 14359 2467 14365
rect 3329 14365 3341 14368
rect 3375 14396 3387 14399
rect 4982 14396 4988 14408
rect 3375 14368 4154 14396
rect 4943 14368 4988 14396
rect 3375 14365 3387 14368
rect 3329 14359 3387 14365
rect 4126 14328 4154 14368
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 10686 14396 10692 14408
rect 10647 14368 10692 14396
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 5166 14328 5172 14340
rect 4126 14300 5172 14328
rect 5166 14288 5172 14300
rect 5224 14288 5230 14340
rect 8662 14288 8668 14340
rect 8720 14328 8726 14340
rect 12342 14328 12348 14340
rect 8720 14300 12348 14328
rect 8720 14288 8726 14300
rect 12342 14288 12348 14300
rect 12400 14328 12406 14340
rect 12452 14337 12480 14436
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 16920 14467 16978 14473
rect 16920 14433 16932 14467
rect 16966 14464 16978 14467
rect 17310 14464 17316 14476
rect 16966 14436 17316 14464
rect 16966 14433 16978 14436
rect 16920 14427 16978 14433
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 17770 14424 17776 14476
rect 17828 14464 17834 14476
rect 17900 14467 17958 14473
rect 17900 14464 17912 14467
rect 17828 14436 17912 14464
rect 17828 14424 17834 14436
rect 17900 14433 17912 14436
rect 17946 14433 17958 14467
rect 17900 14427 17958 14433
rect 12710 14396 12716 14408
rect 12671 14368 12716 14396
rect 12710 14356 12716 14368
rect 12768 14356 12774 14408
rect 15381 14399 15439 14405
rect 15381 14396 15393 14399
rect 15028 14368 15393 14396
rect 12437 14331 12495 14337
rect 12437 14328 12449 14331
rect 12400 14300 12449 14328
rect 12400 14288 12406 14300
rect 12437 14297 12449 14300
rect 12483 14297 12495 14331
rect 12437 14291 12495 14297
rect 15028 14272 15056 14368
rect 15381 14365 15393 14368
rect 15427 14365 15439 14399
rect 15381 14359 15439 14365
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 4430 14260 4436 14272
rect 4212 14232 4436 14260
rect 4212 14220 4218 14232
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 7742 14260 7748 14272
rect 7655 14232 7748 14260
rect 7742 14220 7748 14232
rect 7800 14260 7806 14272
rect 8343 14263 8401 14269
rect 8343 14260 8355 14263
rect 7800 14232 8355 14260
rect 7800 14220 7806 14232
rect 8343 14229 8355 14232
rect 8389 14229 8401 14263
rect 8343 14223 8401 14229
rect 10502 14220 10508 14272
rect 10560 14260 10566 14272
rect 11698 14260 11704 14272
rect 10560 14232 11704 14260
rect 10560 14220 10566 14232
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 13630 14260 13636 14272
rect 13591 14232 13636 14260
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 14553 14263 14611 14269
rect 14553 14229 14565 14263
rect 14599 14260 14611 14263
rect 14734 14260 14740 14272
rect 14599 14232 14740 14260
rect 14599 14229 14611 14232
rect 14553 14223 14611 14229
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 15010 14260 15016 14272
rect 14971 14232 15016 14260
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 15194 14220 15200 14272
rect 15252 14260 15258 14272
rect 16991 14263 17049 14269
rect 16991 14260 17003 14263
rect 15252 14232 17003 14260
rect 15252 14220 15258 14232
rect 16991 14229 17003 14232
rect 17037 14229 17049 14263
rect 16991 14223 17049 14229
rect 17126 14220 17132 14272
rect 17184 14260 17190 14272
rect 18003 14263 18061 14269
rect 18003 14260 18015 14263
rect 17184 14232 18015 14260
rect 17184 14220 17190 14232
rect 18003 14229 18015 14232
rect 18049 14229 18061 14263
rect 18003 14223 18061 14229
rect 1104 14170 20884 14192
rect 1104 14118 4648 14170
rect 4700 14118 4712 14170
rect 4764 14118 4776 14170
rect 4828 14118 4840 14170
rect 4892 14118 11982 14170
rect 12034 14118 12046 14170
rect 12098 14118 12110 14170
rect 12162 14118 12174 14170
rect 12226 14118 19315 14170
rect 19367 14118 19379 14170
rect 19431 14118 19443 14170
rect 19495 14118 19507 14170
rect 19559 14118 20884 14170
rect 1104 14096 20884 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 4430 14056 4436 14068
rect 1452 14028 4436 14056
rect 1452 14016 1458 14028
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 5074 14016 5080 14068
rect 5132 14056 5138 14068
rect 5169 14059 5227 14065
rect 5169 14056 5181 14059
rect 5132 14028 5181 14056
rect 5132 14016 5138 14028
rect 5169 14025 5181 14028
rect 5215 14025 5227 14059
rect 7190 14056 7196 14068
rect 7151 14028 7196 14056
rect 5169 14019 5227 14025
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 8110 14016 8116 14068
rect 8168 14056 8174 14068
rect 8205 14059 8263 14065
rect 8205 14056 8217 14059
rect 8168 14028 8217 14056
rect 8168 14016 8174 14028
rect 8205 14025 8217 14028
rect 8251 14025 8263 14059
rect 8205 14019 8263 14025
rect 11471 14059 11529 14065
rect 11471 14025 11483 14059
rect 11517 14056 11529 14059
rect 15010 14056 15016 14068
rect 11517 14028 15016 14056
rect 11517 14025 11529 14028
rect 11471 14019 11529 14025
rect 15010 14016 15016 14028
rect 15068 14016 15074 14068
rect 15286 14016 15292 14068
rect 15344 14056 15350 14068
rect 18187 14059 18245 14065
rect 18187 14056 18199 14059
rect 15344 14028 18199 14056
rect 15344 14016 15350 14028
rect 18187 14025 18199 14028
rect 18233 14025 18245 14059
rect 18187 14019 18245 14025
rect 1949 13991 2007 13997
rect 1949 13957 1961 13991
rect 1995 13988 2007 13991
rect 2406 13988 2412 14000
rect 1995 13960 2412 13988
rect 1995 13957 2007 13960
rect 1949 13951 2007 13957
rect 1448 13855 1506 13861
rect 1448 13821 1460 13855
rect 1494 13852 1506 13855
rect 1964 13852 1992 13951
rect 2406 13948 2412 13960
rect 2464 13948 2470 14000
rect 2958 13948 2964 14000
rect 3016 13988 3022 14000
rect 3053 13991 3111 13997
rect 3053 13988 3065 13991
rect 3016 13960 3065 13988
rect 3016 13948 3022 13960
rect 3053 13957 3065 13960
rect 3099 13988 3111 13991
rect 4801 13991 4859 13997
rect 4801 13988 4813 13991
rect 3099 13960 4813 13988
rect 3099 13957 3111 13960
rect 3053 13951 3111 13957
rect 4801 13957 4813 13960
rect 4847 13988 4859 13991
rect 4982 13988 4988 14000
rect 4847 13960 4988 13988
rect 4847 13957 4859 13960
rect 4801 13951 4859 13957
rect 4982 13948 4988 13960
rect 5040 13948 5046 14000
rect 10686 13948 10692 14000
rect 10744 13988 10750 14000
rect 11149 13991 11207 13997
rect 11149 13988 11161 13991
rect 10744 13960 11161 13988
rect 10744 13948 10750 13960
rect 11149 13957 11161 13960
rect 11195 13988 11207 13991
rect 17126 13988 17132 14000
rect 11195 13960 17132 13988
rect 11195 13957 11207 13960
rect 11149 13951 11207 13957
rect 17126 13948 17132 13960
rect 17184 13948 17190 14000
rect 19199 13991 19257 13997
rect 19199 13988 19211 13991
rect 17236 13960 19211 13988
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13920 4307 13923
rect 5537 13923 5595 13929
rect 5537 13920 5549 13923
rect 4295 13892 5549 13920
rect 4295 13889 4307 13892
rect 4249 13883 4307 13889
rect 5537 13889 5549 13892
rect 5583 13920 5595 13923
rect 5859 13923 5917 13929
rect 5859 13920 5871 13923
rect 5583 13892 5871 13920
rect 5583 13889 5595 13892
rect 5537 13883 5595 13889
rect 5859 13889 5871 13892
rect 5905 13889 5917 13923
rect 5859 13883 5917 13889
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13920 7435 13923
rect 7742 13920 7748 13932
rect 7423 13892 7748 13920
rect 7423 13889 7435 13892
rect 7377 13883 7435 13889
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 8018 13920 8024 13932
rect 7979 13892 8024 13920
rect 8018 13880 8024 13892
rect 8076 13880 8082 13932
rect 9033 13923 9091 13929
rect 9033 13889 9045 13923
rect 9079 13920 9091 13923
rect 9490 13920 9496 13932
rect 9079 13892 9496 13920
rect 9079 13889 9091 13892
rect 9033 13883 9091 13889
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 10778 13920 10784 13932
rect 10428 13892 10784 13920
rect 5756 13855 5814 13861
rect 5756 13852 5768 13855
rect 1494 13824 1992 13852
rect 1494 13821 1506 13824
rect 1448 13815 1506 13821
rect 5736 13821 5768 13852
rect 5802 13821 5814 13855
rect 5736 13815 5814 13821
rect 1535 13787 1593 13793
rect 1535 13753 1547 13787
rect 1581 13784 1593 13787
rect 2498 13784 2504 13796
rect 1581 13756 2504 13784
rect 1581 13753 1593 13756
rect 1535 13747 1593 13753
rect 2498 13744 2504 13756
rect 2556 13744 2562 13796
rect 2590 13744 2596 13796
rect 2648 13784 2654 13796
rect 3421 13787 3479 13793
rect 3421 13784 3433 13787
rect 2648 13756 3433 13784
rect 2648 13744 2654 13756
rect 3421 13753 3433 13756
rect 3467 13753 3479 13787
rect 3421 13747 3479 13753
rect 4065 13787 4123 13793
rect 4065 13753 4077 13787
rect 4111 13784 4123 13787
rect 4338 13784 4344 13796
rect 4111 13756 4344 13784
rect 4111 13753 4123 13756
rect 4065 13747 4123 13753
rect 4338 13744 4344 13756
rect 4396 13744 4402 13796
rect 4430 13744 4436 13796
rect 4488 13784 4494 13796
rect 5736 13784 5764 13815
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 10134 13852 10140 13864
rect 8168 13824 10140 13852
rect 8168 13812 8174 13824
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 10428 13861 10456 13892
rect 10778 13880 10784 13892
rect 10836 13920 10842 13932
rect 12526 13920 12532 13932
rect 10836 13892 12296 13920
rect 12487 13892 12532 13920
rect 10836 13880 10842 13892
rect 10413 13855 10471 13861
rect 10413 13821 10425 13855
rect 10459 13821 10471 13855
rect 10413 13815 10471 13821
rect 10870 13812 10876 13864
rect 10928 13852 10934 13864
rect 11368 13855 11426 13861
rect 11368 13852 11380 13855
rect 10928 13824 11380 13852
rect 10928 13812 10934 13824
rect 11368 13821 11380 13824
rect 11414 13852 11426 13855
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 11414 13824 11805 13852
rect 11414 13821 11426 13824
rect 11368 13815 11426 13821
rect 11793 13821 11805 13824
rect 11839 13821 11851 13855
rect 11793 13815 11851 13821
rect 6181 13787 6239 13793
rect 6181 13784 6193 13787
rect 4488 13756 6193 13784
rect 4488 13744 4494 13756
rect 6181 13753 6193 13756
rect 6227 13784 6239 13787
rect 6227 13756 7144 13784
rect 6227 13753 6239 13756
rect 6181 13747 6239 13753
rect 2317 13719 2375 13725
rect 2317 13685 2329 13719
rect 2363 13716 2375 13719
rect 2608 13716 2636 13744
rect 6638 13716 6644 13728
rect 2363 13688 2636 13716
rect 6599 13688 6644 13716
rect 2363 13685 2375 13688
rect 2317 13679 2375 13685
rect 6638 13676 6644 13688
rect 6696 13676 6702 13728
rect 7116 13716 7144 13756
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 7469 13787 7527 13793
rect 7469 13784 7481 13787
rect 7248 13756 7481 13784
rect 7248 13744 7254 13756
rect 7469 13753 7481 13756
rect 7515 13753 7527 13787
rect 7469 13747 7527 13753
rect 9401 13787 9459 13793
rect 9401 13753 9413 13787
rect 9447 13784 9459 13787
rect 9674 13784 9680 13796
rect 9447 13756 9680 13784
rect 9447 13753 9459 13756
rect 9401 13747 9459 13753
rect 9674 13744 9680 13756
rect 9732 13784 9738 13796
rect 12268 13793 12296 13892
rect 12526 13880 12532 13892
rect 12584 13880 12590 13932
rect 12802 13920 12808 13932
rect 12763 13892 12808 13920
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 14090 13920 14096 13932
rect 14051 13892 14096 13920
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 17236 13920 17264 13960
rect 19199 13957 19211 13960
rect 19245 13957 19257 13991
rect 19199 13951 19257 13957
rect 18509 13923 18567 13929
rect 18509 13920 18521 13923
rect 14332 13892 17264 13920
rect 18099 13892 18521 13920
rect 14332 13880 14338 13892
rect 14918 13812 14924 13864
rect 14976 13852 14982 13864
rect 15470 13852 15476 13864
rect 14976 13824 15399 13852
rect 15431 13824 15476 13852
rect 14976 13812 14982 13824
rect 9814 13787 9872 13793
rect 9814 13784 9826 13787
rect 9732 13756 9826 13784
rect 9732 13744 9738 13756
rect 9814 13753 9826 13756
rect 9860 13753 9872 13787
rect 9814 13747 9872 13753
rect 12253 13787 12311 13793
rect 12253 13753 12265 13787
rect 12299 13784 12311 13787
rect 12621 13787 12679 13793
rect 12621 13784 12633 13787
rect 12299 13756 12633 13784
rect 12299 13753 12311 13756
rect 12253 13747 12311 13753
rect 12621 13753 12633 13756
rect 12667 13753 12679 13787
rect 12621 13747 12679 13753
rect 13170 13744 13176 13796
rect 13228 13784 13234 13796
rect 13541 13787 13599 13793
rect 13541 13784 13553 13787
rect 13228 13756 13553 13784
rect 13228 13744 13234 13756
rect 13541 13753 13553 13756
rect 13587 13784 13599 13787
rect 13722 13784 13728 13796
rect 13587 13756 13728 13784
rect 13587 13753 13599 13756
rect 13541 13747 13599 13753
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 13909 13787 13967 13793
rect 13909 13753 13921 13787
rect 13955 13784 13967 13787
rect 14182 13784 14188 13796
rect 13955 13756 14188 13784
rect 13955 13753 13967 13756
rect 13909 13747 13967 13753
rect 8205 13719 8263 13725
rect 8205 13716 8217 13719
rect 7116 13688 8217 13716
rect 8205 13685 8217 13688
rect 8251 13716 8263 13719
rect 8297 13719 8355 13725
rect 8297 13716 8309 13719
rect 8251 13688 8309 13716
rect 8251 13685 8263 13688
rect 8205 13679 8263 13685
rect 8297 13685 8309 13688
rect 8343 13716 8355 13719
rect 8846 13716 8852 13728
rect 8343 13688 8852 13716
rect 8343 13685 8355 13688
rect 8297 13679 8355 13685
rect 8846 13676 8852 13688
rect 8904 13676 8910 13728
rect 9490 13676 9496 13728
rect 9548 13716 9554 13728
rect 11238 13716 11244 13728
rect 9548 13688 11244 13716
rect 9548 13676 9554 13688
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 11606 13676 11612 13728
rect 11664 13716 11670 13728
rect 12802 13716 12808 13728
rect 11664 13688 12808 13716
rect 11664 13676 11670 13688
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 13630 13676 13636 13728
rect 13688 13716 13694 13728
rect 13924 13716 13952 13747
rect 14182 13744 14188 13756
rect 14240 13744 14246 13796
rect 14734 13784 14740 13796
rect 14695 13756 14740 13784
rect 14734 13744 14740 13756
rect 14792 13744 14798 13796
rect 15371 13784 15399 13824
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 15580 13784 15608 13815
rect 15746 13812 15752 13864
rect 15804 13852 15810 13864
rect 16117 13855 16175 13861
rect 16117 13852 16129 13855
rect 15804 13824 16129 13852
rect 15804 13812 15810 13824
rect 16117 13821 16129 13824
rect 16163 13821 16175 13855
rect 16117 13815 16175 13821
rect 14844 13756 15332 13784
rect 15371 13756 15608 13784
rect 16132 13784 16160 13815
rect 17126 13812 17132 13864
rect 17184 13852 17190 13864
rect 18099 13861 18127 13892
rect 18509 13889 18521 13892
rect 18555 13889 18567 13923
rect 19521 13923 19579 13929
rect 19521 13920 19533 13923
rect 18509 13883 18567 13889
rect 19306 13892 19533 13920
rect 18084 13855 18142 13861
rect 18084 13852 18096 13855
rect 17184 13824 18096 13852
rect 17184 13812 17190 13824
rect 18084 13821 18096 13824
rect 18130 13821 18142 13855
rect 19093 13852 19099 13864
rect 19054 13824 19099 13852
rect 18084 13815 18142 13821
rect 19093 13812 19099 13824
rect 19151 13812 19157 13864
rect 17402 13784 17408 13796
rect 16132 13756 17408 13784
rect 13688 13688 13952 13716
rect 13688 13676 13694 13688
rect 14642 13676 14648 13728
rect 14700 13716 14706 13728
rect 14844 13716 14872 13756
rect 14700 13688 14872 13716
rect 14700 13676 14706 13688
rect 14918 13676 14924 13728
rect 14976 13716 14982 13728
rect 15013 13719 15071 13725
rect 15013 13716 15025 13719
rect 14976 13688 15025 13716
rect 14976 13676 14982 13688
rect 15013 13685 15025 13688
rect 15059 13685 15071 13719
rect 15304 13716 15332 13756
rect 17402 13744 17408 13756
rect 17460 13744 17466 13796
rect 17770 13784 17776 13796
rect 17731 13756 17776 13784
rect 17770 13744 17776 13756
rect 17828 13744 17834 13796
rect 15657 13719 15715 13725
rect 15657 13716 15669 13719
rect 15304 13688 15669 13716
rect 15013 13679 15071 13685
rect 15657 13685 15669 13688
rect 15703 13685 15715 13719
rect 15657 13679 15715 13685
rect 16945 13719 17003 13725
rect 16945 13685 16957 13719
rect 16991 13716 17003 13719
rect 17310 13716 17316 13728
rect 16991 13688 17316 13716
rect 16991 13685 17003 13688
rect 16945 13679 17003 13685
rect 17310 13676 17316 13688
rect 17368 13676 17374 13728
rect 19058 13676 19064 13728
rect 19116 13716 19122 13728
rect 19306 13716 19334 13892
rect 19521 13889 19533 13892
rect 19567 13889 19579 13923
rect 19521 13883 19579 13889
rect 19116 13688 19334 13716
rect 19116 13676 19122 13688
rect 1104 13626 20884 13648
rect 1104 13574 8315 13626
rect 8367 13574 8379 13626
rect 8431 13574 8443 13626
rect 8495 13574 8507 13626
rect 8559 13574 15648 13626
rect 15700 13574 15712 13626
rect 15764 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 20884 13626
rect 1104 13552 20884 13574
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 3605 13515 3663 13521
rect 3605 13512 3617 13515
rect 2556 13484 3617 13512
rect 2556 13472 2562 13484
rect 3605 13481 3617 13484
rect 3651 13481 3663 13515
rect 6546 13512 6552 13524
rect 6507 13484 6552 13512
rect 3605 13475 3663 13481
rect 6546 13472 6552 13484
rect 6604 13472 6610 13524
rect 9306 13472 9312 13524
rect 9364 13512 9370 13524
rect 11514 13512 11520 13524
rect 9364 13484 11520 13512
rect 9364 13472 9370 13484
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 12434 13512 12440 13524
rect 12395 13484 12440 13512
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 12710 13512 12716 13524
rect 12671 13484 12716 13512
rect 12710 13472 12716 13484
rect 12768 13512 12774 13524
rect 14642 13512 14648 13524
rect 12768 13484 14648 13512
rect 12768 13472 12774 13484
rect 14642 13472 14648 13484
rect 14700 13472 14706 13524
rect 16945 13515 17003 13521
rect 16945 13512 16957 13515
rect 14844 13484 16957 13512
rect 1854 13404 1860 13456
rect 1912 13444 1918 13456
rect 1994 13447 2052 13453
rect 1994 13444 2006 13447
rect 1912 13416 2006 13444
rect 1912 13404 1918 13416
rect 1994 13413 2006 13416
rect 2040 13413 2052 13447
rect 1994 13407 2052 13413
rect 4338 13404 4344 13456
rect 4396 13444 4402 13456
rect 4801 13447 4859 13453
rect 4801 13444 4813 13447
rect 4396 13416 4813 13444
rect 4396 13404 4402 13416
rect 4801 13413 4813 13416
rect 4847 13413 4859 13447
rect 5350 13444 5356 13456
rect 5311 13416 5356 13444
rect 4801 13407 4859 13413
rect 5350 13404 5356 13416
rect 5408 13404 5414 13456
rect 5994 13404 6000 13456
rect 6052 13444 6058 13456
rect 6822 13444 6828 13456
rect 6052 13416 6828 13444
rect 6052 13404 6058 13416
rect 6822 13404 6828 13416
rect 6880 13404 6886 13456
rect 7282 13444 7288 13456
rect 7243 13416 7288 13444
rect 7282 13404 7288 13416
rect 7340 13404 7346 13456
rect 10870 13444 10876 13456
rect 10831 13416 10876 13444
rect 10870 13404 10876 13416
rect 10928 13404 10934 13456
rect 13259 13447 13317 13453
rect 13259 13413 13271 13447
rect 13305 13444 13317 13447
rect 13722 13444 13728 13456
rect 13305 13416 13728 13444
rect 13305 13413 13317 13416
rect 13259 13407 13317 13413
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 2590 13376 2596 13388
rect 2551 13348 2596 13376
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 9582 13376 9588 13388
rect 9543 13348 9588 13376
rect 9582 13336 9588 13348
rect 9640 13336 9646 13388
rect 14844 13376 14872 13484
rect 16945 13481 16957 13484
rect 16991 13481 17003 13515
rect 16945 13475 17003 13481
rect 18138 13472 18144 13524
rect 18196 13512 18202 13524
rect 18555 13515 18613 13521
rect 18555 13512 18567 13515
rect 18196 13484 18567 13512
rect 18196 13472 18202 13484
rect 18555 13481 18567 13484
rect 18601 13481 18613 13515
rect 18555 13475 18613 13481
rect 15102 13444 15108 13456
rect 15063 13416 15108 13444
rect 15102 13404 15108 13416
rect 15160 13404 15166 13456
rect 15470 13444 15476 13456
rect 15431 13416 15476 13444
rect 15470 13404 15476 13416
rect 15528 13404 15534 13456
rect 12912 13348 14872 13376
rect 17129 13379 17187 13385
rect 12912 13320 12940 13348
rect 17129 13345 17141 13379
rect 17175 13376 17187 13379
rect 17218 13376 17224 13388
rect 17175 13348 17224 13376
rect 17175 13345 17187 13348
rect 17129 13339 17187 13345
rect 17218 13336 17224 13348
rect 17276 13336 17282 13388
rect 17402 13376 17408 13388
rect 17363 13348 17408 13376
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 18484 13379 18542 13385
rect 18484 13345 18496 13379
rect 18530 13376 18542 13379
rect 18782 13376 18788 13388
rect 18530 13348 18788 13376
rect 18530 13345 18542 13348
rect 18484 13339 18542 13345
rect 18782 13336 18788 13348
rect 18840 13336 18846 13388
rect 19496 13379 19554 13385
rect 19496 13345 19508 13379
rect 19542 13376 19554 13379
rect 19610 13376 19616 13388
rect 19542 13348 19616 13376
rect 19542 13345 19554 13348
rect 19496 13339 19554 13345
rect 19610 13336 19616 13348
rect 19668 13336 19674 13388
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 1762 13308 1768 13320
rect 1719 13280 1768 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 1762 13268 1768 13280
rect 1820 13308 1826 13320
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 1820 13280 3249 13308
rect 1820 13268 1826 13280
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 3237 13271 3295 13277
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 5534 13308 5540 13320
rect 4755 13280 5540 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13308 7251 13311
rect 8110 13308 8116 13320
rect 7239 13280 8116 13308
rect 7239 13277 7251 13280
rect 7193 13271 7251 13277
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13277 10839 13311
rect 11054 13308 11060 13320
rect 11015 13280 11060 13308
rect 10781 13271 10839 13277
rect 2222 13200 2228 13252
rect 2280 13240 2286 13252
rect 2869 13243 2927 13249
rect 2869 13240 2881 13243
rect 2280 13212 2881 13240
rect 2280 13200 2286 13212
rect 2869 13209 2881 13212
rect 2915 13209 2927 13243
rect 2869 13203 2927 13209
rect 7745 13243 7803 13249
rect 7745 13209 7757 13243
rect 7791 13240 7803 13243
rect 8018 13240 8024 13252
rect 7791 13212 8024 13240
rect 7791 13209 7803 13212
rect 7745 13203 7803 13209
rect 8018 13200 8024 13212
rect 8076 13240 8082 13252
rect 8754 13240 8760 13252
rect 8076 13212 8760 13240
rect 8076 13200 8082 13212
rect 8754 13200 8760 13212
rect 8812 13200 8818 13252
rect 10796 13240 10824 13271
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 12894 13308 12900 13320
rect 12855 13280 12900 13308
rect 12894 13268 12900 13280
rect 12952 13268 12958 13320
rect 14642 13268 14648 13320
rect 14700 13308 14706 13320
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 14700 13280 15393 13308
rect 14700 13268 14706 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 16022 13308 16028 13320
rect 15983 13280 16028 13308
rect 15381 13271 15439 13277
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 11422 13240 11428 13252
rect 10796 13212 11428 13240
rect 11422 13200 11428 13212
rect 11480 13240 11486 13252
rect 14274 13240 14280 13252
rect 11480 13212 14280 13240
rect 11480 13200 11486 13212
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 4062 13132 4068 13184
rect 4120 13172 4126 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 4120 13144 4261 13172
rect 4120 13132 4126 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 4249 13135 4307 13141
rect 6546 13132 6552 13184
rect 6604 13172 6610 13184
rect 9815 13175 9873 13181
rect 9815 13172 9827 13175
rect 6604 13144 9827 13172
rect 6604 13132 6610 13144
rect 9815 13141 9827 13144
rect 9861 13141 9873 13175
rect 9815 13135 9873 13141
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 13872 13144 13917 13172
rect 13872 13132 13878 13144
rect 14090 13132 14096 13184
rect 14148 13172 14154 13184
rect 14185 13175 14243 13181
rect 14185 13172 14197 13175
rect 14148 13144 14197 13172
rect 14148 13132 14154 13144
rect 14185 13141 14197 13144
rect 14231 13172 14243 13175
rect 17034 13172 17040 13184
rect 14231 13144 17040 13172
rect 14231 13141 14243 13144
rect 14185 13135 14243 13141
rect 17034 13132 17040 13144
rect 17092 13132 17098 13184
rect 17494 13132 17500 13184
rect 17552 13172 17558 13184
rect 19567 13175 19625 13181
rect 19567 13172 19579 13175
rect 17552 13144 19579 13172
rect 17552 13132 17558 13144
rect 19567 13141 19579 13144
rect 19613 13141 19625 13175
rect 19567 13135 19625 13141
rect 1104 13082 20884 13104
rect 1104 13030 4648 13082
rect 4700 13030 4712 13082
rect 4764 13030 4776 13082
rect 4828 13030 4840 13082
rect 4892 13030 11982 13082
rect 12034 13030 12046 13082
rect 12098 13030 12110 13082
rect 12162 13030 12174 13082
rect 12226 13030 19315 13082
rect 19367 13030 19379 13082
rect 19431 13030 19443 13082
rect 19495 13030 19507 13082
rect 19559 13030 20884 13082
rect 1104 13008 20884 13030
rect 4338 12928 4344 12980
rect 4396 12968 4402 12980
rect 4801 12971 4859 12977
rect 4801 12968 4813 12971
rect 4396 12940 4813 12968
rect 4396 12928 4402 12940
rect 4801 12937 4813 12940
rect 4847 12968 4859 12971
rect 5077 12971 5135 12977
rect 5077 12968 5089 12971
rect 4847 12940 5089 12968
rect 4847 12937 4859 12940
rect 4801 12931 4859 12937
rect 5077 12937 5089 12940
rect 5123 12937 5135 12971
rect 5077 12931 5135 12937
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 5767 12971 5825 12977
rect 5767 12968 5779 12971
rect 5224 12940 5779 12968
rect 5224 12928 5230 12940
rect 5767 12937 5779 12940
rect 5813 12937 5825 12971
rect 5767 12931 5825 12937
rect 7282 12928 7288 12980
rect 7340 12968 7346 12980
rect 7745 12971 7803 12977
rect 7745 12968 7757 12971
rect 7340 12940 7757 12968
rect 7340 12928 7346 12940
rect 7745 12937 7757 12940
rect 7791 12937 7803 12971
rect 8110 12968 8116 12980
rect 8071 12940 8116 12968
rect 7745 12931 7803 12937
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 10870 12968 10876 12980
rect 10831 12940 10876 12968
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 12894 12968 12900 12980
rect 12299 12940 12900 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 13909 12971 13967 12977
rect 13909 12968 13921 12971
rect 13872 12940 13921 12968
rect 13872 12928 13878 12940
rect 13909 12937 13921 12940
rect 13955 12968 13967 12971
rect 14182 12968 14188 12980
rect 13955 12940 14188 12968
rect 13955 12937 13967 12940
rect 13909 12931 13967 12937
rect 14182 12928 14188 12940
rect 14240 12968 14246 12980
rect 15105 12971 15163 12977
rect 15105 12968 15117 12971
rect 14240 12940 15117 12968
rect 14240 12928 14246 12940
rect 15105 12937 15117 12940
rect 15151 12968 15163 12971
rect 15470 12968 15476 12980
rect 15151 12940 15476 12968
rect 15151 12937 15163 12940
rect 15105 12931 15163 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 19610 12968 19616 12980
rect 18748 12940 19616 12968
rect 18748 12928 18754 12940
rect 19610 12928 19616 12940
rect 19668 12928 19674 12980
rect 5534 12900 5540 12912
rect 5495 12872 5540 12900
rect 5534 12860 5540 12872
rect 5592 12860 5598 12912
rect 6454 12860 6460 12912
rect 6512 12900 6518 12912
rect 9582 12900 9588 12912
rect 6512 12872 9588 12900
rect 6512 12860 6518 12872
rect 9582 12860 9588 12872
rect 9640 12900 9646 12912
rect 10505 12903 10563 12909
rect 10505 12900 10517 12903
rect 9640 12872 10517 12900
rect 9640 12860 9646 12872
rect 10505 12869 10517 12872
rect 10551 12900 10563 12903
rect 11882 12900 11888 12912
rect 10551 12872 11888 12900
rect 10551 12869 10563 12872
rect 10505 12863 10563 12869
rect 11882 12860 11888 12872
rect 11940 12860 11946 12912
rect 12434 12860 12440 12912
rect 12492 12900 12498 12912
rect 14645 12903 14703 12909
rect 12492 12872 12572 12900
rect 12492 12860 12498 12872
rect 1486 12792 1492 12844
rect 1544 12832 1550 12844
rect 2133 12835 2191 12841
rect 2133 12832 2145 12835
rect 1544 12804 2145 12832
rect 1544 12792 1550 12804
rect 2133 12801 2145 12804
rect 2179 12832 2191 12835
rect 3053 12835 3111 12841
rect 3053 12832 3065 12835
rect 2179 12804 3065 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 3053 12801 3065 12804
rect 3099 12801 3111 12835
rect 6822 12832 6828 12844
rect 6783 12804 6828 12832
rect 3053 12795 3111 12801
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 12544 12841 12572 12872
rect 14645 12869 14657 12903
rect 14691 12900 14703 12903
rect 14826 12900 14832 12912
rect 14691 12872 14832 12900
rect 14691 12869 14703 12872
rect 14645 12863 14703 12869
rect 14826 12860 14832 12872
rect 14884 12900 14890 12912
rect 16209 12903 16267 12909
rect 16209 12900 16221 12903
rect 14884 12872 16221 12900
rect 14884 12860 14890 12872
rect 16209 12869 16221 12872
rect 16255 12869 16267 12903
rect 16209 12863 16267 12869
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12801 12587 12835
rect 12802 12832 12808 12844
rect 12763 12804 12808 12832
rect 12529 12795 12587 12801
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 14090 12832 14096 12844
rect 14051 12804 14096 12832
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 15657 12835 15715 12841
rect 15657 12801 15669 12835
rect 15703 12832 15715 12835
rect 16390 12832 16396 12844
rect 15703 12804 16396 12832
rect 15703 12801 15715 12804
rect 15657 12795 15715 12801
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 16945 12835 17003 12841
rect 16945 12801 16957 12835
rect 16991 12832 17003 12835
rect 17402 12832 17408 12844
rect 16991 12804 17408 12832
rect 16991 12801 17003 12804
rect 16945 12795 17003 12801
rect 17402 12792 17408 12804
rect 17460 12832 17466 12844
rect 18598 12832 18604 12844
rect 17460 12804 18604 12832
rect 17460 12792 17466 12804
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 4062 12764 4068 12776
rect 3927 12736 4068 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 5696 12767 5754 12773
rect 5696 12733 5708 12767
rect 5742 12764 5754 12767
rect 6086 12764 6092 12776
rect 5742 12736 6092 12764
rect 5742 12733 5754 12736
rect 5696 12727 5754 12733
rect 6086 12724 6092 12736
rect 6144 12724 6150 12776
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12764 9367 12767
rect 9398 12764 9404 12776
rect 9355 12736 9404 12764
rect 9355 12733 9367 12736
rect 9309 12727 9367 12733
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 11238 12724 11244 12776
rect 11296 12764 11302 12776
rect 11368 12767 11426 12773
rect 11368 12764 11380 12767
rect 11296 12736 11380 12764
rect 11296 12724 11302 12736
rect 11368 12733 11380 12736
rect 11414 12764 11426 12767
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 11414 12736 11805 12764
rect 11414 12733 11426 12736
rect 11368 12727 11426 12733
rect 11793 12733 11805 12736
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 17126 12724 17132 12776
rect 17184 12764 17190 12776
rect 17678 12764 17684 12776
rect 17184 12736 17684 12764
rect 17184 12724 17190 12736
rect 17678 12724 17684 12736
rect 17736 12724 17742 12776
rect 18084 12767 18142 12773
rect 18084 12733 18096 12767
rect 18130 12733 18142 12767
rect 18084 12727 18142 12733
rect 2222 12656 2228 12708
rect 2280 12696 2286 12708
rect 2774 12696 2780 12708
rect 2280 12668 2325 12696
rect 2735 12668 2780 12696
rect 2280 12656 2286 12668
rect 2774 12656 2780 12668
rect 2832 12656 2838 12708
rect 3786 12696 3792 12708
rect 3699 12668 3792 12696
rect 3786 12656 3792 12668
rect 3844 12696 3850 12708
rect 4243 12699 4301 12705
rect 4243 12696 4255 12699
rect 3844 12668 4255 12696
rect 3844 12656 3850 12668
rect 4243 12665 4255 12668
rect 4289 12696 4301 12699
rect 6638 12696 6644 12708
rect 4289 12668 6644 12696
rect 4289 12665 4301 12668
rect 4243 12659 4301 12665
rect 6638 12656 6644 12668
rect 6696 12696 6702 12708
rect 7187 12699 7245 12705
rect 7187 12696 7199 12699
rect 6696 12668 7199 12696
rect 6696 12656 6702 12668
rect 7187 12665 7199 12668
rect 7233 12696 7245 12699
rect 9217 12699 9275 12705
rect 9217 12696 9229 12699
rect 7233 12668 9229 12696
rect 7233 12665 7245 12668
rect 7187 12659 7245 12665
rect 9217 12665 9229 12668
rect 9263 12696 9275 12699
rect 12618 12696 12624 12708
rect 9263 12668 9674 12696
rect 12579 12668 12624 12696
rect 9263 12665 9275 12668
rect 9217 12659 9275 12665
rect 9646 12640 9674 12668
rect 12618 12656 12624 12668
rect 12676 12656 12682 12708
rect 14182 12656 14188 12708
rect 14240 12696 14246 12708
rect 15749 12699 15807 12705
rect 14240 12668 14285 12696
rect 14240 12656 14246 12668
rect 15749 12665 15761 12699
rect 15795 12665 15807 12699
rect 15749 12659 15807 12665
rect 1765 12631 1823 12637
rect 1765 12597 1777 12631
rect 1811 12628 1823 12631
rect 1854 12628 1860 12640
rect 1811 12600 1860 12628
rect 1811 12597 1823 12600
rect 1765 12591 1823 12597
rect 1854 12588 1860 12600
rect 1912 12628 1918 12640
rect 2958 12628 2964 12640
rect 1912 12600 2964 12628
rect 1912 12588 1918 12600
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 9646 12628 9680 12640
rect 9635 12600 9680 12628
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 10229 12631 10287 12637
rect 10229 12597 10241 12631
rect 10275 12628 10287 12631
rect 10318 12628 10324 12640
rect 10275 12600 10324 12628
rect 10275 12597 10287 12600
rect 10229 12591 10287 12597
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 11471 12631 11529 12637
rect 11471 12597 11483 12631
rect 11517 12628 11529 12631
rect 13446 12628 13452 12640
rect 11517 12600 13452 12628
rect 11517 12597 11529 12600
rect 11471 12591 11529 12597
rect 13446 12588 13452 12600
rect 13504 12588 13510 12640
rect 13541 12631 13599 12637
rect 13541 12597 13553 12631
rect 13587 12628 13599 12631
rect 13722 12628 13728 12640
rect 13587 12600 13728 12628
rect 13587 12597 13599 12600
rect 13541 12591 13599 12597
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 15470 12628 15476 12640
rect 15431 12600 15476 12628
rect 15470 12588 15476 12600
rect 15528 12628 15534 12640
rect 15764 12628 15792 12659
rect 16114 12656 16120 12708
rect 16172 12696 16178 12708
rect 18099 12696 18127 12727
rect 18966 12724 18972 12776
rect 19024 12764 19030 12776
rect 19128 12767 19186 12773
rect 19128 12764 19140 12767
rect 19024 12736 19140 12764
rect 19024 12724 19030 12736
rect 19128 12733 19140 12736
rect 19174 12764 19186 12767
rect 19174 12736 19932 12764
rect 19174 12733 19186 12736
rect 19128 12727 19186 12733
rect 18506 12696 18512 12708
rect 16172 12668 18512 12696
rect 16172 12656 16178 12668
rect 18506 12656 18512 12668
rect 18564 12656 18570 12708
rect 19904 12640 19932 12736
rect 17218 12628 17224 12640
rect 15528 12600 15792 12628
rect 17179 12600 17224 12628
rect 15528 12588 15534 12600
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 18187 12631 18245 12637
rect 18187 12628 18199 12631
rect 17460 12600 18199 12628
rect 17460 12588 17466 12600
rect 18187 12597 18199 12600
rect 18233 12597 18245 12631
rect 18187 12591 18245 12597
rect 18782 12588 18788 12640
rect 18840 12628 18846 12640
rect 18877 12631 18935 12637
rect 18877 12628 18889 12631
rect 18840 12600 18889 12628
rect 18840 12588 18846 12600
rect 18877 12597 18889 12600
rect 18923 12597 18935 12631
rect 18877 12591 18935 12597
rect 18966 12588 18972 12640
rect 19024 12628 19030 12640
rect 19199 12631 19257 12637
rect 19199 12628 19211 12631
rect 19024 12600 19211 12628
rect 19024 12588 19030 12600
rect 19199 12597 19211 12600
rect 19245 12597 19257 12631
rect 19886 12628 19892 12640
rect 19847 12600 19892 12628
rect 19199 12591 19257 12597
rect 19886 12588 19892 12600
rect 19944 12588 19950 12640
rect 1104 12538 20884 12560
rect 1104 12486 8315 12538
rect 8367 12486 8379 12538
rect 8431 12486 8443 12538
rect 8495 12486 8507 12538
rect 8559 12486 15648 12538
rect 15700 12486 15712 12538
rect 15764 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 20884 12538
rect 1104 12464 20884 12486
rect 1854 12424 1860 12436
rect 1815 12396 1860 12424
rect 1854 12384 1860 12396
rect 1912 12384 1918 12436
rect 2222 12384 2228 12436
rect 2280 12424 2286 12436
rect 2409 12427 2467 12433
rect 2409 12424 2421 12427
rect 2280 12396 2421 12424
rect 2280 12384 2286 12396
rect 2409 12393 2421 12396
rect 2455 12393 2467 12427
rect 2409 12387 2467 12393
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 2958 12424 2964 12436
rect 2823 12396 2964 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 2958 12384 2964 12396
rect 3016 12424 3022 12436
rect 3786 12424 3792 12436
rect 3016 12396 3792 12424
rect 3016 12384 3022 12396
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 4157 12427 4215 12433
rect 4157 12424 4169 12427
rect 4120 12396 4169 12424
rect 4120 12384 4126 12396
rect 4157 12393 4169 12396
rect 4203 12393 4215 12427
rect 6638 12424 6644 12436
rect 6599 12396 6644 12424
rect 4157 12387 4215 12393
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 7469 12427 7527 12433
rect 7469 12424 7481 12427
rect 7340 12396 7481 12424
rect 7340 12384 7346 12396
rect 7469 12393 7481 12396
rect 7515 12393 7527 12427
rect 7469 12387 7527 12393
rect 10689 12427 10747 12433
rect 10689 12393 10701 12427
rect 10735 12424 10747 12427
rect 10870 12424 10876 12436
rect 10735 12396 10876 12424
rect 10735 12393 10747 12396
rect 10689 12387 10747 12393
rect 10870 12384 10876 12396
rect 10928 12424 10934 12436
rect 12345 12427 12403 12433
rect 12345 12424 12357 12427
rect 10928 12396 12357 12424
rect 10928 12384 10934 12396
rect 12345 12393 12357 12396
rect 12391 12424 12403 12427
rect 12618 12424 12624 12436
rect 12391 12396 12624 12424
rect 12391 12393 12403 12396
rect 12345 12387 12403 12393
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 12805 12427 12863 12433
rect 12805 12393 12817 12427
rect 12851 12424 12863 12427
rect 18509 12427 18567 12433
rect 18509 12424 18521 12427
rect 12851 12396 18521 12424
rect 12851 12393 12863 12396
rect 12805 12387 12863 12393
rect 8110 12356 8116 12368
rect 7852 12328 8116 12356
rect 4062 12288 4068 12300
rect 4023 12260 4068 12288
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 4525 12291 4583 12297
rect 4525 12288 4537 12291
rect 4212 12260 4537 12288
rect 4212 12248 4218 12260
rect 4525 12257 4537 12260
rect 4571 12257 4583 12291
rect 4525 12251 4583 12257
rect 5994 12248 6000 12300
rect 6052 12288 6058 12300
rect 6273 12291 6331 12297
rect 6273 12288 6285 12291
rect 6052 12260 6285 12288
rect 6052 12248 6058 12260
rect 6273 12257 6285 12260
rect 6319 12288 6331 12291
rect 6730 12288 6736 12300
rect 6319 12260 6736 12288
rect 6319 12257 6331 12260
rect 6273 12251 6331 12257
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 7193 12291 7251 12297
rect 7193 12257 7205 12291
rect 7239 12288 7251 12291
rect 7852 12288 7880 12328
rect 8110 12316 8116 12328
rect 8168 12356 8174 12368
rect 8205 12359 8263 12365
rect 8205 12356 8217 12359
rect 8168 12328 8217 12356
rect 8168 12316 8174 12328
rect 8205 12325 8217 12328
rect 8251 12325 8263 12359
rect 8754 12356 8760 12368
rect 8715 12328 8760 12356
rect 8205 12319 8263 12325
rect 8754 12316 8760 12328
rect 8812 12316 8818 12368
rect 9674 12316 9680 12368
rect 9732 12356 9738 12368
rect 10090 12359 10148 12365
rect 10090 12356 10102 12359
rect 9732 12328 10102 12356
rect 9732 12316 9738 12328
rect 10090 12325 10102 12328
rect 10136 12325 10148 12359
rect 10090 12319 10148 12325
rect 11057 12359 11115 12365
rect 11057 12325 11069 12359
rect 11103 12356 11115 12359
rect 11146 12356 11152 12368
rect 11103 12328 11152 12356
rect 11103 12325 11115 12328
rect 11057 12319 11115 12325
rect 11146 12316 11152 12328
rect 11204 12316 11210 12368
rect 11422 12356 11428 12368
rect 11383 12328 11428 12356
rect 11422 12316 11428 12328
rect 11480 12316 11486 12368
rect 11882 12288 11888 12300
rect 7239 12260 7880 12288
rect 11843 12260 11888 12288
rect 7239 12257 7251 12260
rect 7193 12251 7251 12257
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 12912 12297 12940 12396
rect 18509 12393 18521 12396
rect 18555 12393 18567 12427
rect 18509 12387 18567 12393
rect 13259 12359 13317 12365
rect 13259 12325 13271 12359
rect 13305 12356 13317 12359
rect 13722 12356 13728 12368
rect 13305 12328 13728 12356
rect 13305 12325 13317 12328
rect 13259 12319 13317 12325
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 15470 12356 15476 12368
rect 13832 12328 15476 12356
rect 13832 12297 13860 12328
rect 15470 12316 15476 12328
rect 15528 12316 15534 12368
rect 16022 12356 16028 12368
rect 15983 12328 16028 12356
rect 16022 12316 16028 12328
rect 16080 12316 16086 12368
rect 16390 12356 16396 12368
rect 16303 12328 16396 12356
rect 16390 12316 16396 12328
rect 16448 12356 16454 12368
rect 17402 12356 17408 12368
rect 16448 12328 17408 12356
rect 16448 12316 16454 12328
rect 17402 12316 17408 12328
rect 17460 12316 17466 12368
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12257 12955 12291
rect 12897 12251 12955 12257
rect 13817 12291 13875 12297
rect 13817 12257 13829 12291
rect 13863 12257 13875 12291
rect 17126 12288 17132 12300
rect 17087 12260 17132 12288
rect 13817 12251 13875 12257
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 17313 12291 17371 12297
rect 17313 12288 17325 12291
rect 17276 12260 17325 12288
rect 17276 12248 17282 12260
rect 17313 12257 17325 12260
rect 17359 12257 17371 12291
rect 18414 12288 18420 12300
rect 18375 12260 18420 12288
rect 17313 12251 17371 12257
rect 18414 12248 18420 12260
rect 18472 12248 18478 12300
rect 18598 12248 18604 12300
rect 18656 12288 18662 12300
rect 18877 12291 18935 12297
rect 18877 12288 18889 12291
rect 18656 12260 18889 12288
rect 18656 12248 18662 12260
rect 18877 12257 18889 12260
rect 18923 12257 18935 12291
rect 18877 12251 18935 12257
rect 1489 12223 1547 12229
rect 1489 12189 1501 12223
rect 1535 12220 1547 12223
rect 2130 12220 2136 12232
rect 1535 12192 2136 12220
rect 1535 12189 1547 12192
rect 1489 12183 1547 12189
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12220 8171 12223
rect 8202 12220 8208 12232
rect 8159 12192 8208 12220
rect 8159 12189 8171 12192
rect 8113 12183 8171 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 9769 12223 9827 12229
rect 9769 12189 9781 12223
rect 9815 12220 9827 12223
rect 11238 12220 11244 12232
rect 9815 12192 11244 12220
rect 9815 12189 9827 12192
rect 9769 12183 9827 12189
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 13446 12180 13452 12232
rect 13504 12220 13510 12232
rect 14642 12220 14648 12232
rect 13504 12192 14648 12220
rect 13504 12180 13510 12192
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 15028 12192 15393 12220
rect 7190 12112 7196 12164
rect 7248 12152 7254 12164
rect 7929 12155 7987 12161
rect 7929 12152 7941 12155
rect 7248 12124 7941 12152
rect 7248 12112 7254 12124
rect 7929 12121 7941 12124
rect 7975 12152 7987 12155
rect 10962 12152 10968 12164
rect 7975 12124 10968 12152
rect 7975 12121 7987 12124
rect 7929 12115 7987 12121
rect 10962 12112 10968 12124
rect 11020 12112 11026 12164
rect 15028 12161 15056 12192
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 17402 12220 17408 12232
rect 17363 12192 17408 12220
rect 15381 12183 15439 12189
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 12023 12155 12081 12161
rect 12023 12121 12035 12155
rect 12069 12152 12081 12155
rect 15013 12155 15071 12161
rect 15013 12152 15025 12155
rect 12069 12124 15025 12152
rect 12069 12121 12081 12124
rect 12023 12115 12081 12121
rect 15013 12121 15025 12124
rect 15059 12121 15071 12155
rect 15013 12115 15071 12121
rect 2866 12044 2872 12096
rect 2924 12084 2930 12096
rect 3053 12087 3111 12093
rect 3053 12084 3065 12087
rect 2924 12056 3065 12084
rect 2924 12044 2930 12056
rect 3053 12053 3065 12056
rect 3099 12053 3111 12087
rect 3053 12047 3111 12053
rect 4522 12044 4528 12096
rect 4580 12084 4586 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 4580 12056 5089 12084
rect 4580 12044 4586 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 9398 12084 9404 12096
rect 9359 12056 9404 12084
rect 5077 12047 5135 12053
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 13722 12044 13728 12096
rect 13780 12084 13786 12096
rect 14093 12087 14151 12093
rect 14093 12084 14105 12087
rect 13780 12056 14105 12084
rect 13780 12044 13786 12056
rect 14093 12053 14105 12056
rect 14139 12053 14151 12087
rect 14093 12047 14151 12053
rect 14826 12044 14832 12096
rect 14884 12084 14890 12096
rect 18782 12084 18788 12096
rect 14884 12056 18788 12084
rect 14884 12044 14890 12056
rect 18782 12044 18788 12056
rect 18840 12044 18846 12096
rect 1104 11994 20884 12016
rect 1104 11942 4648 11994
rect 4700 11942 4712 11994
rect 4764 11942 4776 11994
rect 4828 11942 4840 11994
rect 4892 11942 11982 11994
rect 12034 11942 12046 11994
rect 12098 11942 12110 11994
rect 12162 11942 12174 11994
rect 12226 11942 19315 11994
rect 19367 11942 19379 11994
rect 19431 11942 19443 11994
rect 19495 11942 19507 11994
rect 19559 11942 20884 11994
rect 1104 11920 20884 11942
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 5994 11880 6000 11892
rect 4212 11852 4257 11880
rect 5955 11852 6000 11880
rect 4212 11840 4218 11852
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 6365 11883 6423 11889
rect 6365 11849 6377 11883
rect 6411 11880 6423 11883
rect 6638 11880 6644 11892
rect 6411 11852 6644 11880
rect 6411 11849 6423 11852
rect 6365 11843 6423 11849
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 8110 11880 8116 11892
rect 8071 11852 8116 11880
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 8202 11840 8208 11892
rect 8260 11880 8266 11892
rect 8481 11883 8539 11889
rect 8481 11880 8493 11883
rect 8260 11852 8493 11880
rect 8260 11840 8266 11852
rect 8481 11849 8493 11852
rect 8527 11849 8539 11883
rect 8481 11843 8539 11849
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 15286 11880 15292 11892
rect 9824 11852 15292 11880
rect 9824 11840 9830 11852
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 16209 11883 16267 11889
rect 16209 11880 16221 11883
rect 15528 11852 16221 11880
rect 15528 11840 15534 11852
rect 16209 11849 16221 11852
rect 16255 11849 16267 11883
rect 16209 11843 16267 11849
rect 16899 11883 16957 11889
rect 16899 11849 16911 11883
rect 16945 11880 16957 11883
rect 17862 11880 17868 11892
rect 16945 11852 17868 11880
rect 16945 11849 16957 11852
rect 16899 11843 16957 11849
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 18598 11880 18604 11892
rect 18559 11852 18604 11880
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 19245 11883 19303 11889
rect 19245 11849 19257 11883
rect 19291 11880 19303 11883
rect 20070 11880 20076 11892
rect 19291 11852 20076 11880
rect 19291 11849 19303 11852
rect 19245 11843 19303 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 11146 11812 11152 11824
rect 10244 11784 11152 11812
rect 4982 11744 4988 11756
rect 4943 11716 4988 11744
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 7190 11744 7196 11756
rect 7151 11716 7196 11744
rect 7190 11704 7196 11716
rect 7248 11704 7254 11756
rect 7834 11744 7840 11756
rect 7795 11716 7840 11744
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 10244 11753 10272 11784
rect 11146 11772 11152 11784
rect 11204 11772 11210 11824
rect 11238 11772 11244 11824
rect 11296 11812 11302 11824
rect 17402 11812 17408 11824
rect 11296 11784 17408 11812
rect 11296 11772 11302 11784
rect 17402 11772 17408 11784
rect 17460 11772 17466 11824
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11744 10931 11747
rect 11054 11744 11060 11756
rect 10919 11716 11060 11744
rect 10919 11713 10931 11716
rect 10873 11707 10931 11713
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 11882 11744 11888 11756
rect 11843 11716 11888 11744
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 15286 11744 15292 11756
rect 12912 11716 15292 11744
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11676 1458 11688
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1452 11648 1961 11676
rect 1452 11636 1458 11648
rect 1949 11645 1961 11648
rect 1995 11645 2007 11679
rect 1949 11639 2007 11645
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 2866 11676 2872 11688
rect 2731 11648 2872 11676
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 8700 11679 8758 11685
rect 8700 11676 8712 11679
rect 8260 11648 8712 11676
rect 8260 11636 8266 11648
rect 8700 11645 8712 11648
rect 8746 11676 8758 11679
rect 9125 11679 9183 11685
rect 9125 11676 9137 11679
rect 8746 11648 9137 11676
rect 8746 11645 8758 11648
rect 8700 11639 8758 11645
rect 9125 11645 9137 11648
rect 9171 11676 9183 11679
rect 9490 11676 9496 11688
rect 9171 11648 9496 11676
rect 9171 11645 9183 11648
rect 9125 11639 9183 11645
rect 9490 11636 9496 11648
rect 9548 11636 9554 11688
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 12912 11685 12940 11716
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 15378 11704 15384 11756
rect 15436 11744 15442 11756
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 15436 11716 18061 11744
rect 15436 11704 15442 11716
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 12472 11679 12530 11685
rect 12472 11676 12484 11679
rect 12400 11648 12484 11676
rect 12400 11636 12406 11648
rect 12472 11645 12484 11648
rect 12518 11676 12530 11679
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12518 11648 12909 11676
rect 12518 11645 12530 11648
rect 12472 11639 12530 11645
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 13446 11676 13452 11688
rect 13407 11648 13452 11676
rect 12897 11639 12955 11645
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 15105 11679 15163 11685
rect 15105 11676 15117 11679
rect 13556 11648 15117 11676
rect 4522 11608 4528 11620
rect 4483 11580 4528 11608
rect 4522 11568 4528 11580
rect 4580 11568 4586 11620
rect 4617 11611 4675 11617
rect 4617 11577 4629 11611
rect 4663 11577 4675 11611
rect 4617 11571 4675 11577
rect 14 11500 20 11552
rect 72 11540 78 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 72 11512 1593 11540
rect 72 11500 78 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 1581 11503 1639 11509
rect 2409 11543 2467 11549
rect 2409 11509 2421 11543
rect 2455 11540 2467 11543
rect 2498 11540 2504 11552
rect 2455 11512 2504 11540
rect 2455 11509 2467 11512
rect 2409 11503 2467 11509
rect 2498 11500 2504 11512
rect 2556 11540 2562 11552
rect 2958 11540 2964 11552
rect 2556 11512 2964 11540
rect 2556 11500 2562 11512
rect 2958 11500 2964 11512
rect 3016 11540 3022 11552
rect 3053 11543 3111 11549
rect 3053 11540 3065 11543
rect 3016 11512 3065 11540
rect 3016 11500 3022 11512
rect 3053 11509 3065 11512
rect 3099 11509 3111 11543
rect 3053 11503 3111 11509
rect 3605 11543 3663 11549
rect 3605 11509 3617 11543
rect 3651 11540 3663 11543
rect 4632 11540 4660 11571
rect 7282 11568 7288 11620
rect 7340 11608 7346 11620
rect 7340 11580 7385 11608
rect 7340 11568 7346 11580
rect 10318 11568 10324 11620
rect 10376 11608 10382 11620
rect 10376 11580 10421 11608
rect 10376 11568 10382 11580
rect 10502 11568 10508 11620
rect 10560 11608 10566 11620
rect 12575 11611 12633 11617
rect 12575 11608 12587 11611
rect 10560 11580 12587 11608
rect 10560 11568 10566 11580
rect 12575 11577 12587 11580
rect 12621 11577 12633 11611
rect 13556 11608 13584 11648
rect 15105 11645 15117 11648
rect 15151 11676 15163 11679
rect 15194 11676 15200 11688
rect 15151 11648 15200 11676
rect 15151 11645 15163 11648
rect 15105 11639 15163 11645
rect 15194 11636 15200 11648
rect 15252 11636 15258 11688
rect 15657 11679 15715 11685
rect 15657 11676 15669 11679
rect 15304 11648 15669 11676
rect 13722 11608 13728 11620
rect 12575 11571 12633 11577
rect 12728 11580 13584 11608
rect 13680 11580 13728 11608
rect 5445 11543 5503 11549
rect 5445 11540 5457 11543
rect 3651 11512 5457 11540
rect 3651 11509 3663 11512
rect 3605 11503 3663 11509
rect 5445 11509 5457 11512
rect 5491 11509 5503 11543
rect 5445 11503 5503 11509
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 8803 11543 8861 11549
rect 8803 11540 8815 11543
rect 6420 11512 8815 11540
rect 6420 11500 6426 11512
rect 8803 11509 8815 11512
rect 8849 11509 8861 11543
rect 8803 11503 8861 11509
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 9732 11512 9781 11540
rect 9732 11500 9738 11512
rect 9769 11509 9781 11512
rect 9815 11509 9827 11543
rect 9769 11503 9827 11509
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 12728 11540 12756 11580
rect 13722 11568 13728 11580
rect 13780 11617 13786 11620
rect 13780 11611 13828 11617
rect 13780 11577 13782 11611
rect 13816 11577 13828 11611
rect 15304 11608 15332 11648
rect 15657 11645 15669 11648
rect 15703 11645 15715 11679
rect 16796 11679 16854 11685
rect 16796 11676 16808 11679
rect 15657 11639 15715 11645
rect 16592 11648 16808 11676
rect 13780 11571 13828 11577
rect 14660 11580 15332 11608
rect 13780 11568 13813 11571
rect 13262 11540 13268 11552
rect 10652 11512 12756 11540
rect 13223 11512 13268 11540
rect 10652 11500 10658 11512
rect 13262 11500 13268 11512
rect 13320 11540 13326 11552
rect 13785 11540 13813 11568
rect 14660 11552 14688 11580
rect 16022 11568 16028 11620
rect 16080 11608 16086 11620
rect 16592 11617 16620 11648
rect 16796 11645 16808 11648
rect 16842 11645 16854 11679
rect 16796 11639 16854 11645
rect 17034 11636 17040 11688
rect 17092 11676 17098 11688
rect 17218 11676 17224 11688
rect 17092 11648 17224 11676
rect 17092 11636 17098 11648
rect 17218 11636 17224 11648
rect 17276 11676 17282 11688
rect 17589 11679 17647 11685
rect 17589 11676 17601 11679
rect 17276 11648 17601 11676
rect 17276 11636 17282 11648
rect 17589 11645 17601 11648
rect 17635 11645 17647 11679
rect 17589 11639 17647 11645
rect 18506 11636 18512 11688
rect 18564 11676 18570 11688
rect 19061 11679 19119 11685
rect 19061 11676 19073 11679
rect 18564 11648 19073 11676
rect 18564 11636 18570 11648
rect 19061 11645 19073 11648
rect 19107 11676 19119 11679
rect 19613 11679 19671 11685
rect 19613 11676 19625 11679
rect 19107 11648 19625 11676
rect 19107 11645 19119 11648
rect 19061 11639 19119 11645
rect 19613 11645 19625 11648
rect 19659 11645 19671 11679
rect 19613 11639 19671 11645
rect 16577 11611 16635 11617
rect 16577 11608 16589 11611
rect 16080 11580 16589 11608
rect 16080 11568 16086 11580
rect 16577 11577 16589 11580
rect 16623 11577 16635 11611
rect 16577 11571 16635 11577
rect 17126 11568 17132 11620
rect 17184 11608 17190 11620
rect 17313 11611 17371 11617
rect 17313 11608 17325 11611
rect 17184 11580 17325 11608
rect 17184 11568 17190 11580
rect 17313 11577 17325 11580
rect 17359 11608 17371 11611
rect 18230 11608 18236 11620
rect 17359 11580 18236 11608
rect 17359 11577 17371 11580
rect 17313 11571 17371 11577
rect 18230 11568 18236 11580
rect 18288 11568 18294 11620
rect 14366 11540 14372 11552
rect 13320 11512 13813 11540
rect 14327 11512 14372 11540
rect 13320 11500 13326 11512
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 14642 11540 14648 11552
rect 14603 11512 14648 11540
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 15289 11543 15347 11549
rect 15289 11540 15301 11543
rect 15160 11512 15301 11540
rect 15160 11500 15166 11512
rect 15289 11509 15301 11512
rect 15335 11509 15347 11543
rect 15289 11503 15347 11509
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18414 11540 18420 11552
rect 18104 11512 18420 11540
rect 18104 11500 18110 11512
rect 18414 11500 18420 11512
rect 18472 11540 18478 11552
rect 18877 11543 18935 11549
rect 18877 11540 18889 11543
rect 18472 11512 18889 11540
rect 18472 11500 18478 11512
rect 18877 11509 18889 11512
rect 18923 11509 18935 11543
rect 18877 11503 18935 11509
rect 1104 11450 20884 11472
rect 1104 11398 8315 11450
rect 8367 11398 8379 11450
rect 8431 11398 8443 11450
rect 8495 11398 8507 11450
rect 8559 11398 15648 11450
rect 15700 11398 15712 11450
rect 15764 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 20884 11450
rect 1104 11376 20884 11398
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4157 11339 4215 11345
rect 4157 11336 4169 11339
rect 4120 11308 4169 11336
rect 4120 11296 4126 11308
rect 4157 11305 4169 11308
rect 4203 11305 4215 11339
rect 5074 11336 5080 11348
rect 5035 11308 5080 11336
rect 4157 11299 4215 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 7469 11339 7527 11345
rect 7469 11336 7481 11339
rect 7340 11308 7481 11336
rect 7340 11296 7346 11308
rect 7469 11305 7481 11308
rect 7515 11305 7527 11339
rect 7469 11299 7527 11305
rect 7834 11296 7840 11348
rect 7892 11336 7898 11348
rect 10229 11339 10287 11345
rect 7892 11308 8800 11336
rect 7892 11296 7898 11308
rect 2403 11271 2461 11277
rect 2403 11237 2415 11271
rect 2449 11268 2461 11271
rect 2498 11268 2504 11280
rect 2449 11240 2504 11268
rect 2449 11237 2461 11240
rect 2403 11231 2461 11237
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 6638 11268 6644 11280
rect 5644 11240 6644 11268
rect 5350 11160 5356 11212
rect 5408 11200 5414 11212
rect 5644 11209 5672 11240
rect 6638 11228 6644 11240
rect 6696 11228 6702 11280
rect 8110 11228 8116 11280
rect 8168 11268 8174 11280
rect 8772 11277 8800 11308
rect 10229 11305 10241 11339
rect 10275 11336 10287 11339
rect 10318 11336 10324 11348
rect 10275 11308 10324 11336
rect 10275 11305 10287 11308
rect 10229 11299 10287 11305
rect 10318 11296 10324 11308
rect 10376 11336 10382 11348
rect 12802 11336 12808 11348
rect 10376 11308 10548 11336
rect 10376 11296 10382 11308
rect 8205 11271 8263 11277
rect 8205 11268 8217 11271
rect 8168 11240 8217 11268
rect 8168 11228 8174 11240
rect 8205 11237 8217 11240
rect 8251 11237 8263 11271
rect 8205 11231 8263 11237
rect 8757 11271 8815 11277
rect 8757 11237 8769 11271
rect 8803 11237 8815 11271
rect 10410 11268 10416 11280
rect 10371 11240 10416 11268
rect 8757 11231 8815 11237
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 10520 11277 10548 11308
rect 11415 11308 12808 11336
rect 10505 11271 10563 11277
rect 10505 11237 10517 11271
rect 10551 11237 10563 11271
rect 10505 11231 10563 11237
rect 11057 11271 11115 11277
rect 11057 11237 11069 11271
rect 11103 11268 11115 11271
rect 11415 11268 11443 11308
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 13446 11336 13452 11348
rect 13035 11308 13452 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 13446 11296 13452 11308
rect 13504 11336 13510 11348
rect 16945 11339 17003 11345
rect 16945 11336 16957 11339
rect 13504 11308 16957 11336
rect 13504 11296 13510 11308
rect 16945 11305 16957 11308
rect 16991 11305 17003 11339
rect 16945 11299 17003 11305
rect 11103 11240 11443 11268
rect 11103 11237 11115 11240
rect 11057 11231 11115 11237
rect 11790 11228 11796 11280
rect 11848 11268 11854 11280
rect 12069 11271 12127 11277
rect 12069 11268 12081 11271
rect 11848 11240 12081 11268
rect 11848 11228 11854 11240
rect 12069 11237 12081 11240
rect 12115 11237 12127 11271
rect 12069 11231 12127 11237
rect 13262 11228 13268 11280
rect 13320 11268 13326 11280
rect 13770 11271 13828 11277
rect 13770 11268 13782 11271
rect 13320 11240 13782 11268
rect 13320 11228 13326 11240
rect 13770 11237 13782 11240
rect 13816 11237 13828 11271
rect 13770 11231 13828 11237
rect 14366 11228 14372 11280
rect 14424 11268 14430 11280
rect 15010 11268 15016 11280
rect 14424 11240 15016 11268
rect 14424 11228 14430 11240
rect 15010 11228 15016 11240
rect 15068 11268 15074 11280
rect 15473 11271 15531 11277
rect 15473 11268 15485 11271
rect 15068 11240 15485 11268
rect 15068 11228 15074 11240
rect 15473 11237 15485 11240
rect 15519 11237 15531 11271
rect 15473 11231 15531 11237
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 5408 11172 5641 11200
rect 5408 11160 5414 11172
rect 5629 11169 5641 11172
rect 5675 11169 5687 11203
rect 5629 11163 5687 11169
rect 16114 11160 16120 11212
rect 16172 11200 16178 11212
rect 16482 11200 16488 11212
rect 16172 11172 16488 11200
rect 16172 11160 16178 11172
rect 16482 11160 16488 11172
rect 16540 11200 16546 11212
rect 16853 11203 16911 11209
rect 16853 11200 16865 11203
rect 16540 11172 16865 11200
rect 16540 11160 16546 11172
rect 16853 11169 16865 11172
rect 16899 11169 16911 11203
rect 17310 11200 17316 11212
rect 17271 11172 17316 11200
rect 16853 11163 16911 11169
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 19061 11203 19119 11209
rect 19061 11169 19073 11203
rect 19107 11169 19119 11203
rect 19061 11163 19119 11169
rect 2041 11135 2099 11141
rect 2041 11132 2053 11135
rect 1872 11104 2053 11132
rect 1670 10956 1676 11008
rect 1728 10996 1734 11008
rect 1872 11005 1900 11104
rect 2041 11101 2053 11104
rect 2087 11101 2099 11135
rect 2041 11095 2099 11101
rect 2314 11092 2320 11144
rect 2372 11132 2378 11144
rect 2774 11132 2780 11144
rect 2372 11104 2780 11132
rect 2372 11092 2378 11104
rect 2774 11092 2780 11104
rect 2832 11132 2838 11144
rect 3605 11135 3663 11141
rect 3605 11132 3617 11135
rect 2832 11104 3617 11132
rect 2832 11092 2838 11104
rect 3605 11101 3617 11104
rect 3651 11101 3663 11135
rect 3605 11095 3663 11101
rect 2130 11024 2136 11076
rect 2188 11064 2194 11076
rect 3237 11067 3295 11073
rect 3237 11064 3249 11067
rect 2188 11036 3249 11064
rect 2188 11024 2194 11036
rect 3237 11033 3249 11036
rect 3283 11033 3295 11067
rect 3620 11064 3648 11095
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4709 11135 4767 11141
rect 4709 11132 4721 11135
rect 4120 11104 4721 11132
rect 4120 11092 4126 11104
rect 4709 11101 4721 11104
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 6365 11135 6423 11141
rect 6365 11101 6377 11135
rect 6411 11132 6423 11135
rect 6546 11132 6552 11144
rect 6411 11104 6552 11132
rect 6411 11101 6423 11104
rect 6365 11095 6423 11101
rect 6546 11092 6552 11104
rect 6604 11092 6610 11144
rect 6822 11132 6828 11144
rect 6783 11104 6828 11132
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11132 7987 11135
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 7975 11104 8125 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8113 11101 8125 11104
rect 8159 11132 8171 11135
rect 8754 11132 8760 11144
rect 8159 11104 8760 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 8754 11092 8760 11104
rect 8812 11092 8818 11144
rect 11977 11135 12035 11141
rect 11977 11101 11989 11135
rect 12023 11132 12035 11135
rect 12434 11132 12440 11144
rect 12023 11104 12440 11132
rect 12023 11101 12035 11104
rect 11977 11095 12035 11101
rect 12434 11092 12440 11104
rect 12492 11132 12498 11144
rect 13446 11132 13452 11144
rect 12492 11104 12756 11132
rect 13407 11104 13452 11132
rect 12492 11092 12498 11104
rect 4982 11064 4988 11076
rect 3620 11036 4988 11064
rect 3237 11027 3295 11033
rect 4982 11024 4988 11036
rect 5040 11024 5046 11076
rect 6914 11064 6920 11076
rect 5276 11036 6920 11064
rect 1857 10999 1915 11005
rect 1857 10996 1869 10999
rect 1728 10968 1869 10996
rect 1728 10956 1734 10968
rect 1857 10965 1869 10968
rect 1903 10965 1915 10999
rect 2958 10996 2964 11008
rect 2919 10968 2964 10996
rect 1857 10959 1915 10965
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 4157 10999 4215 11005
rect 4157 10965 4169 10999
rect 4203 10996 4215 10999
rect 4341 10999 4399 11005
rect 4341 10996 4353 10999
rect 4203 10968 4353 10996
rect 4203 10965 4215 10968
rect 4157 10959 4215 10965
rect 4341 10965 4353 10968
rect 4387 10996 4399 10999
rect 5276 10996 5304 11036
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 11514 11024 11520 11076
rect 11572 11064 11578 11076
rect 12529 11067 12587 11073
rect 12529 11064 12541 11067
rect 11572 11036 12541 11064
rect 11572 11024 11578 11036
rect 12529 11033 12541 11036
rect 12575 11033 12587 11067
rect 12728 11064 12756 11104
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 15378 11132 15384 11144
rect 15339 11104 15384 11132
rect 15378 11092 15384 11104
rect 15436 11092 15442 11144
rect 16022 11132 16028 11144
rect 15983 11104 16028 11132
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 14458 11064 14464 11076
rect 12728 11036 14464 11064
rect 12529 11027 12587 11033
rect 14458 11024 14464 11036
rect 14516 11024 14522 11076
rect 15286 11024 15292 11076
rect 15344 11064 15350 11076
rect 19076 11064 19104 11163
rect 19150 11064 19156 11076
rect 15344 11036 19156 11064
rect 15344 11024 15350 11036
rect 19150 11024 19156 11036
rect 19208 11024 19214 11076
rect 5902 10996 5908 11008
rect 4387 10968 5304 10996
rect 5863 10968 5908 10996
rect 4387 10965 4399 10968
rect 4341 10959 4399 10965
rect 5902 10956 5908 10968
rect 5960 10956 5966 11008
rect 13354 10996 13360 11008
rect 13315 10968 13360 10996
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 14366 10996 14372 11008
rect 14327 10968 14372 10996
rect 14366 10956 14372 10968
rect 14424 10956 14430 11008
rect 15105 10999 15163 11005
rect 15105 10965 15117 10999
rect 15151 10996 15163 10999
rect 15194 10996 15200 11008
rect 15151 10968 15200 10996
rect 15151 10965 15163 10968
rect 15105 10959 15163 10965
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 19245 10999 19303 11005
rect 19245 10965 19257 10999
rect 19291 10996 19303 10999
rect 20438 10996 20444 11008
rect 19291 10968 20444 10996
rect 19291 10965 19303 10968
rect 19245 10959 19303 10965
rect 20438 10956 20444 10968
rect 20496 10956 20502 11008
rect 1104 10906 20884 10928
rect 1104 10854 4648 10906
rect 4700 10854 4712 10906
rect 4764 10854 4776 10906
rect 4828 10854 4840 10906
rect 4892 10854 11982 10906
rect 12034 10854 12046 10906
rect 12098 10854 12110 10906
rect 12162 10854 12174 10906
rect 12226 10854 19315 10906
rect 19367 10854 19379 10906
rect 19431 10854 19443 10906
rect 19495 10854 19507 10906
rect 19559 10854 20884 10906
rect 1104 10832 20884 10854
rect 2409 10795 2467 10801
rect 2409 10761 2421 10795
rect 2455 10792 2467 10795
rect 2498 10792 2504 10804
rect 2455 10764 2504 10792
rect 2455 10761 2467 10764
rect 2409 10755 2467 10761
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 4433 10795 4491 10801
rect 4433 10761 4445 10795
rect 4479 10792 4491 10795
rect 4709 10795 4767 10801
rect 4709 10792 4721 10795
rect 4479 10764 4721 10792
rect 4479 10761 4491 10764
rect 4433 10755 4491 10761
rect 4709 10761 4721 10764
rect 4755 10792 4767 10795
rect 5626 10792 5632 10804
rect 4755 10764 5632 10792
rect 4755 10761 4767 10764
rect 4709 10755 4767 10761
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 6273 10795 6331 10801
rect 6273 10761 6285 10795
rect 6319 10792 6331 10795
rect 6638 10792 6644 10804
rect 6319 10764 6644 10792
rect 6319 10761 6331 10764
rect 6273 10755 6331 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 8110 10752 8116 10804
rect 8168 10792 8174 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 8168 10764 8217 10792
rect 8168 10752 8174 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 10318 10792 10324 10804
rect 10279 10764 10324 10792
rect 8205 10755 8263 10761
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 11885 10795 11943 10801
rect 11885 10792 11897 10795
rect 11848 10764 11897 10792
rect 11848 10752 11854 10764
rect 11885 10761 11897 10764
rect 11931 10761 11943 10795
rect 11885 10755 11943 10761
rect 15013 10795 15071 10801
rect 15013 10761 15025 10795
rect 15059 10792 15071 10795
rect 15378 10792 15384 10804
rect 15059 10764 15384 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 19150 10792 19156 10804
rect 19111 10764 19156 10792
rect 19150 10752 19156 10764
rect 19208 10792 19214 10804
rect 19794 10792 19800 10804
rect 19208 10764 19800 10792
rect 19208 10752 19214 10764
rect 19794 10752 19800 10764
rect 19852 10752 19858 10804
rect 2041 10727 2099 10733
rect 2041 10693 2053 10727
rect 2087 10724 2099 10727
rect 8846 10724 8852 10736
rect 2087 10696 8852 10724
rect 2087 10693 2099 10696
rect 2041 10687 2099 10693
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 2056 10588 2084 10687
rect 8846 10684 8852 10696
rect 8904 10684 8910 10736
rect 12897 10727 12955 10733
rect 12897 10693 12909 10727
rect 12943 10724 12955 10727
rect 13446 10724 13452 10736
rect 12943 10696 13452 10724
rect 12943 10693 12955 10696
rect 12897 10687 12955 10693
rect 13446 10684 13452 10696
rect 13504 10724 13510 10736
rect 16942 10724 16948 10736
rect 13504 10696 16948 10724
rect 13504 10684 13510 10696
rect 16942 10684 16948 10696
rect 17000 10684 17006 10736
rect 4295 10659 4353 10665
rect 4295 10625 4307 10659
rect 4341 10656 4353 10659
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 4341 10628 5273 10656
rect 4341 10625 4353 10628
rect 4295 10619 4353 10625
rect 5261 10625 5273 10628
rect 5307 10656 5319 10659
rect 5902 10656 5908 10668
rect 5307 10628 5908 10656
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10656 7067 10659
rect 7282 10656 7288 10668
rect 7055 10628 7288 10656
rect 7055 10625 7067 10628
rect 7009 10619 7067 10625
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 11057 10659 11115 10665
rect 11057 10656 11069 10659
rect 9916 10628 11069 10656
rect 9916 10616 9922 10628
rect 11057 10625 11069 10628
rect 11103 10656 11115 10659
rect 11790 10656 11796 10668
rect 11103 10628 11796 10656
rect 11103 10625 11115 10628
rect 11057 10619 11115 10625
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 13354 10656 13360 10668
rect 13315 10628 13360 10656
rect 13354 10616 13360 10628
rect 13412 10656 13418 10668
rect 16298 10656 16304 10668
rect 13412 10628 16304 10656
rect 13412 10616 13418 10628
rect 16298 10616 16304 10628
rect 16356 10616 16362 10668
rect 16577 10659 16635 10665
rect 16577 10625 16589 10659
rect 16623 10656 16635 10659
rect 17310 10656 17316 10668
rect 16623 10628 17316 10656
rect 16623 10625 16635 10628
rect 16577 10619 16635 10625
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 4062 10588 4068 10600
rect 1443 10560 2084 10588
rect 4023 10560 4068 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4208 10591 4266 10597
rect 4208 10557 4220 10591
rect 4254 10588 4266 10591
rect 4433 10591 4491 10597
rect 4433 10588 4445 10591
rect 4254 10560 4445 10588
rect 4254 10557 4266 10560
rect 4208 10551 4266 10557
rect 4356 10532 4384 10560
rect 4433 10557 4445 10560
rect 4479 10557 4491 10591
rect 4433 10551 4491 10557
rect 8941 10591 8999 10597
rect 8941 10557 8953 10591
rect 8987 10588 8999 10591
rect 9030 10588 9036 10600
rect 8987 10560 9036 10588
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 9030 10548 9036 10560
rect 9088 10548 9094 10600
rect 16736 10591 16794 10597
rect 16736 10557 16748 10591
rect 16782 10588 16794 10591
rect 17126 10588 17132 10600
rect 16782 10560 17132 10588
rect 16782 10557 16794 10560
rect 16736 10551 16794 10557
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 18012 10560 18061 10588
rect 18012 10548 18018 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10557 18567 10591
rect 18509 10551 18567 10557
rect 2682 10520 2688 10532
rect 2643 10492 2688 10520
rect 2682 10480 2688 10492
rect 2740 10480 2746 10532
rect 2777 10523 2835 10529
rect 2777 10489 2789 10523
rect 2823 10489 2835 10523
rect 2777 10483 2835 10489
rect 3329 10523 3387 10529
rect 3329 10489 3341 10523
rect 3375 10520 3387 10523
rect 3375 10492 4154 10520
rect 3375 10489 3387 10492
rect 3329 10483 3387 10489
rect 106 10412 112 10464
rect 164 10452 170 10464
rect 1581 10455 1639 10461
rect 1581 10452 1593 10455
rect 164 10424 1593 10452
rect 164 10412 170 10424
rect 1581 10421 1593 10424
rect 1627 10421 1639 10455
rect 1581 10415 1639 10421
rect 2590 10412 2596 10464
rect 2648 10452 2654 10464
rect 2792 10452 2820 10483
rect 3605 10455 3663 10461
rect 3605 10452 3617 10455
rect 2648 10424 3617 10452
rect 2648 10412 2654 10424
rect 3605 10421 3617 10424
rect 3651 10421 3663 10455
rect 4126 10452 4154 10492
rect 4338 10480 4344 10532
rect 4396 10480 4402 10532
rect 5350 10520 5356 10532
rect 5311 10492 5356 10520
rect 5350 10480 5356 10492
rect 5408 10480 5414 10532
rect 5902 10520 5908 10532
rect 5863 10492 5908 10520
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 6641 10523 6699 10529
rect 6641 10489 6653 10523
rect 6687 10520 6699 10523
rect 7371 10523 7429 10529
rect 7371 10520 7383 10523
rect 6687 10492 7383 10520
rect 6687 10489 6699 10492
rect 6641 10483 6699 10489
rect 7371 10489 7383 10492
rect 7417 10520 7429 10523
rect 8849 10523 8907 10529
rect 8849 10520 8861 10523
rect 7417 10492 8861 10520
rect 7417 10489 7429 10492
rect 7371 10483 7429 10489
rect 8849 10489 8861 10492
rect 8895 10520 8907 10523
rect 9303 10523 9361 10529
rect 9303 10520 9315 10523
rect 8895 10492 9315 10520
rect 8895 10489 8907 10492
rect 8849 10483 8907 10489
rect 9303 10489 9315 10492
rect 9349 10520 9361 10523
rect 9674 10520 9680 10532
rect 9349 10492 9680 10520
rect 9349 10489 9361 10492
rect 9303 10483 9361 10489
rect 4246 10452 4252 10464
rect 4126 10424 4252 10452
rect 3605 10415 3663 10421
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 5074 10452 5080 10464
rect 4987 10424 5080 10452
rect 5074 10412 5080 10424
rect 5132 10452 5138 10464
rect 6656 10452 6684 10483
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 10778 10520 10784 10532
rect 10739 10492 10784 10520
rect 10778 10480 10784 10492
rect 10836 10480 10842 10532
rect 10870 10480 10876 10532
rect 10928 10520 10934 10532
rect 13678 10523 13736 10529
rect 13678 10520 13690 10523
rect 10928 10492 10973 10520
rect 13464 10492 13690 10520
rect 10928 10480 10934 10492
rect 13464 10464 13492 10492
rect 13678 10489 13690 10492
rect 13724 10489 13736 10523
rect 15194 10520 15200 10532
rect 15155 10492 15200 10520
rect 13678 10483 13736 10489
rect 15194 10480 15200 10492
rect 15252 10480 15258 10532
rect 15289 10523 15347 10529
rect 15289 10489 15301 10523
rect 15335 10489 15347 10523
rect 15289 10483 15347 10489
rect 15841 10523 15899 10529
rect 15841 10489 15853 10523
rect 15887 10520 15899 10523
rect 16022 10520 16028 10532
rect 15887 10492 16028 10520
rect 15887 10489 15899 10492
rect 15841 10483 15899 10489
rect 7926 10452 7932 10464
rect 5132 10424 6684 10452
rect 7887 10424 7932 10452
rect 5132 10412 5138 10424
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 9861 10455 9919 10461
rect 9861 10421 9873 10455
rect 9907 10452 9919 10455
rect 11606 10452 11612 10464
rect 9907 10424 11612 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 13262 10452 13268 10464
rect 13175 10424 13268 10452
rect 13262 10412 13268 10424
rect 13320 10452 13326 10464
rect 13446 10452 13452 10464
rect 13320 10424 13452 10452
rect 13320 10412 13326 10424
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 14277 10455 14335 10461
rect 14277 10421 14289 10455
rect 14323 10452 14335 10455
rect 14553 10455 14611 10461
rect 14553 10452 14565 10455
rect 14323 10424 14565 10452
rect 14323 10421 14335 10424
rect 14277 10415 14335 10421
rect 14553 10421 14565 10424
rect 14599 10452 14611 10455
rect 15304 10452 15332 10483
rect 16022 10480 16028 10492
rect 16080 10480 16086 10532
rect 18524 10520 18552 10551
rect 17880 10492 18552 10520
rect 17880 10464 17908 10492
rect 14599 10424 15332 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 15470 10412 15476 10464
rect 15528 10452 15534 10464
rect 16114 10452 16120 10464
rect 15528 10424 16120 10452
rect 15528 10412 15534 10424
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 16807 10455 16865 10461
rect 16807 10452 16819 10455
rect 16632 10424 16819 10452
rect 16632 10412 16638 10424
rect 16807 10421 16819 10424
rect 16853 10421 16865 10455
rect 17862 10452 17868 10464
rect 17823 10424 17868 10452
rect 16807 10415 16865 10421
rect 17862 10412 17868 10424
rect 17920 10412 17926 10464
rect 18138 10452 18144 10464
rect 18099 10424 18144 10452
rect 18138 10412 18144 10424
rect 18196 10412 18202 10464
rect 19610 10452 19616 10464
rect 19571 10424 19616 10452
rect 19610 10412 19616 10424
rect 19668 10412 19674 10464
rect 1104 10362 20884 10384
rect 1104 10310 8315 10362
rect 8367 10310 8379 10362
rect 8431 10310 8443 10362
rect 8495 10310 8507 10362
rect 8559 10310 15648 10362
rect 15700 10310 15712 10362
rect 15764 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 20884 10362
rect 1104 10288 20884 10310
rect 1210 10208 1216 10260
rect 1268 10248 1274 10260
rect 1535 10251 1593 10257
rect 1535 10248 1547 10251
rect 1268 10220 1547 10248
rect 1268 10208 1274 10220
rect 1535 10217 1547 10220
rect 1581 10217 1593 10251
rect 1535 10211 1593 10217
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2498 10248 2504 10260
rect 1995 10220 2504 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 3418 10248 3424 10260
rect 2740 10220 3424 10248
rect 2740 10208 2746 10220
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 5350 10208 5356 10260
rect 5408 10248 5414 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 5408 10220 5457 10248
rect 5408 10208 5414 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5445 10211 5503 10217
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 10410 10248 10416 10260
rect 9539 10220 10416 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 10410 10208 10416 10220
rect 10468 10208 10474 10260
rect 10597 10251 10655 10257
rect 10597 10217 10609 10251
rect 10643 10248 10655 10251
rect 10870 10248 10876 10260
rect 10643 10220 10876 10248
rect 10643 10217 10655 10220
rect 10597 10211 10655 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 12434 10248 12440 10260
rect 12395 10220 12440 10248
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 14826 10248 14832 10260
rect 13693 10220 14832 10248
rect 2590 10180 2596 10192
rect 2551 10152 2596 10180
rect 2590 10140 2596 10152
rect 2648 10140 2654 10192
rect 2958 10140 2964 10192
rect 3016 10180 3022 10192
rect 4249 10183 4307 10189
rect 4249 10180 4261 10183
rect 3016 10152 4261 10180
rect 3016 10140 3022 10152
rect 4249 10149 4261 10152
rect 4295 10149 4307 10183
rect 4249 10143 4307 10149
rect 4801 10183 4859 10189
rect 4801 10149 4813 10183
rect 4847 10180 4859 10183
rect 4982 10180 4988 10192
rect 4847 10152 4988 10180
rect 4847 10149 4859 10152
rect 4801 10143 4859 10149
rect 4982 10140 4988 10152
rect 5040 10140 5046 10192
rect 5810 10180 5816 10192
rect 5771 10152 5816 10180
rect 5810 10140 5816 10152
rect 5868 10140 5874 10192
rect 7837 10183 7895 10189
rect 7837 10149 7849 10183
rect 7883 10180 7895 10183
rect 7926 10180 7932 10192
rect 7883 10152 7932 10180
rect 7883 10149 7895 10152
rect 7837 10143 7895 10149
rect 7926 10140 7932 10152
rect 7984 10140 7990 10192
rect 8389 10183 8447 10189
rect 8389 10149 8401 10183
rect 8435 10180 8447 10183
rect 9858 10180 9864 10192
rect 8435 10152 9864 10180
rect 8435 10149 8447 10152
rect 8389 10143 8447 10149
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 9998 10183 10056 10189
rect 9998 10149 10010 10183
rect 10044 10149 10056 10183
rect 9998 10143 10056 10149
rect 1464 10115 1522 10121
rect 1464 10081 1476 10115
rect 1510 10112 1522 10115
rect 2314 10112 2320 10124
rect 1510 10084 2320 10112
rect 1510 10081 1522 10084
rect 1464 10075 1522 10081
rect 2314 10072 2320 10084
rect 2372 10072 2378 10124
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 10013 10112 10041 10143
rect 10778 10140 10784 10192
rect 10836 10180 10842 10192
rect 11241 10183 11299 10189
rect 11241 10180 11253 10183
rect 10836 10152 11253 10180
rect 10836 10140 10842 10152
rect 11241 10149 11253 10152
rect 11287 10149 11299 10183
rect 11606 10180 11612 10192
rect 11567 10152 11612 10180
rect 11241 10143 11299 10149
rect 11606 10140 11612 10152
rect 11664 10140 11670 10192
rect 11790 10140 11796 10192
rect 11848 10180 11854 10192
rect 13693 10180 13721 10220
rect 14826 10208 14832 10220
rect 14884 10208 14890 10260
rect 15010 10248 15016 10260
rect 14971 10220 15016 10248
rect 15010 10208 15016 10220
rect 15068 10208 15074 10260
rect 16942 10248 16948 10260
rect 16903 10220 16948 10248
rect 16942 10208 16948 10220
rect 17000 10208 17006 10260
rect 18506 10248 18512 10260
rect 18467 10220 18512 10248
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 11848 10152 13721 10180
rect 11848 10140 11854 10152
rect 13814 10140 13820 10192
rect 13872 10180 13878 10192
rect 13872 10152 13917 10180
rect 13872 10140 13878 10152
rect 14366 10140 14372 10192
rect 14424 10180 14430 10192
rect 15102 10180 15108 10192
rect 14424 10152 15108 10180
rect 14424 10140 14430 10152
rect 15102 10140 15108 10152
rect 15160 10180 15166 10192
rect 15473 10183 15531 10189
rect 15473 10180 15485 10183
rect 15160 10152 15485 10180
rect 15160 10140 15166 10152
rect 15473 10149 15485 10152
rect 15519 10149 15531 10183
rect 16022 10180 16028 10192
rect 15983 10152 16028 10180
rect 15473 10143 15531 10149
rect 16022 10140 16028 10152
rect 16080 10140 16086 10192
rect 16114 10140 16120 10192
rect 16172 10180 16178 10192
rect 16172 10152 18460 10180
rect 16172 10140 16178 10152
rect 18432 10124 18460 10152
rect 9640 10084 10041 10112
rect 9640 10072 9646 10084
rect 16666 10072 16672 10124
rect 16724 10112 16730 10124
rect 16853 10115 16911 10121
rect 16853 10112 16865 10115
rect 16724 10084 16865 10112
rect 16724 10072 16730 10084
rect 16853 10081 16865 10084
rect 16899 10081 16911 10115
rect 17310 10112 17316 10124
rect 17271 10084 17316 10112
rect 16853 10075 16911 10081
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10044 2559 10047
rect 3326 10044 3332 10056
rect 2547 10016 3332 10044
rect 2547 10013 2559 10016
rect 2501 10007 2559 10013
rect 3326 10004 3332 10016
rect 3384 10044 3390 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3384 10016 3801 10044
rect 3384 10004 3390 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4246 10044 4252 10056
rect 4203 10016 4252 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4246 10004 4252 10016
rect 4304 10004 4310 10056
rect 5718 10044 5724 10056
rect 5679 10016 5724 10044
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10013 6055 10047
rect 6914 10044 6920 10056
rect 6875 10016 6920 10044
rect 5997 10007 6055 10013
rect 3053 9979 3111 9985
rect 3053 9945 3065 9979
rect 3099 9976 3111 9979
rect 4522 9976 4528 9988
rect 3099 9948 4528 9976
rect 3099 9945 3111 9948
rect 3053 9939 3111 9945
rect 4522 9936 4528 9948
rect 4580 9976 4586 9988
rect 5902 9976 5908 9988
rect 4580 9948 5908 9976
rect 4580 9936 4586 9948
rect 5902 9936 5908 9948
rect 5960 9976 5966 9988
rect 6012 9976 6040 10007
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10044 7803 10047
rect 8018 10044 8024 10056
rect 7791 10016 8024 10044
rect 7791 10013 7803 10016
rect 7745 10007 7803 10013
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 9490 10004 9496 10056
rect 9548 10044 9554 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9548 10016 9689 10044
rect 9548 10004 9554 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 11514 10044 11520 10056
rect 11475 10016 11520 10044
rect 9677 10007 9735 10013
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 11790 10044 11796 10056
rect 11751 10016 11796 10044
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 13725 10047 13783 10053
rect 13725 10044 13737 10047
rect 13596 10016 13737 10044
rect 13596 10004 13602 10016
rect 13725 10013 13737 10016
rect 13771 10013 13783 10047
rect 14366 10044 14372 10056
rect 14327 10016 14372 10044
rect 13725 10007 13783 10013
rect 14366 10004 14372 10016
rect 14424 10044 14430 10056
rect 15381 10047 15439 10053
rect 15381 10044 15393 10047
rect 14424 10016 15393 10044
rect 14424 10004 14430 10016
rect 15381 10013 15393 10016
rect 15427 10013 15439 10047
rect 16868 10044 16896 10075
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 18414 10112 18420 10124
rect 18327 10084 18420 10112
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 18874 10112 18880 10124
rect 18835 10084 18880 10112
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 17954 10044 17960 10056
rect 16868 10016 17960 10044
rect 15381 10007 15439 10013
rect 17954 10004 17960 10016
rect 18012 10044 18018 10056
rect 18049 10047 18107 10053
rect 18049 10044 18061 10047
rect 18012 10016 18061 10044
rect 18012 10004 18018 10016
rect 18049 10013 18061 10016
rect 18095 10013 18107 10047
rect 18049 10007 18107 10013
rect 5960 9948 6040 9976
rect 5960 9936 5966 9948
rect 2222 9908 2228 9920
rect 2183 9880 2228 9908
rect 2222 9868 2228 9880
rect 2280 9868 2286 9920
rect 5166 9908 5172 9920
rect 5127 9880 5172 9908
rect 5166 9868 5172 9880
rect 5224 9868 5230 9920
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6362 9908 6368 9920
rect 5776 9880 6368 9908
rect 5776 9868 5782 9880
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 7282 9908 7288 9920
rect 7243 9880 7288 9908
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 9030 9908 9036 9920
rect 8991 9880 9036 9908
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 13446 9908 13452 9920
rect 13407 9880 13452 9908
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 14734 9908 14740 9920
rect 14695 9880 14740 9908
rect 14734 9868 14740 9880
rect 14792 9868 14798 9920
rect 1104 9818 20884 9840
rect 1104 9766 4648 9818
rect 4700 9766 4712 9818
rect 4764 9766 4776 9818
rect 4828 9766 4840 9818
rect 4892 9766 11982 9818
rect 12034 9766 12046 9818
rect 12098 9766 12110 9818
rect 12162 9766 12174 9818
rect 12226 9766 19315 9818
rect 19367 9766 19379 9818
rect 19431 9766 19443 9818
rect 19495 9766 19507 9818
rect 19559 9766 20884 9818
rect 1104 9744 20884 9766
rect 2590 9704 2596 9716
rect 2551 9676 2596 9704
rect 2590 9664 2596 9676
rect 2648 9704 2654 9716
rect 2869 9707 2927 9713
rect 2869 9704 2881 9707
rect 2648 9676 2881 9704
rect 2648 9664 2654 9676
rect 2869 9673 2881 9676
rect 2915 9673 2927 9707
rect 2869 9667 2927 9673
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3237 9707 3295 9713
rect 3237 9704 3249 9707
rect 3016 9676 3249 9704
rect 3016 9664 3022 9676
rect 3237 9673 3249 9676
rect 3283 9673 3295 9707
rect 3237 9667 3295 9673
rect 5537 9707 5595 9713
rect 5537 9673 5549 9707
rect 5583 9704 5595 9707
rect 5810 9704 5816 9716
rect 5583 9676 5816 9704
rect 5583 9673 5595 9676
rect 5537 9667 5595 9673
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 6273 9707 6331 9713
rect 6273 9673 6285 9707
rect 6319 9704 6331 9707
rect 6362 9704 6368 9716
rect 6319 9676 6368 9704
rect 6319 9673 6331 9676
rect 6273 9667 6331 9673
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 8110 9704 8116 9716
rect 6610 9676 8116 9704
rect 198 9596 204 9648
rect 256 9636 262 9648
rect 3605 9639 3663 9645
rect 3605 9636 3617 9639
rect 256 9608 3617 9636
rect 256 9596 262 9608
rect 3605 9605 3617 9608
rect 3651 9605 3663 9639
rect 3605 9599 3663 9605
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 6610 9636 6638 9676
rect 8110 9664 8116 9676
rect 8168 9704 8174 9716
rect 8662 9704 8668 9716
rect 8168 9676 8668 9704
rect 8168 9664 8174 9676
rect 8662 9664 8668 9676
rect 8720 9664 8726 9716
rect 11606 9704 11612 9716
rect 11567 9676 11612 9704
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 14093 9707 14151 9713
rect 14093 9704 14105 9707
rect 13872 9676 14105 9704
rect 13872 9664 13878 9676
rect 14093 9673 14105 9676
rect 14139 9704 14151 9707
rect 14461 9707 14519 9713
rect 14461 9704 14473 9707
rect 14139 9676 14473 9704
rect 14139 9673 14151 9676
rect 14093 9667 14151 9673
rect 14461 9673 14473 9676
rect 14507 9704 14519 9707
rect 14826 9704 14832 9716
rect 14507 9676 14832 9704
rect 14507 9673 14519 9676
rect 14461 9667 14519 9673
rect 14826 9664 14832 9676
rect 14884 9664 14890 9716
rect 17310 9704 17316 9716
rect 17271 9676 17316 9704
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 4212 9608 6638 9636
rect 4212 9596 4218 9608
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 10873 9639 10931 9645
rect 9732 9608 9777 9636
rect 9732 9596 9738 9608
rect 10873 9605 10885 9639
rect 10919 9636 10931 9639
rect 11698 9636 11704 9648
rect 10919 9608 11704 9636
rect 10919 9605 10931 9608
rect 10873 9599 10931 9605
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 14918 9596 14924 9648
rect 14976 9636 14982 9648
rect 15194 9636 15200 9648
rect 14976 9608 15200 9636
rect 14976 9596 14982 9608
rect 15194 9596 15200 9608
rect 15252 9636 15258 9648
rect 15289 9639 15347 9645
rect 15289 9636 15301 9639
rect 15252 9608 15301 9636
rect 15252 9596 15258 9608
rect 15289 9605 15301 9608
rect 15335 9605 15347 9639
rect 15289 9599 15347 9605
rect 6641 9571 6699 9577
rect 2700 9540 4568 9568
rect 1486 9460 1492 9512
rect 1544 9500 1550 9512
rect 1673 9503 1731 9509
rect 1673 9500 1685 9503
rect 1544 9472 1685 9500
rect 1544 9460 1550 9472
rect 1673 9469 1685 9472
rect 1719 9500 1731 9503
rect 2222 9500 2228 9512
rect 1719 9472 2228 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 2035 9435 2093 9441
rect 2035 9401 2047 9435
rect 2081 9432 2093 9435
rect 2406 9432 2412 9444
rect 2081 9404 2412 9432
rect 2081 9401 2093 9404
rect 2035 9395 2093 9401
rect 2406 9392 2412 9404
rect 2464 9432 2470 9444
rect 2700 9432 2728 9540
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9500 3479 9503
rect 3467 9472 4108 9500
rect 3467 9469 3479 9472
rect 3421 9463 3479 9469
rect 2464 9404 2728 9432
rect 2464 9392 2470 9404
rect 4080 9373 4108 9472
rect 4540 9441 4568 9540
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 7929 9571 7987 9577
rect 6687 9540 7420 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 7392 9512 7420 9540
rect 7929 9537 7941 9571
rect 7975 9568 7987 9571
rect 8018 9568 8024 9580
rect 7975 9540 8024 9568
rect 7975 9537 7987 9540
rect 7929 9531 7987 9537
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9568 8539 9571
rect 8662 9568 8668 9580
rect 8527 9540 8668 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 8662 9528 8668 9540
rect 8720 9568 8726 9580
rect 9214 9568 9220 9580
rect 8720 9540 9220 9568
rect 8720 9528 8726 9540
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 11514 9568 11520 9580
rect 9876 9540 11520 9568
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9500 4675 9503
rect 4663 9472 5212 9500
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 5184 9444 5212 9472
rect 6730 9460 6736 9512
rect 6788 9500 6794 9512
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6788 9472 6837 9500
rect 6788 9460 6794 9472
rect 6825 9469 6837 9472
rect 6871 9500 6883 9503
rect 6914 9500 6920 9512
rect 6871 9472 6920 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7374 9500 7380 9512
rect 7335 9472 7380 9500
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9500 9183 9503
rect 9876 9500 9904 9540
rect 11514 9528 11520 9540
rect 11572 9568 11578 9580
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 11572 9540 11897 9568
rect 11572 9528 11578 9540
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 14734 9568 14740 9580
rect 14647 9540 14740 9568
rect 11885 9531 11943 9537
rect 14734 9528 14740 9540
rect 14792 9568 14798 9580
rect 19751 9571 19809 9577
rect 19751 9568 19763 9571
rect 14792 9540 19763 9568
rect 14792 9528 14798 9540
rect 19751 9537 19763 9540
rect 19797 9537 19809 9571
rect 19751 9531 19809 9537
rect 9171 9472 9904 9500
rect 9953 9503 10011 9509
rect 9171 9469 9183 9472
rect 9125 9463 9183 9469
rect 9953 9469 9965 9503
rect 9999 9500 10011 9503
rect 10870 9500 10876 9512
rect 9999 9472 10876 9500
rect 9999 9469 10011 9472
rect 9953 9463 10011 9469
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 12894 9500 12900 9512
rect 12855 9472 12900 9500
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 16206 9500 16212 9512
rect 15672 9472 16212 9500
rect 4525 9435 4583 9441
rect 4525 9401 4537 9435
rect 4571 9432 4583 9435
rect 4979 9435 5037 9441
rect 4979 9432 4991 9435
rect 4571 9404 4991 9432
rect 4571 9401 4583 9404
rect 4525 9395 4583 9401
rect 4979 9401 4991 9404
rect 5025 9432 5037 9435
rect 5074 9432 5080 9444
rect 5025 9404 5080 9432
rect 5025 9401 5037 9404
rect 4979 9395 5037 9401
rect 5074 9392 5080 9404
rect 5132 9392 5138 9444
rect 5166 9392 5172 9444
rect 5224 9432 5230 9444
rect 8573 9435 8631 9441
rect 5224 9404 6868 9432
rect 5224 9392 5230 9404
rect 4065 9367 4123 9373
rect 4065 9333 4077 9367
rect 4111 9364 4123 9367
rect 5350 9364 5356 9376
rect 4111 9336 5356 9364
rect 4111 9333 4123 9336
rect 4065 9327 4123 9333
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 6086 9364 6092 9376
rect 5500 9336 6092 9364
rect 5500 9324 5506 9336
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6840 9364 6868 9404
rect 8573 9401 8585 9435
rect 8619 9401 8631 9435
rect 8573 9395 8631 9401
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 6840 9336 6929 9364
rect 6917 9333 6929 9336
rect 6963 9333 6975 9367
rect 6917 9327 6975 9333
rect 8297 9367 8355 9373
rect 8297 9333 8309 9367
rect 8343 9364 8355 9367
rect 8588 9364 8616 9395
rect 9674 9392 9680 9444
rect 9732 9432 9738 9444
rect 10274 9435 10332 9441
rect 10274 9432 10286 9435
rect 9732 9404 10286 9432
rect 9732 9392 9738 9404
rect 10274 9401 10286 9404
rect 10320 9432 10332 9435
rect 11149 9435 11207 9441
rect 11149 9432 11161 9435
rect 10320 9404 11161 9432
rect 10320 9401 10332 9404
rect 10274 9395 10332 9401
rect 11149 9401 11161 9404
rect 11195 9432 11207 9435
rect 12710 9432 12716 9444
rect 11195 9404 12716 9432
rect 11195 9401 11207 9404
rect 11149 9395 11207 9401
rect 12710 9392 12716 9404
rect 12768 9432 12774 9444
rect 13218 9435 13276 9441
rect 13218 9432 13230 9435
rect 12768 9404 13230 9432
rect 12768 9392 12774 9404
rect 13218 9401 13230 9404
rect 13264 9432 13276 9435
rect 13446 9432 13452 9444
rect 13264 9404 13452 9432
rect 13264 9401 13276 9404
rect 13218 9395 13276 9401
rect 13446 9392 13452 9404
rect 13504 9392 13510 9444
rect 14826 9392 14832 9444
rect 14884 9432 14890 9444
rect 14884 9404 14929 9432
rect 14884 9392 14890 9404
rect 9582 9364 9588 9376
rect 8343 9336 9588 9364
rect 8343 9333 8355 9336
rect 8297 9327 8355 9333
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 14550 9324 14556 9376
rect 14608 9364 14614 9376
rect 15672 9373 15700 9472
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 16761 9503 16819 9509
rect 16761 9469 16773 9503
rect 16807 9500 16819 9503
rect 17310 9500 17316 9512
rect 16807 9472 17316 9500
rect 16807 9469 16819 9472
rect 16761 9463 16819 9469
rect 16114 9432 16120 9444
rect 16027 9404 16120 9432
rect 16114 9392 16120 9404
rect 16172 9432 16178 9444
rect 16776 9432 16804 9463
rect 17310 9460 17316 9472
rect 17368 9460 17374 9512
rect 18046 9500 18052 9512
rect 18007 9472 18052 9500
rect 18046 9460 18052 9472
rect 18104 9460 18110 9512
rect 18509 9503 18567 9509
rect 18509 9469 18521 9503
rect 18555 9469 18567 9503
rect 18509 9463 18567 9469
rect 17862 9432 17868 9444
rect 16172 9404 16804 9432
rect 17775 9404 17868 9432
rect 16172 9392 16178 9404
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 14608 9336 15669 9364
rect 14608 9324 14614 9336
rect 15657 9333 15669 9336
rect 15703 9333 15715 9367
rect 16298 9364 16304 9376
rect 16259 9336 16304 9364
rect 15657 9327 15715 9333
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 17310 9324 17316 9376
rect 17368 9364 17374 9376
rect 17788 9373 17816 9404
rect 17862 9392 17868 9404
rect 17920 9432 17926 9444
rect 18524 9432 18552 9463
rect 18598 9460 18604 9512
rect 18656 9500 18662 9512
rect 19648 9503 19706 9509
rect 19648 9500 19660 9503
rect 18656 9472 19660 9500
rect 18656 9460 18662 9472
rect 19648 9469 19660 9472
rect 19694 9500 19706 9503
rect 19886 9500 19892 9512
rect 19694 9472 19892 9500
rect 19694 9469 19706 9472
rect 19648 9463 19706 9469
rect 19886 9460 19892 9472
rect 19944 9500 19950 9512
rect 20073 9503 20131 9509
rect 20073 9500 20085 9503
rect 19944 9472 20085 9500
rect 19944 9460 19950 9472
rect 20073 9469 20085 9472
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 18874 9432 18880 9444
rect 17920 9404 18880 9432
rect 17920 9392 17926 9404
rect 18874 9392 18880 9404
rect 18932 9432 18938 9444
rect 19061 9435 19119 9441
rect 19061 9432 19073 9435
rect 18932 9404 19073 9432
rect 18932 9392 18938 9404
rect 19061 9401 19073 9404
rect 19107 9401 19119 9435
rect 19061 9395 19119 9401
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17368 9336 17785 9364
rect 17368 9324 17374 9336
rect 17773 9333 17785 9336
rect 17819 9333 17831 9367
rect 18138 9364 18144 9376
rect 18099 9336 18144 9364
rect 17773 9327 17831 9333
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 1104 9274 20884 9296
rect 1104 9222 8315 9274
rect 8367 9222 8379 9274
rect 8431 9222 8443 9274
rect 8495 9222 8507 9274
rect 8559 9222 15648 9274
rect 15700 9222 15712 9274
rect 15764 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 20884 9274
rect 1104 9200 20884 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 3050 9120 3056 9172
rect 3108 9120 3114 9172
rect 3234 9120 3240 9172
rect 3292 9160 3298 9172
rect 3513 9163 3571 9169
rect 3513 9160 3525 9163
rect 3292 9132 3525 9160
rect 3292 9120 3298 9132
rect 3513 9129 3525 9132
rect 3559 9160 3571 9163
rect 4154 9160 4160 9172
rect 3559 9132 4160 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 6822 9160 6828 9172
rect 4304 9132 6828 9160
rect 4304 9120 4310 9132
rect 3068 9092 3096 9120
rect 4522 9092 4528 9104
rect 3068 9064 4528 9092
rect 4522 9052 4528 9064
rect 4580 9052 4586 9104
rect 5261 9095 5319 9101
rect 5261 9061 5273 9095
rect 5307 9092 5319 9095
rect 5442 9092 5448 9104
rect 5307 9064 5448 9092
rect 5307 9061 5319 9064
rect 5261 9055 5319 9061
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 5537 9095 5595 9101
rect 5537 9061 5549 9095
rect 5583 9092 5595 9095
rect 5810 9092 5816 9104
rect 5583 9064 5816 9092
rect 5583 9061 5595 9064
rect 5537 9055 5595 9061
rect 5810 9052 5816 9064
rect 5868 9052 5874 9104
rect 6104 9101 6132 9132
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7926 9160 7932 9172
rect 7887 9132 7932 9160
rect 7926 9120 7932 9132
rect 7984 9120 7990 9172
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 8662 9160 8668 9172
rect 8527 9132 8668 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 12894 9160 12900 9172
rect 10796 9132 12020 9160
rect 12855 9132 12900 9160
rect 10796 9104 10824 9132
rect 6089 9095 6147 9101
rect 6089 9061 6101 9095
rect 6135 9061 6147 9095
rect 6089 9055 6147 9061
rect 6638 9052 6644 9104
rect 6696 9092 6702 9104
rect 7101 9095 7159 9101
rect 7101 9092 7113 9095
rect 6696 9064 7113 9092
rect 6696 9052 6702 9064
rect 7101 9061 7113 9064
rect 7147 9061 7159 9095
rect 7101 9055 7159 9061
rect 9582 9052 9588 9104
rect 9640 9092 9646 9104
rect 9861 9095 9919 9101
rect 9861 9092 9873 9095
rect 9640 9064 9873 9092
rect 9640 9052 9646 9064
rect 9861 9061 9873 9064
rect 9907 9061 9919 9095
rect 9861 9055 9919 9061
rect 10413 9095 10471 9101
rect 10413 9061 10425 9095
rect 10459 9092 10471 9095
rect 10778 9092 10784 9104
rect 10459 9064 10784 9092
rect 10459 9061 10471 9064
rect 10413 9055 10471 9061
rect 10778 9052 10784 9064
rect 10836 9052 10842 9104
rect 11330 9092 11336 9104
rect 11291 9064 11336 9092
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 11425 9095 11483 9101
rect 11425 9061 11437 9095
rect 11471 9092 11483 9095
rect 11698 9092 11704 9104
rect 11471 9064 11704 9092
rect 11471 9061 11483 9064
rect 11425 9055 11483 9061
rect 11698 9052 11704 9064
rect 11756 9052 11762 9104
rect 11992 9101 12020 9132
rect 12894 9120 12900 9132
rect 12952 9160 12958 9172
rect 15381 9163 15439 9169
rect 15381 9160 15393 9163
rect 12952 9132 15393 9160
rect 12952 9120 12958 9132
rect 15381 9129 15393 9132
rect 15427 9129 15439 9163
rect 16942 9160 16948 9172
rect 16903 9132 16948 9160
rect 15381 9123 15439 9129
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 18414 9120 18420 9172
rect 18472 9160 18478 9172
rect 18877 9163 18935 9169
rect 18877 9160 18889 9163
rect 18472 9132 18889 9160
rect 18472 9120 18478 9132
rect 18877 9129 18889 9132
rect 18923 9129 18935 9163
rect 18877 9123 18935 9129
rect 11977 9095 12035 9101
rect 11977 9061 11989 9095
rect 12023 9061 12035 9095
rect 13538 9092 13544 9104
rect 13499 9064 13544 9092
rect 11977 9055 12035 9061
rect 13538 9052 13544 9064
rect 13596 9052 13602 9104
rect 13814 9092 13820 9104
rect 13775 9064 13820 9092
rect 13814 9052 13820 9064
rect 13872 9052 13878 9104
rect 14366 9092 14372 9104
rect 14327 9064 14372 9092
rect 14366 9052 14372 9064
rect 14424 9052 14430 9104
rect 15102 9092 15108 9104
rect 15063 9064 15108 9092
rect 15102 9052 15108 9064
rect 15160 9052 15166 9104
rect 18046 9092 18052 9104
rect 15304 9064 18052 9092
rect 1302 8984 1308 9036
rect 1360 9024 1366 9036
rect 1397 9027 1455 9033
rect 1397 9024 1409 9027
rect 1360 8996 1409 9024
rect 1360 8984 1366 8996
rect 1397 8993 1409 8996
rect 1443 8993 1455 9027
rect 1854 9024 1860 9036
rect 1815 8996 1860 9024
rect 1397 8987 1455 8993
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 2038 8984 2044 9036
rect 2096 9024 2102 9036
rect 2774 9024 2780 9036
rect 2096 8996 2780 9024
rect 2096 8984 2102 8996
rect 2774 8984 2780 8996
rect 2832 9024 2838 9036
rect 2996 9027 3054 9033
rect 2996 9024 3008 9027
rect 2832 8996 3008 9024
rect 2832 8984 2838 8996
rect 2996 8993 3008 8996
rect 3042 8993 3054 9027
rect 2996 8987 3054 8993
rect 3237 9027 3295 9033
rect 3237 8993 3249 9027
rect 3283 9024 3295 9027
rect 3326 9024 3332 9036
rect 3283 8996 3332 9024
rect 3283 8993 3295 8996
rect 3237 8987 3295 8993
rect 3326 8984 3332 8996
rect 3384 8984 3390 9036
rect 4338 8984 4344 9036
rect 4396 9033 4402 9036
rect 4396 9027 4434 9033
rect 4422 8993 4434 9027
rect 4396 8987 4434 8993
rect 8640 9027 8698 9033
rect 8640 8993 8652 9027
rect 8686 9024 8698 9027
rect 8846 9024 8852 9036
rect 8686 8996 8852 9024
rect 8686 8993 8698 8996
rect 8640 8987 8698 8993
rect 4396 8984 4402 8987
rect 8846 8984 8852 8996
rect 8904 8984 8910 9036
rect 9490 9024 9496 9036
rect 9451 8996 9496 9024
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 2498 8956 2504 8968
rect 2459 8928 2504 8956
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 4479 8959 4537 8965
rect 4479 8925 4491 8959
rect 4525 8956 4537 8959
rect 7006 8956 7012 8968
rect 4525 8928 7012 8956
rect 4525 8925 4537 8928
rect 4479 8919 4537 8925
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 9766 8956 9772 8968
rect 9727 8928 9772 8956
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 10870 8956 10876 8968
rect 10827 8928 10876 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8925 13783 8959
rect 14384 8956 14412 9052
rect 14458 8984 14464 9036
rect 14516 9024 14522 9036
rect 15304 9033 15332 9064
rect 18046 9052 18052 9064
rect 18104 9052 18110 9104
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 14516 8996 15301 9024
rect 14516 8984 14522 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 15654 8984 15660 9036
rect 15712 9024 15718 9036
rect 15841 9027 15899 9033
rect 15841 9024 15853 9027
rect 15712 8996 15853 9024
rect 15712 8984 15718 8996
rect 15841 8993 15853 8996
rect 15887 9024 15899 9027
rect 16114 9024 16120 9036
rect 15887 8996 16120 9024
rect 15887 8993 15899 8996
rect 15841 8987 15899 8993
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 16206 8984 16212 9036
rect 16264 9024 16270 9036
rect 16758 9024 16764 9036
rect 16264 8996 16764 9024
rect 16264 8984 16270 8996
rect 16758 8984 16764 8996
rect 16816 9024 16822 9036
rect 16853 9027 16911 9033
rect 16853 9024 16865 9027
rect 16816 8996 16865 9024
rect 16816 8984 16822 8996
rect 16853 8993 16865 8996
rect 16899 8993 16911 9027
rect 17310 9024 17316 9036
rect 17271 8996 17316 9024
rect 16853 8987 16911 8993
rect 17310 8984 17316 8996
rect 17368 8984 17374 9036
rect 17678 8984 17684 9036
rect 17736 9024 17742 9036
rect 18484 9027 18542 9033
rect 18484 9024 18496 9027
rect 17736 8996 18496 9024
rect 17736 8984 17742 8996
rect 18484 8993 18496 8996
rect 18530 9024 18542 9027
rect 18874 9024 18880 9036
rect 18530 8996 18880 9024
rect 18530 8993 18542 8996
rect 18484 8987 18542 8993
rect 18874 8984 18880 8996
rect 18932 8984 18938 9036
rect 19150 8984 19156 9036
rect 19208 9024 19214 9036
rect 19464 9027 19522 9033
rect 19464 9024 19476 9027
rect 19208 8996 19476 9024
rect 19208 8984 19214 8996
rect 19464 8993 19476 8996
rect 19510 8993 19522 9027
rect 19464 8987 19522 8993
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 14384 8928 16313 8956
rect 13725 8919 13783 8925
rect 16301 8925 16313 8928
rect 16347 8956 16359 8959
rect 16482 8956 16488 8968
rect 16347 8928 16488 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 7558 8888 7564 8900
rect 7519 8860 7564 8888
rect 7558 8848 7564 8860
rect 7616 8848 7622 8900
rect 9033 8891 9091 8897
rect 9033 8888 9045 8891
rect 8404 8860 9045 8888
rect 2869 8823 2927 8829
rect 2869 8789 2881 8823
rect 2915 8820 2927 8823
rect 2958 8820 2964 8832
rect 2915 8792 2964 8820
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3878 8820 3884 8832
rect 3839 8792 3884 8820
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 4580 8792 4813 8820
rect 4580 8780 4586 8792
rect 4801 8789 4813 8792
rect 4847 8789 4859 8823
rect 4801 8783 4859 8789
rect 5442 8780 5448 8832
rect 5500 8820 5506 8832
rect 6365 8823 6423 8829
rect 6365 8820 6377 8823
rect 5500 8792 6377 8820
rect 5500 8780 5506 8792
rect 6365 8789 6377 8792
rect 6411 8789 6423 8823
rect 6365 8783 6423 8789
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 8404 8820 8432 8860
rect 9033 8857 9045 8860
rect 9079 8857 9091 8891
rect 9033 8851 9091 8857
rect 6972 8792 8432 8820
rect 8711 8823 8769 8829
rect 6972 8780 6978 8792
rect 8711 8789 8723 8823
rect 8757 8820 8769 8823
rect 8938 8820 8944 8832
rect 8757 8792 8944 8820
rect 8757 8789 8769 8792
rect 8711 8783 8769 8789
rect 8938 8780 8944 8792
rect 8996 8780 9002 8832
rect 10686 8780 10692 8832
rect 10744 8820 10750 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 10744 8792 11069 8820
rect 10744 8780 10750 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 13740 8820 13768 8919
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 14274 8848 14280 8900
rect 14332 8888 14338 8900
rect 15930 8888 15936 8900
rect 14332 8860 15936 8888
rect 14332 8848 14338 8860
rect 15930 8848 15936 8860
rect 15988 8848 15994 8900
rect 14734 8820 14740 8832
rect 13740 8792 14740 8820
rect 11057 8783 11115 8789
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 16632 8792 16681 8820
rect 16632 8780 16638 8792
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 16669 8783 16727 8789
rect 16850 8780 16856 8832
rect 16908 8820 16914 8832
rect 18555 8823 18613 8829
rect 18555 8820 18567 8823
rect 16908 8792 18567 8820
rect 16908 8780 16914 8792
rect 18555 8789 18567 8792
rect 18601 8789 18613 8823
rect 18555 8783 18613 8789
rect 18966 8780 18972 8832
rect 19024 8820 19030 8832
rect 19567 8823 19625 8829
rect 19567 8820 19579 8823
rect 19024 8792 19579 8820
rect 19024 8780 19030 8792
rect 19567 8789 19579 8792
rect 19613 8789 19625 8823
rect 19567 8783 19625 8789
rect 1104 8730 20884 8752
rect 1104 8678 4648 8730
rect 4700 8678 4712 8730
rect 4764 8678 4776 8730
rect 4828 8678 4840 8730
rect 4892 8678 11982 8730
rect 12034 8678 12046 8730
rect 12098 8678 12110 8730
rect 12162 8678 12174 8730
rect 12226 8678 19315 8730
rect 19367 8678 19379 8730
rect 19431 8678 19443 8730
rect 19495 8678 19507 8730
rect 19559 8678 20884 8730
rect 1104 8656 20884 8678
rect 2774 8616 2780 8628
rect 2735 8588 2780 8616
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 5810 8616 5816 8628
rect 5675 8588 5816 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 6089 8619 6147 8625
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 7374 8616 7380 8628
rect 6135 8588 7380 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 8846 8616 8852 8628
rect 8619 8588 8852 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9582 8616 9588 8628
rect 9543 8588 9588 8616
rect 9582 8576 9588 8588
rect 9640 8616 9646 8628
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 9640 8588 9873 8616
rect 9640 8576 9646 8588
rect 9861 8585 9873 8588
rect 9907 8585 9919 8619
rect 11698 8616 11704 8628
rect 11659 8588 11704 8616
rect 9861 8579 9919 8585
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 12710 8616 12716 8628
rect 12671 8588 12716 8616
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 13814 8616 13820 8628
rect 13771 8588 13820 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 13814 8576 13820 8588
rect 13872 8616 13878 8628
rect 14001 8619 14059 8625
rect 14001 8616 14013 8619
rect 13872 8588 14013 8616
rect 13872 8576 13878 8588
rect 14001 8585 14013 8588
rect 14047 8585 14059 8619
rect 14001 8579 14059 8585
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 19751 8619 19809 8625
rect 19751 8616 19763 8619
rect 14792 8588 19763 8616
rect 14792 8576 14798 8588
rect 19751 8585 19763 8588
rect 19797 8585 19809 8619
rect 19751 8579 19809 8585
rect 4338 8508 4344 8560
rect 4396 8548 4402 8560
rect 4433 8551 4491 8557
rect 4433 8548 4445 8551
rect 4396 8520 4445 8548
rect 4396 8508 4402 8520
rect 4433 8517 4445 8520
rect 4479 8548 4491 8551
rect 8202 8548 8208 8560
rect 4479 8520 8208 8548
rect 4479 8517 4491 8520
rect 4433 8511 4491 8517
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 13538 8508 13544 8560
rect 13596 8548 13602 8560
rect 18966 8548 18972 8560
rect 13596 8520 18972 8548
rect 13596 8508 13602 8520
rect 18966 8508 18972 8520
rect 19024 8508 19030 8560
rect 2498 8480 2504 8492
rect 1688 8452 2504 8480
rect 1688 8421 1716 8452
rect 2498 8440 2504 8452
rect 2556 8440 2562 8492
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 3476 8452 4077 8480
rect 3476 8440 3482 8452
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8381 1731 8415
rect 1673 8375 1731 8381
rect 1854 8372 1860 8424
rect 1912 8412 1918 8424
rect 1949 8415 2007 8421
rect 1949 8412 1961 8415
rect 1912 8384 1961 8412
rect 1912 8372 1918 8384
rect 1949 8381 1961 8384
rect 1995 8412 2007 8415
rect 3234 8412 3240 8424
rect 1995 8384 2544 8412
rect 3195 8384 3240 8412
rect 1995 8381 2007 8384
rect 1949 8375 2007 8381
rect 2130 8344 2136 8356
rect 2091 8316 2136 8344
rect 2130 8304 2136 8316
rect 2188 8304 2194 8356
rect 2516 8288 2544 8384
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 3528 8421 3556 8452
rect 4065 8449 4077 8452
rect 4111 8480 4123 8483
rect 4111 8452 5120 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 3513 8415 3571 8421
rect 3513 8381 3525 8415
rect 3559 8381 3571 8415
rect 4338 8412 4344 8424
rect 3513 8375 3571 8381
rect 4126 8384 4344 8412
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 4126 8344 4154 8384
rect 4338 8372 4344 8384
rect 4396 8372 4402 8424
rect 4522 8412 4528 8424
rect 4483 8384 4528 8412
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 5092 8421 5120 8452
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 6328 8452 7205 8480
rect 6328 8440 6334 8452
rect 7193 8449 7205 8452
rect 7239 8480 7251 8483
rect 7650 8480 7656 8492
rect 7239 8452 7656 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 10778 8440 10784 8492
rect 10836 8480 10842 8492
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10836 8452 11069 8480
rect 10836 8440 10842 8452
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8480 12311 8483
rect 12805 8483 12863 8489
rect 12805 8480 12817 8483
rect 12299 8452 12817 8480
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 12805 8449 12817 8452
rect 12851 8480 12863 8483
rect 14642 8480 14648 8492
rect 12851 8452 14648 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 14918 8480 14924 8492
rect 14879 8452 14924 8480
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 15654 8480 15660 8492
rect 15615 8452 15660 8480
rect 15654 8440 15660 8452
rect 15712 8480 15718 8492
rect 15930 8480 15936 8492
rect 15712 8452 15936 8480
rect 15712 8440 15718 8452
rect 15930 8440 15936 8452
rect 15988 8440 15994 8492
rect 16025 8483 16083 8489
rect 16025 8449 16037 8483
rect 16071 8480 16083 8483
rect 16206 8480 16212 8492
rect 16071 8452 16212 8480
rect 16071 8449 16083 8452
rect 16025 8443 16083 8449
rect 16206 8440 16212 8452
rect 16264 8440 16270 8492
rect 16942 8440 16948 8492
rect 17000 8480 17006 8492
rect 17770 8480 17776 8492
rect 17000 8452 17776 8480
rect 17000 8440 17006 8452
rect 17770 8440 17776 8452
rect 17828 8480 17834 8492
rect 17828 8452 18184 8480
rect 17828 8440 17834 8452
rect 5077 8415 5135 8421
rect 5077 8381 5089 8415
rect 5123 8412 5135 8415
rect 6089 8415 6147 8421
rect 6089 8412 6101 8415
rect 5123 8384 6101 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 6089 8381 6101 8384
rect 6135 8381 6147 8415
rect 6089 8375 6147 8381
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8662 8412 8668 8424
rect 8251 8384 8668 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 16117 8415 16175 8421
rect 16117 8381 16129 8415
rect 16163 8381 16175 8415
rect 16224 8412 16252 8440
rect 16577 8415 16635 8421
rect 16577 8412 16589 8415
rect 16224 8384 16589 8412
rect 16117 8375 16175 8381
rect 16577 8381 16589 8384
rect 16623 8412 16635 8415
rect 17129 8415 17187 8421
rect 17129 8412 17141 8415
rect 16623 8384 17141 8412
rect 16623 8381 16635 8384
rect 16577 8375 16635 8381
rect 17129 8381 17141 8384
rect 17175 8412 17187 8415
rect 17310 8412 17316 8424
rect 17175 8384 17316 8412
rect 17175 8381 17187 8384
rect 17129 8375 17187 8381
rect 6273 8347 6331 8353
rect 3752 8316 4154 8344
rect 4264 8316 4476 8344
rect 3752 8304 3758 8316
rect 2498 8276 2504 8288
rect 2459 8248 2504 8276
rect 2498 8236 2504 8248
rect 2556 8236 2562 8288
rect 2866 8236 2872 8288
rect 2924 8276 2930 8288
rect 3053 8279 3111 8285
rect 3053 8276 3065 8279
rect 2924 8248 3065 8276
rect 2924 8236 2930 8248
rect 3053 8245 3065 8248
rect 3099 8245 3111 8279
rect 3053 8239 3111 8245
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 4264 8276 4292 8316
rect 4120 8248 4292 8276
rect 4448 8276 4476 8316
rect 6273 8313 6285 8347
rect 6319 8344 6331 8347
rect 6917 8347 6975 8353
rect 6917 8344 6929 8347
rect 6319 8316 6929 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 6917 8313 6929 8316
rect 6963 8313 6975 8347
rect 6917 8307 6975 8313
rect 7009 8347 7067 8353
rect 7009 8313 7021 8347
rect 7055 8344 7067 8347
rect 7190 8344 7196 8356
rect 7055 8316 7196 8344
rect 7055 8313 7067 8316
rect 7009 8307 7067 8313
rect 4617 8279 4675 8285
rect 4617 8276 4629 8279
rect 4448 8248 4629 8276
rect 4120 8236 4126 8248
rect 4617 8245 4629 8248
rect 4663 8245 4675 8279
rect 6638 8276 6644 8288
rect 6599 8248 6644 8276
rect 4617 8239 4675 8245
rect 6638 8236 6644 8248
rect 6696 8236 6702 8288
rect 6932 8276 6960 8307
rect 7190 8304 7196 8316
rect 7248 8304 7254 8356
rect 9027 8347 9085 8353
rect 9027 8313 9039 8347
rect 9073 8344 9085 8347
rect 9674 8344 9680 8356
rect 9073 8316 9680 8344
rect 9073 8313 9085 8316
rect 9027 8307 9085 8313
rect 9674 8304 9680 8316
rect 9732 8304 9738 8356
rect 10778 8344 10784 8356
rect 10739 8316 10784 8344
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 10870 8304 10876 8356
rect 10928 8344 10934 8356
rect 10928 8316 10973 8344
rect 10928 8304 10934 8316
rect 12710 8304 12716 8356
rect 12768 8344 12774 8356
rect 13126 8347 13184 8353
rect 13126 8344 13138 8347
rect 12768 8316 13138 8344
rect 12768 8304 12774 8316
rect 13126 8313 13138 8316
rect 13172 8313 13184 8347
rect 14645 8347 14703 8353
rect 14645 8344 14657 8347
rect 13126 8307 13184 8313
rect 14568 8316 14657 8344
rect 7098 8276 7104 8288
rect 6932 8248 7104 8276
rect 7098 8236 7104 8248
rect 7156 8236 7162 8288
rect 10597 8279 10655 8285
rect 10597 8245 10609 8279
rect 10643 8276 10655 8279
rect 10888 8276 10916 8304
rect 14568 8288 14596 8316
rect 14645 8313 14657 8316
rect 14691 8313 14703 8347
rect 14645 8307 14703 8313
rect 14734 8304 14740 8356
rect 14792 8344 14798 8356
rect 16132 8344 16160 8375
rect 17310 8372 17316 8384
rect 17368 8372 17374 8424
rect 18156 8421 18184 8452
rect 18141 8415 18199 8421
rect 18141 8381 18153 8415
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 19680 8415 19738 8421
rect 19680 8381 19692 8415
rect 19726 8412 19738 8415
rect 19794 8412 19800 8424
rect 19726 8384 19800 8412
rect 19726 8381 19738 8384
rect 19680 8375 19738 8381
rect 19794 8372 19800 8384
rect 19852 8412 19858 8424
rect 20073 8415 20131 8421
rect 20073 8412 20085 8415
rect 19852 8384 20085 8412
rect 19852 8372 19858 8384
rect 20073 8381 20085 8384
rect 20119 8381 20131 8415
rect 20073 8375 20131 8381
rect 16482 8344 16488 8356
rect 14792 8316 14837 8344
rect 16132 8316 16488 8344
rect 14792 8304 14798 8316
rect 16482 8304 16488 8316
rect 16540 8344 16546 8356
rect 17034 8344 17040 8356
rect 16540 8316 17040 8344
rect 16540 8304 16546 8316
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 17218 8304 17224 8356
rect 17276 8344 17282 8356
rect 19150 8344 19156 8356
rect 17276 8316 19156 8344
rect 17276 8304 17282 8316
rect 19150 8304 19156 8316
rect 19208 8344 19214 8356
rect 19429 8347 19487 8353
rect 19429 8344 19441 8347
rect 19208 8316 19441 8344
rect 19208 8304 19214 8316
rect 19429 8313 19441 8316
rect 19475 8313 19487 8347
rect 19429 8307 19487 8313
rect 10643 8248 10916 8276
rect 10643 8245 10655 8248
rect 10597 8239 10655 8245
rect 14182 8236 14188 8288
rect 14240 8276 14246 8288
rect 14366 8276 14372 8288
rect 14240 8248 14372 8276
rect 14240 8236 14246 8248
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 14550 8236 14556 8288
rect 14608 8236 14614 8288
rect 16206 8276 16212 8288
rect 16167 8248 16212 8276
rect 16206 8236 16212 8248
rect 16264 8236 16270 8288
rect 18414 8236 18420 8288
rect 18472 8276 18478 8288
rect 18509 8279 18567 8285
rect 18509 8276 18521 8279
rect 18472 8248 18521 8276
rect 18472 8236 18478 8248
rect 18509 8245 18521 8248
rect 18555 8245 18567 8279
rect 18509 8239 18567 8245
rect 18966 8236 18972 8288
rect 19024 8276 19030 8288
rect 19061 8279 19119 8285
rect 19061 8276 19073 8279
rect 19024 8248 19073 8276
rect 19024 8236 19030 8248
rect 19061 8245 19073 8248
rect 19107 8245 19119 8279
rect 19061 8239 19119 8245
rect 1104 8186 20884 8208
rect 1104 8134 8315 8186
rect 8367 8134 8379 8186
rect 8431 8134 8443 8186
rect 8495 8134 8507 8186
rect 8559 8134 15648 8186
rect 15700 8134 15712 8186
rect 15764 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 20884 8186
rect 1104 8112 20884 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 2498 8072 2504 8084
rect 2411 8044 2504 8072
rect 2498 8032 2504 8044
rect 2556 8072 2562 8084
rect 3418 8072 3424 8084
rect 2556 8044 3424 8072
rect 2556 8032 2562 8044
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 3568 8044 4445 8072
rect 3568 8032 3574 8044
rect 4433 8041 4445 8044
rect 4479 8041 4491 8075
rect 5902 8072 5908 8084
rect 5863 8044 5908 8072
rect 4433 8035 4491 8041
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 7006 8032 7012 8084
rect 7064 8072 7070 8084
rect 11977 8075 12035 8081
rect 11977 8072 11989 8075
rect 7064 8044 11989 8072
rect 7064 8032 7070 8044
rect 11977 8041 11989 8044
rect 12023 8041 12035 8075
rect 11977 8035 12035 8041
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 14553 8075 14611 8081
rect 14553 8072 14565 8075
rect 13872 8044 14565 8072
rect 13872 8032 13878 8044
rect 14553 8041 14565 8044
rect 14599 8072 14611 8075
rect 14734 8072 14740 8084
rect 14599 8044 14740 8072
rect 14599 8041 14611 8044
rect 14553 8035 14611 8041
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 14829 8075 14887 8081
rect 14829 8041 14841 8075
rect 14875 8072 14887 8075
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14875 8044 15025 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 15013 8041 15025 8044
rect 15059 8072 15071 8075
rect 16850 8072 16856 8084
rect 15059 8044 16856 8072
rect 15059 8041 15071 8044
rect 15013 8035 15071 8041
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 18230 8032 18236 8084
rect 18288 8072 18294 8084
rect 19061 8075 19119 8081
rect 19061 8072 19073 8075
rect 18288 8044 19073 8072
rect 18288 8032 18294 8044
rect 19061 8041 19073 8044
rect 19107 8041 19119 8075
rect 19061 8035 19119 8041
rect 1302 7964 1308 8016
rect 1360 8004 1366 8016
rect 2777 8007 2835 8013
rect 2777 8004 2789 8007
rect 1360 7976 2789 8004
rect 1360 7964 1366 7976
rect 2777 7973 2789 7976
rect 2823 7973 2835 8007
rect 2777 7967 2835 7973
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7905 1639 7939
rect 1581 7899 1639 7905
rect 1596 7868 1624 7899
rect 1670 7896 1676 7948
rect 1728 7936 1734 7948
rect 1949 7939 2007 7945
rect 1949 7936 1961 7939
rect 1728 7908 1961 7936
rect 1728 7896 1734 7908
rect 1949 7905 1961 7908
rect 1995 7936 2007 7939
rect 2498 7936 2504 7948
rect 1995 7908 2504 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 1762 7868 1768 7880
rect 1596 7840 1768 7868
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 2792 7800 2820 7967
rect 3878 7964 3884 8016
rect 3936 8004 3942 8016
rect 5353 8007 5411 8013
rect 5353 8004 5365 8007
rect 3936 7976 5365 8004
rect 3936 7964 3942 7976
rect 5353 7973 5365 7976
rect 5399 7973 5411 8007
rect 7469 8007 7527 8013
rect 7469 8004 7481 8007
rect 5353 7967 5411 7973
rect 6472 7976 7481 8004
rect 3028 7939 3086 7945
rect 3028 7905 3040 7939
rect 3074 7936 3086 7939
rect 3142 7936 3148 7948
rect 3074 7908 3148 7936
rect 3074 7905 3086 7908
rect 3028 7899 3086 7905
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 4157 7939 4215 7945
rect 4157 7905 4169 7939
rect 4203 7905 4215 7939
rect 4157 7899 4215 7905
rect 4172 7868 4200 7899
rect 4338 7896 4344 7948
rect 4396 7936 4402 7948
rect 5074 7936 5080 7948
rect 4396 7908 5080 7936
rect 4396 7896 4402 7908
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 6472 7945 6500 7976
rect 7469 7973 7481 7976
rect 7515 8004 7527 8007
rect 8478 8004 8484 8016
rect 7515 7976 8484 8004
rect 7515 7973 7527 7976
rect 7469 7967 7527 7973
rect 8478 7964 8484 7976
rect 8536 7964 8542 8016
rect 9493 8007 9551 8013
rect 9493 7973 9505 8007
rect 9539 8004 9551 8007
rect 9766 8004 9772 8016
rect 9539 7976 9772 8004
rect 9539 7973 9551 7976
rect 9493 7967 9551 7973
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 10090 8007 10148 8013
rect 10090 7973 10102 8007
rect 10136 7973 10148 8007
rect 11330 8004 11336 8016
rect 11291 7976 11336 8004
rect 10090 7967 10148 7973
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7905 6515 7939
rect 6457 7899 6515 7905
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 9674 7936 9680 7948
rect 8803 7908 9680 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 9674 7896 9680 7908
rect 9732 7936 9738 7948
rect 10105 7936 10133 7967
rect 11330 7964 11336 7976
rect 11388 7964 11394 8016
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 13034 8007 13092 8013
rect 13034 8004 13046 8007
rect 12768 7976 13046 8004
rect 12768 7964 12774 7976
rect 13034 7973 13046 7976
rect 13080 8004 13092 8007
rect 13262 8004 13268 8016
rect 13080 7976 13268 8004
rect 13080 7973 13092 7976
rect 13034 7967 13092 7973
rect 13262 7964 13268 7976
rect 13320 7964 13326 8016
rect 13906 8004 13912 8016
rect 13648 7976 13912 8004
rect 11422 7936 11428 7948
rect 9732 7908 10133 7936
rect 11383 7908 11428 7936
rect 9732 7896 9738 7908
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 13648 7945 13676 7976
rect 13906 7964 13912 7976
rect 13964 8004 13970 8016
rect 14001 8007 14059 8013
rect 14001 8004 14013 8007
rect 13964 7976 14013 8004
rect 13964 7964 13970 7976
rect 14001 7973 14013 7976
rect 14047 8004 14059 8007
rect 15473 8007 15531 8013
rect 15473 8004 15485 8007
rect 14047 7976 15485 8004
rect 14047 7973 14059 7976
rect 14001 7967 14059 7973
rect 15473 7973 15485 7976
rect 15519 8004 15531 8007
rect 16298 8004 16304 8016
rect 15519 7976 16304 8004
rect 15519 7973 15531 7976
rect 15473 7967 15531 7973
rect 16298 7964 16304 7976
rect 16356 7964 16362 8016
rect 16758 8004 16764 8016
rect 16719 7976 16764 8004
rect 16758 7964 16764 7976
rect 16816 8004 16822 8016
rect 17218 8004 17224 8016
rect 16816 7976 17224 8004
rect 16816 7964 16822 7976
rect 17218 7964 17224 7976
rect 17276 7964 17282 8016
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 14550 7896 14556 7948
rect 14608 7936 14614 7948
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 14608 7908 14841 7936
rect 14608 7896 14614 7908
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7936 16175 7939
rect 16574 7936 16580 7948
rect 16163 7908 16580 7936
rect 16163 7905 16175 7908
rect 16117 7899 16175 7905
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 16666 7896 16672 7948
rect 16724 7936 16730 7948
rect 16945 7939 17003 7945
rect 16945 7936 16957 7939
rect 16724 7908 16957 7936
rect 16724 7896 16730 7908
rect 16945 7905 16957 7908
rect 16991 7905 17003 7939
rect 16945 7899 17003 7905
rect 18417 7939 18475 7945
rect 18417 7905 18429 7939
rect 18463 7905 18475 7939
rect 18417 7899 18475 7905
rect 4172 7840 5120 7868
rect 4982 7800 4988 7812
rect 2792 7772 4988 7800
rect 4982 7760 4988 7772
rect 5040 7760 5046 7812
rect 3234 7732 3240 7744
rect 3195 7704 3240 7732
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 3881 7735 3939 7741
rect 3881 7701 3893 7735
rect 3927 7732 3939 7735
rect 4430 7732 4436 7744
rect 3927 7704 4436 7732
rect 3927 7701 3939 7704
rect 3881 7695 3939 7701
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 5092 7741 5120 7840
rect 5442 7828 5448 7880
rect 5500 7868 5506 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5500 7840 5549 7868
rect 5500 7828 5506 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7868 7435 7871
rect 7558 7868 7564 7880
rect 7423 7840 7564 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 9766 7868 9772 7880
rect 7708 7840 7753 7868
rect 9727 7840 9772 7868
rect 7708 7828 7714 7840
rect 9766 7828 9772 7840
rect 9824 7828 9830 7880
rect 12710 7868 12716 7880
rect 12671 7840 12716 7868
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15381 7871 15439 7877
rect 15381 7868 15393 7871
rect 15252 7840 15393 7868
rect 15252 7828 15258 7840
rect 15381 7837 15393 7840
rect 15427 7837 15439 7871
rect 15381 7831 15439 7837
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 16853 7871 16911 7877
rect 16853 7868 16865 7871
rect 15528 7840 16865 7868
rect 15528 7828 15534 7840
rect 16853 7837 16865 7840
rect 16899 7837 16911 7871
rect 16853 7831 16911 7837
rect 6917 7803 6975 7809
rect 6917 7769 6929 7803
rect 6963 7800 6975 7803
rect 7190 7800 7196 7812
rect 6963 7772 7196 7800
rect 6963 7769 6975 7772
rect 6917 7763 6975 7769
rect 7190 7760 7196 7772
rect 7248 7800 7254 7812
rect 9122 7800 9128 7812
rect 7248 7772 9128 7800
rect 7248 7760 7254 7772
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 10689 7803 10747 7809
rect 10689 7769 10701 7803
rect 10735 7800 10747 7803
rect 10870 7800 10876 7812
rect 10735 7772 10876 7800
rect 10735 7769 10747 7772
rect 10689 7763 10747 7769
rect 10870 7760 10876 7772
rect 10928 7800 10934 7812
rect 11330 7800 11336 7812
rect 10928 7772 11336 7800
rect 10928 7760 10934 7772
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 15286 7760 15292 7812
rect 15344 7800 15350 7812
rect 18432 7800 18460 7899
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 18874 7868 18880 7880
rect 18831 7840 18880 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 19150 7800 19156 7812
rect 15344 7772 19156 7800
rect 15344 7760 15350 7772
rect 19150 7760 19156 7772
rect 19208 7760 19214 7812
rect 5077 7735 5135 7741
rect 5077 7701 5089 7735
rect 5123 7732 5135 7735
rect 5166 7732 5172 7744
rect 5123 7704 5172 7732
rect 5123 7701 5135 7704
rect 5077 7695 5135 7701
rect 5166 7692 5172 7704
rect 5224 7692 5230 7744
rect 5258 7692 5264 7744
rect 5316 7732 5322 7744
rect 7650 7732 7656 7744
rect 5316 7704 7656 7732
rect 5316 7692 5322 7704
rect 7650 7692 7656 7704
rect 7708 7692 7714 7744
rect 8389 7735 8447 7741
rect 8389 7701 8401 7735
rect 8435 7732 8447 7735
rect 8478 7732 8484 7744
rect 8435 7704 8484 7732
rect 8435 7701 8447 7704
rect 8389 7695 8447 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 9030 7732 9036 7744
rect 8991 7704 9036 7732
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 11514 7692 11520 7744
rect 11572 7732 11578 7744
rect 11655 7735 11713 7741
rect 11655 7732 11667 7735
rect 11572 7704 11667 7732
rect 11572 7692 11578 7704
rect 11655 7701 11667 7704
rect 11701 7701 11713 7735
rect 11655 7695 11713 7701
rect 15010 7692 15016 7744
rect 15068 7732 15074 7744
rect 15562 7732 15568 7744
rect 15068 7704 15568 7732
rect 15068 7692 15074 7704
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 16301 7735 16359 7741
rect 16301 7732 16313 7735
rect 15804 7704 16313 7732
rect 15804 7692 15810 7704
rect 16301 7701 16313 7704
rect 16347 7732 16359 7735
rect 16482 7732 16488 7744
rect 16347 7704 16488 7732
rect 16347 7701 16359 7704
rect 16301 7695 16359 7701
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 18414 7692 18420 7744
rect 18472 7732 18478 7744
rect 18555 7735 18613 7741
rect 18555 7732 18567 7735
rect 18472 7704 18567 7732
rect 18472 7692 18478 7704
rect 18555 7701 18567 7704
rect 18601 7701 18613 7735
rect 18555 7695 18613 7701
rect 18693 7735 18751 7741
rect 18693 7701 18705 7735
rect 18739 7732 18751 7735
rect 18782 7732 18788 7744
rect 18739 7704 18788 7732
rect 18739 7701 18751 7704
rect 18693 7695 18751 7701
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 1104 7642 20884 7664
rect 1104 7590 4648 7642
rect 4700 7590 4712 7642
rect 4764 7590 4776 7642
rect 4828 7590 4840 7642
rect 4892 7590 11982 7642
rect 12034 7590 12046 7642
rect 12098 7590 12110 7642
rect 12162 7590 12174 7642
rect 12226 7590 19315 7642
rect 19367 7590 19379 7642
rect 19431 7590 19443 7642
rect 19495 7590 19507 7642
rect 19559 7590 20884 7642
rect 1104 7568 20884 7590
rect 1670 7528 1676 7540
rect 1631 7500 1676 7528
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 9030 7528 9036 7540
rect 2096 7500 9036 7528
rect 2096 7488 2102 7500
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 9732 7500 9777 7528
rect 9732 7488 9738 7500
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 12713 7531 12771 7537
rect 12713 7528 12725 7531
rect 10284 7500 12725 7528
rect 10284 7488 10290 7500
rect 12713 7497 12725 7500
rect 12759 7528 12771 7531
rect 12897 7531 12955 7537
rect 12897 7528 12909 7531
rect 12759 7500 12909 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 12897 7497 12909 7500
rect 12943 7497 12955 7531
rect 13262 7528 13268 7540
rect 13223 7500 13268 7528
rect 12897 7491 12955 7497
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 16298 7528 16304 7540
rect 16259 7500 16304 7528
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 3053 7463 3111 7469
rect 3053 7429 3065 7463
rect 3099 7460 3111 7463
rect 3142 7460 3148 7472
rect 3099 7432 3148 7460
rect 3099 7429 3111 7432
rect 3053 7423 3111 7429
rect 3142 7420 3148 7432
rect 3200 7420 3206 7472
rect 3786 7420 3792 7472
rect 3844 7460 3850 7472
rect 3973 7463 4031 7469
rect 3973 7460 3985 7463
rect 3844 7432 3985 7460
rect 3844 7420 3850 7432
rect 3973 7429 3985 7432
rect 4019 7460 4031 7463
rect 4062 7460 4068 7472
rect 4019 7432 4068 7460
rect 4019 7429 4031 7432
rect 3973 7423 4031 7429
rect 4062 7420 4068 7432
rect 4120 7460 4126 7472
rect 4203 7463 4261 7469
rect 4203 7460 4215 7463
rect 4120 7432 4215 7460
rect 4120 7420 4126 7432
rect 4203 7429 4215 7432
rect 4249 7429 4261 7463
rect 4203 7423 4261 7429
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7429 4399 7463
rect 5074 7460 5080 7472
rect 5035 7432 5080 7460
rect 4341 7423 4399 7429
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7392 3663 7395
rect 3651 7364 4154 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 2130 7284 2136 7336
rect 2188 7324 2194 7336
rect 2409 7327 2467 7333
rect 2409 7324 2421 7327
rect 2188 7296 2421 7324
rect 2188 7284 2194 7296
rect 2409 7293 2421 7296
rect 2455 7324 2467 7327
rect 3878 7324 3884 7336
rect 2455 7296 3884 7324
rect 2455 7293 2467 7296
rect 2409 7287 2467 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 4126 7324 4154 7364
rect 4246 7324 4252 7336
rect 4126 7296 4252 7324
rect 4246 7284 4252 7296
rect 4304 7324 4310 7336
rect 4356 7324 4384 7423
rect 5074 7420 5080 7432
rect 5132 7420 5138 7472
rect 5629 7463 5687 7469
rect 5629 7429 5641 7463
rect 5675 7460 5687 7463
rect 5902 7460 5908 7472
rect 5675 7432 5908 7460
rect 5675 7429 5687 7432
rect 5629 7423 5687 7429
rect 5902 7420 5908 7432
rect 5960 7420 5966 7472
rect 9766 7420 9772 7472
rect 9824 7460 9830 7472
rect 10965 7463 11023 7469
rect 10965 7460 10977 7463
rect 9824 7432 10977 7460
rect 9824 7420 9830 7432
rect 10965 7429 10977 7432
rect 11011 7460 11023 7463
rect 16022 7460 16028 7472
rect 11011 7432 16028 7460
rect 11011 7429 11023 7432
rect 10965 7423 11023 7429
rect 16022 7420 16028 7432
rect 16080 7420 16086 7472
rect 4430 7352 4436 7404
rect 4488 7392 4494 7404
rect 4801 7395 4859 7401
rect 4488 7364 4533 7392
rect 4488 7352 4494 7364
rect 4801 7361 4813 7395
rect 4847 7392 4859 7395
rect 9214 7392 9220 7404
rect 4847 7364 9220 7392
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 9490 7352 9496 7404
rect 9548 7392 9554 7404
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9548 7364 9965 7392
rect 9548 7352 9554 7364
rect 9953 7361 9965 7364
rect 9999 7392 10011 7395
rect 11514 7392 11520 7404
rect 9999 7364 11520 7392
rect 9999 7361 10011 7364
rect 9953 7355 10011 7361
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 13814 7392 13820 7404
rect 13775 7364 13820 7392
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14918 7392 14924 7404
rect 14507 7364 14924 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 15243 7364 15884 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 5626 7324 5632 7336
rect 4304 7296 5632 7324
rect 4304 7284 4310 7296
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 5772 7327 5830 7333
rect 5772 7293 5784 7327
rect 5818 7324 5830 7327
rect 6181 7327 6239 7333
rect 6181 7324 6193 7327
rect 5818 7296 6193 7324
rect 5818 7293 5830 7296
rect 5772 7287 5830 7293
rect 6181 7293 6193 7296
rect 6227 7324 6239 7327
rect 6454 7324 6460 7336
rect 6227 7296 6460 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 6454 7284 6460 7296
rect 6512 7284 6518 7336
rect 7834 7284 7840 7336
rect 7892 7324 7898 7336
rect 8297 7327 8355 7333
rect 8297 7324 8309 7327
rect 7892 7296 8309 7324
rect 7892 7284 7898 7296
rect 8297 7293 8309 7296
rect 8343 7324 8355 7327
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 8343 7296 8585 7324
rect 8343 7293 8355 7296
rect 8297 7287 8355 7293
rect 8573 7293 8585 7296
rect 8619 7324 8631 7327
rect 8662 7324 8668 7336
rect 8619 7296 8668 7324
rect 8619 7293 8631 7296
rect 8573 7287 8631 7293
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7324 8999 7327
rect 9306 7324 9312 7336
rect 8987 7296 9312 7324
rect 8987 7293 8999 7296
rect 8941 7287 8999 7293
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 12504 7327 12562 7333
rect 12504 7293 12516 7327
rect 12550 7324 12562 7327
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 12550 7296 12725 7324
rect 12550 7293 12562 7296
rect 12504 7287 12562 7293
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 15289 7327 15347 7333
rect 15289 7324 15301 7327
rect 12713 7287 12771 7293
rect 14568 7296 15301 7324
rect 1762 7256 1768 7268
rect 1723 7228 1768 7256
rect 1762 7216 1768 7228
rect 1820 7216 1826 7268
rect 4065 7259 4123 7265
rect 4065 7225 4077 7259
rect 4111 7225 4123 7259
rect 4065 7219 4123 7225
rect 5859 7259 5917 7265
rect 5859 7225 5871 7259
rect 5905 7256 5917 7259
rect 6914 7256 6920 7268
rect 5905 7228 6920 7256
rect 5905 7225 5917 7228
rect 5859 7219 5917 7225
rect 3970 7148 3976 7200
rect 4028 7188 4034 7200
rect 4080 7188 4108 7219
rect 6914 7216 6920 7228
rect 6972 7216 6978 7268
rect 7006 7216 7012 7268
rect 7064 7256 7070 7268
rect 7558 7256 7564 7268
rect 7064 7228 7109 7256
rect 7519 7228 7564 7256
rect 7064 7216 7070 7228
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 7742 7216 7748 7268
rect 7800 7256 7806 7268
rect 8389 7259 8447 7265
rect 8389 7256 8401 7259
rect 7800 7228 8401 7256
rect 7800 7216 7806 7228
rect 8389 7225 8401 7228
rect 8435 7225 8447 7259
rect 8389 7219 8447 7225
rect 4338 7188 4344 7200
rect 4028 7160 4344 7188
rect 4028 7148 4034 7160
rect 4338 7148 4344 7160
rect 4396 7148 4402 7200
rect 6546 7188 6552 7200
rect 6507 7160 6552 7188
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 6638 7148 6644 7200
rect 6696 7188 6702 7200
rect 7837 7191 7895 7197
rect 7837 7188 7849 7191
rect 6696 7160 7849 7188
rect 6696 7148 6702 7160
rect 7837 7157 7849 7160
rect 7883 7157 7895 7191
rect 8404 7188 8432 7219
rect 8478 7216 8484 7268
rect 8536 7256 8542 7268
rect 9030 7256 9036 7268
rect 8536 7228 9036 7256
rect 8536 7216 8542 7228
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 10042 7256 10048 7268
rect 10003 7228 10048 7256
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 10594 7256 10600 7268
rect 10555 7228 10600 7256
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 11422 7216 11428 7268
rect 11480 7256 11486 7268
rect 11609 7259 11667 7265
rect 11609 7256 11621 7259
rect 11480 7228 11621 7256
rect 11480 7216 11486 7228
rect 11609 7225 11621 7228
rect 11655 7256 11667 7259
rect 13906 7256 13912 7268
rect 11655 7228 13400 7256
rect 13867 7228 13912 7256
rect 11655 7225 11667 7228
rect 11609 7219 11667 7225
rect 9309 7191 9367 7197
rect 9309 7188 9321 7191
rect 8404 7160 9321 7188
rect 7837 7151 7895 7157
rect 9309 7157 9321 7160
rect 9355 7188 9367 7191
rect 9398 7188 9404 7200
rect 9355 7160 9404 7188
rect 9355 7157 9367 7160
rect 9309 7151 9367 7157
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 12575 7191 12633 7197
rect 12575 7188 12587 7191
rect 9824 7160 12587 7188
rect 9824 7148 9830 7160
rect 12575 7157 12587 7160
rect 12621 7157 12633 7191
rect 13372 7188 13400 7228
rect 13906 7216 13912 7228
rect 13964 7216 13970 7268
rect 14568 7200 14596 7296
rect 15289 7293 15301 7296
rect 15335 7324 15347 7327
rect 15746 7324 15752 7336
rect 15335 7296 15752 7324
rect 15335 7293 15347 7296
rect 15289 7287 15347 7293
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 15856 7333 15884 7364
rect 16390 7352 16396 7404
rect 16448 7392 16454 7404
rect 18049 7395 18107 7401
rect 18049 7392 18061 7395
rect 16448 7364 18061 7392
rect 16448 7352 16454 7364
rect 18049 7361 18061 7364
rect 18095 7392 18107 7395
rect 18782 7392 18788 7404
rect 18095 7364 18788 7392
rect 18095 7361 18107 7364
rect 18049 7355 18107 7361
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 15841 7327 15899 7333
rect 15841 7293 15853 7327
rect 15887 7324 15899 7327
rect 15930 7324 15936 7336
rect 15887 7296 15936 7324
rect 15887 7293 15899 7296
rect 15841 7287 15899 7293
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 16574 7284 16580 7336
rect 16632 7324 16638 7336
rect 16888 7327 16946 7333
rect 16888 7324 16900 7327
rect 16632 7296 16900 7324
rect 16632 7284 16638 7296
rect 16888 7293 16900 7296
rect 16934 7324 16946 7327
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 16934 7296 17325 7324
rect 16934 7293 16946 7296
rect 16888 7287 16946 7293
rect 17313 7293 17325 7296
rect 17359 7293 17371 7327
rect 17770 7324 17776 7336
rect 17731 7296 17776 7324
rect 17313 7287 17371 7293
rect 17770 7284 17776 7296
rect 17828 7324 17834 7336
rect 18141 7327 18199 7333
rect 18141 7324 18153 7327
rect 17828 7296 18153 7324
rect 17828 7284 17834 7296
rect 18141 7293 18153 7296
rect 18187 7293 18199 7327
rect 18141 7287 18199 7293
rect 18414 7284 18420 7336
rect 18472 7324 18478 7336
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 18472 7296 19441 7324
rect 18472 7284 18478 7296
rect 19429 7293 19441 7296
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 14642 7216 14648 7268
rect 14700 7256 14706 7268
rect 14700 7228 15332 7256
rect 14700 7216 14706 7228
rect 14274 7188 14280 7200
rect 13372 7160 14280 7188
rect 12575 7151 12633 7157
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 14550 7148 14556 7200
rect 14608 7188 14614 7200
rect 14737 7191 14795 7197
rect 14737 7188 14749 7191
rect 14608 7160 14749 7188
rect 14608 7148 14614 7160
rect 14737 7157 14749 7160
rect 14783 7157 14795 7191
rect 15304 7188 15332 7228
rect 16758 7216 16764 7268
rect 16816 7256 16822 7268
rect 19613 7259 19671 7265
rect 19613 7256 19625 7259
rect 16816 7228 19625 7256
rect 16816 7216 16822 7228
rect 19613 7225 19625 7228
rect 19659 7225 19671 7259
rect 19613 7219 19671 7225
rect 15381 7191 15439 7197
rect 15381 7188 15393 7191
rect 15304 7160 15393 7188
rect 14737 7151 14795 7157
rect 15381 7157 15393 7160
rect 15427 7157 15439 7191
rect 16666 7188 16672 7200
rect 16627 7160 16672 7188
rect 15381 7151 15439 7157
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 16850 7148 16856 7200
rect 16908 7188 16914 7200
rect 16991 7191 17049 7197
rect 16991 7188 17003 7191
rect 16908 7160 17003 7188
rect 16908 7148 16914 7160
rect 16991 7157 17003 7160
rect 17037 7157 17049 7191
rect 16991 7151 17049 7157
rect 17126 7148 17132 7200
rect 17184 7188 17190 7200
rect 18874 7188 18880 7200
rect 17184 7160 18880 7188
rect 17184 7148 17190 7160
rect 18874 7148 18880 7160
rect 18932 7188 18938 7200
rect 19061 7191 19119 7197
rect 19061 7188 19073 7191
rect 18932 7160 19073 7188
rect 18932 7148 18938 7160
rect 19061 7157 19073 7160
rect 19107 7157 19119 7191
rect 19061 7151 19119 7157
rect 1104 7098 20884 7120
rect 1104 7046 8315 7098
rect 8367 7046 8379 7098
rect 8431 7046 8443 7098
rect 8495 7046 8507 7098
rect 8559 7046 15648 7098
rect 15700 7046 15712 7098
rect 15764 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 20884 7098
rect 1104 7024 20884 7046
rect 1854 6944 1860 6996
rect 1912 6984 1918 6996
rect 2961 6987 3019 6993
rect 2961 6984 2973 6987
rect 1912 6956 2973 6984
rect 1912 6944 1918 6956
rect 2961 6953 2973 6956
rect 3007 6984 3019 6987
rect 4982 6984 4988 6996
rect 3007 6956 4988 6984
rect 3007 6953 3019 6956
rect 2961 6947 3019 6953
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 5166 6984 5172 6996
rect 5079 6956 5172 6984
rect 5166 6944 5172 6956
rect 5224 6984 5230 6996
rect 7742 6984 7748 6996
rect 5224 6956 7748 6984
rect 5224 6944 5230 6956
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 9490 6984 9496 6996
rect 9451 6956 9496 6984
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 10042 6944 10048 6996
rect 10100 6984 10106 6996
rect 10689 6987 10747 6993
rect 10689 6984 10701 6987
rect 10100 6956 10701 6984
rect 10100 6944 10106 6956
rect 10689 6953 10701 6956
rect 10735 6953 10747 6987
rect 12710 6984 12716 6996
rect 12671 6956 12716 6984
rect 10689 6947 10747 6953
rect 12710 6944 12716 6956
rect 12768 6944 12774 6996
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14645 6987 14703 6993
rect 14645 6984 14657 6987
rect 13872 6956 14657 6984
rect 13872 6944 13878 6956
rect 14645 6953 14657 6956
rect 14691 6984 14703 6987
rect 16850 6984 16856 6996
rect 14691 6956 16856 6984
rect 14691 6953 14703 6956
rect 14645 6947 14703 6953
rect 16850 6944 16856 6956
rect 16908 6944 16914 6996
rect 18782 6944 18788 6996
rect 18840 6984 18846 6996
rect 18877 6987 18935 6993
rect 18877 6984 18889 6987
rect 18840 6956 18889 6984
rect 18840 6944 18846 6956
rect 18877 6953 18889 6956
rect 18923 6953 18935 6987
rect 18877 6947 18935 6953
rect 19150 6944 19156 6996
rect 19208 6984 19214 6996
rect 19245 6987 19303 6993
rect 19245 6984 19257 6987
rect 19208 6956 19257 6984
rect 19208 6944 19214 6956
rect 19245 6953 19257 6956
rect 19291 6953 19303 6987
rect 19245 6947 19303 6953
rect 1762 6916 1768 6928
rect 1723 6888 1768 6916
rect 1762 6876 1768 6888
rect 1820 6876 1826 6928
rect 5902 6916 5908 6928
rect 5863 6888 5908 6916
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 6730 6876 6736 6928
rect 6788 6916 6794 6928
rect 7098 6916 7104 6928
rect 6788 6888 7104 6916
rect 6788 6876 6794 6888
rect 7098 6876 7104 6888
rect 7156 6876 7162 6928
rect 8754 6916 8760 6928
rect 7208 6888 8760 6916
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 5350 6848 5356 6860
rect 4111 6820 5356 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 5350 6808 5356 6820
rect 5408 6848 5414 6860
rect 5445 6851 5503 6857
rect 5445 6848 5457 6851
rect 5408 6820 5457 6848
rect 5408 6808 5414 6820
rect 5445 6817 5457 6820
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 5718 6848 5724 6860
rect 5675 6820 5724 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 5718 6808 5724 6820
rect 5776 6848 5782 6860
rect 6638 6848 6644 6860
rect 5776 6820 6644 6848
rect 5776 6808 5782 6820
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1719 6752 3464 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 1118 6672 1124 6724
rect 1176 6712 1182 6724
rect 2225 6715 2283 6721
rect 2225 6712 2237 6715
rect 1176 6684 2237 6712
rect 1176 6672 1182 6684
rect 2225 6681 2237 6684
rect 2271 6712 2283 6715
rect 2314 6712 2320 6724
rect 2271 6684 2320 6712
rect 2271 6681 2283 6684
rect 2225 6675 2283 6681
rect 2314 6672 2320 6684
rect 2372 6672 2378 6724
rect 3436 6656 3464 6752
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4212 6783 4270 6789
rect 4212 6780 4224 6783
rect 4028 6752 4224 6780
rect 4028 6740 4034 6752
rect 4212 6749 4224 6752
rect 4258 6749 4270 6783
rect 4430 6780 4436 6792
rect 4343 6752 4436 6780
rect 4212 6743 4270 6749
rect 4430 6740 4436 6752
rect 4488 6780 4494 6792
rect 7208 6780 7236 6888
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 9858 6916 9864 6928
rect 9819 6888 9864 6916
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 10413 6919 10471 6925
rect 10413 6885 10425 6919
rect 10459 6916 10471 6919
rect 10594 6916 10600 6928
rect 10459 6888 10600 6916
rect 10459 6885 10471 6888
rect 10413 6879 10471 6885
rect 10594 6876 10600 6888
rect 10652 6876 10658 6928
rect 11330 6876 11336 6928
rect 11388 6916 11394 6928
rect 11425 6919 11483 6925
rect 11425 6916 11437 6919
rect 11388 6888 11437 6916
rect 11388 6876 11394 6888
rect 11425 6885 11437 6888
rect 11471 6885 11483 6919
rect 13722 6916 13728 6928
rect 13683 6888 13728 6916
rect 11425 6879 11483 6885
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 15105 6919 15163 6925
rect 15105 6885 15117 6919
rect 15151 6916 15163 6919
rect 15194 6916 15200 6928
rect 15151 6888 15200 6916
rect 15151 6885 15163 6888
rect 15105 6879 15163 6885
rect 15194 6876 15200 6888
rect 15252 6916 15258 6928
rect 18555 6919 18613 6925
rect 18555 6916 18567 6919
rect 15252 6888 18567 6916
rect 15252 6876 15258 6888
rect 18555 6885 18567 6888
rect 18601 6885 18613 6919
rect 18555 6879 18613 6885
rect 7469 6851 7527 6857
rect 7469 6848 7481 6851
rect 4488 6752 7236 6780
rect 7300 6820 7481 6848
rect 4488 6740 4494 6752
rect 4062 6672 4068 6724
rect 4120 6712 4126 6724
rect 4525 6715 4583 6721
rect 4525 6712 4537 6715
rect 4120 6684 4537 6712
rect 4120 6672 4126 6684
rect 4525 6681 4537 6684
rect 4571 6681 4583 6715
rect 4525 6675 4583 6681
rect 5074 6672 5080 6724
rect 5132 6712 5138 6724
rect 5132 6684 6960 6712
rect 5132 6672 5138 6684
rect 6932 6656 6960 6684
rect 2682 6644 2688 6656
rect 2643 6616 2688 6644
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 3418 6644 3424 6656
rect 3379 6616 3424 6644
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3878 6644 3884 6656
rect 3839 6616 3884 6644
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 4341 6647 4399 6653
rect 4341 6644 4353 6647
rect 4304 6616 4353 6644
rect 4304 6604 4310 6616
rect 4341 6613 4353 6616
rect 4387 6613 4399 6647
rect 6546 6644 6552 6656
rect 6507 6616 6552 6644
rect 4341 6607 4399 6613
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 6822 6644 6828 6656
rect 6783 6616 6828 6644
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7300 6653 7328 6820
rect 7469 6817 7481 6820
rect 7515 6817 7527 6851
rect 7926 6848 7932 6860
rect 7887 6820 7932 6848
rect 7469 6811 7527 6817
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 15010 6808 15016 6860
rect 15068 6848 15074 6860
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 15068 6820 15301 6848
rect 15068 6808 15074 6820
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 15749 6851 15807 6857
rect 15749 6817 15761 6851
rect 15795 6848 15807 6851
rect 15930 6848 15936 6860
rect 15795 6820 15936 6848
rect 15795 6817 15807 6820
rect 15749 6811 15807 6817
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 16850 6848 16856 6860
rect 16811 6820 16856 6848
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 17126 6848 17132 6860
rect 17087 6820 17132 6848
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 18468 6851 18526 6857
rect 18468 6817 18480 6851
rect 18514 6848 18526 6851
rect 18690 6848 18696 6860
rect 18514 6820 18696 6848
rect 18514 6817 18526 6820
rect 18468 6811 18526 6817
rect 18690 6808 18696 6820
rect 18748 6808 18754 6860
rect 19496 6851 19554 6857
rect 19496 6817 19508 6851
rect 19542 6848 19554 6851
rect 19702 6848 19708 6860
rect 19542 6820 19708 6848
rect 19542 6817 19554 6820
rect 19496 6811 19554 6817
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 9214 6780 9220 6792
rect 8251 6752 9220 6780
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 11333 6783 11391 6789
rect 11333 6749 11345 6783
rect 11379 6780 11391 6783
rect 11422 6780 11428 6792
rect 11379 6752 11428 6780
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11606 6780 11612 6792
rect 11567 6752 11612 6780
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6780 13691 6783
rect 13814 6780 13820 6792
rect 13679 6752 13820 6780
rect 13679 6749 13691 6752
rect 13633 6743 13691 6749
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 13924 6752 15853 6780
rect 7558 6672 7564 6724
rect 7616 6712 7622 6724
rect 11057 6715 11115 6721
rect 11057 6712 11069 6715
rect 7616 6684 11069 6712
rect 7616 6672 7622 6684
rect 11057 6681 11069 6684
rect 11103 6681 11115 6715
rect 11057 6675 11115 6681
rect 12710 6672 12716 6724
rect 12768 6712 12774 6724
rect 13924 6712 13952 6752
rect 15841 6749 15853 6752
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 16942 6780 16948 6792
rect 16448 6752 16948 6780
rect 16448 6740 16454 6752
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 17310 6780 17316 6792
rect 17271 6752 17316 6780
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 12768 6684 13952 6712
rect 14185 6715 14243 6721
rect 12768 6672 12774 6684
rect 14185 6681 14197 6715
rect 14231 6712 14243 6715
rect 14458 6712 14464 6724
rect 14231 6684 14464 6712
rect 14231 6681 14243 6684
rect 14185 6675 14243 6681
rect 14458 6672 14464 6684
rect 14516 6672 14522 6724
rect 17034 6672 17040 6724
rect 17092 6712 17098 6724
rect 19567 6715 19625 6721
rect 19567 6712 19579 6715
rect 17092 6684 19579 6712
rect 17092 6672 17098 6684
rect 19567 6681 19579 6684
rect 19613 6681 19625 6715
rect 19567 6675 19625 6681
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 6972 6616 7297 6644
rect 6972 6604 6978 6616
rect 7285 6613 7297 6616
rect 7331 6613 7343 6647
rect 7285 6607 7343 6613
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 8662 6644 8668 6656
rect 8619 6616 8668 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 8846 6644 8852 6656
rect 8807 6616 8852 6644
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 18782 6644 18788 6656
rect 10836 6616 18788 6644
rect 10836 6604 10842 6616
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 1104 6554 20884 6576
rect 1104 6502 4648 6554
rect 4700 6502 4712 6554
rect 4764 6502 4776 6554
rect 4828 6502 4840 6554
rect 4892 6502 11982 6554
rect 12034 6502 12046 6554
rect 12098 6502 12110 6554
rect 12162 6502 12174 6554
rect 12226 6502 19315 6554
rect 19367 6502 19379 6554
rect 19431 6502 19443 6554
rect 19495 6502 19507 6554
rect 19559 6502 20884 6554
rect 1104 6480 20884 6502
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6440 1731 6443
rect 1762 6440 1768 6452
rect 1719 6412 1768 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 1762 6400 1768 6412
rect 1820 6400 1826 6452
rect 3694 6440 3700 6452
rect 3655 6412 3700 6440
rect 3694 6400 3700 6412
rect 3752 6400 3758 6452
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 5776 6412 5821 6440
rect 5776 6400 5782 6412
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5960 6412 6009 6440
rect 5960 6400 5966 6412
rect 5997 6409 6009 6412
rect 6043 6440 6055 6443
rect 8018 6440 8024 6452
rect 6043 6412 8024 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 11330 6440 11336 6452
rect 11291 6412 11336 6440
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 13262 6440 13268 6452
rect 12299 6412 13268 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 3421 6375 3479 6381
rect 3421 6341 3433 6375
rect 3467 6372 3479 6375
rect 3602 6372 3608 6384
rect 3467 6344 3608 6372
rect 3467 6341 3479 6344
rect 3421 6335 3479 6341
rect 2038 6304 2044 6316
rect 1999 6276 2044 6304
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 2314 6304 2320 6316
rect 2275 6276 2320 6304
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 3528 6245 3556 6344
rect 3602 6332 3608 6344
rect 3660 6332 3666 6384
rect 9125 6375 9183 6381
rect 9125 6341 9137 6375
rect 9171 6372 9183 6375
rect 9950 6372 9956 6384
rect 9171 6344 9956 6372
rect 9171 6341 9183 6344
rect 9125 6335 9183 6341
rect 9950 6332 9956 6344
rect 10008 6332 10014 6384
rect 5350 6304 5356 6316
rect 5311 6276 5356 6304
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 7374 6304 7380 6316
rect 7335 6276 7380 6304
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 10192 6276 10333 6304
rect 10192 6264 10198 6276
rect 10321 6273 10333 6276
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 3513 6239 3571 6245
rect 3513 6205 3525 6239
rect 3559 6205 3571 6239
rect 3513 6199 3571 6205
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6236 4951 6239
rect 5166 6236 5172 6248
rect 4939 6208 5172 6236
rect 4939 6205 4951 6208
rect 4893 6199 4951 6205
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6205 5503 6239
rect 5445 6199 5503 6205
rect 6549 6239 6607 6245
rect 6549 6205 6561 6239
rect 6595 6236 6607 6239
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6595 6208 7021 6236
rect 6595 6205 6607 6208
rect 6549 6199 6607 6205
rect 7009 6205 7021 6208
rect 7055 6236 7067 6239
rect 7190 6236 7196 6248
rect 7055 6208 7196 6236
rect 7055 6205 7067 6208
rect 7009 6199 7067 6205
rect 2130 6168 2136 6180
rect 2091 6140 2136 6168
rect 2130 6128 2136 6140
rect 2188 6128 2194 6180
rect 3050 6168 3056 6180
rect 2963 6140 3056 6168
rect 3050 6128 3056 6140
rect 3108 6168 3114 6180
rect 4430 6168 4436 6180
rect 3108 6140 4436 6168
rect 3108 6128 3114 6140
rect 4430 6128 4436 6140
rect 4488 6128 4494 6180
rect 4525 6171 4583 6177
rect 4525 6137 4537 6171
rect 4571 6168 4583 6171
rect 4982 6168 4988 6180
rect 4571 6140 4988 6168
rect 4571 6137 4583 6140
rect 4525 6131 4583 6137
rect 4982 6128 4988 6140
rect 5040 6168 5046 6180
rect 5460 6168 5488 6199
rect 7190 6196 7196 6208
rect 7248 6236 7254 6248
rect 7834 6236 7840 6248
rect 7248 6208 7840 6236
rect 7248 6196 7254 6208
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6236 8263 6239
rect 8662 6236 8668 6248
rect 8251 6208 8668 6236
rect 8251 6205 8263 6208
rect 8205 6199 8263 6205
rect 8662 6196 8668 6208
rect 8720 6236 8726 6248
rect 9306 6236 9312 6248
rect 8720 6208 9312 6236
rect 8720 6196 8726 6208
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6236 11943 6239
rect 12434 6236 12440 6248
rect 11931 6208 12440 6236
rect 11931 6205 11943 6208
rect 11885 6199 11943 6205
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 5040 6140 5488 6168
rect 5040 6128 5046 6140
rect 6638 6128 6644 6180
rect 6696 6168 6702 6180
rect 6825 6171 6883 6177
rect 6825 6168 6837 6171
rect 6696 6140 6837 6168
rect 6696 6128 6702 6140
rect 6825 6137 6837 6140
rect 6871 6168 6883 6171
rect 7653 6171 7711 6177
rect 7653 6168 7665 6171
rect 6871 6140 7665 6168
rect 6871 6137 6883 6140
rect 6825 6131 6883 6137
rect 7653 6137 7665 6140
rect 7699 6137 7711 6171
rect 7653 6131 7711 6137
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 8526 6171 8584 6177
rect 8526 6168 8538 6171
rect 8076 6140 8538 6168
rect 8076 6128 8082 6140
rect 8526 6137 8538 6140
rect 8572 6137 8584 6171
rect 10042 6168 10048 6180
rect 10003 6140 10048 6168
rect 8526 6131 8584 6137
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 10137 6171 10195 6177
rect 10137 6137 10149 6171
rect 10183 6137 10195 6171
rect 10137 6131 10195 6137
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4065 6103 4123 6109
rect 4065 6100 4077 6103
rect 4028 6072 4077 6100
rect 4028 6060 4034 6072
rect 4065 6069 4077 6072
rect 4111 6069 4123 6103
rect 9398 6100 9404 6112
rect 9359 6072 9404 6100
rect 4065 6063 4123 6069
rect 9398 6060 9404 6072
rect 9456 6100 9462 6112
rect 9769 6103 9827 6109
rect 9769 6100 9781 6103
rect 9456 6072 9781 6100
rect 9456 6060 9462 6072
rect 9769 6069 9781 6072
rect 9815 6100 9827 6103
rect 9858 6100 9864 6112
rect 9815 6072 9864 6100
rect 9815 6069 9827 6072
rect 9769 6063 9827 6069
rect 9858 6060 9864 6072
rect 9916 6100 9922 6112
rect 10152 6100 10180 6131
rect 9916 6072 10180 6100
rect 9916 6060 9922 6072
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 12820 6109 12848 6412
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 13722 6440 13728 6452
rect 13403 6412 13728 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 13722 6400 13728 6412
rect 13780 6440 13786 6452
rect 14001 6443 14059 6449
rect 14001 6440 14013 6443
rect 13780 6412 14013 6440
rect 13780 6400 13786 6412
rect 14001 6409 14013 6412
rect 14047 6440 14059 6443
rect 14366 6440 14372 6452
rect 14047 6412 14372 6440
rect 14047 6409 14059 6412
rect 14001 6403 14059 6409
rect 14366 6400 14372 6412
rect 14424 6400 14430 6452
rect 15289 6443 15347 6449
rect 15289 6409 15301 6443
rect 15335 6440 15347 6443
rect 15930 6440 15936 6452
rect 15335 6412 15936 6440
rect 15335 6409 15347 6412
rect 15289 6403 15347 6409
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 16850 6440 16856 6452
rect 16811 6412 16856 6440
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 17589 6443 17647 6449
rect 17589 6440 17601 6443
rect 17000 6412 17601 6440
rect 17000 6400 17006 6412
rect 17589 6409 17601 6412
rect 17635 6409 17647 6443
rect 17589 6403 17647 6409
rect 18601 6443 18659 6449
rect 18601 6409 18613 6443
rect 18647 6440 18659 6443
rect 18690 6440 18696 6452
rect 18647 6412 18696 6440
rect 18647 6409 18659 6412
rect 18601 6403 18659 6409
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 19613 6443 19671 6449
rect 19613 6409 19625 6443
rect 19659 6440 19671 6443
rect 19702 6440 19708 6452
rect 19659 6412 19708 6440
rect 19659 6409 19671 6412
rect 19613 6403 19671 6409
rect 19702 6400 19708 6412
rect 19760 6400 19766 6452
rect 19794 6400 19800 6452
rect 19852 6440 19858 6452
rect 19889 6443 19947 6449
rect 19889 6440 19901 6443
rect 19852 6412 19901 6440
rect 19852 6400 19858 6412
rect 19889 6409 19901 6412
rect 19935 6409 19947 6443
rect 19889 6403 19947 6409
rect 13814 6332 13820 6384
rect 13872 6372 13878 6384
rect 19199 6375 19257 6381
rect 19199 6372 19211 6375
rect 13872 6344 19211 6372
rect 13872 6332 13878 6344
rect 19199 6341 19211 6344
rect 19245 6341 19257 6375
rect 19199 6335 19257 6341
rect 14274 6304 14280 6316
rect 14187 6276 14280 6304
rect 14274 6264 14280 6276
rect 14332 6304 14338 6316
rect 17034 6304 17040 6316
rect 14332 6276 17040 6304
rect 14332 6264 14338 6276
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 15102 6196 15108 6248
rect 15160 6236 15166 6248
rect 15749 6239 15807 6245
rect 15749 6236 15761 6239
rect 15160 6208 15761 6236
rect 15160 6196 15166 6208
rect 15749 6205 15761 6208
rect 15795 6236 15807 6239
rect 16114 6236 16120 6248
rect 15795 6208 16120 6236
rect 15795 6205 15807 6208
rect 15749 6199 15807 6205
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 16206 6196 16212 6248
rect 16264 6236 16270 6248
rect 19128 6239 19186 6245
rect 16264 6208 16309 6236
rect 16264 6196 16270 6208
rect 19128 6205 19140 6239
rect 19174 6236 19186 6239
rect 19794 6236 19800 6248
rect 19174 6208 19800 6236
rect 19174 6205 19186 6208
rect 19128 6199 19186 6205
rect 19794 6196 19800 6208
rect 19852 6196 19858 6248
rect 14366 6128 14372 6180
rect 14424 6168 14430 6180
rect 14921 6171 14979 6177
rect 14424 6140 14469 6168
rect 14424 6128 14430 6140
rect 14921 6137 14933 6171
rect 14967 6168 14979 6171
rect 15470 6168 15476 6180
rect 14967 6140 15476 6168
rect 14967 6137 14979 6140
rect 14921 6131 14979 6137
rect 15470 6128 15476 6140
rect 15528 6128 15534 6180
rect 15654 6128 15660 6180
rect 15712 6168 15718 6180
rect 17126 6168 17132 6180
rect 15712 6140 17132 6168
rect 15712 6128 15718 6140
rect 17126 6128 17132 6140
rect 17184 6168 17190 6180
rect 17221 6171 17279 6177
rect 17221 6168 17233 6171
rect 17184 6140 17233 6168
rect 17184 6128 17190 6140
rect 17221 6137 17233 6140
rect 17267 6137 17279 6171
rect 17221 6131 17279 6137
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 12768 6072 12817 6100
rect 12768 6060 12774 6072
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 12805 6063 12863 6069
rect 14182 6060 14188 6112
rect 14240 6100 14246 6112
rect 14550 6100 14556 6112
rect 14240 6072 14556 6100
rect 14240 6060 14246 6072
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 14826 6060 14832 6112
rect 14884 6100 14890 6112
rect 15565 6103 15623 6109
rect 15565 6100 15577 6103
rect 14884 6072 15577 6100
rect 14884 6060 14890 6072
rect 15565 6069 15577 6072
rect 15611 6069 15623 6103
rect 16022 6100 16028 6112
rect 15983 6072 16028 6100
rect 15565 6063 15623 6069
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 18046 6100 18052 6112
rect 18007 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 1104 6010 20884 6032
rect 1104 5958 8315 6010
rect 8367 5958 8379 6010
rect 8431 5958 8443 6010
rect 8495 5958 8507 6010
rect 8559 5958 15648 6010
rect 15700 5958 15712 6010
rect 15764 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 20884 6010
rect 1104 5936 20884 5958
rect 2130 5856 2136 5908
rect 2188 5896 2194 5908
rect 2869 5899 2927 5905
rect 2869 5896 2881 5899
rect 2188 5868 2881 5896
rect 2188 5856 2194 5868
rect 2869 5865 2881 5868
rect 2915 5865 2927 5899
rect 2869 5859 2927 5865
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 4246 5896 4252 5908
rect 3568 5868 4252 5896
rect 3568 5856 3574 5868
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 5442 5896 5448 5908
rect 5403 5868 5448 5896
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 8757 5899 8815 5905
rect 8757 5865 8769 5899
rect 8803 5896 8815 5899
rect 9398 5896 9404 5908
rect 8803 5868 9404 5896
rect 8803 5865 8815 5868
rect 8757 5859 8815 5865
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 9493 5899 9551 5905
rect 9493 5865 9505 5899
rect 9539 5896 9551 5899
rect 9674 5896 9680 5908
rect 9539 5868 9680 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 10042 5856 10048 5908
rect 10100 5896 10106 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10100 5868 10701 5896
rect 10100 5856 10106 5868
rect 10689 5865 10701 5868
rect 10735 5896 10747 5899
rect 11379 5899 11437 5905
rect 11379 5896 11391 5899
rect 10735 5868 11391 5896
rect 10735 5865 10747 5868
rect 10689 5859 10747 5865
rect 11379 5865 11391 5868
rect 11425 5865 11437 5899
rect 11379 5859 11437 5865
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 16945 5899 17003 5905
rect 16945 5896 16957 5899
rect 12492 5868 16957 5896
rect 12492 5856 12498 5868
rect 16945 5865 16957 5868
rect 16991 5865 17003 5899
rect 16945 5859 17003 5865
rect 2311 5831 2369 5837
rect 2311 5797 2323 5831
rect 2357 5828 2369 5831
rect 2406 5828 2412 5840
rect 2357 5800 2412 5828
rect 2357 5797 2369 5800
rect 2311 5791 2369 5797
rect 2406 5788 2412 5800
rect 2464 5788 2470 5840
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 7469 5831 7527 5837
rect 7469 5828 7481 5831
rect 4120 5800 7481 5828
rect 4120 5788 4126 5800
rect 7469 5797 7481 5800
rect 7515 5828 7527 5831
rect 7926 5828 7932 5840
rect 7515 5800 7932 5828
rect 7515 5797 7527 5800
rect 7469 5791 7527 5797
rect 7926 5788 7932 5800
rect 7984 5788 7990 5840
rect 8018 5788 8024 5840
rect 8076 5828 8082 5840
rect 8158 5831 8216 5837
rect 8158 5828 8170 5831
rect 8076 5800 8170 5828
rect 8076 5788 8082 5800
rect 8158 5797 8170 5800
rect 8204 5797 8216 5831
rect 8158 5791 8216 5797
rect 8938 5788 8944 5840
rect 8996 5828 9002 5840
rect 9033 5831 9091 5837
rect 9033 5828 9045 5831
rect 8996 5800 9045 5828
rect 8996 5788 9002 5800
rect 9033 5797 9045 5800
rect 9079 5828 9091 5831
rect 9769 5831 9827 5837
rect 9769 5828 9781 5831
rect 9079 5800 9781 5828
rect 9079 5797 9091 5800
rect 9033 5791 9091 5797
rect 9769 5797 9781 5800
rect 9815 5797 9827 5831
rect 9769 5791 9827 5797
rect 9861 5831 9919 5837
rect 9861 5797 9873 5831
rect 9907 5828 9919 5831
rect 9950 5828 9956 5840
rect 9907 5800 9956 5828
rect 9907 5797 9919 5800
rect 9861 5791 9919 5797
rect 9950 5788 9956 5800
rect 10008 5788 10014 5840
rect 12710 5788 12716 5840
rect 12768 5828 12774 5840
rect 12850 5831 12908 5837
rect 12850 5828 12862 5831
rect 12768 5800 12862 5828
rect 12768 5788 12774 5800
rect 12850 5797 12862 5800
rect 12896 5797 12908 5831
rect 15378 5828 15384 5840
rect 12850 5791 12908 5797
rect 13464 5800 15384 5828
rect 4801 5763 4859 5769
rect 4801 5729 4813 5763
rect 4847 5760 4859 5763
rect 5166 5760 5172 5772
rect 4847 5732 5172 5760
rect 4847 5729 4859 5732
rect 4801 5723 4859 5729
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5760 5411 5763
rect 5442 5760 5448 5772
rect 5399 5732 5448 5760
rect 5399 5729 5411 5732
rect 5353 5723 5411 5729
rect 5442 5720 5448 5732
rect 5500 5720 5506 5772
rect 6454 5760 6460 5772
rect 6415 5732 6460 5760
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 11276 5763 11334 5769
rect 11276 5760 11288 5763
rect 11256 5729 11288 5760
rect 11322 5729 11334 5763
rect 11256 5723 11334 5729
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5692 2007 5695
rect 4430 5692 4436 5704
rect 1995 5664 4436 5692
rect 1995 5661 2007 5664
rect 1949 5655 2007 5661
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 5258 5692 5264 5704
rect 5219 5664 5264 5692
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 7834 5692 7840 5704
rect 5592 5664 5672 5692
rect 7795 5664 7840 5692
rect 5592 5652 5598 5664
rect 3421 5627 3479 5633
rect 3421 5593 3433 5627
rect 3467 5624 3479 5627
rect 3694 5624 3700 5636
rect 3467 5596 3700 5624
rect 3467 5593 3479 5596
rect 3421 5587 3479 5593
rect 3694 5584 3700 5596
rect 3752 5584 3758 5636
rect 5644 5624 5672 5664
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 11256 5636 11284 5723
rect 11422 5720 11428 5772
rect 11480 5760 11486 5772
rect 11701 5763 11759 5769
rect 11701 5760 11713 5763
rect 11480 5732 11713 5760
rect 11480 5720 11486 5732
rect 11701 5729 11713 5732
rect 11747 5729 11759 5763
rect 11701 5723 11759 5729
rect 12986 5720 12992 5772
rect 13044 5760 13050 5772
rect 13464 5769 13492 5800
rect 15378 5788 15384 5800
rect 15436 5828 15442 5840
rect 15473 5831 15531 5837
rect 15473 5828 15485 5831
rect 15436 5800 15485 5828
rect 15436 5788 15442 5800
rect 15473 5797 15485 5800
rect 15519 5797 15531 5831
rect 15473 5791 15531 5797
rect 16114 5788 16120 5840
rect 16172 5828 16178 5840
rect 16298 5828 16304 5840
rect 16172 5800 16304 5828
rect 16172 5788 16178 5800
rect 16298 5788 16304 5800
rect 16356 5788 16362 5840
rect 13449 5763 13507 5769
rect 13449 5760 13461 5763
rect 13044 5732 13461 5760
rect 13044 5720 13050 5732
rect 13449 5729 13461 5732
rect 13495 5729 13507 5763
rect 13449 5723 13507 5729
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 14274 5760 14280 5772
rect 13872 5732 13917 5760
rect 14235 5732 14280 5760
rect 13872 5720 13878 5732
rect 14274 5720 14280 5732
rect 14332 5720 14338 5772
rect 15102 5760 15108 5772
rect 15063 5732 15108 5760
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 16482 5720 16488 5772
rect 16540 5760 16546 5772
rect 16853 5763 16911 5769
rect 16853 5760 16865 5763
rect 16540 5732 16865 5760
rect 16540 5720 16546 5732
rect 16853 5729 16865 5732
rect 16899 5760 16911 5763
rect 17126 5760 17132 5772
rect 16899 5732 17132 5760
rect 16899 5729 16911 5732
rect 16853 5723 16911 5729
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 17310 5760 17316 5772
rect 17271 5732 17316 5760
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 18417 5763 18475 5769
rect 18417 5729 18429 5763
rect 18463 5760 18475 5763
rect 18506 5760 18512 5772
rect 18463 5732 18512 5760
rect 18463 5729 18475 5732
rect 18417 5723 18475 5729
rect 18506 5720 18512 5732
rect 18564 5720 18570 5772
rect 19058 5720 19064 5772
rect 19116 5760 19122 5772
rect 19464 5763 19522 5769
rect 19464 5760 19476 5763
rect 19116 5732 19476 5760
rect 19116 5720 19122 5732
rect 19464 5729 19476 5732
rect 19510 5729 19522 5763
rect 19464 5723 19522 5729
rect 12526 5692 12532 5704
rect 12487 5664 12532 5692
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 11238 5624 11244 5636
rect 5644 5596 11244 5624
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 15194 5584 15200 5636
rect 15252 5624 15258 5636
rect 15396 5624 15424 5655
rect 15470 5652 15476 5704
rect 15528 5692 15534 5704
rect 15657 5695 15715 5701
rect 15657 5692 15669 5695
rect 15528 5664 15669 5692
rect 15528 5652 15534 5664
rect 15657 5661 15669 5664
rect 15703 5661 15715 5695
rect 15657 5655 15715 5661
rect 15746 5652 15752 5704
rect 15804 5692 15810 5704
rect 19567 5695 19625 5701
rect 19567 5692 19579 5695
rect 15804 5664 19579 5692
rect 15804 5652 15810 5664
rect 19567 5661 19579 5664
rect 19613 5661 19625 5695
rect 19567 5655 19625 5661
rect 18555 5627 18613 5633
rect 18555 5624 18567 5627
rect 15252 5596 18567 5624
rect 15252 5584 15258 5596
rect 18555 5593 18567 5596
rect 18601 5593 18613 5627
rect 18555 5587 18613 5593
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 3786 5556 3792 5568
rect 3747 5528 3792 5556
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 5994 5556 6000 5568
rect 5955 5528 6000 5556
rect 5994 5516 6000 5528
rect 6052 5516 6058 5568
rect 6362 5556 6368 5568
rect 6323 5528 6368 5556
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 6595 5559 6653 5565
rect 6595 5525 6607 5559
rect 6641 5556 6653 5559
rect 6730 5556 6736 5568
rect 6641 5528 6736 5556
rect 6641 5525 6653 5528
rect 6595 5519 6653 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 7006 5556 7012 5568
rect 6967 5528 7012 5556
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 11054 5556 11060 5568
rect 11015 5528 11060 5556
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 1104 5466 20884 5488
rect 1104 5414 4648 5466
rect 4700 5414 4712 5466
rect 4764 5414 4776 5466
rect 4828 5414 4840 5466
rect 4892 5414 11982 5466
rect 12034 5414 12046 5466
rect 12098 5414 12110 5466
rect 12162 5414 12174 5466
rect 12226 5414 19315 5466
rect 19367 5414 19379 5466
rect 19431 5414 19443 5466
rect 19495 5414 19507 5466
rect 19559 5414 20884 5466
rect 1104 5392 20884 5414
rect 2406 5312 2412 5364
rect 2464 5352 2470 5364
rect 2501 5355 2559 5361
rect 2501 5352 2513 5355
rect 2464 5324 2513 5352
rect 2464 5312 2470 5324
rect 2501 5321 2513 5324
rect 2547 5321 2559 5355
rect 2501 5315 2559 5321
rect 4430 5312 4436 5364
rect 4488 5352 4494 5364
rect 6822 5352 6828 5364
rect 4488 5324 6828 5352
rect 4488 5312 4494 5324
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 8018 5352 8024 5364
rect 7979 5324 8024 5352
rect 8018 5312 8024 5324
rect 8076 5352 8082 5364
rect 9309 5355 9367 5361
rect 9309 5352 9321 5355
rect 8076 5324 9321 5352
rect 8076 5312 8082 5324
rect 9309 5321 9321 5324
rect 9355 5352 9367 5355
rect 9398 5352 9404 5364
rect 9355 5324 9404 5352
rect 9355 5321 9367 5324
rect 9309 5315 9367 5321
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 9950 5352 9956 5364
rect 9815 5324 9956 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 11238 5352 11244 5364
rect 11199 5324 11244 5352
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12526 5352 12532 5364
rect 12299 5324 12532 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 12526 5312 12532 5324
rect 12584 5352 12590 5364
rect 13998 5352 14004 5364
rect 12584 5324 14004 5352
rect 12584 5312 12590 5324
rect 13998 5312 14004 5324
rect 14056 5312 14062 5364
rect 15378 5352 15384 5364
rect 15339 5324 15384 5352
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17313 5355 17371 5361
rect 17313 5352 17325 5355
rect 17184 5324 17325 5352
rect 17184 5312 17190 5324
rect 17313 5321 17325 5324
rect 17359 5321 17371 5355
rect 17313 5315 17371 5321
rect 18782 5312 18788 5364
rect 18840 5352 18846 5364
rect 19199 5355 19257 5361
rect 19199 5352 19211 5355
rect 18840 5324 19211 5352
rect 18840 5312 18846 5324
rect 19199 5321 19211 5324
rect 19245 5321 19257 5355
rect 19199 5315 19257 5321
rect 4246 5284 4252 5296
rect 4126 5256 4252 5284
rect 2038 5216 2044 5228
rect 1999 5188 2044 5216
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 3786 5176 3792 5228
rect 3844 5216 3850 5228
rect 4126 5216 4154 5256
rect 4246 5244 4252 5256
rect 4304 5244 4310 5296
rect 7558 5284 7564 5296
rect 7208 5256 7564 5284
rect 5166 5216 5172 5228
rect 3844 5188 4154 5216
rect 5127 5188 5172 5216
rect 3844 5176 3850 5188
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5994 5216 6000 5228
rect 5276 5188 6000 5216
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5148 3295 5151
rect 3602 5148 3608 5160
rect 3283 5120 3608 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 3602 5108 3608 5120
rect 3660 5108 3666 5160
rect 3694 5108 3700 5160
rect 3752 5148 3758 5160
rect 4111 5151 4169 5157
rect 4111 5148 4123 5151
rect 3752 5120 4123 5148
rect 3752 5108 3758 5120
rect 4111 5117 4123 5120
rect 4157 5117 4169 5151
rect 4111 5111 4169 5117
rect 4338 5108 4344 5160
rect 4396 5148 4402 5160
rect 5184 5148 5212 5176
rect 5276 5157 5304 5188
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 7208 5157 7236 5256
rect 7558 5244 7564 5256
rect 7616 5244 7622 5296
rect 10505 5287 10563 5293
rect 10505 5253 10517 5287
rect 10551 5284 10563 5287
rect 10594 5284 10600 5296
rect 10551 5256 10600 5284
rect 10551 5253 10563 5256
rect 10505 5247 10563 5253
rect 10594 5244 10600 5256
rect 10652 5284 10658 5296
rect 11609 5287 11667 5293
rect 11609 5284 11621 5287
rect 10652 5256 11621 5284
rect 10652 5244 10658 5256
rect 11609 5253 11621 5256
rect 11655 5253 11667 5287
rect 12710 5284 12716 5296
rect 12671 5256 12716 5284
rect 11609 5247 11667 5253
rect 12710 5244 12716 5256
rect 12768 5244 12774 5296
rect 13909 5287 13967 5293
rect 13909 5284 13921 5287
rect 13464 5256 13921 5284
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 7423 5188 9965 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 9953 5185 9965 5188
rect 9999 5216 10011 5219
rect 10686 5216 10692 5228
rect 9999 5188 10692 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 12897 5219 12955 5225
rect 12897 5185 12909 5219
rect 12943 5216 12955 5219
rect 13464 5216 13492 5256
rect 13909 5253 13921 5256
rect 13955 5284 13967 5287
rect 15746 5284 15752 5296
rect 13955 5256 15752 5284
rect 13955 5253 13967 5256
rect 13909 5247 13967 5253
rect 15746 5244 15752 5256
rect 15804 5244 15810 5296
rect 19058 5244 19064 5296
rect 19116 5284 19122 5296
rect 19521 5287 19579 5293
rect 19521 5284 19533 5287
rect 19116 5256 19533 5284
rect 19116 5244 19122 5256
rect 19521 5253 19533 5256
rect 19567 5253 19579 5287
rect 19521 5247 19579 5253
rect 12943 5188 13492 5216
rect 13541 5219 13599 5225
rect 12943 5185 12955 5188
rect 12897 5179 12955 5185
rect 13541 5185 13553 5219
rect 13587 5216 13599 5219
rect 15930 5216 15936 5228
rect 13587 5188 13814 5216
rect 15891 5188 15936 5216
rect 13587 5185 13599 5188
rect 13541 5179 13599 5185
rect 4396 5120 5212 5148
rect 5261 5151 5319 5157
rect 4396 5108 4402 5120
rect 5261 5117 5273 5151
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 7168 5151 7236 5157
rect 7168 5117 7180 5151
rect 7214 5120 7236 5151
rect 7214 5117 7226 5120
rect 7168 5111 7226 5117
rect 1578 5080 1584 5092
rect 1539 5052 1584 5080
rect 1578 5040 1584 5052
rect 1636 5040 1642 5092
rect 1670 5040 1676 5092
rect 1728 5080 1734 5092
rect 1728 5052 1773 5080
rect 1728 5040 1734 5052
rect 2866 5040 2872 5092
rect 2924 5080 2930 5092
rect 5276 5080 5304 5111
rect 2924 5052 5304 5080
rect 5460 5080 5488 5111
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 7340 5120 8125 5148
rect 7340 5108 7346 5120
rect 8113 5117 8125 5120
rect 8159 5148 8171 5151
rect 8938 5148 8944 5160
rect 8159 5120 8944 5148
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 8938 5108 8944 5120
rect 8996 5108 9002 5160
rect 13786 5092 13814 5188
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16574 5176 16580 5228
rect 16632 5216 16638 5228
rect 19889 5219 19947 5225
rect 19889 5216 19901 5219
rect 16632 5188 19901 5216
rect 16632 5176 16638 5188
rect 15657 5151 15715 5157
rect 15657 5117 15669 5151
rect 15703 5148 15715 5151
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15703 5120 16037 5148
rect 15703 5117 15715 5120
rect 15657 5111 15715 5117
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 16025 5111 16083 5117
rect 17954 5108 17960 5160
rect 18012 5148 18018 5160
rect 19143 5157 19171 5188
rect 19889 5185 19901 5188
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 18116 5151 18174 5157
rect 18116 5148 18128 5151
rect 18012 5120 18128 5148
rect 18012 5108 18018 5120
rect 18116 5117 18128 5120
rect 18162 5148 18174 5151
rect 18877 5151 18935 5157
rect 18877 5148 18889 5151
rect 18162 5120 18889 5148
rect 18162 5117 18174 5120
rect 18116 5111 18174 5117
rect 18877 5117 18889 5120
rect 18923 5117 18935 5151
rect 18877 5111 18935 5117
rect 19128 5151 19186 5157
rect 19128 5117 19140 5151
rect 19174 5117 19186 5151
rect 19128 5111 19186 5117
rect 6181 5083 6239 5089
rect 6181 5080 6193 5083
rect 5460 5052 6193 5080
rect 2924 5040 2930 5052
rect 6181 5049 6193 5052
rect 6227 5080 6239 5083
rect 6822 5080 6828 5092
rect 6227 5052 6828 5080
rect 6227 5049 6239 5052
rect 6181 5043 6239 5049
rect 6822 5040 6828 5052
rect 6880 5040 6886 5092
rect 8018 5040 8024 5092
rect 8076 5080 8082 5092
rect 8434 5083 8492 5089
rect 8434 5080 8446 5083
rect 8076 5052 8446 5080
rect 8076 5040 8082 5052
rect 8434 5049 8446 5052
rect 8480 5049 8492 5083
rect 10045 5083 10103 5089
rect 8434 5043 8492 5049
rect 9048 5052 9904 5080
rect 4801 5015 4859 5021
rect 4801 4981 4813 5015
rect 4847 5012 4859 5015
rect 5074 5012 5080 5024
rect 4847 4984 5080 5012
rect 4847 4981 4859 4984
rect 4801 4975 4859 4981
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 5258 4972 5264 5024
rect 5316 5012 5322 5024
rect 5537 5015 5595 5021
rect 5537 5012 5549 5015
rect 5316 4984 5549 5012
rect 5316 4972 5322 4984
rect 5537 4981 5549 4984
rect 5583 4981 5595 5015
rect 6454 5012 6460 5024
rect 6415 4984 6460 5012
rect 5537 4975 5595 4981
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 9048 5021 9076 5052
rect 9876 5024 9904 5052
rect 10045 5049 10057 5083
rect 10091 5049 10103 5083
rect 12986 5080 12992 5092
rect 12947 5052 12992 5080
rect 10045 5043 10103 5049
rect 9033 5015 9091 5021
rect 9033 4981 9045 5015
rect 9079 4981 9091 5015
rect 9033 4975 9091 4981
rect 9858 4972 9864 5024
rect 9916 5012 9922 5024
rect 10060 5012 10088 5043
rect 12986 5040 12992 5052
rect 13044 5040 13050 5092
rect 13786 5052 13820 5092
rect 13814 5040 13820 5052
rect 13872 5080 13878 5092
rect 14458 5080 14464 5092
rect 13872 5052 14464 5080
rect 13872 5040 13878 5052
rect 14458 5040 14464 5052
rect 14516 5040 14522 5092
rect 14553 5083 14611 5089
rect 14553 5049 14565 5083
rect 14599 5049 14611 5083
rect 14553 5043 14611 5049
rect 15105 5083 15163 5089
rect 15105 5049 15117 5083
rect 15151 5080 15163 5083
rect 16114 5080 16120 5092
rect 15151 5052 16120 5080
rect 15151 5049 15163 5052
rect 15105 5043 15163 5049
rect 10873 5015 10931 5021
rect 10873 5012 10885 5015
rect 9916 4984 10885 5012
rect 9916 4972 9922 4984
rect 10873 4981 10885 4984
rect 10919 4981 10931 5015
rect 10873 4975 10931 4981
rect 14277 5015 14335 5021
rect 14277 4981 14289 5015
rect 14323 5012 14335 5015
rect 14366 5012 14372 5024
rect 14323 4984 14372 5012
rect 14323 4981 14335 4984
rect 14277 4975 14335 4981
rect 14366 4972 14372 4984
rect 14424 5012 14430 5024
rect 14568 5012 14596 5043
rect 16114 5040 16120 5052
rect 16172 5040 16178 5092
rect 14424 4984 14596 5012
rect 14424 4972 14430 4984
rect 15470 4972 15476 5024
rect 15528 5012 15534 5024
rect 15657 5015 15715 5021
rect 15657 5012 15669 5015
rect 15528 4984 15669 5012
rect 15528 4972 15534 4984
rect 15657 4981 15669 4984
rect 15703 5012 15715 5015
rect 15749 5015 15807 5021
rect 15749 5012 15761 5015
rect 15703 4984 15761 5012
rect 15703 4981 15715 4984
rect 15657 4975 15715 4981
rect 15749 4981 15761 4984
rect 15795 4981 15807 5015
rect 15749 4975 15807 4981
rect 17037 5015 17095 5021
rect 17037 4981 17049 5015
rect 17083 5012 17095 5015
rect 17310 5012 17316 5024
rect 17083 4984 17316 5012
rect 17083 4981 17095 4984
rect 17037 4975 17095 4981
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 17402 4972 17408 5024
rect 17460 5012 17466 5024
rect 18187 5015 18245 5021
rect 18187 5012 18199 5015
rect 17460 4984 18199 5012
rect 17460 4972 17466 4984
rect 18187 4981 18199 4984
rect 18233 4981 18245 5015
rect 18506 5012 18512 5024
rect 18467 4984 18512 5012
rect 18187 4975 18245 4981
rect 18506 4972 18512 4984
rect 18564 4972 18570 5024
rect 1104 4922 20884 4944
rect 1104 4870 8315 4922
rect 8367 4870 8379 4922
rect 8431 4870 8443 4922
rect 8495 4870 8507 4922
rect 8559 4870 15648 4922
rect 15700 4870 15712 4922
rect 15764 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 20884 4922
rect 1104 4848 20884 4870
rect 2866 4808 2872 4820
rect 1596 4780 2544 4808
rect 2827 4780 2872 4808
rect 1596 4681 1624 4780
rect 1943 4743 2001 4749
rect 1943 4709 1955 4743
rect 1989 4740 2001 4743
rect 2406 4740 2412 4752
rect 1989 4712 2412 4740
rect 1989 4709 2001 4712
rect 1943 4703 2001 4709
rect 2406 4700 2412 4712
rect 2464 4700 2470 4752
rect 2516 4740 2544 4780
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 3421 4811 3479 4817
rect 3421 4777 3433 4811
rect 3467 4808 3479 4811
rect 3786 4808 3792 4820
rect 3467 4780 3792 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 4080 4780 4169 4808
rect 2958 4740 2964 4752
rect 2516 4712 2964 4740
rect 2958 4700 2964 4712
rect 3016 4740 3022 4752
rect 4080 4740 4108 4780
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 4157 4771 4215 4777
rect 4522 4768 4528 4820
rect 4580 4808 4586 4820
rect 7009 4811 7067 4817
rect 7009 4808 7021 4811
rect 4580 4780 7021 4808
rect 4580 4768 4586 4780
rect 7009 4777 7021 4780
rect 7055 4777 7067 4811
rect 7466 4808 7472 4820
rect 7427 4780 7472 4808
rect 7009 4771 7067 4777
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 7834 4808 7840 4820
rect 7795 4780 7840 4808
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 8938 4808 8944 4820
rect 8899 4780 8944 4808
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 9272 4780 9321 4808
rect 9272 4768 9278 4780
rect 9309 4777 9321 4780
rect 9355 4777 9367 4811
rect 9309 4771 9367 4777
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 10686 4808 10692 4820
rect 9456 4780 9996 4808
rect 10647 4780 10692 4808
rect 9456 4768 9462 4780
rect 6362 4740 6368 4752
rect 3016 4712 4108 4740
rect 4816 4712 6368 4740
rect 3016 4700 3022 4712
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4641 1639 4675
rect 1581 4635 1639 4641
rect 3694 4632 3700 4684
rect 3752 4672 3758 4684
rect 3881 4675 3939 4681
rect 3881 4672 3893 4675
rect 3752 4644 3893 4672
rect 3752 4632 3758 4644
rect 3881 4641 3893 4644
rect 3927 4672 3939 4675
rect 4154 4672 4160 4684
rect 3927 4644 4160 4672
rect 3927 4641 3939 4644
rect 3881 4635 3939 4641
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 4338 4672 4344 4684
rect 4299 4644 4344 4672
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 4816 4604 4844 4712
rect 6362 4700 6368 4712
rect 6420 4700 6426 4752
rect 8110 4740 8116 4752
rect 7944 4712 8116 4740
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 4982 4672 4988 4684
rect 4939 4644 4988 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 5258 4672 5264 4684
rect 5132 4644 5264 4672
rect 5132 4632 5138 4644
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 6178 4672 6184 4684
rect 6043 4644 6184 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4672 6331 4675
rect 6546 4672 6552 4684
rect 6319 4644 6552 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 7834 4632 7840 4684
rect 7892 4672 7898 4684
rect 7944 4681 7972 4712
rect 8110 4700 8116 4712
rect 8168 4700 8174 4752
rect 8202 4700 8208 4752
rect 8260 4740 8266 4752
rect 9232 4740 9260 4768
rect 9858 4740 9864 4752
rect 8260 4712 9260 4740
rect 9819 4712 9864 4740
rect 8260 4700 8266 4712
rect 9858 4700 9864 4712
rect 9916 4700 9922 4752
rect 9968 4740 9996 4780
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 12161 4811 12219 4817
rect 12161 4777 12173 4811
rect 12207 4808 12219 4811
rect 13078 4808 13084 4820
rect 12207 4780 13084 4808
rect 12207 4777 12219 4780
rect 12161 4771 12219 4777
rect 13078 4768 13084 4780
rect 13136 4808 13142 4820
rect 13814 4808 13820 4820
rect 13136 4780 13216 4808
rect 13136 4768 13142 4780
rect 11330 4740 11336 4752
rect 9968 4712 11336 4740
rect 11330 4700 11336 4712
rect 11388 4740 11394 4752
rect 11603 4743 11661 4749
rect 11603 4740 11615 4743
rect 11388 4712 11615 4740
rect 11388 4700 11394 4712
rect 11603 4709 11615 4712
rect 11649 4740 11661 4743
rect 12710 4740 12716 4752
rect 11649 4712 12716 4740
rect 11649 4709 11661 4712
rect 11603 4703 11661 4709
rect 12710 4700 12716 4712
rect 12768 4700 12774 4752
rect 12894 4740 12900 4752
rect 12855 4712 12900 4740
rect 12894 4700 12900 4712
rect 12952 4700 12958 4752
rect 13188 4749 13216 4780
rect 13740 4780 13820 4808
rect 13740 4749 13768 4780
rect 13814 4768 13820 4780
rect 13872 4808 13878 4820
rect 14369 4811 14427 4817
rect 14369 4808 14381 4811
rect 13872 4780 14381 4808
rect 13872 4768 13878 4780
rect 14369 4777 14381 4780
rect 14415 4777 14427 4811
rect 14369 4771 14427 4777
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 16945 4811 17003 4817
rect 16945 4808 16957 4811
rect 14700 4780 16957 4808
rect 14700 4768 14706 4780
rect 16945 4777 16957 4780
rect 16991 4777 17003 4811
rect 16945 4771 17003 4777
rect 13173 4743 13231 4749
rect 13173 4709 13185 4743
rect 13219 4709 13231 4743
rect 13173 4703 13231 4709
rect 13725 4743 13783 4749
rect 13725 4709 13737 4743
rect 13771 4709 13783 4743
rect 13725 4703 13783 4709
rect 15102 4700 15108 4752
rect 15160 4740 15166 4752
rect 15160 4712 15792 4740
rect 15160 4700 15166 4712
rect 7929 4675 7987 4681
rect 7929 4672 7941 4675
rect 7892 4644 7941 4672
rect 7892 4632 7898 4644
rect 7929 4641 7941 4644
rect 7975 4641 7987 4675
rect 7929 4635 7987 4641
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8389 4675 8447 4681
rect 8389 4672 8401 4675
rect 8076 4644 8401 4672
rect 8076 4632 8082 4644
rect 8389 4641 8401 4644
rect 8435 4641 8447 4675
rect 8389 4635 8447 4641
rect 12342 4632 12348 4684
rect 12400 4672 12406 4684
rect 15013 4675 15071 4681
rect 12400 4644 12940 4672
rect 12400 4632 12406 4644
rect 2516 4576 4844 4604
rect 6733 4607 6791 4613
rect 1762 4496 1768 4548
rect 1820 4536 1826 4548
rect 2516 4545 2544 4576
rect 6733 4573 6745 4607
rect 6779 4604 6791 4607
rect 6914 4604 6920 4616
rect 6779 4576 6920 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 6914 4564 6920 4576
rect 6972 4564 6978 4616
rect 8662 4604 8668 4616
rect 8623 4576 8668 4604
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 9122 4564 9128 4616
rect 9180 4604 9186 4616
rect 9582 4604 9588 4616
rect 9180 4576 9588 4604
rect 9180 4564 9186 4576
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4604 9827 4607
rect 10134 4604 10140 4616
rect 9815 4576 10041 4604
rect 10095 4576 10140 4604
rect 9815 4573 9827 4576
rect 9769 4567 9827 4573
rect 2501 4539 2559 4545
rect 2501 4536 2513 4539
rect 1820 4508 2513 4536
rect 1820 4496 1826 4508
rect 2501 4505 2513 4508
rect 2547 4505 2559 4539
rect 2501 4499 2559 4505
rect 5258 4496 5264 4548
rect 5316 4536 5322 4548
rect 5537 4539 5595 4545
rect 5537 4536 5549 4539
rect 5316 4508 5549 4536
rect 5316 4496 5322 4508
rect 5537 4505 5549 4508
rect 5583 4536 5595 4539
rect 6089 4539 6147 4545
rect 6089 4536 6101 4539
rect 5583 4508 6101 4536
rect 5583 4505 5595 4508
rect 5537 4499 5595 4505
rect 6089 4505 6101 4508
rect 6135 4536 6147 4539
rect 6362 4536 6368 4548
rect 6135 4508 6368 4536
rect 6135 4505 6147 4508
rect 6089 4499 6147 4505
rect 6362 4496 6368 4508
rect 6420 4496 6426 4548
rect 10013 4536 10041 4576
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4604 11299 4607
rect 11698 4604 11704 4616
rect 11287 4576 11704 4604
rect 11287 4573 11299 4576
rect 11241 4567 11299 4573
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 12912 4604 12940 4644
rect 15013 4641 15025 4675
rect 15059 4672 15071 4675
rect 15194 4672 15200 4684
rect 15059 4644 15200 4672
rect 15059 4641 15071 4644
rect 15013 4635 15071 4641
rect 15194 4632 15200 4644
rect 15252 4632 15258 4684
rect 15378 4672 15384 4684
rect 15339 4644 15384 4672
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 15764 4681 15792 4712
rect 15749 4675 15807 4681
rect 15749 4641 15761 4675
rect 15795 4641 15807 4675
rect 15749 4635 15807 4641
rect 16298 4632 16304 4684
rect 16356 4672 16362 4684
rect 16666 4672 16672 4684
rect 16356 4644 16672 4672
rect 16356 4632 16362 4644
rect 16666 4632 16672 4644
rect 16724 4672 16730 4684
rect 16853 4675 16911 4681
rect 16853 4672 16865 4675
rect 16724 4644 16865 4672
rect 16724 4632 16730 4644
rect 16853 4641 16865 4644
rect 16899 4641 16911 4675
rect 17310 4672 17316 4684
rect 17271 4644 17316 4672
rect 16853 4635 16911 4641
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 18417 4675 18475 4681
rect 18417 4641 18429 4675
rect 18463 4672 18475 4675
rect 18690 4672 18696 4684
rect 18463 4644 18696 4672
rect 18463 4641 18475 4644
rect 18417 4635 18475 4641
rect 18690 4632 18696 4644
rect 18748 4672 18754 4684
rect 19150 4672 19156 4684
rect 18748 4644 19156 4672
rect 18748 4632 18754 4644
rect 19150 4632 19156 4644
rect 19208 4672 19214 4684
rect 19556 4675 19614 4681
rect 19556 4672 19568 4675
rect 19208 4644 19568 4672
rect 19208 4632 19214 4644
rect 19556 4641 19568 4644
rect 19602 4641 19614 4675
rect 19556 4635 19614 4641
rect 13081 4607 13139 4613
rect 13081 4604 13093 4607
rect 12912 4576 13093 4604
rect 13081 4573 13093 4576
rect 13127 4604 13139 4607
rect 13127 4576 13952 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 11054 4536 11060 4548
rect 10013 4508 11060 4536
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 12437 4539 12495 4545
rect 12437 4536 12449 4539
rect 11256 4508 12449 4536
rect 11256 4480 11284 4508
rect 12437 4505 12449 4508
rect 12483 4505 12495 4539
rect 13924 4536 13952 4576
rect 13998 4564 14004 4616
rect 14056 4604 14062 4616
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 14056 4576 15853 4604
rect 14056 4564 14062 4576
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 19659 4539 19717 4545
rect 19659 4536 19671 4539
rect 13924 4508 19671 4536
rect 12437 4499 12495 4505
rect 19659 4505 19671 4508
rect 19705 4505 19717 4539
rect 19659 4499 19717 4505
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 5442 4468 5448 4480
rect 5224 4440 5448 4468
rect 5224 4428 5230 4440
rect 5442 4428 5448 4440
rect 5500 4468 5506 4480
rect 5905 4471 5963 4477
rect 5905 4468 5917 4471
rect 5500 4440 5917 4468
rect 5500 4428 5506 4440
rect 5905 4437 5917 4440
rect 5951 4468 5963 4471
rect 6178 4468 6184 4480
rect 5951 4440 6184 4468
rect 5951 4437 5963 4440
rect 5905 4431 5963 4437
rect 6178 4428 6184 4440
rect 6236 4428 6242 4480
rect 11238 4428 11244 4480
rect 11296 4428 11302 4480
rect 13538 4428 13544 4480
rect 13596 4468 13602 4480
rect 14093 4471 14151 4477
rect 14093 4468 14105 4471
rect 13596 4440 14105 4468
rect 13596 4428 13602 4440
rect 14093 4437 14105 4440
rect 14139 4468 14151 4471
rect 16574 4468 16580 4480
rect 14139 4440 16580 4468
rect 14139 4437 14151 4440
rect 14093 4431 14151 4437
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 18601 4471 18659 4477
rect 18601 4437 18613 4471
rect 18647 4468 18659 4471
rect 18874 4468 18880 4480
rect 18647 4440 18880 4468
rect 18647 4437 18659 4440
rect 18601 4431 18659 4437
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 1104 4378 20884 4400
rect 1104 4326 4648 4378
rect 4700 4326 4712 4378
rect 4764 4326 4776 4378
rect 4828 4326 4840 4378
rect 4892 4326 11982 4378
rect 12034 4326 12046 4378
rect 12098 4326 12110 4378
rect 12162 4326 12174 4378
rect 12226 4326 19315 4378
rect 19367 4326 19379 4378
rect 19431 4326 19443 4378
rect 19495 4326 19507 4378
rect 19559 4326 20884 4378
rect 1104 4304 20884 4326
rect 2130 4224 2136 4276
rect 2188 4264 2194 4276
rect 2685 4267 2743 4273
rect 2685 4264 2697 4267
rect 2188 4236 2697 4264
rect 2188 4224 2194 4236
rect 2685 4233 2697 4236
rect 2731 4264 2743 4267
rect 3050 4264 3056 4276
rect 2731 4236 3056 4264
rect 2731 4233 2743 4236
rect 2685 4227 2743 4233
rect 3050 4224 3056 4236
rect 3108 4224 3114 4276
rect 3513 4267 3571 4273
rect 3513 4233 3525 4267
rect 3559 4264 3571 4267
rect 3602 4264 3608 4276
rect 3559 4236 3608 4264
rect 3559 4233 3571 4236
rect 3513 4227 3571 4233
rect 3602 4224 3608 4236
rect 3660 4264 3666 4276
rect 4338 4264 4344 4276
rect 3660 4236 4344 4264
rect 3660 4224 3666 4236
rect 4338 4224 4344 4236
rect 4396 4264 4402 4276
rect 6638 4264 6644 4276
rect 4396 4236 6644 4264
rect 4396 4224 4402 4236
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 7466 4264 7472 4276
rect 6840 4236 7472 4264
rect 5258 4196 5264 4208
rect 5219 4168 5264 4196
rect 5258 4156 5264 4168
rect 5316 4156 5322 4208
rect 5442 4156 5448 4208
rect 5500 4196 5506 4208
rect 6840 4196 6868 4236
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 7558 4224 7564 4276
rect 7616 4264 7622 4276
rect 8205 4267 8263 4273
rect 8205 4264 8217 4267
rect 7616 4236 8217 4264
rect 7616 4224 7622 4236
rect 8205 4233 8217 4236
rect 8251 4264 8263 4267
rect 9398 4264 9404 4276
rect 8251 4236 9404 4264
rect 8251 4233 8263 4236
rect 8205 4227 8263 4233
rect 5500 4168 6868 4196
rect 5500 4156 5506 4168
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 1854 4128 1860 4140
rect 1719 4100 1860 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 4246 4128 4252 4140
rect 4126 4100 4252 4128
rect 4126 4072 4154 4100
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4128 4399 4131
rect 7282 4128 7288 4140
rect 4387 4100 7288 4128
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8260 4100 8309 4128
rect 8260 4088 8266 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4029 3939 4063
rect 4062 4060 4068 4072
rect 4023 4032 4068 4060
rect 3881 4023 3939 4029
rect 1762 3992 1768 4004
rect 1723 3964 1768 3992
rect 1762 3952 1768 3964
rect 1820 3952 1826 4004
rect 3896 3992 3924 4023
rect 4062 4020 4068 4032
rect 4120 4032 4154 4072
rect 4522 4060 4528 4072
rect 4264 4032 4528 4060
rect 4120 4020 4126 4032
rect 4264 4004 4292 4032
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 5166 4060 5172 4072
rect 5127 4032 5172 4060
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 5445 4063 5503 4069
rect 5445 4060 5457 4063
rect 5316 4032 5457 4060
rect 5316 4020 5322 4032
rect 5445 4029 5457 4032
rect 5491 4060 5503 4063
rect 5534 4060 5540 4072
rect 5491 4032 5540 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6696 4032 6837 4060
rect 6696 4020 6702 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4029 7067 4063
rect 7009 4023 7067 4029
rect 7377 4063 7435 4069
rect 7377 4029 7389 4063
rect 7423 4060 7435 4063
rect 8110 4060 8116 4072
rect 7423 4032 8116 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 4246 3992 4252 4004
rect 3896 3964 4252 3992
rect 4246 3952 4252 3964
rect 4304 3952 4310 4004
rect 4430 3952 4436 4004
rect 4488 3992 4494 4004
rect 7024 3992 7052 4023
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 8655 4001 8683 4236
rect 9398 4224 9404 4236
rect 9456 4224 9462 4276
rect 9858 4264 9864 4276
rect 9819 4236 9864 4264
rect 9858 4224 9864 4236
rect 9916 4224 9922 4276
rect 11054 4224 11060 4276
rect 11112 4264 11118 4276
rect 12575 4267 12633 4273
rect 12575 4264 12587 4267
rect 11112 4236 12587 4264
rect 11112 4224 11118 4236
rect 12575 4233 12587 4236
rect 12621 4233 12633 4267
rect 12575 4227 12633 4233
rect 12710 4224 12716 4276
rect 12768 4264 12774 4276
rect 13357 4267 13415 4273
rect 13357 4264 13369 4267
rect 12768 4236 13369 4264
rect 12768 4224 12774 4236
rect 13357 4233 13369 4236
rect 13403 4264 13415 4267
rect 13906 4264 13912 4276
rect 13403 4236 13912 4264
rect 13403 4233 13415 4236
rect 13357 4227 13415 4233
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 14366 4224 14372 4276
rect 14424 4264 14430 4276
rect 14461 4267 14519 4273
rect 14461 4264 14473 4267
rect 14424 4236 14473 4264
rect 14424 4224 14430 4236
rect 14461 4233 14473 4236
rect 14507 4233 14519 4267
rect 14461 4227 14519 4233
rect 14550 4224 14556 4276
rect 14608 4264 14614 4276
rect 14737 4267 14795 4273
rect 14737 4264 14749 4267
rect 14608 4236 14749 4264
rect 14608 4224 14614 4236
rect 14737 4233 14749 4236
rect 14783 4264 14795 4267
rect 15378 4264 15384 4276
rect 14783 4236 15384 4264
rect 14783 4233 14795 4236
rect 14737 4227 14795 4233
rect 15378 4224 15384 4236
rect 15436 4224 15442 4276
rect 16666 4264 16672 4276
rect 16627 4236 16672 4264
rect 16666 4224 16672 4236
rect 16724 4224 16730 4276
rect 19150 4264 19156 4276
rect 19111 4236 19156 4264
rect 19150 4224 19156 4236
rect 19208 4264 19214 4276
rect 20073 4267 20131 4273
rect 20073 4264 20085 4267
rect 19208 4236 20085 4264
rect 19208 4224 19214 4236
rect 20073 4233 20085 4236
rect 20119 4233 20131 4267
rect 20073 4227 20131 4233
rect 10594 4196 10600 4208
rect 10152 4168 10600 4196
rect 10152 4137 10180 4168
rect 10594 4156 10600 4168
rect 10652 4156 10658 4208
rect 11330 4196 11336 4208
rect 11291 4168 11336 4196
rect 11330 4156 11336 4168
rect 11388 4156 11394 4208
rect 11698 4196 11704 4208
rect 11611 4168 11704 4196
rect 11698 4156 11704 4168
rect 11756 4196 11762 4208
rect 14642 4196 14648 4208
rect 11756 4168 14648 4196
rect 11756 4156 11762 4168
rect 14642 4156 14648 4168
rect 14700 4156 14706 4208
rect 18322 4196 18328 4208
rect 18283 4168 18328 4196
rect 18322 4156 18328 4168
rect 18380 4156 18386 4208
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 10115 4100 10149 4128
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10410 4128 10416 4140
rect 10371 4100 10416 4128
rect 10137 4091 10195 4097
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12342 4128 12348 4140
rect 12299 4100 12348 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 13538 4128 13544 4140
rect 13499 4100 13544 4128
rect 13538 4088 13544 4100
rect 13596 4088 13602 4140
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 21542 4128 21548 4140
rect 17552 4100 21548 4128
rect 17552 4088 17558 4100
rect 21542 4088 21548 4100
rect 21600 4088 21606 4140
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4060 9275 4063
rect 12504 4063 12562 4069
rect 9263 4032 9904 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 7653 3995 7711 4001
rect 7653 3992 7665 3995
rect 4488 3964 7665 3992
rect 4488 3952 4494 3964
rect 7653 3961 7665 3964
rect 7699 3961 7711 3995
rect 7653 3955 7711 3961
rect 8638 3995 8696 4001
rect 8638 3961 8650 3995
rect 8684 3992 8696 3995
rect 8754 3992 8760 4004
rect 8684 3964 8760 3992
rect 8684 3961 8696 3964
rect 8638 3955 8696 3961
rect 8754 3952 8760 3964
rect 8812 3952 8818 4004
rect 9876 3992 9904 4032
rect 12504 4029 12516 4063
rect 12550 4060 12562 4063
rect 12550 4029 12572 4060
rect 12504 4023 12572 4029
rect 10226 3992 10232 4004
rect 9876 3964 10232 3992
rect 10226 3952 10232 3964
rect 10284 3952 10290 4004
rect 12544 3992 12572 4023
rect 16758 4020 16764 4072
rect 16816 4060 16822 4072
rect 17773 4063 17831 4069
rect 17773 4060 17785 4063
rect 16816 4032 17785 4060
rect 16816 4020 16822 4032
rect 17773 4029 17785 4032
rect 17819 4060 17831 4063
rect 18046 4060 18052 4072
rect 17819 4032 18052 4060
rect 17819 4029 17831 4032
rect 17773 4023 17831 4029
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 18230 4020 18236 4072
rect 18288 4060 18294 4072
rect 18325 4063 18383 4069
rect 18325 4060 18337 4063
rect 18288 4032 18337 4060
rect 18288 4020 18294 4032
rect 18325 4029 18337 4032
rect 18371 4029 18383 4063
rect 19648 4063 19706 4069
rect 19648 4060 19660 4063
rect 18325 4023 18383 4029
rect 19306 4032 19660 4060
rect 12989 3995 13047 4001
rect 12989 3992 13001 3995
rect 12544 3964 13001 3992
rect 12989 3961 13001 3964
rect 13035 3992 13047 3995
rect 13722 3992 13728 4004
rect 13035 3964 13728 3992
rect 13035 3961 13047 3964
rect 12989 3955 13047 3961
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 15010 3952 15016 4004
rect 15068 3992 15074 4004
rect 15381 3995 15439 4001
rect 15381 3992 15393 3995
rect 15068 3964 15393 3992
rect 15068 3952 15074 3964
rect 15304 3936 15332 3964
rect 15381 3961 15393 3964
rect 15427 3961 15439 3995
rect 15381 3955 15439 3961
rect 15470 3952 15476 4004
rect 15528 3992 15534 4004
rect 15528 3964 15573 3992
rect 15528 3952 15534 3964
rect 15838 3952 15844 4004
rect 15896 3992 15902 4004
rect 16025 3995 16083 4001
rect 16025 3992 16037 3995
rect 15896 3964 16037 3992
rect 15896 3952 15902 3964
rect 16025 3961 16037 3964
rect 16071 3992 16083 3995
rect 16114 3992 16120 4004
rect 16071 3964 16120 3992
rect 16071 3961 16083 3964
rect 16025 3955 16083 3961
rect 16114 3952 16120 3964
rect 16172 3992 16178 4004
rect 16172 3964 17908 3992
rect 16172 3952 16178 3964
rect 3145 3927 3203 3933
rect 3145 3893 3157 3927
rect 3191 3924 3203 3927
rect 3878 3924 3884 3936
rect 3191 3896 3884 3924
rect 3191 3893 3203 3896
rect 3145 3887 3203 3893
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 4709 3927 4767 3933
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 4982 3924 4988 3936
rect 4755 3896 4988 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5077 3927 5135 3933
rect 5077 3893 5089 3927
rect 5123 3924 5135 3927
rect 5258 3924 5264 3936
rect 5123 3896 5264 3924
rect 5123 3893 5135 3896
rect 5077 3887 5135 3893
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 5442 3884 5448 3936
rect 5500 3924 5506 3936
rect 5629 3927 5687 3933
rect 5629 3924 5641 3927
rect 5500 3896 5641 3924
rect 5500 3884 5506 3896
rect 5629 3893 5641 3896
rect 5675 3893 5687 3927
rect 5629 3887 5687 3893
rect 5810 3884 5816 3936
rect 5868 3924 5874 3936
rect 6181 3927 6239 3933
rect 6181 3924 6193 3927
rect 5868 3896 6193 3924
rect 5868 3884 5874 3896
rect 6181 3893 6193 3896
rect 6227 3924 6239 3927
rect 6362 3924 6368 3936
rect 6227 3896 6368 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 9490 3924 9496 3936
rect 9451 3896 9496 3924
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 13906 3924 13912 3936
rect 13867 3896 13912 3924
rect 13906 3884 13912 3896
rect 13964 3884 13970 3936
rect 15102 3924 15108 3936
rect 15063 3896 15108 3924
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15286 3884 15292 3936
rect 15344 3884 15350 3936
rect 15488 3924 15516 3952
rect 16301 3927 16359 3933
rect 16301 3924 16313 3927
rect 15488 3896 16313 3924
rect 16301 3893 16313 3896
rect 16347 3893 16359 3927
rect 16850 3924 16856 3936
rect 16811 3896 16856 3924
rect 16301 3887 16359 3893
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 17310 3924 17316 3936
rect 17271 3896 17316 3924
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 17880 3924 17908 3964
rect 19306 3924 19334 4032
rect 19648 4029 19660 4032
rect 19694 4060 19706 4063
rect 20441 4063 20499 4069
rect 20441 4060 20453 4063
rect 19694 4032 20453 4060
rect 19694 4029 19706 4032
rect 19648 4023 19706 4029
rect 20441 4029 20453 4032
rect 20487 4029 20499 4063
rect 20441 4023 20499 4029
rect 19751 3995 19809 4001
rect 19751 3961 19763 3995
rect 19797 3992 19809 3995
rect 21082 3992 21088 4004
rect 19797 3964 21088 3992
rect 19797 3961 19809 3964
rect 19751 3955 19809 3961
rect 21082 3952 21088 3964
rect 21140 3952 21146 4004
rect 17880 3896 19334 3924
rect 1104 3834 20884 3856
rect 1104 3782 8315 3834
rect 8367 3782 8379 3834
rect 8431 3782 8443 3834
rect 8495 3782 8507 3834
rect 8559 3782 15648 3834
rect 15700 3782 15712 3834
rect 15764 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 20884 3834
rect 1104 3760 20884 3782
rect 2130 3720 2136 3732
rect 2091 3692 2136 3720
rect 2130 3680 2136 3692
rect 2188 3680 2194 3732
rect 3697 3723 3755 3729
rect 3697 3689 3709 3723
rect 3743 3720 3755 3723
rect 4062 3720 4068 3732
rect 3743 3692 4068 3720
rect 3743 3689 3755 3692
rect 3697 3683 3755 3689
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 4617 3723 4675 3729
rect 4617 3689 4629 3723
rect 4663 3720 4675 3723
rect 5074 3720 5080 3732
rect 4663 3692 5080 3720
rect 4663 3689 4675 3692
rect 4617 3683 4675 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 7558 3720 7564 3732
rect 7519 3692 7564 3720
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 8662 3680 8668 3732
rect 8720 3720 8726 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 8720 3692 9413 3720
rect 8720 3680 8726 3692
rect 9401 3689 9413 3692
rect 9447 3689 9459 3723
rect 9401 3683 9459 3689
rect 10226 3680 10232 3732
rect 10284 3720 10290 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10284 3692 10701 3720
rect 10284 3680 10290 3692
rect 10689 3689 10701 3692
rect 10735 3689 10747 3723
rect 12434 3720 12440 3732
rect 10689 3683 10747 3689
rect 12084 3692 12440 3720
rect 2958 3652 2964 3664
rect 2608 3624 2964 3652
rect 2608 3593 2636 3624
rect 2958 3612 2964 3624
rect 3016 3612 3022 3664
rect 7190 3652 7196 3664
rect 4126 3624 7052 3652
rect 7151 3624 7196 3652
rect 2593 3587 2651 3593
rect 2593 3553 2605 3587
rect 2639 3553 2651 3587
rect 3050 3584 3056 3596
rect 3011 3556 3056 3584
rect 2593 3547 2651 3553
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 4126 3593 4154 3624
rect 4111 3587 4169 3593
rect 4111 3553 4123 3587
rect 4157 3553 4169 3587
rect 4111 3547 4169 3553
rect 4338 3544 4344 3596
rect 4396 3584 4402 3596
rect 4893 3587 4951 3593
rect 4893 3584 4905 3587
rect 4396 3556 4905 3584
rect 4396 3544 4402 3556
rect 4893 3553 4905 3556
rect 4939 3553 4951 3587
rect 5074 3584 5080 3596
rect 5035 3556 5080 3584
rect 4893 3547 4951 3553
rect 4908 3516 4936 3547
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 5353 3587 5411 3593
rect 5353 3553 5365 3587
rect 5399 3584 5411 3587
rect 5534 3584 5540 3596
rect 5399 3556 5540 3584
rect 5399 3553 5411 3556
rect 5353 3547 5411 3553
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 6638 3584 6644 3596
rect 6599 3556 6644 3584
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 6822 3584 6828 3596
rect 6783 3556 6828 3584
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 7024 3584 7052 3624
rect 7190 3612 7196 3624
rect 7248 3612 7254 3664
rect 8202 3652 8208 3664
rect 8163 3624 8208 3652
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 9858 3652 9864 3664
rect 9819 3624 9864 3652
rect 9858 3612 9864 3624
rect 9916 3612 9922 3664
rect 12084 3661 12112 3692
rect 12434 3680 12440 3692
rect 12492 3720 12498 3732
rect 13078 3720 13084 3732
rect 12492 3692 13084 3720
rect 12492 3680 12498 3692
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 14369 3723 14427 3729
rect 14369 3689 14381 3723
rect 14415 3720 14427 3723
rect 15470 3720 15476 3732
rect 14415 3692 15476 3720
rect 14415 3689 14427 3692
rect 14369 3683 14427 3689
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 16298 3720 16304 3732
rect 16259 3692 16304 3720
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 16942 3720 16948 3732
rect 16903 3692 16948 3720
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 12069 3655 12127 3661
rect 12069 3621 12081 3655
rect 12115 3621 12127 3655
rect 12069 3615 12127 3621
rect 13811 3655 13869 3661
rect 13811 3621 13823 3655
rect 13857 3652 13869 3655
rect 13906 3652 13912 3664
rect 13857 3624 13912 3652
rect 13857 3621 13869 3624
rect 13811 3615 13869 3621
rect 13906 3612 13912 3624
rect 13964 3612 13970 3664
rect 12621 3587 12679 3593
rect 7024 3556 7972 3584
rect 5626 3516 5632 3528
rect 4908 3488 5632 3516
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3516 5871 3519
rect 7834 3516 7840 3528
rect 5859 3488 7840 3516
rect 5859 3485 5871 3488
rect 5813 3479 5871 3485
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 106 3408 112 3460
rect 164 3448 170 3460
rect 4203 3451 4261 3457
rect 4203 3448 4215 3451
rect 164 3420 4215 3448
rect 164 3408 170 3420
rect 4203 3417 4215 3420
rect 4249 3417 4261 3451
rect 4203 3411 4261 3417
rect 5169 3451 5227 3457
rect 5169 3417 5181 3451
rect 5215 3448 5227 3451
rect 6270 3448 6276 3460
rect 5215 3420 6276 3448
rect 5215 3417 5227 3420
rect 5169 3411 5227 3417
rect 6270 3408 6276 3420
rect 6328 3408 6334 3460
rect 6546 3448 6552 3460
rect 6507 3420 6552 3448
rect 6546 3408 6552 3420
rect 6604 3408 6610 3460
rect 7944 3448 7972 3556
rect 12621 3553 12633 3587
rect 12667 3584 12679 3587
rect 15010 3584 15016 3596
rect 12667 3556 15016 3584
rect 12667 3553 12679 3556
rect 12621 3547 12679 3553
rect 15010 3544 15016 3556
rect 15068 3544 15074 3596
rect 15562 3584 15568 3596
rect 15523 3556 15568 3584
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 17126 3584 17132 3596
rect 17087 3556 17132 3584
rect 17126 3544 17132 3556
rect 17184 3544 17190 3596
rect 17310 3584 17316 3596
rect 17271 3556 17316 3584
rect 17310 3544 17316 3556
rect 17368 3544 17374 3596
rect 19058 3584 19064 3596
rect 19019 3556 19064 3584
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8159 3488 9137 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 9125 3485 9137 3488
rect 9171 3516 9183 3519
rect 9398 3516 9404 3528
rect 9171 3488 9404 3516
rect 9171 3485 9183 3488
rect 9125 3479 9183 3485
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3516 9827 3519
rect 10134 3516 10140 3528
rect 9815 3488 10140 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 10134 3476 10140 3488
rect 10192 3516 10198 3528
rect 11146 3516 11152 3528
rect 10192 3488 11152 3516
rect 10192 3476 10198 3488
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 11977 3519 12035 3525
rect 11977 3485 11989 3519
rect 12023 3485 12035 3519
rect 13446 3516 13452 3528
rect 13407 3488 13452 3516
rect 11977 3479 12035 3485
rect 8665 3451 8723 3457
rect 8665 3448 8677 3451
rect 7944 3420 8677 3448
rect 8665 3417 8677 3420
rect 8711 3448 8723 3451
rect 8846 3448 8852 3460
rect 8711 3420 8852 3448
rect 8711 3417 8723 3420
rect 8665 3411 8723 3417
rect 8846 3408 8852 3420
rect 8904 3448 8910 3460
rect 10321 3451 10379 3457
rect 10321 3448 10333 3451
rect 8904 3420 10333 3448
rect 8904 3408 8910 3420
rect 10321 3417 10333 3420
rect 10367 3448 10379 3451
rect 10410 3448 10416 3460
rect 10367 3420 10416 3448
rect 10367 3417 10379 3420
rect 10321 3411 10379 3417
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 11793 3451 11851 3457
rect 11793 3417 11805 3451
rect 11839 3448 11851 3451
rect 11992 3448 12020 3479
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 15286 3516 15292 3528
rect 15247 3488 15292 3516
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 18417 3519 18475 3525
rect 18417 3516 18429 3519
rect 16632 3488 18429 3516
rect 16632 3476 16638 3488
rect 18417 3485 18429 3488
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 17402 3448 17408 3460
rect 11839 3420 17408 3448
rect 11839 3417 11851 3420
rect 11793 3411 11851 3417
rect 17402 3408 17408 3420
rect 17460 3408 17466 3460
rect 1673 3383 1731 3389
rect 1673 3349 1685 3383
rect 1719 3380 1731 3383
rect 2222 3380 2228 3392
rect 1719 3352 2228 3380
rect 1719 3349 1731 3352
rect 1673 3343 1731 3349
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 2409 3383 2467 3389
rect 2409 3349 2421 3383
rect 2455 3380 2467 3383
rect 3786 3380 3792 3392
rect 2455 3352 3792 3380
rect 2455 3349 2467 3352
rect 2409 3343 2467 3349
rect 3786 3340 3792 3352
rect 3844 3380 3850 3392
rect 4430 3380 4436 3392
rect 3844 3352 4436 3380
rect 3844 3340 3850 3352
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 6178 3380 6184 3392
rect 6139 3352 6184 3380
rect 6178 3340 6184 3352
rect 6236 3340 6242 3392
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 10594 3380 10600 3392
rect 9180 3352 10600 3380
rect 9180 3340 9186 3352
rect 10594 3340 10600 3352
rect 10652 3380 10658 3392
rect 11057 3383 11115 3389
rect 11057 3380 11069 3383
rect 10652 3352 11069 3380
rect 10652 3340 10658 3352
rect 11057 3349 11069 3352
rect 11103 3349 11115 3383
rect 14642 3380 14648 3392
rect 14603 3352 14648 3380
rect 11057 3343 11115 3349
rect 14642 3340 14648 3352
rect 14700 3340 14706 3392
rect 1104 3290 20884 3312
rect 1104 3238 4648 3290
rect 4700 3238 4712 3290
rect 4764 3238 4776 3290
rect 4828 3238 4840 3290
rect 4892 3238 11982 3290
rect 12034 3238 12046 3290
rect 12098 3238 12110 3290
rect 12162 3238 12174 3290
rect 12226 3238 19315 3290
rect 19367 3238 19379 3290
rect 19431 3238 19443 3290
rect 19495 3238 19507 3290
rect 19559 3238 20884 3290
rect 1104 3216 20884 3238
rect 1949 3179 2007 3185
rect 1949 3145 1961 3179
rect 1995 3176 2007 3179
rect 2179 3179 2237 3185
rect 2179 3176 2191 3179
rect 1995 3148 2191 3176
rect 1995 3145 2007 3148
rect 1949 3139 2007 3145
rect 2179 3145 2191 3148
rect 2225 3176 2237 3179
rect 3970 3176 3976 3188
rect 2225 3148 3976 3176
rect 2225 3145 2237 3148
rect 2179 3139 2237 3145
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 4120 3148 6193 3176
rect 4120 3136 4126 3148
rect 6181 3145 6193 3148
rect 6227 3176 6239 3179
rect 6638 3176 6644 3188
rect 6227 3148 6644 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 8665 3179 8723 3185
rect 8665 3145 8677 3179
rect 8711 3176 8723 3179
rect 8754 3176 8760 3188
rect 8711 3148 8760 3176
rect 8711 3145 8723 3148
rect 8665 3139 8723 3145
rect 8754 3136 8760 3148
rect 8812 3136 8818 3188
rect 9677 3179 9735 3185
rect 9677 3145 9689 3179
rect 9723 3176 9735 3179
rect 9858 3176 9864 3188
rect 9723 3148 9864 3176
rect 9723 3145 9735 3148
rect 9677 3139 9735 3145
rect 9858 3136 9864 3148
rect 9916 3176 9922 3188
rect 9953 3179 10011 3185
rect 9953 3176 9965 3179
rect 9916 3148 9965 3176
rect 9916 3136 9922 3148
rect 9953 3145 9965 3148
rect 9999 3145 10011 3179
rect 9953 3139 10011 3145
rect 13446 3136 13452 3188
rect 13504 3176 13510 3188
rect 13909 3179 13967 3185
rect 13909 3176 13921 3179
rect 13504 3148 13921 3176
rect 13504 3136 13510 3148
rect 13909 3145 13921 3148
rect 13955 3176 13967 3179
rect 16942 3176 16948 3188
rect 13955 3148 16948 3176
rect 13955 3145 13967 3148
rect 13909 3139 13967 3145
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 17313 3179 17371 3185
rect 17313 3176 17325 3179
rect 17184 3148 17325 3176
rect 17184 3136 17190 3148
rect 17313 3145 17325 3148
rect 17359 3145 17371 3179
rect 17313 3139 17371 3145
rect 2314 3108 2320 3120
rect 2275 3080 2320 3108
rect 2314 3068 2320 3080
rect 2372 3108 2378 3120
rect 3326 3108 3332 3120
rect 2372 3080 3332 3108
rect 2372 3068 2378 3080
rect 3326 3068 3332 3080
rect 3384 3068 3390 3120
rect 3513 3111 3571 3117
rect 3513 3077 3525 3111
rect 3559 3108 3571 3111
rect 5074 3108 5080 3120
rect 3559 3080 5080 3108
rect 3559 3077 3571 3080
rect 3513 3071 3571 3077
rect 2130 3000 2136 3052
rect 2188 3040 2194 3052
rect 2409 3043 2467 3049
rect 2409 3040 2421 3043
rect 2188 3012 2421 3040
rect 2188 3000 2194 3012
rect 2409 3009 2421 3012
rect 2455 3040 2467 3043
rect 2498 3040 2504 3052
rect 2455 3012 2504 3040
rect 2455 3009 2467 3012
rect 2409 3003 2467 3009
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 2774 3040 2780 3052
rect 2735 3012 2780 3040
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2972 2099 2975
rect 2590 2972 2596 2984
rect 2087 2944 2596 2972
rect 2087 2941 2099 2944
rect 2041 2935 2099 2941
rect 2590 2932 2596 2944
rect 2648 2932 2654 2984
rect 3620 2981 3648 3080
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 7929 3111 7987 3117
rect 7929 3077 7941 3111
rect 7975 3108 7987 3111
rect 8202 3108 8208 3120
rect 7975 3080 8208 3108
rect 7975 3077 7987 3080
rect 7929 3071 7987 3077
rect 8202 3068 8208 3080
rect 8260 3108 8266 3120
rect 10321 3111 10379 3117
rect 10321 3108 10333 3111
rect 8260 3080 10333 3108
rect 8260 3068 8266 3080
rect 10321 3077 10333 3080
rect 10367 3077 10379 3111
rect 10321 3071 10379 3077
rect 14277 3111 14335 3117
rect 14277 3077 14289 3111
rect 14323 3108 14335 3111
rect 16850 3108 16856 3120
rect 14323 3080 16856 3108
rect 14323 3077 14335 3080
rect 14277 3071 14335 3077
rect 4246 3040 4252 3052
rect 4207 3012 4252 3040
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 6546 3040 6552 3052
rect 5092 3012 6552 3040
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2941 3663 2975
rect 3605 2935 3663 2941
rect 3694 2932 3700 2984
rect 3752 2972 3758 2984
rect 3878 2972 3884 2984
rect 3752 2944 3797 2972
rect 3839 2944 3884 2972
rect 3752 2932 3758 2944
rect 3878 2932 3884 2944
rect 3936 2972 3942 2984
rect 5092 2972 5120 3012
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 7006 3040 7012 3052
rect 6967 3012 7012 3040
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 8662 3000 8668 3052
rect 8720 3040 8726 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 8720 3012 8769 3040
rect 8720 3000 8726 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 9214 3000 9220 3052
rect 9272 3040 9278 3052
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 9272 3012 10517 3040
rect 9272 3000 9278 3012
rect 10505 3009 10517 3012
rect 10551 3009 10563 3043
rect 14182 3040 14188 3052
rect 10505 3003 10563 3009
rect 12452 3012 14188 3040
rect 5442 2972 5448 2984
rect 3936 2944 5120 2972
rect 5403 2944 5448 2972
rect 3936 2932 3942 2944
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 5626 2972 5632 2984
rect 5587 2944 5632 2972
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 5905 2975 5963 2981
rect 5905 2941 5917 2975
rect 5951 2972 5963 2975
rect 7742 2972 7748 2984
rect 5951 2944 7748 2972
rect 5951 2941 5963 2944
rect 5905 2935 5963 2941
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 8110 2932 8116 2984
rect 8168 2972 8174 2984
rect 10594 2972 10600 2984
rect 8168 2944 9674 2972
rect 10555 2944 10600 2972
rect 8168 2932 8174 2944
rect 106 2864 112 2916
rect 164 2904 170 2916
rect 3970 2904 3976 2916
rect 164 2876 3976 2904
rect 164 2864 170 2876
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 6549 2907 6607 2913
rect 6549 2904 6561 2907
rect 4126 2876 6561 2904
rect 3050 2836 3056 2848
rect 3011 2808 3056 2836
rect 3050 2796 3056 2808
rect 3108 2836 3114 2848
rect 4126 2836 4154 2876
rect 6549 2873 6561 2876
rect 6595 2904 6607 2907
rect 6822 2904 6828 2916
rect 6595 2876 6828 2904
rect 6595 2873 6607 2876
rect 6549 2867 6607 2873
rect 6822 2864 6828 2876
rect 6880 2864 6886 2916
rect 7371 2907 7429 2913
rect 7371 2873 7383 2907
rect 7417 2904 7429 2907
rect 7558 2904 7564 2916
rect 7417 2876 7564 2904
rect 7417 2873 7429 2876
rect 7371 2867 7429 2873
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 8754 2864 8760 2916
rect 8812 2904 8818 2916
rect 9078 2907 9136 2913
rect 9078 2904 9090 2907
rect 8812 2876 9090 2904
rect 8812 2864 8818 2876
rect 9078 2873 9090 2876
rect 9124 2873 9136 2907
rect 9646 2904 9674 2944
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 12452 2981 12480 3012
rect 14182 3000 14188 3012
rect 14240 3000 14246 3052
rect 14476 3049 14504 3080
rect 16850 3068 16856 3080
rect 16908 3068 16914 3120
rect 14461 3043 14519 3049
rect 14461 3009 14473 3043
rect 14507 3009 14519 3043
rect 15562 3040 15568 3052
rect 15523 3012 15568 3040
rect 14461 3003 14519 3009
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 16114 3000 16120 3052
rect 16172 3040 16178 3052
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 16172 3012 18061 3040
rect 16172 3000 16178 3012
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 12069 2975 12127 2981
rect 12069 2941 12081 2975
rect 12115 2972 12127 2975
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12115 2944 12449 2972
rect 12115 2941 12127 2944
rect 12069 2935 12127 2941
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12897 2975 12955 2981
rect 12897 2941 12909 2975
rect 12943 2941 12955 2975
rect 12897 2935 12955 2941
rect 12161 2907 12219 2913
rect 12161 2904 12173 2907
rect 9646 2876 12173 2904
rect 9078 2867 9136 2873
rect 12161 2873 12173 2876
rect 12207 2904 12219 2907
rect 12912 2904 12940 2935
rect 13262 2932 13268 2984
rect 13320 2972 13326 2984
rect 13541 2975 13599 2981
rect 13541 2972 13553 2975
rect 13320 2944 13553 2972
rect 13320 2932 13326 2944
rect 13541 2941 13553 2944
rect 13587 2972 13599 2975
rect 13906 2972 13912 2984
rect 13587 2944 13912 2972
rect 13587 2941 13599 2944
rect 13541 2935 13599 2941
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 15105 2975 15163 2981
rect 15105 2941 15117 2975
rect 15151 2972 15163 2975
rect 15930 2972 15936 2984
rect 15151 2944 15936 2972
rect 15151 2941 15163 2944
rect 15105 2935 15163 2941
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 16209 2975 16267 2981
rect 16209 2941 16221 2975
rect 16255 2972 16267 2975
rect 16298 2972 16304 2984
rect 16255 2944 16304 2972
rect 16255 2941 16267 2944
rect 16209 2935 16267 2941
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 16393 2975 16451 2981
rect 16393 2941 16405 2975
rect 16439 2972 16451 2975
rect 16945 2975 17003 2981
rect 16945 2972 16957 2975
rect 16439 2944 16957 2972
rect 16439 2941 16451 2944
rect 16393 2935 16451 2941
rect 16945 2941 16957 2944
rect 16991 2972 17003 2975
rect 17310 2972 17316 2984
rect 16991 2944 17316 2972
rect 16991 2941 17003 2944
rect 16945 2935 17003 2941
rect 12207 2876 12940 2904
rect 12207 2873 12219 2876
rect 12161 2867 12219 2873
rect 4706 2836 4712 2848
rect 3108 2808 4154 2836
rect 4667 2808 4712 2836
rect 3108 2796 3114 2808
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 5074 2836 5080 2848
rect 5035 2808 5080 2836
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 6270 2796 6276 2848
rect 6328 2836 6334 2848
rect 8297 2839 8355 2845
rect 8297 2836 8309 2839
rect 6328 2808 8309 2836
rect 6328 2796 6334 2808
rect 8297 2805 8309 2808
rect 8343 2836 8355 2839
rect 8662 2836 8668 2848
rect 8343 2808 8668 2836
rect 8343 2805 8355 2808
rect 8297 2799 8355 2805
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 9214 2796 9220 2848
rect 9272 2836 9278 2848
rect 11793 2839 11851 2845
rect 11793 2836 11805 2839
rect 9272 2808 11805 2836
rect 9272 2796 9278 2808
rect 11793 2805 11805 2808
rect 11839 2836 11851 2839
rect 12069 2839 12127 2845
rect 12069 2836 12081 2839
rect 11839 2808 12081 2836
rect 11839 2805 11851 2808
rect 11793 2799 11851 2805
rect 12069 2805 12081 2808
rect 12115 2805 12127 2839
rect 12710 2836 12716 2848
rect 12671 2808 12716 2836
rect 12069 2799 12127 2805
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 12912 2836 12940 2876
rect 14553 2907 14611 2913
rect 14553 2873 14565 2907
rect 14599 2904 14611 2907
rect 14642 2904 14648 2916
rect 14599 2876 14648 2904
rect 14599 2873 14611 2876
rect 14553 2867 14611 2873
rect 14642 2864 14648 2876
rect 14700 2864 14706 2916
rect 15749 2907 15807 2913
rect 15749 2904 15761 2907
rect 15120 2876 15761 2904
rect 15120 2848 15148 2876
rect 15749 2873 15761 2876
rect 15795 2904 15807 2907
rect 15795 2876 15976 2904
rect 15795 2873 15807 2876
rect 15749 2867 15807 2873
rect 15948 2848 15976 2876
rect 15102 2836 15108 2848
rect 12912 2808 15108 2836
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 15381 2839 15439 2845
rect 15381 2836 15393 2839
rect 15252 2808 15393 2836
rect 15252 2796 15258 2808
rect 15381 2805 15393 2808
rect 15427 2836 15439 2839
rect 15565 2839 15623 2845
rect 15565 2836 15577 2839
rect 15427 2808 15577 2836
rect 15427 2805 15439 2808
rect 15381 2799 15439 2805
rect 15565 2805 15577 2808
rect 15611 2805 15623 2839
rect 15565 2799 15623 2805
rect 15930 2796 15936 2848
rect 15988 2796 15994 2848
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 16408 2836 16436 2935
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 17770 2932 17776 2984
rect 17828 2972 17834 2984
rect 18141 2975 18199 2981
rect 18141 2972 18153 2975
rect 17828 2944 18153 2972
rect 17828 2932 17834 2944
rect 18141 2941 18153 2944
rect 18187 2941 18199 2975
rect 18141 2935 18199 2941
rect 16482 2864 16488 2916
rect 16540 2904 16546 2916
rect 19613 2907 19671 2913
rect 19613 2904 19625 2907
rect 16540 2876 19625 2904
rect 16540 2864 16546 2876
rect 19613 2873 19625 2876
rect 19659 2873 19671 2907
rect 19613 2867 19671 2873
rect 16172 2808 16436 2836
rect 16172 2796 16178 2808
rect 16666 2796 16672 2848
rect 16724 2836 16730 2848
rect 16761 2839 16819 2845
rect 16761 2836 16773 2839
rect 16724 2808 16773 2836
rect 16724 2796 16730 2808
rect 16761 2805 16773 2808
rect 16807 2805 16819 2839
rect 17770 2836 17776 2848
rect 17731 2808 17776 2836
rect 16761 2799 16819 2805
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 19058 2836 19064 2848
rect 19019 2808 19064 2836
rect 19058 2796 19064 2808
rect 19116 2796 19122 2848
rect 1104 2746 20884 2768
rect 1104 2694 8315 2746
rect 8367 2694 8379 2746
rect 8431 2694 8443 2746
rect 8495 2694 8507 2746
rect 8559 2694 15648 2746
rect 15700 2694 15712 2746
rect 15764 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 20884 2746
rect 1104 2672 20884 2694
rect 3694 2632 3700 2644
rect 3655 2604 3700 2632
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 4341 2635 4399 2641
rect 4341 2601 4353 2635
rect 4387 2632 4399 2635
rect 8202 2632 8208 2644
rect 4387 2604 8208 2632
rect 4387 2601 4399 2604
rect 4341 2595 4399 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 9214 2632 9220 2644
rect 8527 2604 9220 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9306 2592 9312 2644
rect 9364 2632 9370 2644
rect 9861 2635 9919 2641
rect 9861 2632 9873 2635
rect 9364 2604 9873 2632
rect 9364 2592 9370 2604
rect 9861 2601 9873 2604
rect 9907 2601 9919 2635
rect 9861 2595 9919 2601
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 10781 2635 10839 2641
rect 10781 2632 10793 2635
rect 10192 2604 10793 2632
rect 10192 2592 10198 2604
rect 10781 2601 10793 2604
rect 10827 2601 10839 2635
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 10781 2595 10839 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 12805 2635 12863 2641
rect 12805 2632 12817 2635
rect 12768 2604 12817 2632
rect 12768 2592 12774 2604
rect 12805 2601 12817 2604
rect 12851 2601 12863 2635
rect 13262 2632 13268 2644
rect 13223 2604 13268 2632
rect 12805 2595 12863 2601
rect 2961 2567 3019 2573
rect 2961 2533 2973 2567
rect 3007 2564 3019 2567
rect 3602 2564 3608 2576
rect 3007 2536 3608 2564
rect 3007 2533 3019 2536
rect 2961 2527 3019 2533
rect 3602 2524 3608 2536
rect 3660 2524 3666 2576
rect 4706 2524 4712 2576
rect 4764 2564 4770 2576
rect 4801 2567 4859 2573
rect 4801 2564 4813 2567
rect 4764 2536 4813 2564
rect 4764 2524 4770 2536
rect 4801 2533 4813 2536
rect 4847 2564 4859 2567
rect 4847 2536 5580 2564
rect 4847 2533 4859 2536
rect 4801 2527 4859 2533
rect 5552 2508 5580 2536
rect 5626 2524 5632 2576
rect 5684 2564 5690 2576
rect 6641 2567 6699 2573
rect 6641 2564 6653 2567
rect 5684 2536 6653 2564
rect 5684 2524 5690 2536
rect 6641 2533 6653 2536
rect 6687 2564 6699 2567
rect 9490 2564 9496 2576
rect 6687 2536 9496 2564
rect 6687 2533 6699 2536
rect 6641 2527 6699 2533
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2496 2283 2499
rect 2271 2468 2452 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 2314 2360 2320 2372
rect 2056 2332 2320 2360
rect 1670 2292 1676 2304
rect 1631 2264 1676 2292
rect 1670 2252 1676 2264
rect 1728 2292 1734 2304
rect 2056 2301 2084 2332
rect 2314 2320 2320 2332
rect 2372 2320 2378 2372
rect 2424 2360 2452 2468
rect 2498 2456 2504 2508
rect 2556 2496 2562 2508
rect 3329 2499 3387 2505
rect 2556 2468 2601 2496
rect 2556 2456 2562 2468
rect 3329 2465 3341 2499
rect 3375 2496 3387 2499
rect 4157 2499 4215 2505
rect 4157 2496 4169 2499
rect 3375 2468 4169 2496
rect 3375 2465 3387 2468
rect 3329 2459 3387 2465
rect 4157 2465 4169 2468
rect 4203 2496 4215 2499
rect 4522 2496 4528 2508
rect 4203 2468 4528 2496
rect 4203 2465 4215 2468
rect 4157 2459 4215 2465
rect 4522 2456 4528 2468
rect 4580 2496 4586 2508
rect 4580 2468 5120 2496
rect 4580 2456 4586 2468
rect 5092 2428 5120 2468
rect 5166 2456 5172 2508
rect 5224 2496 5230 2508
rect 5261 2499 5319 2505
rect 5261 2496 5273 2499
rect 5224 2468 5273 2496
rect 5224 2456 5230 2468
rect 5261 2465 5273 2468
rect 5307 2465 5319 2499
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 5261 2459 5319 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 7193 2499 7251 2505
rect 5868 2468 6408 2496
rect 5868 2456 5874 2468
rect 5718 2428 5724 2440
rect 3160 2400 5028 2428
rect 5092 2400 5724 2428
rect 3160 2360 3188 2400
rect 2424 2332 3188 2360
rect 3694 2320 3700 2372
rect 3752 2360 3758 2372
rect 4522 2360 4528 2372
rect 3752 2332 4528 2360
rect 3752 2320 3758 2332
rect 4522 2320 4528 2332
rect 4580 2320 4586 2372
rect 5000 2360 5028 2400
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 6380 2437 6408 2468
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 7282 2496 7288 2508
rect 7239 2468 7288 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 7392 2505 7420 2536
rect 9490 2524 9496 2536
rect 9548 2564 9554 2576
rect 12069 2567 12127 2573
rect 9548 2536 10272 2564
rect 9548 2524 9554 2536
rect 7377 2499 7435 2505
rect 7377 2465 7389 2499
rect 7423 2465 7435 2499
rect 7377 2459 7435 2465
rect 7558 2456 7564 2508
rect 7616 2496 7622 2508
rect 8297 2499 8355 2505
rect 8297 2496 8309 2499
rect 7616 2468 8309 2496
rect 7616 2456 7622 2468
rect 8297 2465 8309 2468
rect 8343 2496 8355 2499
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 8343 2468 8493 2496
rect 8343 2465 8355 2468
rect 8297 2459 8355 2465
rect 8481 2465 8493 2468
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8619 2468 9137 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 9309 2499 9367 2505
rect 9309 2465 9321 2499
rect 9355 2496 9367 2499
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9355 2468 9781 2496
rect 9355 2465 9367 2468
rect 9309 2459 9367 2465
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 10134 2496 10140 2508
rect 9815 2468 10140 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2397 6055 2431
rect 5997 2391 6055 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 6454 2428 6460 2440
rect 6411 2400 6460 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 5350 2360 5356 2372
rect 5000 2332 5212 2360
rect 5263 2332 5356 2360
rect 2041 2295 2099 2301
rect 2041 2292 2053 2295
rect 1728 2264 2053 2292
rect 1728 2252 1734 2264
rect 2041 2261 2053 2264
rect 2087 2261 2099 2295
rect 5074 2292 5080 2304
rect 5035 2264 5080 2292
rect 2041 2255 2099 2261
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 5184 2292 5212 2332
rect 5350 2320 5356 2332
rect 5408 2360 5414 2372
rect 5810 2360 5816 2372
rect 5408 2332 5816 2360
rect 5408 2320 5414 2332
rect 5810 2320 5816 2332
rect 5868 2320 5874 2372
rect 6012 2360 6040 2391
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7064 2400 7481 2428
rect 7064 2388 7070 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 9140 2428 9168 2459
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 10244 2505 10272 2536
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 12618 2564 12624 2576
rect 12115 2536 12624 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2465 10287 2499
rect 10229 2459 10287 2465
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 12084 2496 12112 2527
rect 12618 2524 12624 2536
rect 12676 2524 12682 2576
rect 11471 2468 12112 2496
rect 12820 2496 12848 2595
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 14642 2632 14648 2644
rect 14323 2604 14648 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 14642 2592 14648 2604
rect 14700 2592 14706 2644
rect 16574 2632 16580 2644
rect 15580 2604 16580 2632
rect 13280 2564 13308 2592
rect 13678 2567 13736 2573
rect 13678 2564 13690 2567
rect 13280 2536 13690 2564
rect 13678 2533 13690 2536
rect 13724 2533 13736 2567
rect 13678 2527 13736 2533
rect 15580 2508 15608 2604
rect 16574 2592 16580 2604
rect 16632 2592 16638 2644
rect 17494 2592 17500 2644
rect 17552 2632 17558 2644
rect 17589 2635 17647 2641
rect 17589 2632 17601 2635
rect 17552 2604 17601 2632
rect 17552 2592 17558 2604
rect 17589 2601 17601 2604
rect 17635 2601 17647 2635
rect 18782 2632 18788 2644
rect 18743 2604 18788 2632
rect 17589 2595 17647 2601
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 13357 2499 13415 2505
rect 13357 2496 13369 2499
rect 12820 2468 13369 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 13357 2465 13369 2468
rect 13403 2465 13415 2499
rect 13357 2459 13415 2465
rect 14826 2456 14832 2508
rect 14884 2496 14890 2508
rect 15286 2496 15292 2508
rect 14884 2468 15292 2496
rect 14884 2456 14890 2468
rect 15286 2456 15292 2468
rect 15344 2496 15350 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15344 2468 15485 2496
rect 15344 2456 15350 2468
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 15562 2456 15568 2508
rect 15620 2496 15626 2508
rect 15620 2468 15713 2496
rect 15620 2456 15626 2468
rect 15746 2456 15752 2508
rect 15804 2496 15810 2508
rect 16758 2496 16764 2508
rect 15804 2468 16764 2496
rect 15804 2456 15810 2468
rect 16758 2456 16764 2468
rect 16816 2456 16822 2508
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2496 17095 2499
rect 17512 2496 17540 2592
rect 17083 2468 17540 2496
rect 17083 2465 17095 2468
rect 17037 2459 17095 2465
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 18417 2499 18475 2505
rect 18417 2496 18429 2499
rect 18104 2468 18429 2496
rect 18104 2456 18110 2468
rect 18417 2465 18429 2468
rect 18463 2465 18475 2499
rect 18417 2459 18475 2465
rect 13630 2428 13636 2440
rect 9140 2400 13636 2428
rect 7469 2391 7527 2397
rect 13630 2388 13636 2400
rect 13688 2388 13694 2440
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 14918 2428 14924 2440
rect 14240 2400 14924 2428
rect 14240 2388 14246 2400
rect 14918 2388 14924 2400
rect 14976 2428 14982 2440
rect 15933 2431 15991 2437
rect 15933 2428 15945 2431
rect 14976 2400 15945 2428
rect 14976 2388 14982 2400
rect 15933 2397 15945 2400
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 7098 2360 7104 2372
rect 6012 2332 7104 2360
rect 7098 2320 7104 2332
rect 7156 2360 7162 2372
rect 8757 2363 8815 2369
rect 7156 2332 8156 2360
rect 7156 2320 7162 2332
rect 7650 2292 7656 2304
rect 5184 2264 7656 2292
rect 7650 2252 7656 2264
rect 7708 2292 7714 2304
rect 8018 2292 8024 2304
rect 7708 2264 8024 2292
rect 7708 2252 7714 2264
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 8128 2292 8156 2332
rect 8757 2329 8769 2363
rect 8803 2360 8815 2363
rect 10042 2360 10048 2372
rect 8803 2332 10048 2360
rect 8803 2329 8815 2332
rect 8757 2323 8815 2329
rect 10042 2320 10048 2332
rect 10100 2320 10106 2372
rect 11609 2363 11667 2369
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 15378 2360 15384 2372
rect 11655 2332 15384 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 15378 2320 15384 2332
rect 15436 2320 15442 2372
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 8128 2264 9321 2292
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 14826 2292 14832 2304
rect 14787 2264 14832 2292
rect 9309 2255 9367 2261
rect 14826 2252 14832 2264
rect 14884 2252 14890 2304
rect 15102 2252 15108 2304
rect 15160 2292 15166 2304
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 15160 2264 15209 2292
rect 15160 2252 15166 2264
rect 15197 2261 15209 2264
rect 15243 2292 15255 2295
rect 15746 2292 15752 2304
rect 15243 2264 15752 2292
rect 15243 2261 15255 2264
rect 15197 2255 15255 2261
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 17218 2292 17224 2304
rect 17179 2264 17224 2292
rect 17218 2252 17224 2264
rect 17276 2252 17282 2304
rect 18046 2292 18052 2304
rect 18007 2264 18052 2292
rect 18046 2252 18052 2264
rect 18104 2252 18110 2304
rect 1104 2202 20884 2224
rect 1104 2150 4648 2202
rect 4700 2150 4712 2202
rect 4764 2150 4776 2202
rect 4828 2150 4840 2202
rect 4892 2150 11982 2202
rect 12034 2150 12046 2202
rect 12098 2150 12110 2202
rect 12162 2150 12174 2202
rect 12226 2150 19315 2202
rect 19367 2150 19379 2202
rect 19431 2150 19443 2202
rect 19495 2150 19507 2202
rect 19559 2150 20884 2202
rect 1104 2128 20884 2150
rect 4522 2048 4528 2100
rect 4580 2088 4586 2100
rect 5350 2088 5356 2100
rect 4580 2060 5356 2088
rect 4580 2048 4586 2060
rect 5350 2048 5356 2060
rect 5408 2048 5414 2100
rect 8018 1980 8024 2032
rect 8076 2020 8082 2032
rect 18414 2020 18420 2032
rect 8076 1992 18420 2020
rect 8076 1980 8082 1992
rect 18414 1980 18420 1992
rect 18472 1980 18478 2032
rect 12066 1912 12072 1964
rect 12124 1952 12130 1964
rect 18506 1952 18512 1964
rect 12124 1924 18512 1952
rect 12124 1912 12130 1924
rect 18506 1912 18512 1924
rect 18564 1912 18570 1964
<< via1 >>
rect 4648 19558 4700 19610
rect 4712 19558 4764 19610
rect 4776 19558 4828 19610
rect 4840 19558 4892 19610
rect 11982 19558 12034 19610
rect 12046 19558 12098 19610
rect 12110 19558 12162 19610
rect 12174 19558 12226 19610
rect 19315 19558 19367 19610
rect 19379 19558 19431 19610
rect 19443 19558 19495 19610
rect 19507 19558 19559 19610
rect 2872 19456 2924 19508
rect 1124 19252 1176 19304
rect 5264 19295 5316 19304
rect 5264 19261 5273 19295
rect 5273 19261 5307 19295
rect 5307 19261 5316 19295
rect 5264 19252 5316 19261
rect 1308 19184 1360 19236
rect 6276 19252 6328 19304
rect 6000 19227 6052 19236
rect 6000 19193 6009 19227
rect 6009 19193 6043 19227
rect 6043 19193 6052 19227
rect 6000 19184 6052 19193
rect 1492 19116 1544 19168
rect 4068 19159 4120 19168
rect 4068 19125 4077 19159
rect 4077 19125 4111 19159
rect 4111 19125 4120 19159
rect 4068 19116 4120 19125
rect 5632 19116 5684 19168
rect 6920 19159 6972 19168
rect 6920 19125 6929 19159
rect 6929 19125 6963 19159
rect 6963 19125 6972 19159
rect 6920 19116 6972 19125
rect 8208 19116 8260 19168
rect 9220 19116 9272 19168
rect 10324 19159 10376 19168
rect 10324 19125 10333 19159
rect 10333 19125 10367 19159
rect 10367 19125 10376 19159
rect 10324 19116 10376 19125
rect 11152 19116 11204 19168
rect 8315 19014 8367 19066
rect 8379 19014 8431 19066
rect 8443 19014 8495 19066
rect 8507 19014 8559 19066
rect 15648 19014 15700 19066
rect 15712 19014 15764 19066
rect 15776 19014 15828 19066
rect 15840 19014 15892 19066
rect 2228 18955 2280 18964
rect 2228 18921 2237 18955
rect 2237 18921 2271 18955
rect 2271 18921 2280 18955
rect 2228 18912 2280 18921
rect 5080 18912 5132 18964
rect 5264 18955 5316 18964
rect 5264 18921 5273 18955
rect 5273 18921 5307 18955
rect 5307 18921 5316 18955
rect 5264 18912 5316 18921
rect 6552 18912 6604 18964
rect 21548 18912 21600 18964
rect 2320 18776 2372 18828
rect 5080 18776 5132 18828
rect 6092 18776 6144 18828
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 7564 18819 7616 18828
rect 7564 18785 7573 18819
rect 7573 18785 7607 18819
rect 7607 18785 7616 18819
rect 7564 18776 7616 18785
rect 7840 18819 7892 18828
rect 7840 18785 7849 18819
rect 7849 18785 7883 18819
rect 7883 18785 7892 18819
rect 7840 18776 7892 18785
rect 9680 18776 9732 18828
rect 11428 18819 11480 18828
rect 11428 18785 11437 18819
rect 11437 18785 11471 18819
rect 11471 18785 11480 18819
rect 11428 18776 11480 18785
rect 6368 18751 6420 18760
rect 6368 18717 6377 18751
rect 6377 18717 6411 18751
rect 6411 18717 6420 18751
rect 6368 18708 6420 18717
rect 2688 18640 2740 18692
rect 5264 18640 5316 18692
rect 1860 18572 1912 18624
rect 3056 18615 3108 18624
rect 3056 18581 3065 18615
rect 3065 18581 3099 18615
rect 3099 18581 3108 18615
rect 3056 18572 3108 18581
rect 8944 18572 8996 18624
rect 4648 18470 4700 18522
rect 4712 18470 4764 18522
rect 4776 18470 4828 18522
rect 4840 18470 4892 18522
rect 11982 18470 12034 18522
rect 12046 18470 12098 18522
rect 12110 18470 12162 18522
rect 12174 18470 12226 18522
rect 19315 18470 19367 18522
rect 19379 18470 19431 18522
rect 19443 18470 19495 18522
rect 19507 18470 19559 18522
rect 7840 18411 7892 18420
rect 3516 18300 3568 18352
rect 7840 18377 7849 18411
rect 7849 18377 7883 18411
rect 7883 18377 7892 18411
rect 7840 18368 7892 18377
rect 14280 18368 14332 18420
rect 16028 18368 16080 18420
rect 18328 18368 18380 18420
rect 1308 18164 1360 18216
rect 3056 18207 3108 18216
rect 1860 18096 1912 18148
rect 3056 18173 3065 18207
rect 3065 18173 3099 18207
rect 3099 18173 3108 18207
rect 3056 18164 3108 18173
rect 4344 18164 4396 18216
rect 8116 18300 8168 18352
rect 5264 18275 5316 18284
rect 5264 18241 5273 18275
rect 5273 18241 5307 18275
rect 5307 18241 5316 18275
rect 5264 18232 5316 18241
rect 6276 18232 6328 18284
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 7840 18164 7892 18216
rect 6092 18096 6144 18148
rect 7656 18096 7708 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 3056 18071 3108 18080
rect 3056 18037 3065 18071
rect 3065 18037 3099 18071
rect 3099 18037 3108 18071
rect 3056 18028 3108 18037
rect 3148 18028 3200 18080
rect 6736 18028 6788 18080
rect 8668 18028 8720 18080
rect 9404 18164 9456 18216
rect 10692 18164 10744 18216
rect 13636 18207 13688 18216
rect 13636 18173 13645 18207
rect 13645 18173 13679 18207
rect 13679 18173 13688 18207
rect 13636 18164 13688 18173
rect 16856 18207 16908 18216
rect 9772 18139 9824 18148
rect 9772 18105 9781 18139
rect 9781 18105 9815 18139
rect 9815 18105 9824 18139
rect 9772 18096 9824 18105
rect 16856 18173 16865 18207
rect 16865 18173 16899 18207
rect 16899 18173 16908 18207
rect 16856 18164 16908 18173
rect 9680 18028 9732 18080
rect 10600 18071 10652 18080
rect 10600 18037 10609 18071
rect 10609 18037 10643 18071
rect 10643 18037 10652 18071
rect 10600 18028 10652 18037
rect 10876 18028 10928 18080
rect 11428 18071 11480 18080
rect 11428 18037 11437 18071
rect 11437 18037 11471 18071
rect 11471 18037 11480 18071
rect 11428 18028 11480 18037
rect 15936 18028 15988 18080
rect 8315 17926 8367 17978
rect 8379 17926 8431 17978
rect 8443 17926 8495 17978
rect 8507 17926 8559 17978
rect 15648 17926 15700 17978
rect 15712 17926 15764 17978
rect 15776 17926 15828 17978
rect 15840 17926 15892 17978
rect 2320 17824 2372 17876
rect 3148 17824 3200 17876
rect 2688 17756 2740 17808
rect 3976 17756 4028 17808
rect 7564 17824 7616 17876
rect 9496 17824 9548 17876
rect 10600 17824 10652 17876
rect 20444 17824 20496 17876
rect 9404 17756 9456 17808
rect 16856 17756 16908 17808
rect 1584 17731 1636 17740
rect 1584 17697 1593 17731
rect 1593 17697 1627 17731
rect 1627 17697 1636 17731
rect 1584 17688 1636 17697
rect 1860 17731 1912 17740
rect 1860 17697 1869 17731
rect 1869 17697 1903 17731
rect 1903 17697 1912 17731
rect 1860 17688 1912 17697
rect 1768 17620 1820 17672
rect 2964 17552 3016 17604
rect 2780 17527 2832 17536
rect 2780 17493 2789 17527
rect 2789 17493 2823 17527
rect 2823 17493 2832 17527
rect 2780 17484 2832 17493
rect 3884 17688 3936 17740
rect 4160 17688 4212 17740
rect 5724 17731 5776 17740
rect 5724 17697 5733 17731
rect 5733 17697 5767 17731
rect 5767 17697 5776 17731
rect 5724 17688 5776 17697
rect 6276 17731 6328 17740
rect 6276 17697 6285 17731
rect 6285 17697 6319 17731
rect 6319 17697 6328 17731
rect 6276 17688 6328 17697
rect 8116 17731 8168 17740
rect 8116 17697 8125 17731
rect 8125 17697 8159 17731
rect 8159 17697 8168 17731
rect 8116 17688 8168 17697
rect 8576 17731 8628 17740
rect 8576 17697 8585 17731
rect 8585 17697 8619 17731
rect 8619 17697 8628 17731
rect 8576 17688 8628 17697
rect 9956 17731 10008 17740
rect 9956 17697 9965 17731
rect 9965 17697 9999 17731
rect 9999 17697 10008 17731
rect 9956 17688 10008 17697
rect 3608 17484 3660 17536
rect 4528 17620 4580 17672
rect 6460 17663 6512 17672
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 8760 17663 8812 17672
rect 8760 17629 8769 17663
rect 8769 17629 8803 17663
rect 8803 17629 8812 17663
rect 8760 17620 8812 17629
rect 11336 17688 11388 17740
rect 12348 17731 12400 17740
rect 12348 17697 12366 17731
rect 12366 17697 12400 17731
rect 12348 17688 12400 17697
rect 13452 17688 13504 17740
rect 15292 17688 15344 17740
rect 5172 17552 5224 17604
rect 7564 17552 7616 17604
rect 10048 17552 10100 17604
rect 10140 17552 10192 17604
rect 4436 17484 4488 17536
rect 5080 17527 5132 17536
rect 5080 17493 5089 17527
rect 5089 17493 5123 17527
rect 5123 17493 5132 17527
rect 5080 17484 5132 17493
rect 6184 17484 6236 17536
rect 6828 17527 6880 17536
rect 6828 17493 6837 17527
rect 6837 17493 6871 17527
rect 6871 17493 6880 17527
rect 6828 17484 6880 17493
rect 7380 17484 7432 17536
rect 10968 17484 11020 17536
rect 12532 17484 12584 17536
rect 4648 17382 4700 17434
rect 4712 17382 4764 17434
rect 4776 17382 4828 17434
rect 4840 17382 4892 17434
rect 11982 17382 12034 17434
rect 12046 17382 12098 17434
rect 12110 17382 12162 17434
rect 12174 17382 12226 17434
rect 19315 17382 19367 17434
rect 19379 17382 19431 17434
rect 19443 17382 19495 17434
rect 19507 17382 19559 17434
rect 1860 17280 1912 17332
rect 20 17212 72 17264
rect 6276 17323 6328 17332
rect 6276 17289 6285 17323
rect 6285 17289 6319 17323
rect 6319 17289 6328 17323
rect 6276 17280 6328 17289
rect 6644 17280 6696 17332
rect 12348 17280 12400 17332
rect 13452 17323 13504 17332
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 15936 17280 15988 17332
rect 4344 17212 4396 17264
rect 3884 17144 3936 17196
rect 3608 17076 3660 17128
rect 3976 17119 4028 17128
rect 3976 17085 3985 17119
rect 3985 17085 4019 17119
rect 4019 17085 4028 17119
rect 3976 17076 4028 17085
rect 4344 17119 4396 17128
rect 4344 17085 4353 17119
rect 4353 17085 4387 17119
rect 4387 17085 4396 17119
rect 4344 17076 4396 17085
rect 6920 17187 6972 17196
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 1584 16940 1636 16992
rect 1860 16940 1912 16992
rect 2780 17008 2832 17060
rect 4436 17008 4488 17060
rect 6276 17008 6328 17060
rect 7380 17008 7432 17060
rect 9404 17212 9456 17264
rect 7656 17144 7708 17196
rect 10600 17144 10652 17196
rect 8576 17076 8628 17128
rect 9036 17119 9088 17128
rect 7932 17008 7984 17060
rect 2872 16940 2924 16992
rect 3884 16983 3936 16992
rect 3884 16949 3893 16983
rect 3893 16949 3927 16983
rect 3927 16949 3936 16983
rect 3884 16940 3936 16949
rect 4160 16940 4212 16992
rect 5356 16940 5408 16992
rect 5724 16940 5776 16992
rect 8116 16983 8168 16992
rect 8116 16949 8125 16983
rect 8125 16949 8159 16983
rect 8159 16949 8168 16983
rect 8116 16940 8168 16949
rect 9036 17085 9045 17119
rect 9045 17085 9079 17119
rect 9079 17085 9088 17119
rect 9036 17076 9088 17085
rect 12624 17076 12676 17128
rect 9312 17051 9364 17060
rect 9312 17017 9321 17051
rect 9321 17017 9355 17051
rect 9355 17017 9364 17051
rect 9312 17008 9364 17017
rect 10600 17008 10652 17060
rect 10876 17051 10928 17060
rect 10876 17017 10885 17051
rect 10885 17017 10919 17051
rect 10919 17017 10928 17051
rect 10876 17008 10928 17017
rect 9956 16940 10008 16992
rect 10508 16940 10560 16992
rect 11336 16983 11388 16992
rect 11336 16949 11345 16983
rect 11345 16949 11379 16983
rect 11379 16949 11388 16983
rect 11336 16940 11388 16949
rect 11520 16940 11572 16992
rect 13452 17008 13504 17060
rect 14556 17051 14608 17060
rect 14556 17017 14565 17051
rect 14565 17017 14599 17051
rect 14599 17017 14608 17051
rect 14556 17008 14608 17017
rect 15292 16940 15344 16992
rect 8315 16838 8367 16890
rect 8379 16838 8431 16890
rect 8443 16838 8495 16890
rect 8507 16838 8559 16890
rect 15648 16838 15700 16890
rect 15712 16838 15764 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 1952 16779 2004 16788
rect 1952 16745 1961 16779
rect 1961 16745 1995 16779
rect 1995 16745 2004 16779
rect 1952 16736 2004 16745
rect 2780 16736 2832 16788
rect 2872 16779 2924 16788
rect 2872 16745 2881 16779
rect 2881 16745 2915 16779
rect 2915 16745 2924 16779
rect 2872 16736 2924 16745
rect 4068 16736 4120 16788
rect 6276 16736 6328 16788
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 8668 16736 8720 16788
rect 9956 16736 10008 16788
rect 10600 16779 10652 16788
rect 10600 16745 10609 16779
rect 10609 16745 10643 16779
rect 10643 16745 10652 16779
rect 10600 16736 10652 16745
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 14556 16736 14608 16788
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 5724 16668 5776 16720
rect 7472 16711 7524 16720
rect 7472 16677 7481 16711
rect 7481 16677 7515 16711
rect 7515 16677 7524 16711
rect 7472 16668 7524 16677
rect 7656 16668 7708 16720
rect 8116 16668 8168 16720
rect 13268 16668 13320 16720
rect 2136 16600 2188 16652
rect 3056 16600 3108 16652
rect 5264 16643 5316 16652
rect 5264 16609 5273 16643
rect 5273 16609 5307 16643
rect 5307 16609 5316 16643
rect 5264 16600 5316 16609
rect 8760 16600 8812 16652
rect 11244 16600 11296 16652
rect 11796 16643 11848 16652
rect 11796 16609 11805 16643
rect 11805 16609 11839 16643
rect 11839 16609 11848 16643
rect 11796 16600 11848 16609
rect 4252 16532 4304 16584
rect 5448 16532 5500 16584
rect 6644 16532 6696 16584
rect 8024 16532 8076 16584
rect 8392 16532 8444 16584
rect 11520 16532 11572 16584
rect 3056 16464 3108 16516
rect 3976 16464 4028 16516
rect 4528 16464 4580 16516
rect 7932 16507 7984 16516
rect 7932 16473 7941 16507
rect 7941 16473 7975 16507
rect 7975 16473 7984 16507
rect 7932 16464 7984 16473
rect 10048 16464 10100 16516
rect 14924 16600 14976 16652
rect 16120 16600 16172 16652
rect 19064 16643 19116 16652
rect 19064 16609 19073 16643
rect 19073 16609 19107 16643
rect 19107 16609 19116 16643
rect 19064 16600 19116 16609
rect 13176 16575 13228 16584
rect 13176 16541 13185 16575
rect 13185 16541 13219 16575
rect 13219 16541 13228 16575
rect 13176 16532 13228 16541
rect 12440 16464 12492 16516
rect 2964 16396 3016 16448
rect 5172 16396 5224 16448
rect 8668 16439 8720 16448
rect 8668 16405 8677 16439
rect 8677 16405 8711 16439
rect 8711 16405 8720 16439
rect 8668 16396 8720 16405
rect 9036 16396 9088 16448
rect 12624 16396 12676 16448
rect 16672 16396 16724 16448
rect 4648 16294 4700 16346
rect 4712 16294 4764 16346
rect 4776 16294 4828 16346
rect 4840 16294 4892 16346
rect 11982 16294 12034 16346
rect 12046 16294 12098 16346
rect 12110 16294 12162 16346
rect 12174 16294 12226 16346
rect 19315 16294 19367 16346
rect 19379 16294 19431 16346
rect 19443 16294 19495 16346
rect 19507 16294 19559 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 1952 16192 2004 16244
rect 4252 16235 4304 16244
rect 4252 16201 4261 16235
rect 4261 16201 4295 16235
rect 4295 16201 4304 16235
rect 4252 16192 4304 16201
rect 6368 16192 6420 16244
rect 7472 16192 7524 16244
rect 8392 16235 8444 16244
rect 8392 16201 8401 16235
rect 8401 16201 8435 16235
rect 8435 16201 8444 16235
rect 8392 16192 8444 16201
rect 9864 16192 9916 16244
rect 11244 16235 11296 16244
rect 11244 16201 11253 16235
rect 11253 16201 11287 16235
rect 11287 16201 11296 16235
rect 11244 16192 11296 16201
rect 11796 16192 11848 16244
rect 16488 16192 16540 16244
rect 4436 16124 4488 16176
rect 4620 16124 4672 16176
rect 4528 16056 4580 16108
rect 10416 16124 10468 16176
rect 9772 16056 9824 16108
rect 13636 16056 13688 16108
rect 3608 16031 3660 16040
rect 3608 15997 3617 16031
rect 3617 15997 3651 16031
rect 3651 15997 3660 16031
rect 3608 15988 3660 15997
rect 4436 15988 4488 16040
rect 13360 16031 13412 16040
rect 2964 15963 3016 15972
rect 2964 15929 2973 15963
rect 2973 15929 3007 15963
rect 3007 15929 3016 15963
rect 2964 15920 3016 15929
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 5080 15920 5132 15972
rect 5356 15963 5408 15972
rect 5356 15929 5365 15963
rect 5365 15929 5399 15963
rect 5399 15929 5408 15963
rect 5356 15920 5408 15929
rect 13360 15997 13369 16031
rect 13369 15997 13403 16031
rect 13403 15997 13412 16031
rect 13360 15988 13412 15997
rect 3148 15852 3200 15904
rect 5724 15895 5776 15904
rect 5724 15861 5733 15895
rect 5733 15861 5767 15895
rect 5767 15861 5776 15895
rect 6644 15895 6696 15904
rect 5724 15852 5776 15861
rect 6644 15861 6653 15895
rect 6653 15861 6687 15895
rect 6687 15861 6696 15895
rect 6644 15852 6696 15861
rect 9588 15920 9640 15972
rect 13268 15920 13320 15972
rect 9864 15852 9916 15904
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 11520 15852 11572 15904
rect 14280 15895 14332 15904
rect 14280 15861 14289 15895
rect 14289 15861 14323 15895
rect 14323 15861 14332 15895
rect 14280 15852 14332 15861
rect 14464 15852 14516 15904
rect 15936 15852 15988 15904
rect 16120 15852 16172 15904
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 8315 15750 8367 15802
rect 8379 15750 8431 15802
rect 8443 15750 8495 15802
rect 8507 15750 8559 15802
rect 15648 15750 15700 15802
rect 15712 15750 15764 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 3148 15691 3200 15700
rect 3148 15657 3157 15691
rect 3157 15657 3191 15691
rect 3191 15657 3200 15691
rect 3148 15648 3200 15657
rect 5264 15691 5316 15700
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 6460 15691 6512 15700
rect 6460 15657 6469 15691
rect 6469 15657 6503 15691
rect 6503 15657 6512 15691
rect 9864 15691 9916 15700
rect 6460 15648 6512 15657
rect 1952 15580 2004 15632
rect 4252 15623 4304 15632
rect 4252 15589 4261 15623
rect 4261 15589 4295 15623
rect 4295 15589 4304 15623
rect 4252 15580 4304 15589
rect 2228 15555 2280 15564
rect 2228 15521 2237 15555
rect 2237 15521 2271 15555
rect 2271 15521 2280 15555
rect 2228 15512 2280 15521
rect 9864 15657 9873 15691
rect 9873 15657 9907 15691
rect 9907 15657 9916 15691
rect 9864 15648 9916 15657
rect 11796 15648 11848 15700
rect 13176 15691 13228 15700
rect 6644 15580 6696 15632
rect 13176 15657 13185 15691
rect 13185 15657 13219 15691
rect 13219 15657 13228 15691
rect 13176 15648 13228 15657
rect 13268 15580 13320 15632
rect 15476 15623 15528 15632
rect 15476 15589 15485 15623
rect 15485 15589 15519 15623
rect 15519 15589 15528 15623
rect 15476 15580 15528 15589
rect 7748 15512 7800 15564
rect 8300 15555 8352 15564
rect 8300 15521 8344 15555
rect 8344 15521 8352 15555
rect 8300 15512 8352 15521
rect 9312 15512 9364 15564
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 13452 15555 13504 15564
rect 13452 15521 13461 15555
rect 13461 15521 13495 15555
rect 13495 15521 13504 15555
rect 13452 15512 13504 15521
rect 16948 15512 17000 15564
rect 3792 15444 3844 15496
rect 4436 15487 4488 15496
rect 4436 15453 4445 15487
rect 4445 15453 4479 15487
rect 4479 15453 4488 15487
rect 4436 15444 4488 15453
rect 5540 15444 5592 15496
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 15660 15487 15712 15496
rect 15660 15453 15669 15487
rect 15669 15453 15703 15487
rect 15703 15453 15712 15487
rect 15660 15444 15712 15453
rect 7380 15376 7432 15428
rect 7840 15419 7892 15428
rect 7840 15385 7849 15419
rect 7849 15385 7883 15419
rect 7883 15385 7892 15419
rect 7840 15376 7892 15385
rect 9036 15376 9088 15428
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 11612 15308 11664 15360
rect 14096 15308 14148 15360
rect 4648 15206 4700 15258
rect 4712 15206 4764 15258
rect 4776 15206 4828 15258
rect 4840 15206 4892 15258
rect 11982 15206 12034 15258
rect 12046 15206 12098 15258
rect 12110 15206 12162 15258
rect 12174 15206 12226 15258
rect 19315 15206 19367 15258
rect 19379 15206 19431 15258
rect 19443 15206 19495 15258
rect 19507 15206 19559 15258
rect 4252 15104 4304 15156
rect 5356 15104 5408 15156
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 8300 15104 8352 15113
rect 9864 15104 9916 15156
rect 10600 15147 10652 15156
rect 10600 15113 10609 15147
rect 10609 15113 10643 15147
rect 10643 15113 10652 15147
rect 10600 15104 10652 15113
rect 11796 15147 11848 15156
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 11796 15104 11848 15113
rect 13452 15104 13504 15156
rect 14280 15147 14332 15156
rect 14280 15113 14289 15147
rect 14289 15113 14323 15147
rect 14323 15113 14332 15147
rect 14280 15104 14332 15113
rect 15476 15147 15528 15156
rect 15476 15113 15485 15147
rect 15485 15113 15519 15147
rect 15519 15113 15528 15147
rect 15476 15104 15528 15113
rect 4712 15036 4764 15088
rect 7932 15079 7984 15088
rect 7932 15045 7941 15079
rect 7941 15045 7975 15079
rect 7975 15045 7984 15079
rect 7932 15036 7984 15045
rect 10692 15036 10744 15088
rect 10876 15036 10928 15088
rect 12348 15036 12400 15088
rect 15384 15036 15436 15088
rect 16028 15036 16080 15088
rect 21548 15036 21600 15088
rect 1676 15011 1728 15020
rect 1676 14977 1685 15011
rect 1685 14977 1719 15011
rect 1719 14977 1728 15011
rect 1676 14968 1728 14977
rect 3884 15011 3936 15020
rect 3884 14977 3893 15011
rect 3893 14977 3927 15011
rect 3927 14977 3936 15011
rect 3884 14968 3936 14977
rect 6644 14968 6696 15020
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 8944 15011 8996 15020
rect 8944 14977 8953 15011
rect 8953 14977 8987 15011
rect 8987 14977 8996 15011
rect 8944 14968 8996 14977
rect 9036 14968 9088 15020
rect 11612 14968 11664 15020
rect 13360 14968 13412 15020
rect 14740 14968 14792 15020
rect 15292 14968 15344 15020
rect 15660 14968 15712 15020
rect 1952 14764 2004 14816
rect 4344 14832 4396 14884
rect 3792 14764 3844 14816
rect 4712 14764 4764 14816
rect 5080 14764 5132 14816
rect 12348 14900 12400 14952
rect 7472 14875 7524 14884
rect 7472 14841 7481 14875
rect 7481 14841 7515 14875
rect 7515 14841 7524 14875
rect 8760 14875 8812 14884
rect 7472 14832 7524 14841
rect 8760 14841 8769 14875
rect 8769 14841 8803 14875
rect 8803 14841 8812 14875
rect 8760 14832 8812 14841
rect 6460 14764 6512 14816
rect 10600 14764 10652 14816
rect 11520 14764 11572 14816
rect 13268 14832 13320 14884
rect 14280 14832 14332 14884
rect 16856 14900 16908 14952
rect 18972 14832 19024 14884
rect 15476 14764 15528 14816
rect 16948 14807 17000 14816
rect 16948 14773 16957 14807
rect 16957 14773 16991 14807
rect 16991 14773 17000 14807
rect 16948 14764 17000 14773
rect 17040 14764 17092 14816
rect 8315 14662 8367 14714
rect 8379 14662 8431 14714
rect 8443 14662 8495 14714
rect 8507 14662 8559 14714
rect 15648 14662 15700 14714
rect 15712 14662 15764 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 1952 14560 2004 14612
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 7196 14560 7248 14612
rect 8760 14560 8812 14612
rect 8944 14603 8996 14612
rect 8944 14569 8953 14603
rect 8953 14569 8987 14603
rect 8987 14569 8996 14603
rect 8944 14560 8996 14569
rect 10048 14603 10100 14612
rect 10048 14569 10057 14603
rect 10057 14569 10091 14603
rect 10091 14569 10100 14603
rect 10048 14560 10100 14569
rect 2596 14492 2648 14544
rect 3792 14492 3844 14544
rect 4344 14535 4396 14544
rect 4344 14501 4353 14535
rect 4353 14501 4387 14535
rect 4387 14501 4396 14535
rect 4344 14492 4396 14501
rect 5080 14492 5132 14544
rect 6644 14492 6696 14544
rect 10784 14535 10836 14544
rect 10784 14501 10793 14535
rect 10793 14501 10827 14535
rect 10827 14501 10836 14535
rect 10784 14492 10836 14501
rect 11060 14492 11112 14544
rect 11888 14560 11940 14612
rect 12532 14560 12584 14612
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 13268 14492 13320 14544
rect 15108 14492 15160 14544
rect 16028 14535 16080 14544
rect 16028 14501 16037 14535
rect 16037 14501 16071 14535
rect 16071 14501 16080 14535
rect 16028 14492 16080 14501
rect 6552 14424 6604 14476
rect 8116 14424 8168 14476
rect 4988 14399 5040 14408
rect 4988 14365 4997 14399
rect 4997 14365 5031 14399
rect 5031 14365 5040 14399
rect 4988 14356 5040 14365
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 5172 14288 5224 14340
rect 8668 14288 8720 14340
rect 12348 14288 12400 14340
rect 14556 14424 14608 14476
rect 17316 14424 17368 14476
rect 17776 14424 17828 14476
rect 12716 14399 12768 14408
rect 12716 14365 12725 14399
rect 12725 14365 12759 14399
rect 12759 14365 12768 14399
rect 12716 14356 12768 14365
rect 4160 14220 4212 14272
rect 4436 14220 4488 14272
rect 7748 14263 7800 14272
rect 7748 14229 7757 14263
rect 7757 14229 7791 14263
rect 7791 14229 7800 14263
rect 7748 14220 7800 14229
rect 10508 14220 10560 14272
rect 11704 14220 11756 14272
rect 13636 14263 13688 14272
rect 13636 14229 13645 14263
rect 13645 14229 13679 14263
rect 13679 14229 13688 14263
rect 13636 14220 13688 14229
rect 14740 14220 14792 14272
rect 15016 14263 15068 14272
rect 15016 14229 15025 14263
rect 15025 14229 15059 14263
rect 15059 14229 15068 14263
rect 15016 14220 15068 14229
rect 15200 14220 15252 14272
rect 17132 14220 17184 14272
rect 4648 14118 4700 14170
rect 4712 14118 4764 14170
rect 4776 14118 4828 14170
rect 4840 14118 4892 14170
rect 11982 14118 12034 14170
rect 12046 14118 12098 14170
rect 12110 14118 12162 14170
rect 12174 14118 12226 14170
rect 19315 14118 19367 14170
rect 19379 14118 19431 14170
rect 19443 14118 19495 14170
rect 19507 14118 19559 14170
rect 1400 14016 1452 14068
rect 4436 14016 4488 14068
rect 5080 14016 5132 14068
rect 7196 14059 7248 14068
rect 7196 14025 7205 14059
rect 7205 14025 7239 14059
rect 7239 14025 7248 14059
rect 7196 14016 7248 14025
rect 8116 14016 8168 14068
rect 15016 14016 15068 14068
rect 15292 14016 15344 14068
rect 2412 13948 2464 14000
rect 2964 13948 3016 14000
rect 4988 13948 5040 14000
rect 10692 13948 10744 14000
rect 17132 13948 17184 14000
rect 7748 13880 7800 13932
rect 8024 13923 8076 13932
rect 8024 13889 8033 13923
rect 8033 13889 8067 13923
rect 8067 13889 8076 13923
rect 8024 13880 8076 13889
rect 9496 13923 9548 13932
rect 9496 13889 9505 13923
rect 9505 13889 9539 13923
rect 9539 13889 9548 13923
rect 9496 13880 9548 13889
rect 10784 13923 10836 13932
rect 2504 13787 2556 13796
rect 2504 13753 2513 13787
rect 2513 13753 2547 13787
rect 2547 13753 2556 13787
rect 2504 13744 2556 13753
rect 2596 13787 2648 13796
rect 2596 13753 2605 13787
rect 2605 13753 2639 13787
rect 2639 13753 2648 13787
rect 2596 13744 2648 13753
rect 4344 13787 4396 13796
rect 4344 13753 4353 13787
rect 4353 13753 4387 13787
rect 4387 13753 4396 13787
rect 4344 13744 4396 13753
rect 4436 13744 4488 13796
rect 8116 13812 8168 13864
rect 10140 13812 10192 13864
rect 10784 13889 10793 13923
rect 10793 13889 10827 13923
rect 10827 13889 10836 13923
rect 12532 13923 12584 13932
rect 10784 13880 10836 13889
rect 10876 13812 10928 13864
rect 6644 13719 6696 13728
rect 6644 13685 6653 13719
rect 6653 13685 6687 13719
rect 6687 13685 6696 13719
rect 6644 13676 6696 13685
rect 7196 13744 7248 13796
rect 9680 13744 9732 13796
rect 12532 13889 12541 13923
rect 12541 13889 12575 13923
rect 12575 13889 12584 13923
rect 12532 13880 12584 13889
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 14280 13880 14332 13932
rect 14924 13812 14976 13864
rect 15476 13855 15528 13864
rect 13176 13744 13228 13796
rect 13728 13744 13780 13796
rect 14188 13787 14240 13796
rect 8852 13676 8904 13728
rect 9496 13676 9548 13728
rect 11244 13676 11296 13728
rect 11612 13676 11664 13728
rect 12808 13676 12860 13728
rect 13636 13676 13688 13728
rect 14188 13753 14197 13787
rect 14197 13753 14231 13787
rect 14231 13753 14240 13787
rect 14188 13744 14240 13753
rect 14740 13787 14792 13796
rect 14740 13753 14749 13787
rect 14749 13753 14783 13787
rect 14783 13753 14792 13787
rect 14740 13744 14792 13753
rect 15476 13821 15485 13855
rect 15485 13821 15519 13855
rect 15519 13821 15528 13855
rect 15476 13812 15528 13821
rect 15752 13812 15804 13864
rect 17132 13812 17184 13864
rect 19099 13855 19151 13864
rect 19099 13821 19108 13855
rect 19108 13821 19142 13855
rect 19142 13821 19151 13855
rect 19099 13812 19151 13821
rect 14648 13676 14700 13728
rect 14924 13676 14976 13728
rect 17408 13744 17460 13796
rect 17776 13787 17828 13796
rect 17776 13753 17785 13787
rect 17785 13753 17819 13787
rect 17819 13753 17828 13787
rect 17776 13744 17828 13753
rect 17316 13676 17368 13728
rect 19064 13676 19116 13728
rect 8315 13574 8367 13626
rect 8379 13574 8431 13626
rect 8443 13574 8495 13626
rect 8507 13574 8559 13626
rect 15648 13574 15700 13626
rect 15712 13574 15764 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 2504 13472 2556 13524
rect 6552 13515 6604 13524
rect 6552 13481 6561 13515
rect 6561 13481 6595 13515
rect 6595 13481 6604 13515
rect 6552 13472 6604 13481
rect 9312 13472 9364 13524
rect 11520 13472 11572 13524
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 12716 13515 12768 13524
rect 12716 13481 12725 13515
rect 12725 13481 12759 13515
rect 12759 13481 12768 13515
rect 12716 13472 12768 13481
rect 14648 13472 14700 13524
rect 1860 13404 1912 13456
rect 4344 13404 4396 13456
rect 5356 13447 5408 13456
rect 5356 13413 5365 13447
rect 5365 13413 5399 13447
rect 5399 13413 5408 13447
rect 5356 13404 5408 13413
rect 6000 13404 6052 13456
rect 6828 13447 6880 13456
rect 6828 13413 6837 13447
rect 6837 13413 6871 13447
rect 6871 13413 6880 13447
rect 6828 13404 6880 13413
rect 7288 13447 7340 13456
rect 7288 13413 7297 13447
rect 7297 13413 7331 13447
rect 7331 13413 7340 13447
rect 7288 13404 7340 13413
rect 10876 13447 10928 13456
rect 10876 13413 10885 13447
rect 10885 13413 10919 13447
rect 10919 13413 10928 13447
rect 10876 13404 10928 13413
rect 13728 13404 13780 13456
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 9588 13379 9640 13388
rect 9588 13345 9597 13379
rect 9597 13345 9631 13379
rect 9631 13345 9640 13379
rect 9588 13336 9640 13345
rect 18144 13472 18196 13524
rect 15108 13447 15160 13456
rect 15108 13413 15117 13447
rect 15117 13413 15151 13447
rect 15151 13413 15160 13447
rect 15108 13404 15160 13413
rect 15476 13447 15528 13456
rect 15476 13413 15485 13447
rect 15485 13413 15519 13447
rect 15519 13413 15528 13447
rect 15476 13404 15528 13413
rect 17224 13336 17276 13388
rect 17408 13379 17460 13388
rect 17408 13345 17417 13379
rect 17417 13345 17451 13379
rect 17451 13345 17460 13379
rect 17408 13336 17460 13345
rect 18788 13336 18840 13388
rect 19616 13336 19668 13388
rect 1768 13268 1820 13320
rect 5540 13268 5592 13320
rect 8116 13268 8168 13320
rect 11060 13311 11112 13320
rect 2228 13200 2280 13252
rect 8024 13200 8076 13252
rect 8760 13200 8812 13252
rect 11060 13277 11069 13311
rect 11069 13277 11103 13311
rect 11103 13277 11112 13311
rect 11060 13268 11112 13277
rect 12900 13311 12952 13320
rect 12900 13277 12909 13311
rect 12909 13277 12943 13311
rect 12943 13277 12952 13311
rect 12900 13268 12952 13277
rect 14648 13268 14700 13320
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 11428 13200 11480 13252
rect 14280 13200 14332 13252
rect 4068 13132 4120 13184
rect 6552 13132 6604 13184
rect 13820 13175 13872 13184
rect 13820 13141 13829 13175
rect 13829 13141 13863 13175
rect 13863 13141 13872 13175
rect 13820 13132 13872 13141
rect 14096 13132 14148 13184
rect 17040 13132 17092 13184
rect 17500 13132 17552 13184
rect 4648 13030 4700 13082
rect 4712 13030 4764 13082
rect 4776 13030 4828 13082
rect 4840 13030 4892 13082
rect 11982 13030 12034 13082
rect 12046 13030 12098 13082
rect 12110 13030 12162 13082
rect 12174 13030 12226 13082
rect 19315 13030 19367 13082
rect 19379 13030 19431 13082
rect 19443 13030 19495 13082
rect 19507 13030 19559 13082
rect 4344 12928 4396 12980
rect 5172 12928 5224 12980
rect 7288 12928 7340 12980
rect 8116 12971 8168 12980
rect 8116 12937 8125 12971
rect 8125 12937 8159 12971
rect 8159 12937 8168 12971
rect 8116 12928 8168 12937
rect 10876 12971 10928 12980
rect 10876 12937 10885 12971
rect 10885 12937 10919 12971
rect 10919 12937 10928 12971
rect 10876 12928 10928 12937
rect 12900 12928 12952 12980
rect 13820 12928 13872 12980
rect 14188 12928 14240 12980
rect 15476 12928 15528 12980
rect 18696 12928 18748 12980
rect 19616 12971 19668 12980
rect 19616 12937 19625 12971
rect 19625 12937 19659 12971
rect 19659 12937 19668 12971
rect 19616 12928 19668 12937
rect 5540 12903 5592 12912
rect 5540 12869 5549 12903
rect 5549 12869 5583 12903
rect 5583 12869 5592 12903
rect 5540 12860 5592 12869
rect 6460 12860 6512 12912
rect 9588 12860 9640 12912
rect 11888 12860 11940 12912
rect 12440 12860 12492 12912
rect 1492 12792 1544 12844
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 6828 12792 6880 12801
rect 14832 12860 14884 12912
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 16396 12792 16448 12844
rect 17408 12792 17460 12844
rect 18604 12792 18656 12844
rect 4068 12724 4120 12776
rect 6092 12767 6144 12776
rect 6092 12733 6101 12767
rect 6101 12733 6135 12767
rect 6135 12733 6144 12767
rect 6092 12724 6144 12733
rect 9404 12724 9456 12776
rect 11244 12724 11296 12776
rect 17132 12724 17184 12776
rect 17684 12724 17736 12776
rect 2228 12699 2280 12708
rect 2228 12665 2237 12699
rect 2237 12665 2271 12699
rect 2271 12665 2280 12699
rect 2780 12699 2832 12708
rect 2228 12656 2280 12665
rect 2780 12665 2789 12699
rect 2789 12665 2823 12699
rect 2823 12665 2832 12699
rect 2780 12656 2832 12665
rect 3792 12699 3844 12708
rect 3792 12665 3801 12699
rect 3801 12665 3835 12699
rect 3835 12665 3844 12699
rect 3792 12656 3844 12665
rect 6644 12699 6696 12708
rect 6644 12665 6653 12699
rect 6653 12665 6687 12699
rect 6687 12665 6696 12699
rect 6644 12656 6696 12665
rect 12624 12699 12676 12708
rect 12624 12665 12633 12699
rect 12633 12665 12667 12699
rect 12667 12665 12676 12699
rect 12624 12656 12676 12665
rect 14188 12699 14240 12708
rect 14188 12665 14197 12699
rect 14197 12665 14231 12699
rect 14231 12665 14240 12699
rect 14188 12656 14240 12665
rect 1860 12588 1912 12640
rect 2964 12588 3016 12640
rect 9680 12631 9732 12640
rect 9680 12597 9689 12631
rect 9689 12597 9723 12631
rect 9723 12597 9732 12631
rect 9680 12588 9732 12597
rect 10324 12588 10376 12640
rect 13452 12588 13504 12640
rect 13728 12588 13780 12640
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 16120 12656 16172 12708
rect 18972 12724 19024 12776
rect 18512 12699 18564 12708
rect 18512 12665 18521 12699
rect 18521 12665 18555 12699
rect 18555 12665 18564 12699
rect 18512 12656 18564 12665
rect 17224 12631 17276 12640
rect 15476 12588 15528 12597
rect 17224 12597 17233 12631
rect 17233 12597 17267 12631
rect 17267 12597 17276 12631
rect 17224 12588 17276 12597
rect 17408 12588 17460 12640
rect 18788 12588 18840 12640
rect 18972 12588 19024 12640
rect 19892 12631 19944 12640
rect 19892 12597 19901 12631
rect 19901 12597 19935 12631
rect 19935 12597 19944 12631
rect 19892 12588 19944 12597
rect 8315 12486 8367 12538
rect 8379 12486 8431 12538
rect 8443 12486 8495 12538
rect 8507 12486 8559 12538
rect 15648 12486 15700 12538
rect 15712 12486 15764 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 1860 12427 1912 12436
rect 1860 12393 1869 12427
rect 1869 12393 1903 12427
rect 1903 12393 1912 12427
rect 1860 12384 1912 12393
rect 2228 12384 2280 12436
rect 2964 12384 3016 12436
rect 3792 12384 3844 12436
rect 4068 12384 4120 12436
rect 6644 12427 6696 12436
rect 6644 12393 6653 12427
rect 6653 12393 6687 12427
rect 6687 12393 6696 12427
rect 6644 12384 6696 12393
rect 7288 12384 7340 12436
rect 10876 12384 10928 12436
rect 12624 12384 12676 12436
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 4160 12248 4212 12300
rect 6000 12248 6052 12300
rect 6736 12248 6788 12300
rect 8116 12316 8168 12368
rect 8760 12359 8812 12368
rect 8760 12325 8769 12359
rect 8769 12325 8803 12359
rect 8803 12325 8812 12359
rect 8760 12316 8812 12325
rect 9680 12316 9732 12368
rect 11152 12316 11204 12368
rect 11428 12359 11480 12368
rect 11428 12325 11437 12359
rect 11437 12325 11471 12359
rect 11471 12325 11480 12359
rect 11428 12316 11480 12325
rect 11888 12291 11940 12300
rect 11888 12257 11897 12291
rect 11897 12257 11931 12291
rect 11931 12257 11940 12291
rect 11888 12248 11940 12257
rect 13728 12316 13780 12368
rect 15476 12359 15528 12368
rect 15476 12325 15485 12359
rect 15485 12325 15519 12359
rect 15519 12325 15528 12359
rect 15476 12316 15528 12325
rect 16028 12359 16080 12368
rect 16028 12325 16037 12359
rect 16037 12325 16071 12359
rect 16071 12325 16080 12359
rect 16028 12316 16080 12325
rect 16396 12359 16448 12368
rect 16396 12325 16405 12359
rect 16405 12325 16439 12359
rect 16439 12325 16448 12359
rect 16396 12316 16448 12325
rect 17408 12316 17460 12368
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 17224 12248 17276 12300
rect 18420 12291 18472 12300
rect 18420 12257 18429 12291
rect 18429 12257 18463 12291
rect 18463 12257 18472 12291
rect 18420 12248 18472 12257
rect 18604 12248 18656 12300
rect 2136 12180 2188 12232
rect 8208 12180 8260 12232
rect 11244 12180 11296 12232
rect 13452 12180 13504 12232
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 7196 12112 7248 12164
rect 10968 12112 11020 12164
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17408 12180 17460 12189
rect 2872 12044 2924 12096
rect 4528 12044 4580 12096
rect 9404 12087 9456 12096
rect 9404 12053 9413 12087
rect 9413 12053 9447 12087
rect 9447 12053 9456 12087
rect 9404 12044 9456 12053
rect 13728 12044 13780 12096
rect 14832 12044 14884 12096
rect 18788 12044 18840 12096
rect 4648 11942 4700 11994
rect 4712 11942 4764 11994
rect 4776 11942 4828 11994
rect 4840 11942 4892 11994
rect 11982 11942 12034 11994
rect 12046 11942 12098 11994
rect 12110 11942 12162 11994
rect 12174 11942 12226 11994
rect 19315 11942 19367 11994
rect 19379 11942 19431 11994
rect 19443 11942 19495 11994
rect 19507 11942 19559 11994
rect 4160 11883 4212 11892
rect 4160 11849 4169 11883
rect 4169 11849 4203 11883
rect 4203 11849 4212 11883
rect 6000 11883 6052 11892
rect 4160 11840 4212 11849
rect 6000 11849 6009 11883
rect 6009 11849 6043 11883
rect 6043 11849 6052 11883
rect 6000 11840 6052 11849
rect 6644 11840 6696 11892
rect 8116 11883 8168 11892
rect 8116 11849 8125 11883
rect 8125 11849 8159 11883
rect 8159 11849 8168 11883
rect 8116 11840 8168 11849
rect 8208 11840 8260 11892
rect 9772 11840 9824 11892
rect 15292 11840 15344 11892
rect 15476 11840 15528 11892
rect 17868 11840 17920 11892
rect 18604 11883 18656 11892
rect 18604 11849 18613 11883
rect 18613 11849 18647 11883
rect 18647 11849 18656 11883
rect 18604 11840 18656 11849
rect 20076 11840 20128 11892
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 7196 11747 7248 11756
rect 7196 11713 7205 11747
rect 7205 11713 7239 11747
rect 7239 11713 7248 11747
rect 7196 11704 7248 11713
rect 7840 11747 7892 11756
rect 7840 11713 7849 11747
rect 7849 11713 7883 11747
rect 7883 11713 7892 11747
rect 7840 11704 7892 11713
rect 11152 11772 11204 11824
rect 11244 11815 11296 11824
rect 11244 11781 11253 11815
rect 11253 11781 11287 11815
rect 11287 11781 11296 11815
rect 11244 11772 11296 11781
rect 17408 11772 17460 11824
rect 11060 11704 11112 11756
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 2872 11636 2924 11688
rect 8208 11636 8260 11688
rect 9496 11636 9548 11688
rect 12348 11636 12400 11688
rect 15292 11704 15344 11756
rect 15384 11704 15436 11756
rect 13452 11679 13504 11688
rect 13452 11645 13461 11679
rect 13461 11645 13495 11679
rect 13495 11645 13504 11679
rect 13452 11636 13504 11645
rect 4528 11611 4580 11620
rect 4528 11577 4537 11611
rect 4537 11577 4571 11611
rect 4571 11577 4580 11611
rect 4528 11568 4580 11577
rect 20 11500 72 11552
rect 2504 11500 2556 11552
rect 2964 11500 3016 11552
rect 7288 11611 7340 11620
rect 7288 11577 7297 11611
rect 7297 11577 7331 11611
rect 7331 11577 7340 11611
rect 7288 11568 7340 11577
rect 10324 11611 10376 11620
rect 10324 11577 10333 11611
rect 10333 11577 10367 11611
rect 10367 11577 10376 11611
rect 10324 11568 10376 11577
rect 10508 11568 10560 11620
rect 15200 11679 15252 11688
rect 15200 11645 15209 11679
rect 15209 11645 15243 11679
rect 15243 11645 15252 11679
rect 15200 11636 15252 11645
rect 6368 11500 6420 11552
rect 9680 11500 9732 11552
rect 10600 11500 10652 11552
rect 13728 11568 13780 11620
rect 13268 11543 13320 11552
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 16028 11568 16080 11620
rect 17040 11636 17092 11688
rect 17224 11636 17276 11688
rect 18512 11636 18564 11688
rect 17132 11568 17184 11620
rect 18236 11568 18288 11620
rect 14372 11543 14424 11552
rect 13268 11500 13320 11509
rect 14372 11509 14381 11543
rect 14381 11509 14415 11543
rect 14415 11509 14424 11543
rect 14372 11500 14424 11509
rect 14648 11543 14700 11552
rect 14648 11509 14657 11543
rect 14657 11509 14691 11543
rect 14691 11509 14700 11543
rect 14648 11500 14700 11509
rect 15108 11500 15160 11552
rect 18052 11500 18104 11552
rect 18420 11500 18472 11552
rect 8315 11398 8367 11450
rect 8379 11398 8431 11450
rect 8443 11398 8495 11450
rect 8507 11398 8559 11450
rect 15648 11398 15700 11450
rect 15712 11398 15764 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 4068 11296 4120 11348
rect 5080 11339 5132 11348
rect 5080 11305 5089 11339
rect 5089 11305 5123 11339
rect 5123 11305 5132 11339
rect 5080 11296 5132 11305
rect 7288 11296 7340 11348
rect 7840 11296 7892 11348
rect 2504 11228 2556 11280
rect 6644 11271 6696 11280
rect 5356 11160 5408 11212
rect 6644 11237 6653 11271
rect 6653 11237 6687 11271
rect 6687 11237 6696 11271
rect 6644 11228 6696 11237
rect 8116 11228 8168 11280
rect 10324 11296 10376 11348
rect 10416 11271 10468 11280
rect 10416 11237 10425 11271
rect 10425 11237 10459 11271
rect 10459 11237 10468 11271
rect 10416 11228 10468 11237
rect 12808 11296 12860 11348
rect 13452 11296 13504 11348
rect 11796 11228 11848 11280
rect 13268 11228 13320 11280
rect 14372 11228 14424 11280
rect 15016 11228 15068 11280
rect 16120 11160 16172 11212
rect 16488 11160 16540 11212
rect 17316 11203 17368 11212
rect 17316 11169 17325 11203
rect 17325 11169 17359 11203
rect 17359 11169 17368 11203
rect 17316 11160 17368 11169
rect 1676 10956 1728 11008
rect 2320 11092 2372 11144
rect 2780 11092 2832 11144
rect 2136 11024 2188 11076
rect 4068 11092 4120 11144
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 8760 11092 8812 11144
rect 12440 11092 12492 11144
rect 13452 11135 13504 11144
rect 4988 11024 5040 11076
rect 2964 10999 3016 11008
rect 2964 10965 2973 10999
rect 2973 10965 3007 10999
rect 3007 10965 3016 10999
rect 2964 10956 3016 10965
rect 6920 11024 6972 11076
rect 11520 11024 11572 11076
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 14464 11024 14516 11076
rect 15292 11024 15344 11076
rect 19156 11024 19208 11076
rect 5908 10999 5960 11008
rect 5908 10965 5917 10999
rect 5917 10965 5951 10999
rect 5951 10965 5960 10999
rect 5908 10956 5960 10965
rect 13360 10999 13412 11008
rect 13360 10965 13369 10999
rect 13369 10965 13403 10999
rect 13403 10965 13412 10999
rect 13360 10956 13412 10965
rect 14372 10999 14424 11008
rect 14372 10965 14381 10999
rect 14381 10965 14415 10999
rect 14415 10965 14424 10999
rect 14372 10956 14424 10965
rect 15200 10956 15252 11008
rect 20444 10956 20496 11008
rect 4648 10854 4700 10906
rect 4712 10854 4764 10906
rect 4776 10854 4828 10906
rect 4840 10854 4892 10906
rect 11982 10854 12034 10906
rect 12046 10854 12098 10906
rect 12110 10854 12162 10906
rect 12174 10854 12226 10906
rect 19315 10854 19367 10906
rect 19379 10854 19431 10906
rect 19443 10854 19495 10906
rect 19507 10854 19559 10906
rect 2504 10752 2556 10804
rect 5632 10752 5684 10804
rect 6644 10752 6696 10804
rect 8116 10752 8168 10804
rect 10324 10795 10376 10804
rect 10324 10761 10333 10795
rect 10333 10761 10367 10795
rect 10367 10761 10376 10795
rect 10324 10752 10376 10761
rect 11796 10752 11848 10804
rect 15384 10752 15436 10804
rect 19156 10795 19208 10804
rect 19156 10761 19165 10795
rect 19165 10761 19199 10795
rect 19199 10761 19208 10795
rect 19156 10752 19208 10761
rect 19800 10752 19852 10804
rect 8852 10684 8904 10736
rect 13452 10684 13504 10736
rect 16948 10684 17000 10736
rect 5908 10616 5960 10668
rect 7288 10616 7340 10668
rect 9864 10616 9916 10668
rect 11796 10616 11848 10668
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 16304 10616 16356 10668
rect 17316 10616 17368 10668
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 9036 10548 9088 10600
rect 17132 10591 17184 10600
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 17960 10548 18012 10600
rect 2688 10523 2740 10532
rect 2688 10489 2697 10523
rect 2697 10489 2731 10523
rect 2731 10489 2740 10523
rect 2688 10480 2740 10489
rect 112 10412 164 10464
rect 2596 10412 2648 10464
rect 4344 10480 4396 10532
rect 5356 10523 5408 10532
rect 5356 10489 5365 10523
rect 5365 10489 5399 10523
rect 5399 10489 5408 10523
rect 5356 10480 5408 10489
rect 5908 10523 5960 10532
rect 5908 10489 5917 10523
rect 5917 10489 5951 10523
rect 5951 10489 5960 10523
rect 5908 10480 5960 10489
rect 4252 10412 4304 10464
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 9680 10480 9732 10532
rect 10784 10523 10836 10532
rect 10784 10489 10793 10523
rect 10793 10489 10827 10523
rect 10827 10489 10836 10523
rect 10784 10480 10836 10489
rect 10876 10523 10928 10532
rect 10876 10489 10885 10523
rect 10885 10489 10919 10523
rect 10919 10489 10928 10523
rect 10876 10480 10928 10489
rect 15200 10523 15252 10532
rect 15200 10489 15209 10523
rect 15209 10489 15243 10523
rect 15243 10489 15252 10523
rect 15200 10480 15252 10489
rect 7932 10455 7984 10464
rect 5080 10412 5132 10421
rect 7932 10421 7941 10455
rect 7941 10421 7975 10455
rect 7975 10421 7984 10455
rect 7932 10412 7984 10421
rect 11612 10412 11664 10464
rect 13268 10455 13320 10464
rect 13268 10421 13277 10455
rect 13277 10421 13311 10455
rect 13311 10421 13320 10455
rect 13268 10412 13320 10421
rect 13452 10412 13504 10464
rect 16028 10480 16080 10532
rect 15476 10412 15528 10464
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 16580 10412 16632 10464
rect 17868 10455 17920 10464
rect 17868 10421 17877 10455
rect 17877 10421 17911 10455
rect 17911 10421 17920 10455
rect 17868 10412 17920 10421
rect 18144 10455 18196 10464
rect 18144 10421 18153 10455
rect 18153 10421 18187 10455
rect 18187 10421 18196 10455
rect 18144 10412 18196 10421
rect 19616 10455 19668 10464
rect 19616 10421 19625 10455
rect 19625 10421 19659 10455
rect 19659 10421 19668 10455
rect 19616 10412 19668 10421
rect 8315 10310 8367 10362
rect 8379 10310 8431 10362
rect 8443 10310 8495 10362
rect 8507 10310 8559 10362
rect 15648 10310 15700 10362
rect 15712 10310 15764 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 1216 10208 1268 10260
rect 2504 10208 2556 10260
rect 2688 10208 2740 10260
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 5356 10208 5408 10260
rect 10416 10208 10468 10260
rect 10876 10251 10928 10260
rect 10876 10217 10885 10251
rect 10885 10217 10919 10251
rect 10919 10217 10928 10251
rect 10876 10208 10928 10217
rect 12440 10251 12492 10260
rect 12440 10217 12449 10251
rect 12449 10217 12483 10251
rect 12483 10217 12492 10251
rect 12440 10208 12492 10217
rect 2596 10183 2648 10192
rect 2596 10149 2605 10183
rect 2605 10149 2639 10183
rect 2639 10149 2648 10183
rect 2596 10140 2648 10149
rect 2964 10140 3016 10192
rect 4988 10140 5040 10192
rect 5816 10183 5868 10192
rect 5816 10149 5825 10183
rect 5825 10149 5859 10183
rect 5859 10149 5868 10183
rect 5816 10140 5868 10149
rect 7932 10140 7984 10192
rect 9864 10140 9916 10192
rect 2320 10072 2372 10124
rect 9588 10072 9640 10124
rect 10784 10140 10836 10192
rect 11612 10183 11664 10192
rect 11612 10149 11621 10183
rect 11621 10149 11655 10183
rect 11655 10149 11664 10183
rect 11612 10140 11664 10149
rect 11796 10140 11848 10192
rect 14832 10208 14884 10260
rect 15016 10251 15068 10260
rect 15016 10217 15025 10251
rect 15025 10217 15059 10251
rect 15059 10217 15068 10251
rect 15016 10208 15068 10217
rect 16948 10251 17000 10260
rect 16948 10217 16957 10251
rect 16957 10217 16991 10251
rect 16991 10217 17000 10251
rect 16948 10208 17000 10217
rect 18512 10251 18564 10260
rect 18512 10217 18521 10251
rect 18521 10217 18555 10251
rect 18555 10217 18564 10251
rect 18512 10208 18564 10217
rect 13820 10183 13872 10192
rect 13820 10149 13829 10183
rect 13829 10149 13863 10183
rect 13863 10149 13872 10183
rect 13820 10140 13872 10149
rect 14372 10140 14424 10192
rect 15108 10140 15160 10192
rect 16028 10183 16080 10192
rect 16028 10149 16037 10183
rect 16037 10149 16071 10183
rect 16071 10149 16080 10183
rect 16028 10140 16080 10149
rect 16120 10140 16172 10192
rect 16672 10072 16724 10124
rect 17316 10115 17368 10124
rect 3332 10004 3384 10056
rect 4252 10004 4304 10056
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 6920 10047 6972 10056
rect 4528 9936 4580 9988
rect 5908 9936 5960 9988
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 8024 10004 8076 10056
rect 9496 10004 9548 10056
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 13544 10004 13596 10056
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 17316 10081 17325 10115
rect 17325 10081 17359 10115
rect 17359 10081 17368 10115
rect 17316 10072 17368 10081
rect 18420 10115 18472 10124
rect 18420 10081 18429 10115
rect 18429 10081 18463 10115
rect 18463 10081 18472 10115
rect 18420 10072 18472 10081
rect 18880 10115 18932 10124
rect 18880 10081 18889 10115
rect 18889 10081 18923 10115
rect 18923 10081 18932 10115
rect 18880 10072 18932 10081
rect 17960 10004 18012 10056
rect 2228 9911 2280 9920
rect 2228 9877 2237 9911
rect 2237 9877 2271 9911
rect 2271 9877 2280 9911
rect 2228 9868 2280 9877
rect 5172 9911 5224 9920
rect 5172 9877 5181 9911
rect 5181 9877 5215 9911
rect 5215 9877 5224 9911
rect 5172 9868 5224 9877
rect 5724 9868 5776 9920
rect 6368 9868 6420 9920
rect 7288 9911 7340 9920
rect 7288 9877 7297 9911
rect 7297 9877 7331 9911
rect 7331 9877 7340 9911
rect 7288 9868 7340 9877
rect 9036 9911 9088 9920
rect 9036 9877 9045 9911
rect 9045 9877 9079 9911
rect 9079 9877 9088 9911
rect 9036 9868 9088 9877
rect 13452 9911 13504 9920
rect 13452 9877 13461 9911
rect 13461 9877 13495 9911
rect 13495 9877 13504 9911
rect 13452 9868 13504 9877
rect 14740 9911 14792 9920
rect 14740 9877 14749 9911
rect 14749 9877 14783 9911
rect 14783 9877 14792 9911
rect 14740 9868 14792 9877
rect 4648 9766 4700 9818
rect 4712 9766 4764 9818
rect 4776 9766 4828 9818
rect 4840 9766 4892 9818
rect 11982 9766 12034 9818
rect 12046 9766 12098 9818
rect 12110 9766 12162 9818
rect 12174 9766 12226 9818
rect 19315 9766 19367 9818
rect 19379 9766 19431 9818
rect 19443 9766 19495 9818
rect 19507 9766 19559 9818
rect 2596 9707 2648 9716
rect 2596 9673 2605 9707
rect 2605 9673 2639 9707
rect 2639 9673 2648 9707
rect 2596 9664 2648 9673
rect 2964 9664 3016 9716
rect 5816 9707 5868 9716
rect 5816 9673 5825 9707
rect 5825 9673 5859 9707
rect 5859 9673 5868 9707
rect 5816 9664 5868 9673
rect 6368 9664 6420 9716
rect 204 9596 256 9648
rect 4160 9596 4212 9648
rect 8116 9664 8168 9716
rect 8668 9664 8720 9716
rect 11612 9707 11664 9716
rect 11612 9673 11621 9707
rect 11621 9673 11655 9707
rect 11655 9673 11664 9707
rect 11612 9664 11664 9673
rect 13820 9707 13872 9716
rect 13820 9673 13829 9707
rect 13829 9673 13863 9707
rect 13863 9673 13872 9707
rect 13820 9664 13872 9673
rect 14832 9664 14884 9716
rect 17316 9707 17368 9716
rect 17316 9673 17325 9707
rect 17325 9673 17359 9707
rect 17359 9673 17368 9707
rect 17316 9664 17368 9673
rect 9680 9639 9732 9648
rect 9680 9605 9689 9639
rect 9689 9605 9723 9639
rect 9723 9605 9732 9639
rect 9680 9596 9732 9605
rect 11704 9596 11756 9648
rect 14924 9596 14976 9648
rect 15200 9596 15252 9648
rect 1492 9460 1544 9512
rect 2228 9460 2280 9512
rect 2412 9392 2464 9444
rect 8024 9528 8076 9580
rect 8668 9528 8720 9580
rect 9220 9528 9272 9580
rect 6736 9460 6788 9512
rect 6920 9460 6972 9512
rect 7380 9503 7432 9512
rect 7380 9469 7389 9503
rect 7389 9469 7423 9503
rect 7423 9469 7432 9503
rect 7380 9460 7432 9469
rect 11520 9528 11572 9580
rect 14740 9571 14792 9580
rect 14740 9537 14749 9571
rect 14749 9537 14783 9571
rect 14783 9537 14792 9571
rect 14740 9528 14792 9537
rect 10876 9460 10928 9512
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 16212 9503 16264 9512
rect 5080 9392 5132 9444
rect 5172 9392 5224 9444
rect 5356 9324 5408 9376
rect 5448 9324 5500 9376
rect 6092 9324 6144 9376
rect 9680 9392 9732 9444
rect 12716 9435 12768 9444
rect 12716 9401 12725 9435
rect 12725 9401 12759 9435
rect 12759 9401 12768 9435
rect 12716 9392 12768 9401
rect 13452 9392 13504 9444
rect 14832 9435 14884 9444
rect 14832 9401 14841 9435
rect 14841 9401 14875 9435
rect 14875 9401 14884 9435
rect 14832 9392 14884 9401
rect 9588 9324 9640 9376
rect 14556 9324 14608 9376
rect 16212 9469 16221 9503
rect 16221 9469 16255 9503
rect 16255 9469 16264 9503
rect 16212 9460 16264 9469
rect 16120 9435 16172 9444
rect 16120 9401 16129 9435
rect 16129 9401 16163 9435
rect 16163 9401 16172 9435
rect 17316 9460 17368 9512
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 16120 9392 16172 9401
rect 16304 9367 16356 9376
rect 16304 9333 16313 9367
rect 16313 9333 16347 9367
rect 16347 9333 16356 9367
rect 16304 9324 16356 9333
rect 17316 9324 17368 9376
rect 17868 9392 17920 9444
rect 18604 9460 18656 9512
rect 19892 9460 19944 9512
rect 18880 9392 18932 9444
rect 18144 9367 18196 9376
rect 18144 9333 18153 9367
rect 18153 9333 18187 9367
rect 18187 9333 18196 9367
rect 18144 9324 18196 9333
rect 8315 9222 8367 9274
rect 8379 9222 8431 9274
rect 8443 9222 8495 9274
rect 8507 9222 8559 9274
rect 15648 9222 15700 9274
rect 15712 9222 15764 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 3056 9120 3108 9172
rect 3240 9120 3292 9172
rect 4160 9120 4212 9172
rect 4252 9120 4304 9172
rect 6828 9163 6880 9172
rect 4528 9052 4580 9104
rect 5448 9095 5500 9104
rect 5448 9061 5457 9095
rect 5457 9061 5491 9095
rect 5491 9061 5500 9095
rect 5448 9052 5500 9061
rect 5816 9052 5868 9104
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 7932 9163 7984 9172
rect 7932 9129 7941 9163
rect 7941 9129 7975 9163
rect 7975 9129 7984 9163
rect 7932 9120 7984 9129
rect 8668 9120 8720 9172
rect 12900 9163 12952 9172
rect 6644 9052 6696 9104
rect 9588 9052 9640 9104
rect 10784 9052 10836 9104
rect 11336 9095 11388 9104
rect 11336 9061 11345 9095
rect 11345 9061 11379 9095
rect 11379 9061 11388 9095
rect 11336 9052 11388 9061
rect 11704 9052 11756 9104
rect 12900 9129 12909 9163
rect 12909 9129 12943 9163
rect 12943 9129 12952 9163
rect 12900 9120 12952 9129
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 18420 9120 18472 9172
rect 13544 9095 13596 9104
rect 13544 9061 13553 9095
rect 13553 9061 13587 9095
rect 13587 9061 13596 9095
rect 13544 9052 13596 9061
rect 13820 9095 13872 9104
rect 13820 9061 13829 9095
rect 13829 9061 13863 9095
rect 13863 9061 13872 9095
rect 13820 9052 13872 9061
rect 14372 9095 14424 9104
rect 14372 9061 14381 9095
rect 14381 9061 14415 9095
rect 14415 9061 14424 9095
rect 14372 9052 14424 9061
rect 15108 9095 15160 9104
rect 15108 9061 15117 9095
rect 15117 9061 15151 9095
rect 15151 9061 15160 9095
rect 15108 9052 15160 9061
rect 18052 9095 18104 9104
rect 1308 8984 1360 9036
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 2044 8984 2096 9036
rect 2780 8984 2832 9036
rect 3332 8984 3384 9036
rect 4344 9027 4396 9036
rect 4344 8993 4388 9027
rect 4388 8993 4396 9027
rect 4344 8984 4396 8993
rect 8852 8984 8904 9036
rect 9496 9027 9548 9036
rect 9496 8993 9505 9027
rect 9505 8993 9539 9027
rect 9539 8993 9548 9027
rect 9496 8984 9548 8993
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 9772 8959 9824 8968
rect 9772 8925 9781 8959
rect 9781 8925 9815 8959
rect 9815 8925 9824 8959
rect 9772 8916 9824 8925
rect 10876 8916 10928 8968
rect 14464 8984 14516 9036
rect 18052 9061 18061 9095
rect 18061 9061 18095 9095
rect 18095 9061 18104 9095
rect 18052 9052 18104 9061
rect 15660 8984 15712 9036
rect 16120 8984 16172 9036
rect 16212 8984 16264 9036
rect 16764 8984 16816 9036
rect 17316 9027 17368 9036
rect 17316 8993 17325 9027
rect 17325 8993 17359 9027
rect 17359 8993 17368 9027
rect 17316 8984 17368 8993
rect 17684 8984 17736 9036
rect 18880 8984 18932 9036
rect 19156 8984 19208 9036
rect 7564 8891 7616 8900
rect 7564 8857 7573 8891
rect 7573 8857 7607 8891
rect 7607 8857 7616 8891
rect 7564 8848 7616 8857
rect 2964 8780 3016 8832
rect 3884 8823 3936 8832
rect 3884 8789 3893 8823
rect 3893 8789 3927 8823
rect 3927 8789 3936 8823
rect 3884 8780 3936 8789
rect 4528 8780 4580 8832
rect 5448 8780 5500 8832
rect 6920 8780 6972 8832
rect 8944 8780 8996 8832
rect 10692 8780 10744 8832
rect 16488 8916 16540 8968
rect 14280 8848 14332 8900
rect 15936 8848 15988 8900
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 16580 8780 16632 8832
rect 16856 8780 16908 8832
rect 18972 8780 19024 8832
rect 4648 8678 4700 8730
rect 4712 8678 4764 8730
rect 4776 8678 4828 8730
rect 4840 8678 4892 8730
rect 11982 8678 12034 8730
rect 12046 8678 12098 8730
rect 12110 8678 12162 8730
rect 12174 8678 12226 8730
rect 19315 8678 19367 8730
rect 19379 8678 19431 8730
rect 19443 8678 19495 8730
rect 19507 8678 19559 8730
rect 2780 8619 2832 8628
rect 2780 8585 2789 8619
rect 2789 8585 2823 8619
rect 2823 8585 2832 8619
rect 2780 8576 2832 8585
rect 5816 8576 5868 8628
rect 7380 8576 7432 8628
rect 8852 8576 8904 8628
rect 9588 8619 9640 8628
rect 9588 8585 9597 8619
rect 9597 8585 9631 8619
rect 9631 8585 9640 8619
rect 9588 8576 9640 8585
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 12716 8619 12768 8628
rect 12716 8585 12725 8619
rect 12725 8585 12759 8619
rect 12759 8585 12768 8619
rect 12716 8576 12768 8585
rect 13820 8576 13872 8628
rect 14740 8576 14792 8628
rect 4344 8508 4396 8560
rect 8208 8508 8260 8560
rect 13544 8508 13596 8560
rect 18972 8508 19024 8560
rect 2504 8440 2556 8492
rect 3424 8440 3476 8492
rect 1860 8372 1912 8424
rect 3240 8415 3292 8424
rect 2136 8347 2188 8356
rect 2136 8313 2145 8347
rect 2145 8313 2179 8347
rect 2179 8313 2188 8347
rect 2136 8304 2188 8313
rect 3240 8381 3249 8415
rect 3249 8381 3283 8415
rect 3283 8381 3292 8415
rect 3240 8372 3292 8381
rect 3700 8304 3752 8356
rect 4344 8372 4396 8424
rect 4528 8415 4580 8424
rect 4528 8381 4537 8415
rect 4537 8381 4571 8415
rect 4571 8381 4580 8415
rect 4528 8372 4580 8381
rect 6276 8440 6328 8492
rect 7656 8440 7708 8492
rect 10784 8440 10836 8492
rect 14648 8440 14700 8492
rect 14924 8483 14976 8492
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 15660 8483 15712 8492
rect 15660 8449 15669 8483
rect 15669 8449 15703 8483
rect 15703 8449 15712 8483
rect 15660 8440 15712 8449
rect 15936 8440 15988 8492
rect 16212 8440 16264 8492
rect 16948 8440 17000 8492
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 2504 8279 2556 8288
rect 2504 8245 2513 8279
rect 2513 8245 2547 8279
rect 2547 8245 2556 8279
rect 2504 8236 2556 8245
rect 2872 8236 2924 8288
rect 4068 8236 4120 8288
rect 6644 8279 6696 8288
rect 6644 8245 6653 8279
rect 6653 8245 6687 8279
rect 6687 8245 6696 8279
rect 6644 8236 6696 8245
rect 7196 8304 7248 8356
rect 9680 8304 9732 8356
rect 10784 8347 10836 8356
rect 10784 8313 10793 8347
rect 10793 8313 10827 8347
rect 10827 8313 10836 8347
rect 10784 8304 10836 8313
rect 10876 8347 10928 8356
rect 10876 8313 10885 8347
rect 10885 8313 10919 8347
rect 10919 8313 10928 8347
rect 10876 8304 10928 8313
rect 12716 8304 12768 8356
rect 7104 8236 7156 8288
rect 14740 8347 14792 8356
rect 14740 8313 14749 8347
rect 14749 8313 14783 8347
rect 14783 8313 14792 8347
rect 17316 8372 17368 8424
rect 19800 8372 19852 8424
rect 14740 8304 14792 8313
rect 16488 8304 16540 8356
rect 17040 8304 17092 8356
rect 17224 8304 17276 8356
rect 19156 8304 19208 8356
rect 14188 8236 14240 8288
rect 14372 8279 14424 8288
rect 14372 8245 14381 8279
rect 14381 8245 14415 8279
rect 14415 8245 14424 8279
rect 14372 8236 14424 8245
rect 14556 8236 14608 8288
rect 16212 8279 16264 8288
rect 16212 8245 16221 8279
rect 16221 8245 16255 8279
rect 16255 8245 16264 8279
rect 16212 8236 16264 8245
rect 18420 8236 18472 8288
rect 18972 8236 19024 8288
rect 8315 8134 8367 8186
rect 8379 8134 8431 8186
rect 8443 8134 8495 8186
rect 8507 8134 8559 8186
rect 15648 8134 15700 8186
rect 15712 8134 15764 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 2504 8075 2556 8084
rect 2504 8041 2513 8075
rect 2513 8041 2547 8075
rect 2547 8041 2556 8075
rect 3424 8075 3476 8084
rect 2504 8032 2556 8041
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 3516 8032 3568 8084
rect 5908 8075 5960 8084
rect 5908 8041 5917 8075
rect 5917 8041 5951 8075
rect 5951 8041 5960 8075
rect 5908 8032 5960 8041
rect 7012 8032 7064 8084
rect 13820 8032 13872 8084
rect 14740 8032 14792 8084
rect 16856 8032 16908 8084
rect 18236 8032 18288 8084
rect 1308 7964 1360 8016
rect 1676 7896 1728 7948
rect 2504 7896 2556 7948
rect 1768 7828 1820 7880
rect 3884 7964 3936 8016
rect 3148 7896 3200 7948
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 5080 7896 5132 7948
rect 8484 7964 8536 8016
rect 9772 7964 9824 8016
rect 11336 8007 11388 8016
rect 9680 7896 9732 7948
rect 11336 7973 11345 8007
rect 11345 7973 11379 8007
rect 11379 7973 11388 8007
rect 11336 7964 11388 7973
rect 12716 7964 12768 8016
rect 13268 7964 13320 8016
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 13912 7964 13964 8016
rect 16304 7964 16356 8016
rect 16764 8007 16816 8016
rect 16764 7973 16773 8007
rect 16773 7973 16807 8007
rect 16807 7973 16816 8007
rect 16764 7964 16816 7973
rect 17224 7964 17276 8016
rect 14556 7896 14608 7948
rect 16580 7896 16632 7948
rect 16672 7896 16724 7948
rect 4988 7760 5040 7812
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 4436 7692 4488 7744
rect 5448 7828 5500 7880
rect 7564 7828 7616 7880
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 9772 7871 9824 7880
rect 7656 7828 7708 7837
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12716 7828 12768 7837
rect 15200 7828 15252 7880
rect 15476 7828 15528 7880
rect 7196 7760 7248 7812
rect 9128 7760 9180 7812
rect 10876 7760 10928 7812
rect 11336 7760 11388 7812
rect 15292 7760 15344 7812
rect 18880 7828 18932 7880
rect 19156 7760 19208 7812
rect 5172 7692 5224 7744
rect 5264 7692 5316 7744
rect 7656 7692 7708 7744
rect 8484 7692 8536 7744
rect 9036 7735 9088 7744
rect 9036 7701 9045 7735
rect 9045 7701 9079 7735
rect 9079 7701 9088 7735
rect 9036 7692 9088 7701
rect 11520 7692 11572 7744
rect 15016 7692 15068 7744
rect 15568 7692 15620 7744
rect 15752 7692 15804 7744
rect 16488 7692 16540 7744
rect 18420 7692 18472 7744
rect 18788 7692 18840 7744
rect 4648 7590 4700 7642
rect 4712 7590 4764 7642
rect 4776 7590 4828 7642
rect 4840 7590 4892 7642
rect 11982 7590 12034 7642
rect 12046 7590 12098 7642
rect 12110 7590 12162 7642
rect 12174 7590 12226 7642
rect 19315 7590 19367 7642
rect 19379 7590 19431 7642
rect 19443 7590 19495 7642
rect 19507 7590 19559 7642
rect 1676 7531 1728 7540
rect 1676 7497 1685 7531
rect 1685 7497 1719 7531
rect 1719 7497 1728 7531
rect 1676 7488 1728 7497
rect 2044 7488 2096 7540
rect 9036 7488 9088 7540
rect 9680 7531 9732 7540
rect 9680 7497 9689 7531
rect 9689 7497 9723 7531
rect 9723 7497 9732 7531
rect 9680 7488 9732 7497
rect 10232 7488 10284 7540
rect 13268 7531 13320 7540
rect 13268 7497 13277 7531
rect 13277 7497 13311 7531
rect 13311 7497 13320 7531
rect 13268 7488 13320 7497
rect 16304 7531 16356 7540
rect 16304 7497 16313 7531
rect 16313 7497 16347 7531
rect 16347 7497 16356 7531
rect 16304 7488 16356 7497
rect 3148 7420 3200 7472
rect 3792 7420 3844 7472
rect 4068 7420 4120 7472
rect 5080 7463 5132 7472
rect 2136 7284 2188 7336
rect 3884 7284 3936 7336
rect 4252 7284 4304 7336
rect 5080 7429 5089 7463
rect 5089 7429 5123 7463
rect 5123 7429 5132 7463
rect 5080 7420 5132 7429
rect 5908 7420 5960 7472
rect 9772 7420 9824 7472
rect 16028 7420 16080 7472
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 9220 7352 9272 7404
rect 9496 7352 9548 7404
rect 11520 7352 11572 7404
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 14924 7352 14976 7404
rect 5632 7284 5684 7336
rect 6460 7284 6512 7336
rect 7840 7284 7892 7336
rect 8668 7284 8720 7336
rect 9312 7284 9364 7336
rect 1768 7259 1820 7268
rect 1768 7225 1777 7259
rect 1777 7225 1811 7259
rect 1811 7225 1820 7259
rect 1768 7216 1820 7225
rect 6920 7259 6972 7268
rect 3976 7148 4028 7200
rect 6920 7225 6929 7259
rect 6929 7225 6963 7259
rect 6963 7225 6972 7259
rect 6920 7216 6972 7225
rect 7012 7259 7064 7268
rect 7012 7225 7021 7259
rect 7021 7225 7055 7259
rect 7055 7225 7064 7259
rect 7564 7259 7616 7268
rect 7012 7216 7064 7225
rect 7564 7225 7573 7259
rect 7573 7225 7607 7259
rect 7607 7225 7616 7259
rect 7564 7216 7616 7225
rect 7748 7216 7800 7268
rect 4344 7148 4396 7200
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 6552 7148 6604 7157
rect 6644 7148 6696 7200
rect 8484 7216 8536 7268
rect 9036 7216 9088 7268
rect 10048 7259 10100 7268
rect 10048 7225 10057 7259
rect 10057 7225 10091 7259
rect 10091 7225 10100 7259
rect 10048 7216 10100 7225
rect 10600 7259 10652 7268
rect 10600 7225 10609 7259
rect 10609 7225 10643 7259
rect 10643 7225 10652 7259
rect 10600 7216 10652 7225
rect 11428 7216 11480 7268
rect 13912 7259 13964 7268
rect 9404 7148 9456 7200
rect 9772 7148 9824 7200
rect 13912 7225 13921 7259
rect 13921 7225 13955 7259
rect 13955 7225 13964 7259
rect 13912 7216 13964 7225
rect 15752 7284 15804 7336
rect 16396 7352 16448 7404
rect 18788 7352 18840 7404
rect 15936 7284 15988 7336
rect 16580 7284 16632 7336
rect 17776 7327 17828 7336
rect 17776 7293 17785 7327
rect 17785 7293 17819 7327
rect 17819 7293 17828 7327
rect 17776 7284 17828 7293
rect 18420 7284 18472 7336
rect 14648 7216 14700 7268
rect 14280 7148 14332 7200
rect 14556 7148 14608 7200
rect 16764 7216 16816 7268
rect 16672 7191 16724 7200
rect 16672 7157 16681 7191
rect 16681 7157 16715 7191
rect 16715 7157 16724 7191
rect 16672 7148 16724 7157
rect 16856 7148 16908 7200
rect 17132 7148 17184 7200
rect 18880 7148 18932 7200
rect 8315 7046 8367 7098
rect 8379 7046 8431 7098
rect 8443 7046 8495 7098
rect 8507 7046 8559 7098
rect 15648 7046 15700 7098
rect 15712 7046 15764 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 1860 6944 1912 6996
rect 4988 6944 5040 6996
rect 5172 6987 5224 6996
rect 5172 6953 5181 6987
rect 5181 6953 5215 6987
rect 5215 6953 5224 6987
rect 5172 6944 5224 6953
rect 7748 6944 7800 6996
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 10048 6944 10100 6996
rect 12716 6987 12768 6996
rect 12716 6953 12725 6987
rect 12725 6953 12759 6987
rect 12759 6953 12768 6987
rect 12716 6944 12768 6953
rect 13820 6944 13872 6996
rect 16856 6944 16908 6996
rect 18788 6944 18840 6996
rect 19156 6944 19208 6996
rect 1768 6919 1820 6928
rect 1768 6885 1777 6919
rect 1777 6885 1811 6919
rect 1811 6885 1820 6919
rect 1768 6876 1820 6885
rect 5908 6919 5960 6928
rect 5908 6885 5917 6919
rect 5917 6885 5951 6919
rect 5951 6885 5960 6919
rect 5908 6876 5960 6885
rect 6736 6876 6788 6928
rect 7104 6876 7156 6928
rect 5356 6808 5408 6860
rect 5724 6808 5776 6860
rect 6644 6808 6696 6860
rect 1124 6672 1176 6724
rect 2320 6672 2372 6724
rect 3976 6740 4028 6792
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 8760 6876 8812 6928
rect 9864 6919 9916 6928
rect 9864 6885 9873 6919
rect 9873 6885 9907 6919
rect 9907 6885 9916 6919
rect 9864 6876 9916 6885
rect 10600 6876 10652 6928
rect 11336 6876 11388 6928
rect 13728 6919 13780 6928
rect 13728 6885 13737 6919
rect 13737 6885 13771 6919
rect 13771 6885 13780 6919
rect 13728 6876 13780 6885
rect 15200 6876 15252 6928
rect 4436 6740 4488 6749
rect 4068 6672 4120 6724
rect 5080 6672 5132 6724
rect 2688 6647 2740 6656
rect 2688 6613 2697 6647
rect 2697 6613 2731 6647
rect 2731 6613 2740 6647
rect 2688 6604 2740 6613
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 4252 6604 4304 6656
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 6552 6604 6604 6613
rect 6828 6647 6880 6656
rect 6828 6613 6837 6647
rect 6837 6613 6871 6647
rect 6871 6613 6880 6647
rect 6828 6604 6880 6613
rect 6920 6604 6972 6656
rect 7932 6851 7984 6860
rect 7932 6817 7941 6851
rect 7941 6817 7975 6851
rect 7975 6817 7984 6851
rect 7932 6808 7984 6817
rect 15016 6808 15068 6860
rect 15936 6808 15988 6860
rect 16856 6851 16908 6860
rect 16856 6817 16865 6851
rect 16865 6817 16899 6851
rect 16899 6817 16908 6851
rect 16856 6808 16908 6817
rect 17132 6851 17184 6860
rect 17132 6817 17141 6851
rect 17141 6817 17175 6851
rect 17175 6817 17184 6851
rect 17132 6808 17184 6817
rect 18696 6808 18748 6860
rect 19708 6808 19760 6860
rect 9220 6740 9272 6792
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 11428 6740 11480 6792
rect 11612 6783 11664 6792
rect 11612 6749 11621 6783
rect 11621 6749 11655 6783
rect 11655 6749 11664 6783
rect 11612 6740 11664 6749
rect 13820 6740 13872 6792
rect 7564 6672 7616 6724
rect 12716 6672 12768 6724
rect 16396 6740 16448 6792
rect 16948 6783 17000 6792
rect 16948 6749 16957 6783
rect 16957 6749 16991 6783
rect 16991 6749 17000 6783
rect 16948 6740 17000 6749
rect 17316 6783 17368 6792
rect 17316 6749 17325 6783
rect 17325 6749 17359 6783
rect 17359 6749 17368 6783
rect 17316 6740 17368 6749
rect 14464 6672 14516 6724
rect 17040 6672 17092 6724
rect 8668 6604 8720 6656
rect 8852 6647 8904 6656
rect 8852 6613 8861 6647
rect 8861 6613 8895 6647
rect 8895 6613 8904 6647
rect 8852 6604 8904 6613
rect 10784 6604 10836 6656
rect 18788 6604 18840 6656
rect 4648 6502 4700 6554
rect 4712 6502 4764 6554
rect 4776 6502 4828 6554
rect 4840 6502 4892 6554
rect 11982 6502 12034 6554
rect 12046 6502 12098 6554
rect 12110 6502 12162 6554
rect 12174 6502 12226 6554
rect 19315 6502 19367 6554
rect 19379 6502 19431 6554
rect 19443 6502 19495 6554
rect 19507 6502 19559 6554
rect 1768 6400 1820 6452
rect 3700 6443 3752 6452
rect 3700 6409 3709 6443
rect 3709 6409 3743 6443
rect 3743 6409 3752 6443
rect 3700 6400 3752 6409
rect 5724 6443 5776 6452
rect 5724 6409 5733 6443
rect 5733 6409 5767 6443
rect 5767 6409 5776 6443
rect 5724 6400 5776 6409
rect 5908 6400 5960 6452
rect 8024 6443 8076 6452
rect 8024 6409 8033 6443
rect 8033 6409 8067 6443
rect 8067 6409 8076 6443
rect 8024 6400 8076 6409
rect 11336 6443 11388 6452
rect 11336 6409 11345 6443
rect 11345 6409 11379 6443
rect 11379 6409 11388 6443
rect 11336 6400 11388 6409
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 3608 6332 3660 6384
rect 9956 6332 10008 6384
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5356 6264 5408 6273
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 10140 6264 10192 6316
rect 5172 6196 5224 6248
rect 2136 6171 2188 6180
rect 2136 6137 2145 6171
rect 2145 6137 2179 6171
rect 2179 6137 2188 6171
rect 2136 6128 2188 6137
rect 3056 6171 3108 6180
rect 3056 6137 3065 6171
rect 3065 6137 3099 6171
rect 3099 6137 3108 6171
rect 3056 6128 3108 6137
rect 4436 6128 4488 6180
rect 4988 6128 5040 6180
rect 7196 6196 7248 6248
rect 7840 6196 7892 6248
rect 8668 6196 8720 6248
rect 9312 6196 9364 6248
rect 12440 6239 12492 6248
rect 12440 6205 12449 6239
rect 12449 6205 12483 6239
rect 12483 6205 12492 6239
rect 12440 6196 12492 6205
rect 6644 6128 6696 6180
rect 8024 6128 8076 6180
rect 10048 6171 10100 6180
rect 10048 6137 10057 6171
rect 10057 6137 10091 6171
rect 10091 6137 10100 6171
rect 10048 6128 10100 6137
rect 3976 6060 4028 6112
rect 9404 6103 9456 6112
rect 9404 6069 9413 6103
rect 9413 6069 9447 6103
rect 9447 6069 9456 6103
rect 9404 6060 9456 6069
rect 9864 6060 9916 6112
rect 12716 6060 12768 6112
rect 13268 6400 13320 6452
rect 13728 6443 13780 6452
rect 13728 6409 13737 6443
rect 13737 6409 13771 6443
rect 13771 6409 13780 6443
rect 13728 6400 13780 6409
rect 14372 6400 14424 6452
rect 15936 6400 15988 6452
rect 16856 6443 16908 6452
rect 16856 6409 16865 6443
rect 16865 6409 16899 6443
rect 16899 6409 16908 6443
rect 16856 6400 16908 6409
rect 16948 6400 17000 6452
rect 18696 6400 18748 6452
rect 19708 6400 19760 6452
rect 19800 6400 19852 6452
rect 13820 6332 13872 6384
rect 14280 6307 14332 6316
rect 14280 6273 14289 6307
rect 14289 6273 14323 6307
rect 14323 6273 14332 6307
rect 14280 6264 14332 6273
rect 17040 6264 17092 6316
rect 15108 6196 15160 6248
rect 16120 6196 16172 6248
rect 16212 6239 16264 6248
rect 16212 6205 16221 6239
rect 16221 6205 16255 6239
rect 16255 6205 16264 6239
rect 16212 6196 16264 6205
rect 19800 6196 19852 6248
rect 14372 6171 14424 6180
rect 14372 6137 14381 6171
rect 14381 6137 14415 6171
rect 14415 6137 14424 6171
rect 14372 6128 14424 6137
rect 15476 6128 15528 6180
rect 15660 6128 15712 6180
rect 17132 6128 17184 6180
rect 14188 6060 14240 6112
rect 14556 6060 14608 6112
rect 14832 6060 14884 6112
rect 16028 6103 16080 6112
rect 16028 6069 16037 6103
rect 16037 6069 16071 6103
rect 16071 6069 16080 6103
rect 16028 6060 16080 6069
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 8315 5958 8367 6010
rect 8379 5958 8431 6010
rect 8443 5958 8495 6010
rect 8507 5958 8559 6010
rect 15648 5958 15700 6010
rect 15712 5958 15764 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 2136 5856 2188 5908
rect 3516 5856 3568 5908
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 5448 5899 5500 5908
rect 5448 5865 5457 5899
rect 5457 5865 5491 5899
rect 5491 5865 5500 5899
rect 5448 5856 5500 5865
rect 9404 5856 9456 5908
rect 9680 5856 9732 5908
rect 10048 5856 10100 5908
rect 12440 5856 12492 5908
rect 2412 5788 2464 5840
rect 4068 5788 4120 5840
rect 7932 5788 7984 5840
rect 8024 5788 8076 5840
rect 8944 5788 8996 5840
rect 9956 5788 10008 5840
rect 12716 5788 12768 5840
rect 5172 5720 5224 5772
rect 5448 5720 5500 5772
rect 6460 5763 6512 5772
rect 6460 5729 6469 5763
rect 6469 5729 6503 5763
rect 6503 5729 6512 5763
rect 6460 5720 6512 5729
rect 4436 5652 4488 5704
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 5540 5652 5592 5704
rect 7840 5695 7892 5704
rect 3700 5584 3752 5636
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 11428 5720 11480 5772
rect 12992 5720 13044 5772
rect 15384 5788 15436 5840
rect 16120 5788 16172 5840
rect 16304 5831 16356 5840
rect 16304 5797 16313 5831
rect 16313 5797 16347 5831
rect 16347 5797 16356 5831
rect 16304 5788 16356 5797
rect 13820 5763 13872 5772
rect 13820 5729 13829 5763
rect 13829 5729 13863 5763
rect 13863 5729 13872 5763
rect 14280 5763 14332 5772
rect 13820 5720 13872 5729
rect 14280 5729 14289 5763
rect 14289 5729 14323 5763
rect 14323 5729 14332 5763
rect 14280 5720 14332 5729
rect 15108 5763 15160 5772
rect 15108 5729 15117 5763
rect 15117 5729 15151 5763
rect 15151 5729 15160 5763
rect 15108 5720 15160 5729
rect 16488 5720 16540 5772
rect 17132 5720 17184 5772
rect 17316 5763 17368 5772
rect 17316 5729 17325 5763
rect 17325 5729 17359 5763
rect 17359 5729 17368 5763
rect 17316 5720 17368 5729
rect 18512 5720 18564 5772
rect 19064 5720 19116 5772
rect 12532 5695 12584 5704
rect 12532 5661 12541 5695
rect 12541 5661 12575 5695
rect 12575 5661 12584 5695
rect 12532 5652 12584 5661
rect 11244 5584 11296 5636
rect 15200 5584 15252 5636
rect 15476 5652 15528 5704
rect 15752 5652 15804 5704
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 6000 5559 6052 5568
rect 6000 5525 6009 5559
rect 6009 5525 6043 5559
rect 6043 5525 6052 5559
rect 6000 5516 6052 5525
rect 6368 5559 6420 5568
rect 6368 5525 6377 5559
rect 6377 5525 6411 5559
rect 6411 5525 6420 5559
rect 6368 5516 6420 5525
rect 6736 5516 6788 5568
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 11060 5559 11112 5568
rect 11060 5525 11069 5559
rect 11069 5525 11103 5559
rect 11103 5525 11112 5559
rect 11060 5516 11112 5525
rect 4648 5414 4700 5466
rect 4712 5414 4764 5466
rect 4776 5414 4828 5466
rect 4840 5414 4892 5466
rect 11982 5414 12034 5466
rect 12046 5414 12098 5466
rect 12110 5414 12162 5466
rect 12174 5414 12226 5466
rect 19315 5414 19367 5466
rect 19379 5414 19431 5466
rect 19443 5414 19495 5466
rect 19507 5414 19559 5466
rect 2412 5312 2464 5364
rect 4436 5355 4488 5364
rect 4436 5321 4445 5355
rect 4445 5321 4479 5355
rect 4479 5321 4488 5355
rect 4436 5312 4488 5321
rect 6828 5312 6880 5364
rect 8024 5355 8076 5364
rect 8024 5321 8033 5355
rect 8033 5321 8067 5355
rect 8067 5321 8076 5355
rect 8024 5312 8076 5321
rect 9404 5312 9456 5364
rect 9956 5312 10008 5364
rect 11244 5355 11296 5364
rect 11244 5321 11253 5355
rect 11253 5321 11287 5355
rect 11287 5321 11296 5355
rect 11244 5312 11296 5321
rect 12532 5312 12584 5364
rect 14004 5312 14056 5364
rect 15384 5355 15436 5364
rect 15384 5321 15393 5355
rect 15393 5321 15427 5355
rect 15427 5321 15436 5355
rect 15384 5312 15436 5321
rect 17132 5312 17184 5364
rect 18788 5312 18840 5364
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 3792 5176 3844 5228
rect 4252 5244 4304 5296
rect 7564 5287 7616 5296
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 3608 5151 3660 5160
rect 3608 5117 3617 5151
rect 3617 5117 3651 5151
rect 3651 5117 3660 5151
rect 3608 5108 3660 5117
rect 3700 5108 3752 5160
rect 4344 5151 4396 5160
rect 4344 5117 4353 5151
rect 4353 5117 4387 5151
rect 4387 5117 4396 5151
rect 6000 5176 6052 5228
rect 7564 5253 7573 5287
rect 7573 5253 7607 5287
rect 7607 5253 7616 5287
rect 7564 5244 7616 5253
rect 10600 5244 10652 5296
rect 12716 5287 12768 5296
rect 12716 5253 12725 5287
rect 12725 5253 12759 5287
rect 12759 5253 12768 5287
rect 12716 5244 12768 5253
rect 10692 5176 10744 5228
rect 15752 5244 15804 5296
rect 19064 5244 19116 5296
rect 15936 5219 15988 5228
rect 4344 5108 4396 5117
rect 1584 5083 1636 5092
rect 1584 5049 1593 5083
rect 1593 5049 1627 5083
rect 1627 5049 1636 5083
rect 1584 5040 1636 5049
rect 1676 5083 1728 5092
rect 1676 5049 1685 5083
rect 1685 5049 1719 5083
rect 1719 5049 1728 5083
rect 1676 5040 1728 5049
rect 2872 5040 2924 5092
rect 7288 5108 7340 5160
rect 8944 5108 8996 5160
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16580 5176 16632 5228
rect 17960 5108 18012 5160
rect 6828 5040 6880 5092
rect 8024 5040 8076 5092
rect 5080 4972 5132 5024
rect 5264 4972 5316 5024
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 12992 5083 13044 5092
rect 9864 4972 9916 5024
rect 12992 5049 13001 5083
rect 13001 5049 13035 5083
rect 13035 5049 13044 5083
rect 12992 5040 13044 5049
rect 13820 5040 13872 5092
rect 14464 5083 14516 5092
rect 14464 5049 14473 5083
rect 14473 5049 14507 5083
rect 14507 5049 14516 5083
rect 14464 5040 14516 5049
rect 14372 4972 14424 5024
rect 16120 5040 16172 5092
rect 15476 4972 15528 5024
rect 17316 4972 17368 5024
rect 17408 4972 17460 5024
rect 18512 5015 18564 5024
rect 18512 4981 18521 5015
rect 18521 4981 18555 5015
rect 18555 4981 18564 5015
rect 18512 4972 18564 4981
rect 8315 4870 8367 4922
rect 8379 4870 8431 4922
rect 8443 4870 8495 4922
rect 8507 4870 8559 4922
rect 15648 4870 15700 4922
rect 15712 4870 15764 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 2872 4811 2924 4820
rect 2412 4700 2464 4752
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 3792 4768 3844 4820
rect 2964 4700 3016 4752
rect 4528 4768 4580 4820
rect 7472 4811 7524 4820
rect 7472 4777 7481 4811
rect 7481 4777 7515 4811
rect 7515 4777 7524 4811
rect 7472 4768 7524 4777
rect 7840 4811 7892 4820
rect 7840 4777 7849 4811
rect 7849 4777 7883 4811
rect 7883 4777 7892 4811
rect 7840 4768 7892 4777
rect 8944 4811 8996 4820
rect 8944 4777 8953 4811
rect 8953 4777 8987 4811
rect 8987 4777 8996 4811
rect 8944 4768 8996 4777
rect 9220 4768 9272 4820
rect 9404 4768 9456 4820
rect 10692 4811 10744 4820
rect 3700 4632 3752 4684
rect 4160 4632 4212 4684
rect 4344 4675 4396 4684
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 6368 4700 6420 4752
rect 4988 4632 5040 4684
rect 5080 4675 5132 4684
rect 5080 4641 5089 4675
rect 5089 4641 5123 4675
rect 5123 4641 5132 4675
rect 5080 4632 5132 4641
rect 5264 4632 5316 4684
rect 6184 4632 6236 4684
rect 6552 4632 6604 4684
rect 7840 4632 7892 4684
rect 8116 4700 8168 4752
rect 8208 4700 8260 4752
rect 9864 4743 9916 4752
rect 9864 4709 9873 4743
rect 9873 4709 9907 4743
rect 9907 4709 9916 4743
rect 9864 4700 9916 4709
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 13084 4768 13136 4820
rect 11336 4700 11388 4752
rect 12716 4700 12768 4752
rect 12900 4743 12952 4752
rect 12900 4709 12909 4743
rect 12909 4709 12943 4743
rect 12943 4709 12952 4743
rect 12900 4700 12952 4709
rect 13820 4768 13872 4820
rect 14648 4768 14700 4820
rect 15108 4700 15160 4752
rect 8024 4632 8076 4684
rect 12348 4632 12400 4684
rect 1768 4496 1820 4548
rect 6920 4564 6972 4616
rect 8668 4607 8720 4616
rect 8668 4573 8677 4607
rect 8677 4573 8711 4607
rect 8711 4573 8720 4607
rect 8668 4564 8720 4573
rect 9128 4564 9180 4616
rect 9588 4564 9640 4616
rect 10140 4607 10192 4616
rect 5264 4496 5316 4548
rect 6368 4496 6420 4548
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 11704 4564 11756 4616
rect 15200 4632 15252 4684
rect 15384 4675 15436 4684
rect 15384 4641 15393 4675
rect 15393 4641 15427 4675
rect 15427 4641 15436 4675
rect 15384 4632 15436 4641
rect 16304 4632 16356 4684
rect 16672 4632 16724 4684
rect 17316 4675 17368 4684
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 18696 4632 18748 4684
rect 19156 4632 19208 4684
rect 11060 4539 11112 4548
rect 11060 4505 11069 4539
rect 11069 4505 11103 4539
rect 11103 4505 11112 4539
rect 11060 4496 11112 4505
rect 14004 4564 14056 4616
rect 5172 4428 5224 4480
rect 5448 4428 5500 4480
rect 6184 4428 6236 4480
rect 11244 4428 11296 4480
rect 13544 4428 13596 4480
rect 16580 4428 16632 4480
rect 18880 4428 18932 4480
rect 4648 4326 4700 4378
rect 4712 4326 4764 4378
rect 4776 4326 4828 4378
rect 4840 4326 4892 4378
rect 11982 4326 12034 4378
rect 12046 4326 12098 4378
rect 12110 4326 12162 4378
rect 12174 4326 12226 4378
rect 19315 4326 19367 4378
rect 19379 4326 19431 4378
rect 19443 4326 19495 4378
rect 19507 4326 19559 4378
rect 2136 4224 2188 4276
rect 3056 4224 3108 4276
rect 3608 4224 3660 4276
rect 4344 4224 4396 4276
rect 6644 4267 6696 4276
rect 6644 4233 6653 4267
rect 6653 4233 6687 4267
rect 6687 4233 6696 4267
rect 6644 4224 6696 4233
rect 5264 4199 5316 4208
rect 5264 4165 5273 4199
rect 5273 4165 5307 4199
rect 5307 4165 5316 4199
rect 5264 4156 5316 4165
rect 5448 4156 5500 4208
rect 7472 4224 7524 4276
rect 7564 4224 7616 4276
rect 1860 4088 1912 4140
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 4252 4088 4304 4140
rect 7288 4088 7340 4140
rect 8208 4088 8260 4140
rect 4068 4063 4120 4072
rect 1768 3995 1820 4004
rect 1768 3961 1777 3995
rect 1777 3961 1811 3995
rect 1811 3961 1820 3995
rect 1768 3952 1820 3961
rect 4068 4029 4077 4063
rect 4077 4029 4111 4063
rect 4111 4029 4120 4063
rect 4068 4020 4120 4029
rect 4528 4020 4580 4072
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 5264 4020 5316 4072
rect 5540 4020 5592 4072
rect 6644 4020 6696 4072
rect 4252 3952 4304 4004
rect 4436 3952 4488 4004
rect 8116 4020 8168 4072
rect 9404 4224 9456 4276
rect 9864 4267 9916 4276
rect 9864 4233 9873 4267
rect 9873 4233 9907 4267
rect 9907 4233 9916 4267
rect 9864 4224 9916 4233
rect 11060 4224 11112 4276
rect 12716 4224 12768 4276
rect 13912 4224 13964 4276
rect 14372 4224 14424 4276
rect 14556 4224 14608 4276
rect 15384 4224 15436 4276
rect 16672 4267 16724 4276
rect 16672 4233 16681 4267
rect 16681 4233 16715 4267
rect 16715 4233 16724 4267
rect 16672 4224 16724 4233
rect 19156 4267 19208 4276
rect 19156 4233 19165 4267
rect 19165 4233 19199 4267
rect 19199 4233 19208 4267
rect 19156 4224 19208 4233
rect 10600 4156 10652 4208
rect 11336 4199 11388 4208
rect 11336 4165 11345 4199
rect 11345 4165 11379 4199
rect 11379 4165 11388 4199
rect 11336 4156 11388 4165
rect 11704 4199 11756 4208
rect 11704 4165 11713 4199
rect 11713 4165 11747 4199
rect 11747 4165 11756 4199
rect 11704 4156 11756 4165
rect 14648 4156 14700 4208
rect 18328 4199 18380 4208
rect 18328 4165 18337 4199
rect 18337 4165 18371 4199
rect 18371 4165 18380 4199
rect 18328 4156 18380 4165
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 12348 4088 12400 4140
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 17500 4088 17552 4140
rect 21548 4088 21600 4140
rect 8760 3952 8812 4004
rect 10232 3995 10284 4004
rect 10232 3961 10241 3995
rect 10241 3961 10275 3995
rect 10275 3961 10284 3995
rect 10232 3952 10284 3961
rect 16764 4020 16816 4072
rect 18052 4020 18104 4072
rect 18236 4020 18288 4072
rect 13728 3952 13780 4004
rect 15016 3952 15068 4004
rect 15476 3995 15528 4004
rect 15476 3961 15485 3995
rect 15485 3961 15519 3995
rect 15519 3961 15528 3995
rect 15476 3952 15528 3961
rect 15844 3952 15896 4004
rect 16120 3952 16172 4004
rect 3884 3884 3936 3936
rect 4988 3884 5040 3936
rect 5264 3884 5316 3936
rect 5448 3884 5500 3936
rect 5816 3884 5868 3936
rect 6368 3884 6420 3936
rect 9496 3927 9548 3936
rect 9496 3893 9505 3927
rect 9505 3893 9539 3927
rect 9539 3893 9548 3927
rect 9496 3884 9548 3893
rect 13912 3927 13964 3936
rect 13912 3893 13921 3927
rect 13921 3893 13955 3927
rect 13955 3893 13964 3927
rect 13912 3884 13964 3893
rect 15108 3927 15160 3936
rect 15108 3893 15117 3927
rect 15117 3893 15151 3927
rect 15151 3893 15160 3927
rect 15108 3884 15160 3893
rect 15292 3884 15344 3936
rect 16856 3927 16908 3936
rect 16856 3893 16865 3927
rect 16865 3893 16899 3927
rect 16899 3893 16908 3927
rect 16856 3884 16908 3893
rect 17316 3927 17368 3936
rect 17316 3893 17325 3927
rect 17325 3893 17359 3927
rect 17359 3893 17368 3927
rect 17316 3884 17368 3893
rect 21088 3952 21140 4004
rect 8315 3782 8367 3834
rect 8379 3782 8431 3834
rect 8443 3782 8495 3834
rect 8507 3782 8559 3834
rect 15648 3782 15700 3834
rect 15712 3782 15764 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 2136 3723 2188 3732
rect 2136 3689 2145 3723
rect 2145 3689 2179 3723
rect 2179 3689 2188 3723
rect 2136 3680 2188 3689
rect 4068 3680 4120 3732
rect 5080 3680 5132 3732
rect 7564 3723 7616 3732
rect 7564 3689 7573 3723
rect 7573 3689 7607 3723
rect 7607 3689 7616 3723
rect 7564 3680 7616 3689
rect 8668 3680 8720 3732
rect 10232 3680 10284 3732
rect 2964 3612 3016 3664
rect 7196 3655 7248 3664
rect 3056 3587 3108 3596
rect 3056 3553 3065 3587
rect 3065 3553 3099 3587
rect 3099 3553 3108 3587
rect 3056 3544 3108 3553
rect 4344 3544 4396 3596
rect 5080 3587 5132 3596
rect 5080 3553 5089 3587
rect 5089 3553 5123 3587
rect 5123 3553 5132 3587
rect 5080 3544 5132 3553
rect 5540 3544 5592 3596
rect 6644 3587 6696 3596
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 6828 3587 6880 3596
rect 6828 3553 6837 3587
rect 6837 3553 6871 3587
rect 6871 3553 6880 3587
rect 6828 3544 6880 3553
rect 7196 3621 7205 3655
rect 7205 3621 7239 3655
rect 7239 3621 7248 3655
rect 7196 3612 7248 3621
rect 8208 3655 8260 3664
rect 8208 3621 8217 3655
rect 8217 3621 8251 3655
rect 8251 3621 8260 3655
rect 8208 3612 8260 3621
rect 9864 3655 9916 3664
rect 9864 3621 9873 3655
rect 9873 3621 9907 3655
rect 9907 3621 9916 3655
rect 9864 3612 9916 3621
rect 12440 3680 12492 3732
rect 13084 3723 13136 3732
rect 13084 3689 13093 3723
rect 13093 3689 13127 3723
rect 13127 3689 13136 3723
rect 13084 3680 13136 3689
rect 15476 3680 15528 3732
rect 16304 3723 16356 3732
rect 16304 3689 16313 3723
rect 16313 3689 16347 3723
rect 16347 3689 16356 3723
rect 16304 3680 16356 3689
rect 16948 3723 17000 3732
rect 16948 3689 16957 3723
rect 16957 3689 16991 3723
rect 16991 3689 17000 3723
rect 16948 3680 17000 3689
rect 13912 3612 13964 3664
rect 5632 3476 5684 3528
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 112 3408 164 3460
rect 6276 3408 6328 3460
rect 6552 3451 6604 3460
rect 6552 3417 6561 3451
rect 6561 3417 6595 3451
rect 6595 3417 6604 3451
rect 6552 3408 6604 3417
rect 15016 3587 15068 3596
rect 15016 3553 15025 3587
rect 15025 3553 15059 3587
rect 15059 3553 15068 3587
rect 15016 3544 15068 3553
rect 15568 3587 15620 3596
rect 15568 3553 15577 3587
rect 15577 3553 15611 3587
rect 15611 3553 15620 3587
rect 15568 3544 15620 3553
rect 17132 3587 17184 3596
rect 17132 3553 17141 3587
rect 17141 3553 17175 3587
rect 17175 3553 17184 3587
rect 17132 3544 17184 3553
rect 17316 3587 17368 3596
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 19064 3587 19116 3596
rect 19064 3553 19073 3587
rect 19073 3553 19107 3587
rect 19107 3553 19116 3587
rect 19064 3544 19116 3553
rect 9404 3476 9456 3528
rect 10140 3476 10192 3528
rect 11152 3476 11204 3528
rect 13452 3519 13504 3528
rect 8852 3408 8904 3460
rect 10416 3408 10468 3460
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 16580 3476 16632 3528
rect 17408 3408 17460 3460
rect 2228 3340 2280 3392
rect 3792 3340 3844 3392
rect 4436 3340 4488 3392
rect 6184 3383 6236 3392
rect 6184 3349 6193 3383
rect 6193 3349 6227 3383
rect 6227 3349 6236 3383
rect 6184 3340 6236 3349
rect 9128 3340 9180 3392
rect 10600 3340 10652 3392
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 14648 3340 14700 3349
rect 4648 3238 4700 3290
rect 4712 3238 4764 3290
rect 4776 3238 4828 3290
rect 4840 3238 4892 3290
rect 11982 3238 12034 3290
rect 12046 3238 12098 3290
rect 12110 3238 12162 3290
rect 12174 3238 12226 3290
rect 19315 3238 19367 3290
rect 19379 3238 19431 3290
rect 19443 3238 19495 3290
rect 19507 3238 19559 3290
rect 3976 3136 4028 3188
rect 4068 3136 4120 3188
rect 6644 3136 6696 3188
rect 8760 3136 8812 3188
rect 9864 3136 9916 3188
rect 13452 3136 13504 3188
rect 16948 3136 17000 3188
rect 17132 3136 17184 3188
rect 2320 3111 2372 3120
rect 2320 3077 2329 3111
rect 2329 3077 2363 3111
rect 2363 3077 2372 3111
rect 2320 3068 2372 3077
rect 3332 3068 3384 3120
rect 2136 3000 2188 3052
rect 2504 3000 2556 3052
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 2596 2932 2648 2984
rect 5080 3068 5132 3120
rect 8208 3068 8260 3120
rect 4252 3043 4304 3052
rect 4252 3009 4261 3043
rect 4261 3009 4295 3043
rect 4295 3009 4304 3043
rect 4252 3000 4304 3009
rect 3700 2975 3752 2984
rect 3700 2941 3709 2975
rect 3709 2941 3743 2975
rect 3743 2941 3752 2975
rect 3884 2975 3936 2984
rect 3700 2932 3752 2941
rect 3884 2941 3893 2975
rect 3893 2941 3927 2975
rect 3927 2941 3936 2975
rect 6552 3000 6604 3052
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 8668 3000 8720 3052
rect 9220 3000 9272 3052
rect 5448 2975 5500 2984
rect 3884 2932 3936 2941
rect 5448 2941 5457 2975
rect 5457 2941 5491 2975
rect 5491 2941 5500 2975
rect 5448 2932 5500 2941
rect 5632 2975 5684 2984
rect 5632 2941 5641 2975
rect 5641 2941 5675 2975
rect 5675 2941 5684 2975
rect 5632 2932 5684 2941
rect 7748 2932 7800 2984
rect 8116 2932 8168 2984
rect 10600 2975 10652 2984
rect 112 2864 164 2916
rect 3976 2864 4028 2916
rect 3056 2839 3108 2848
rect 3056 2805 3065 2839
rect 3065 2805 3099 2839
rect 3099 2805 3108 2839
rect 6828 2864 6880 2916
rect 7564 2864 7616 2916
rect 8760 2864 8812 2916
rect 10600 2941 10609 2975
rect 10609 2941 10643 2975
rect 10643 2941 10652 2975
rect 10600 2932 10652 2941
rect 14188 3000 14240 3052
rect 16856 3068 16908 3120
rect 15568 3043 15620 3052
rect 15568 3009 15577 3043
rect 15577 3009 15611 3043
rect 15611 3009 15620 3043
rect 15568 3000 15620 3009
rect 16120 3000 16172 3052
rect 13268 2932 13320 2984
rect 13912 2932 13964 2984
rect 15936 2932 15988 2984
rect 16304 2932 16356 2984
rect 4712 2839 4764 2848
rect 3056 2796 3108 2805
rect 4712 2805 4721 2839
rect 4721 2805 4755 2839
rect 4755 2805 4764 2839
rect 4712 2796 4764 2805
rect 5080 2839 5132 2848
rect 5080 2805 5089 2839
rect 5089 2805 5123 2839
rect 5123 2805 5132 2839
rect 5080 2796 5132 2805
rect 6276 2796 6328 2848
rect 8668 2796 8720 2848
rect 9220 2796 9272 2848
rect 12716 2839 12768 2848
rect 12716 2805 12725 2839
rect 12725 2805 12759 2839
rect 12759 2805 12768 2839
rect 12716 2796 12768 2805
rect 14648 2864 14700 2916
rect 15108 2796 15160 2848
rect 15200 2796 15252 2848
rect 15936 2796 15988 2848
rect 16120 2796 16172 2848
rect 17316 2932 17368 2984
rect 17776 2932 17828 2984
rect 16488 2864 16540 2916
rect 16672 2796 16724 2848
rect 17776 2839 17828 2848
rect 17776 2805 17785 2839
rect 17785 2805 17819 2839
rect 17819 2805 17828 2839
rect 17776 2796 17828 2805
rect 19064 2839 19116 2848
rect 19064 2805 19073 2839
rect 19073 2805 19107 2839
rect 19107 2805 19116 2839
rect 19064 2796 19116 2805
rect 8315 2694 8367 2746
rect 8379 2694 8431 2746
rect 8443 2694 8495 2746
rect 8507 2694 8559 2746
rect 15648 2694 15700 2746
rect 15712 2694 15764 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 3700 2635 3752 2644
rect 3700 2601 3709 2635
rect 3709 2601 3743 2635
rect 3743 2601 3752 2635
rect 3700 2592 3752 2601
rect 8208 2592 8260 2644
rect 9220 2592 9272 2644
rect 9312 2592 9364 2644
rect 10140 2592 10192 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 12716 2592 12768 2644
rect 13268 2635 13320 2644
rect 3608 2524 3660 2576
rect 4712 2524 4764 2576
rect 5632 2524 5684 2576
rect 9496 2567 9548 2576
rect 2320 2363 2372 2372
rect 1676 2295 1728 2304
rect 1676 2261 1685 2295
rect 1685 2261 1719 2295
rect 1719 2261 1728 2295
rect 2320 2329 2329 2363
rect 2329 2329 2363 2363
rect 2363 2329 2372 2363
rect 2320 2320 2372 2329
rect 2504 2499 2556 2508
rect 2504 2465 2513 2499
rect 2513 2465 2547 2499
rect 2547 2465 2556 2499
rect 2504 2456 2556 2465
rect 4528 2456 4580 2508
rect 5172 2456 5224 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 5816 2456 5868 2508
rect 3700 2320 3752 2372
rect 4528 2320 4580 2372
rect 5724 2388 5776 2440
rect 7288 2456 7340 2508
rect 9496 2533 9505 2567
rect 9505 2533 9539 2567
rect 9539 2533 9548 2567
rect 9496 2524 9548 2533
rect 7564 2456 7616 2508
rect 5356 2363 5408 2372
rect 1676 2252 1728 2261
rect 5080 2295 5132 2304
rect 5080 2261 5089 2295
rect 5089 2261 5123 2295
rect 5123 2261 5132 2295
rect 5080 2252 5132 2261
rect 5356 2329 5365 2363
rect 5365 2329 5399 2363
rect 5399 2329 5408 2363
rect 5356 2320 5408 2329
rect 5816 2320 5868 2372
rect 6460 2388 6512 2440
rect 7012 2388 7064 2440
rect 10140 2456 10192 2508
rect 12624 2524 12676 2576
rect 13268 2601 13277 2635
rect 13277 2601 13311 2635
rect 13311 2601 13320 2635
rect 13268 2592 13320 2601
rect 14648 2592 14700 2644
rect 16580 2635 16632 2644
rect 16580 2601 16589 2635
rect 16589 2601 16623 2635
rect 16623 2601 16632 2635
rect 16580 2592 16632 2601
rect 17500 2592 17552 2644
rect 18788 2635 18840 2644
rect 18788 2601 18797 2635
rect 18797 2601 18831 2635
rect 18831 2601 18840 2635
rect 18788 2592 18840 2601
rect 14832 2456 14884 2508
rect 15292 2456 15344 2508
rect 15568 2499 15620 2508
rect 15568 2465 15577 2499
rect 15577 2465 15611 2499
rect 15611 2465 15620 2499
rect 15568 2456 15620 2465
rect 15752 2499 15804 2508
rect 15752 2465 15761 2499
rect 15761 2465 15795 2499
rect 15795 2465 15804 2499
rect 15752 2456 15804 2465
rect 16764 2456 16816 2508
rect 18052 2456 18104 2508
rect 13636 2388 13688 2440
rect 14188 2388 14240 2440
rect 14924 2388 14976 2440
rect 7104 2320 7156 2372
rect 7656 2252 7708 2304
rect 8024 2295 8076 2304
rect 8024 2261 8033 2295
rect 8033 2261 8067 2295
rect 8067 2261 8076 2295
rect 8024 2252 8076 2261
rect 10048 2320 10100 2372
rect 15384 2320 15436 2372
rect 14832 2295 14884 2304
rect 14832 2261 14841 2295
rect 14841 2261 14875 2295
rect 14875 2261 14884 2295
rect 14832 2252 14884 2261
rect 15108 2252 15160 2304
rect 15752 2252 15804 2304
rect 17224 2295 17276 2304
rect 17224 2261 17233 2295
rect 17233 2261 17267 2295
rect 17267 2261 17276 2295
rect 17224 2252 17276 2261
rect 18052 2295 18104 2304
rect 18052 2261 18061 2295
rect 18061 2261 18095 2295
rect 18095 2261 18104 2295
rect 18052 2252 18104 2261
rect 4648 2150 4700 2202
rect 4712 2150 4764 2202
rect 4776 2150 4828 2202
rect 4840 2150 4892 2202
rect 11982 2150 12034 2202
rect 12046 2150 12098 2202
rect 12110 2150 12162 2202
rect 12174 2150 12226 2202
rect 19315 2150 19367 2202
rect 19379 2150 19431 2202
rect 19443 2150 19495 2202
rect 19507 2150 19559 2202
rect 4528 2048 4580 2100
rect 5356 2048 5408 2100
rect 8024 1980 8076 2032
rect 18420 1980 18472 2032
rect 12072 1912 12124 1964
rect 18512 1912 18564 1964
<< metal2 >>
rect 1030 21584 1086 22000
rect 3146 21570 3202 22000
rect 5354 21570 5410 22000
rect 1030 21519 1086 21528
rect 2884 21542 3202 21570
rect 18 20360 74 20369
rect 18 20295 74 20304
rect 32 17270 60 20295
rect 2884 19514 2912 21542
rect 3146 21520 3202 21542
rect 5092 21542 5410 21570
rect 2962 20904 3018 20913
rect 2962 20839 3018 20848
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 1124 19304 1176 19310
rect 110 19272 166 19281
rect 166 19230 336 19258
rect 1124 19246 1176 19252
rect 110 19207 166 19216
rect 20 17264 72 17270
rect 20 17206 72 17212
rect 110 17232 166 17241
rect 166 17190 244 17218
rect 110 17167 166 17176
rect 20 11552 72 11558
rect 20 11494 72 11500
rect 32 8809 60 11494
rect 112 10464 164 10470
rect 112 10406 164 10412
rect 124 9897 152 10406
rect 110 9888 166 9897
rect 110 9823 166 9832
rect 216 9654 244 17190
rect 308 16697 336 19230
rect 294 16688 350 16697
rect 294 16623 350 16632
rect 204 9648 256 9654
rect 204 9590 256 9596
rect 18 8800 74 8809
rect 18 8735 74 8744
rect 1136 6730 1164 19246
rect 1308 19236 1360 19242
rect 1308 19178 1360 19184
rect 1320 18222 1348 19178
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1308 18216 1360 18222
rect 1308 18158 1360 18164
rect 1214 17776 1270 17785
rect 1214 17711 1270 17720
rect 1228 10266 1256 17711
rect 1320 17649 1348 18158
rect 1306 17640 1362 17649
rect 1306 17575 1362 17584
rect 1216 10260 1268 10266
rect 1216 10202 1268 10208
rect 1320 9042 1348 17575
rect 1398 14648 1454 14657
rect 1398 14583 1454 14592
rect 1412 14074 1440 14583
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1412 11694 1440 14010
rect 1504 12850 1532 19110
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 1860 18624 1912 18630
rect 1860 18566 1912 18572
rect 1872 18154 1900 18566
rect 1860 18148 1912 18154
rect 1860 18090 1912 18096
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1596 16998 1624 17682
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1582 16416 1638 16425
rect 1582 16351 1638 16360
rect 1596 16250 1624 16351
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1688 15706 1716 18022
rect 1872 17746 1900 18090
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1688 15026 1716 15642
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1780 13326 1808 17614
rect 1872 17338 1900 17682
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1872 13814 1900 16934
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1964 16250 1992 16730
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 1964 15638 1992 16186
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 1952 15632 2004 15638
rect 2056 15609 2084 15846
rect 2148 15706 2176 16594
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 1952 15574 2004 15580
rect 2042 15600 2098 15609
rect 1964 14822 1992 15574
rect 2240 15570 2268 18906
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2332 17882 2360 18770
rect 2688 18692 2740 18698
rect 2688 18634 2740 18640
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2700 17814 2728 18634
rect 2688 17808 2740 17814
rect 2688 17750 2740 17756
rect 2976 17610 3004 20839
rect 4622 19612 4918 19632
rect 4678 19610 4702 19612
rect 4758 19610 4782 19612
rect 4838 19610 4862 19612
rect 4700 19558 4702 19610
rect 4764 19558 4776 19610
rect 4838 19558 4840 19610
rect 4678 19556 4702 19558
rect 4758 19556 4782 19558
rect 4838 19556 4862 19558
rect 4622 19536 4918 19556
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 3056 18624 3108 18630
rect 3056 18566 3108 18572
rect 3068 18222 3096 18566
rect 3516 18352 3568 18358
rect 3516 18294 3568 18300
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 2964 17604 3016 17610
rect 2964 17546 3016 17552
rect 2780 17536 2832 17542
rect 2780 17478 2832 17484
rect 2792 17066 2820 17478
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2792 16794 2820 17002
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2884 16794 2912 16934
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 3068 16658 3096 18022
rect 3160 17882 3188 18022
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2976 15978 3004 16390
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2042 15535 2098 15544
rect 2228 15564 2280 15570
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14618 1992 14758
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1872 13786 1992 13814
rect 1860 13456 1912 13462
rect 1860 13398 1912 13404
rect 1768 13320 1820 13326
rect 1768 13262 1820 13268
rect 1492 12844 1544 12850
rect 1492 12786 1544 12792
rect 1872 12646 1900 13398
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 1872 12442 1900 12582
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1964 11370 1992 13786
rect 1780 11342 1992 11370
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1308 9036 1360 9042
rect 1308 8978 1360 8984
rect 1320 8022 1348 8978
rect 1504 8090 1532 9454
rect 1688 9178 1716 10950
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1308 8016 1360 8022
rect 1308 7958 1360 7964
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1688 7546 1716 7890
rect 1780 7886 1808 11342
rect 2056 9042 2084 15535
rect 2228 15506 2280 15512
rect 2240 14618 2268 15506
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 2228 13252 2280 13258
rect 2228 13194 2280 13200
rect 2240 12714 2268 13194
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 2240 12442 2268 12650
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2148 11082 2176 12174
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 1872 8430 1900 8978
rect 1950 8936 2006 8945
rect 1950 8871 2006 8880
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1780 7392 1808 7822
rect 1780 7364 1900 7392
rect 1768 7268 1820 7274
rect 1768 7210 1820 7216
rect 1780 6934 1808 7210
rect 1872 7002 1900 7364
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1768 6928 1820 6934
rect 1768 6870 1820 6876
rect 1124 6724 1176 6730
rect 1124 6666 1176 6672
rect 1780 6458 1808 6870
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1964 6225 1992 8871
rect 2148 8362 2176 11018
rect 2332 10130 2360 11086
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2240 9518 2268 9862
rect 2424 9602 2452 13942
rect 2608 13802 2636 14486
rect 2976 14006 3004 15914
rect 2964 14000 3016 14006
rect 2964 13942 3016 13948
rect 2504 13796 2556 13802
rect 2504 13738 2556 13744
rect 2596 13796 2648 13802
rect 2596 13738 2648 13744
rect 2516 13530 2544 13738
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2608 13394 2636 13738
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11286 2544 11494
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2516 10810 2544 11222
rect 2792 11150 2820 12650
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2976 12442 3004 12582
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11694 2912 12038
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2516 10266 2544 10746
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2608 10198 2636 10406
rect 2700 10266 2728 10474
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2608 9722 2636 10134
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2332 9574 2452 9602
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2332 8945 2360 9574
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 2318 8936 2374 8945
rect 2318 8871 2374 8880
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2056 6322 2084 7482
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1950 6216 2006 6225
rect 1950 6151 2006 6160
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1582 5264 1638 5273
rect 1582 5199 1638 5208
rect 1596 5098 1624 5199
rect 1688 5098 1716 5510
rect 2056 5234 2084 6258
rect 2148 6186 2176 7278
rect 2320 6724 2372 6730
rect 2320 6666 2372 6672
rect 2332 6322 2360 6666
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2136 6180 2188 6186
rect 2136 6122 2188 6128
rect 2148 5914 2176 6122
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2424 5846 2452 9386
rect 2502 9072 2558 9081
rect 2502 9007 2558 9016
rect 2780 9036 2832 9042
rect 2516 8974 2544 9007
rect 2780 8978 2832 8984
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2516 8498 2544 8910
rect 2792 8634 2820 8978
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2884 8294 2912 11630
rect 2976 11558 3004 12378
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2976 10198 3004 10950
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 2976 9722 3004 10134
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 3068 9178 3096 16458
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3160 15706 3188 15846
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3146 10568 3202 10577
rect 3146 10503 3202 10512
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2516 8090 2544 8230
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2516 7954 2544 8026
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6225 2728 6598
rect 2686 6216 2742 6225
rect 2686 6151 2742 6160
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 2424 5370 2452 5782
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 1584 5092 1636 5098
rect 1584 5034 1636 5040
rect 1676 5092 1728 5098
rect 1676 5034 1728 5040
rect 1688 5001 1716 5034
rect 1674 4992 1730 5001
rect 1674 4927 1730 4936
rect 1768 4548 1820 4554
rect 1768 4490 1820 4496
rect 1780 4010 1808 4490
rect 2056 4146 2084 5170
rect 2424 4758 2452 5306
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1872 4049 1900 4082
rect 1858 4040 1914 4049
rect 1768 4004 1820 4010
rect 1858 3975 1914 3984
rect 1768 3946 1820 3952
rect 2148 3738 2176 4218
rect 2424 4154 2452 4694
rect 2700 4154 2728 6151
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2884 4826 2912 5034
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2240 4126 2452 4154
rect 2608 4126 2728 4154
rect 2884 4154 2912 4762
rect 2976 4758 3004 8774
rect 3160 7954 3188 10503
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3332 10056 3384 10062
rect 3436 10033 3464 10202
rect 3332 9998 3384 10004
rect 3422 10024 3478 10033
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3252 8430 3280 9114
rect 3344 9042 3372 9998
rect 3422 9959 3478 9968
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3436 8090 3464 8434
rect 3528 8090 3556 18294
rect 3976 17808 4028 17814
rect 3976 17750 4028 17756
rect 3884 17740 3936 17746
rect 3884 17682 3936 17688
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3620 17134 3648 17478
rect 3896 17202 3924 17682
rect 3884 17196 3936 17202
rect 3712 17156 3884 17184
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 3620 16046 3648 17070
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3606 13288 3662 13297
rect 3606 13223 3662 13232
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3160 7478 3188 7890
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 3068 4282 3096 6122
rect 3252 5273 3280 7686
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6497 3464 6598
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3620 6390 3648 13223
rect 3712 8362 3740 17156
rect 3884 17138 3936 17144
rect 3988 17134 4016 17750
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3804 14822 3832 15438
rect 3896 15026 3924 16934
rect 3988 16522 4016 17070
rect 4080 16794 4108 19110
rect 5092 18970 5120 21542
rect 5354 21520 5410 21542
rect 7562 21570 7618 22000
rect 9770 21570 9826 22000
rect 11978 21570 12034 22000
rect 7562 21542 7788 21570
rect 7562 21520 7618 21542
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 6276 19304 6328 19310
rect 6276 19246 6328 19252
rect 5276 18970 5304 19246
rect 6000 19236 6052 19242
rect 6000 19178 6052 19184
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 4622 18524 4918 18544
rect 4678 18522 4702 18524
rect 4758 18522 4782 18524
rect 4838 18522 4862 18524
rect 4700 18470 4702 18522
rect 4764 18470 4776 18522
rect 4838 18470 4840 18522
rect 4678 18468 4702 18470
rect 4758 18468 4782 18470
rect 4838 18468 4862 18470
rect 4622 18448 4918 18468
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4172 16998 4200 17682
rect 4356 17524 4384 18158
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 4436 17536 4488 17542
rect 4356 17496 4436 17524
rect 4356 17270 4384 17496
rect 4436 17478 4488 17484
rect 4540 17354 4568 17614
rect 5092 17542 5120 18770
rect 5276 18698 5304 18906
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5172 17604 5224 17610
rect 5172 17546 5224 17552
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 4622 17436 4918 17456
rect 4678 17434 4702 17436
rect 4758 17434 4782 17436
rect 4838 17434 4862 17436
rect 4700 17382 4702 17434
rect 4764 17382 4776 17434
rect 4838 17382 4840 17434
rect 4678 17380 4702 17382
rect 4758 17380 4782 17382
rect 4838 17380 4862 17382
rect 4622 17360 4918 17380
rect 4448 17326 4568 17354
rect 4344 17264 4396 17270
rect 4344 17206 4396 17212
rect 4356 17134 4384 17206
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 4264 16250 4292 16526
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4264 15162 4292 15574
rect 4356 15348 4384 17070
rect 4448 17066 4476 17326
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 4448 16182 4476 17002
rect 4528 16516 4580 16522
rect 4528 16458 4580 16464
rect 4436 16176 4488 16182
rect 4436 16118 4488 16124
rect 4540 16114 4568 16458
rect 5184 16454 5212 17546
rect 5276 16658 5304 18226
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 4622 16348 4918 16368
rect 4678 16346 4702 16348
rect 4758 16346 4782 16348
rect 4838 16346 4862 16348
rect 4700 16294 4702 16346
rect 4764 16294 4776 16346
rect 4838 16294 4840 16346
rect 4678 16292 4702 16294
rect 4758 16292 4782 16294
rect 4838 16292 4862 16294
rect 4622 16272 4918 16292
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4436 16040 4488 16046
rect 4632 15994 4660 16118
rect 4436 15982 4488 15988
rect 4448 15502 4476 15982
rect 4540 15966 4660 15994
rect 5080 15972 5132 15978
rect 4436 15496 4488 15502
rect 4436 15438 4488 15444
rect 4356 15320 4476 15348
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3804 14550 3832 14758
rect 4356 14550 4384 14826
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 4344 14544 4396 14550
rect 4344 14486 4396 14492
rect 4448 14278 4476 15320
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4436 14272 4488 14278
rect 4436 14214 4488 14220
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 4080 12782 4108 13126
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3804 12442 3832 12650
rect 4080 12442 4108 12718
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4172 12306 4200 14214
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4448 13802 4476 14010
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4436 13796 4488 13802
rect 4436 13738 4488 13744
rect 4356 13462 4384 13738
rect 4540 13682 4568 15966
rect 5080 15914 5132 15920
rect 4622 15260 4918 15280
rect 4678 15258 4702 15260
rect 4758 15258 4782 15260
rect 4838 15258 4862 15260
rect 4700 15206 4702 15258
rect 4764 15206 4776 15258
rect 4838 15206 4840 15258
rect 4678 15204 4702 15206
rect 4758 15204 4782 15206
rect 4838 15204 4862 15206
rect 4622 15184 4918 15204
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4724 14822 4752 15030
rect 5092 14822 5120 15914
rect 5184 15586 5212 16390
rect 5276 15706 5304 16594
rect 5368 16153 5396 16934
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5354 16144 5410 16153
rect 5354 16079 5410 16088
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5184 15558 5304 15586
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5092 14550 5120 14758
rect 5080 14544 5132 14550
rect 5080 14486 5132 14492
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 4622 14172 4918 14192
rect 4678 14170 4702 14172
rect 4758 14170 4782 14172
rect 4838 14170 4862 14172
rect 4700 14118 4702 14170
rect 4764 14118 4776 14170
rect 4838 14118 4840 14170
rect 4678 14116 4702 14118
rect 4758 14116 4782 14118
rect 4838 14116 4862 14118
rect 4622 14096 4918 14116
rect 5000 14006 5028 14350
rect 5092 14074 5120 14486
rect 5172 14340 5224 14346
rect 5172 14282 5224 14288
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4988 14000 5040 14006
rect 4988 13942 5040 13948
rect 4448 13654 4568 13682
rect 4344 13456 4396 13462
rect 4344 13398 4396 13404
rect 4356 12986 4384 13398
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4080 11354 4108 12242
rect 4172 11898 4200 12242
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3790 11248 3846 11257
rect 3790 11183 3846 11192
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3804 7478 3832 11183
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4080 10606 4108 11086
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3896 8022 3924 8774
rect 4080 8294 4108 10542
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 4252 10464 4304 10470
rect 4356 10441 4384 10474
rect 4252 10406 4304 10412
rect 4342 10432 4398 10441
rect 4264 10062 4292 10406
rect 4342 10367 4398 10376
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4172 9178 4200 9590
rect 4264 9178 4292 9998
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4356 8566 4384 8978
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3896 7342 3924 7958
rect 4356 7954 4384 8366
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 3884 7336 3936 7342
rect 3698 7304 3754 7313
rect 3884 7278 3936 7284
rect 3698 7239 3754 7248
rect 3712 6458 3740 7239
rect 3976 7200 4028 7206
rect 3896 7160 3976 7188
rect 3896 6662 3924 7160
rect 3976 7142 4028 7148
rect 4080 7018 4108 7414
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 3988 6990 4108 7018
rect 3988 6798 4016 6990
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3238 5264 3294 5273
rect 3238 5199 3294 5208
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 3528 4154 3556 5850
rect 3700 5636 3752 5642
rect 3700 5578 3752 5584
rect 3712 5166 3740 5578
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3804 5234 3832 5510
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3620 4282 3648 5102
rect 3712 4690 3740 5102
rect 3804 4826 3832 5170
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 2884 4126 3004 4154
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 110 3632 166 3641
rect 110 3567 166 3576
rect 124 3466 152 3567
rect 112 3460 164 3466
rect 112 3402 164 3408
rect 2148 3058 2176 3674
rect 2240 3398 2268 4126
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 112 2916 164 2922
rect 112 2858 164 2864
rect 124 2553 152 2858
rect 110 2544 166 2553
rect 110 2479 166 2488
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 1688 1057 1716 2246
rect 1674 1048 1730 1057
rect 1674 983 1730 992
rect 846 96 902 480
rect 2240 82 2268 3334
rect 2320 3120 2372 3126
rect 2320 3062 2372 3068
rect 2332 2378 2360 3062
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2516 2514 2544 2994
rect 2608 2990 2636 4126
rect 2976 3670 3004 4126
rect 3344 4126 3556 4154
rect 2964 3664 3016 3670
rect 2778 3632 2834 3641
rect 2964 3606 3016 3612
rect 2778 3567 2834 3576
rect 3056 3596 3108 3602
rect 2792 3058 2820 3567
rect 3056 3538 3108 3544
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 3068 2854 3096 3538
rect 3344 3126 3372 4126
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2320 2372 2372 2378
rect 2320 2314 2372 2320
rect 3068 2009 3096 2790
rect 3620 2582 3648 4218
rect 3896 4154 3924 6598
rect 3988 6118 4016 6734
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3804 4126 3924 4154
rect 3804 3398 3832 4126
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3896 2990 3924 3878
rect 3988 3194 4016 6054
rect 4080 5846 4108 6666
rect 4264 6662 4292 7278
rect 4356 7206 4384 7890
rect 4448 7750 4476 13654
rect 4622 13084 4918 13104
rect 4678 13082 4702 13084
rect 4758 13082 4782 13084
rect 4838 13082 4862 13084
rect 4700 13030 4702 13082
rect 4764 13030 4776 13082
rect 4838 13030 4840 13082
rect 4678 13028 4702 13030
rect 4758 13028 4782 13030
rect 4838 13028 4862 13030
rect 4622 13008 4918 13028
rect 5184 12986 5212 14282
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4540 11626 4568 12038
rect 4622 11996 4918 12016
rect 4678 11994 4702 11996
rect 4758 11994 4782 11996
rect 4838 11994 4862 11996
rect 4700 11942 4702 11994
rect 4764 11942 4776 11994
rect 4838 11942 4840 11994
rect 4678 11940 4702 11942
rect 4758 11940 4782 11942
rect 4838 11940 4862 11942
rect 4622 11920 4918 11940
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4528 11620 4580 11626
rect 4528 11562 4580 11568
rect 4540 9994 4568 11562
rect 5000 11082 5028 11698
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 4622 10908 4918 10928
rect 4678 10906 4702 10908
rect 4758 10906 4782 10908
rect 4838 10906 4862 10908
rect 4700 10854 4702 10906
rect 4764 10854 4776 10906
rect 4838 10854 4840 10906
rect 4678 10852 4702 10854
rect 4758 10852 4782 10854
rect 4838 10852 4862 10854
rect 4622 10832 4918 10852
rect 5000 10198 5028 11018
rect 5092 10470 5120 11290
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4622 9820 4918 9840
rect 4678 9818 4702 9820
rect 4758 9818 4782 9820
rect 4838 9818 4862 9820
rect 4700 9766 4702 9818
rect 4764 9766 4776 9818
rect 4838 9766 4840 9818
rect 4678 9764 4702 9766
rect 4758 9764 4782 9766
rect 4838 9764 4862 9766
rect 4622 9744 4918 9764
rect 5092 9450 5120 10406
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5184 9450 5212 9862
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4540 8838 4568 9046
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4540 8430 4568 8774
rect 4622 8732 4918 8752
rect 4678 8730 4702 8732
rect 4758 8730 4782 8732
rect 4838 8730 4862 8732
rect 4700 8678 4702 8730
rect 4764 8678 4776 8730
rect 4838 8678 4840 8730
rect 4678 8676 4702 8678
rect 4758 8676 4782 8678
rect 4838 8676 4862 8678
rect 4622 8656 4918 8676
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7410 4476 7686
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4448 6798 4476 7346
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4264 5914 4292 6598
rect 4448 6186 4476 6734
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4080 4078 4108 5782
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4448 5370 4476 5646
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4252 5296 4304 5302
rect 4304 5256 4384 5284
rect 4252 5238 4304 5244
rect 4356 5166 4384 5256
rect 4344 5160 4396 5166
rect 4344 5102 4396 5108
rect 4540 4826 4568 8366
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 4622 7644 4918 7664
rect 4678 7642 4702 7644
rect 4758 7642 4782 7644
rect 4838 7642 4862 7644
rect 4700 7590 4702 7642
rect 4764 7590 4776 7642
rect 4838 7590 4840 7642
rect 4678 7588 4702 7590
rect 4758 7588 4782 7590
rect 4838 7588 4862 7590
rect 4622 7568 4918 7588
rect 5000 7324 5028 7754
rect 5092 7478 5120 7890
rect 5276 7750 5304 15558
rect 5368 15162 5396 15914
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5368 13462 5396 15098
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5368 10538 5396 11154
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5368 10266 5396 10474
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5460 9382 5488 16526
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5552 13326 5580 15438
rect 5644 13841 5672 19110
rect 5724 17740 5776 17746
rect 5724 17682 5776 17688
rect 5736 17649 5764 17682
rect 5722 17640 5778 17649
rect 5722 17575 5778 17584
rect 5736 16998 5764 17575
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 5736 15910 5764 16662
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5630 13832 5686 13841
rect 5630 13767 5686 13776
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 12918 5580 13262
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5644 10810 5672 13767
rect 6012 13462 6040 19178
rect 6288 18834 6316 19246
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6104 18154 6132 18770
rect 6288 18290 6316 18770
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6276 18284 6328 18290
rect 6276 18226 6328 18232
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 6288 17746 6316 18226
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6000 13456 6052 13462
rect 6000 13398 6052 13404
rect 6196 12968 6224 17478
rect 6288 17338 6316 17682
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 6288 16794 6316 17002
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6380 16250 6408 18702
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6472 15706 6500 17614
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 13297 6500 14758
rect 6564 14482 6592 18906
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6656 16590 6684 17274
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6656 15638 6684 15846
rect 6644 15632 6696 15638
rect 6644 15574 6696 15580
rect 6656 15026 6684 15574
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6656 14550 6684 14962
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6564 13530 6592 14418
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6458 13288 6514 13297
rect 6458 13223 6514 13232
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6196 12940 6316 12968
rect 6090 12880 6146 12889
rect 6090 12815 6146 12824
rect 6104 12782 6132 12815
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6104 12481 6132 12718
rect 6090 12472 6146 12481
rect 6090 12407 6146 12416
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6012 11898 6040 12242
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5920 10674 5948 10950
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5736 9926 5764 9998
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5828 9722 5856 10134
rect 5920 9994 5948 10474
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5368 8956 5396 9318
rect 5446 9208 5502 9217
rect 5446 9143 5502 9152
rect 5460 9110 5488 9143
rect 5828 9110 5856 9658
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5368 8928 5580 8956
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 7886 5488 8774
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 5000 7296 5120 7324
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 4622 6556 4918 6576
rect 4678 6554 4702 6556
rect 4758 6554 4782 6556
rect 4838 6554 4862 6556
rect 4700 6502 4702 6554
rect 4764 6502 4776 6554
rect 4838 6502 4840 6554
rect 4678 6500 4702 6502
rect 4758 6500 4782 6502
rect 4838 6500 4862 6502
rect 4622 6480 4918 6500
rect 5000 6361 5028 6938
rect 5092 6730 5120 7296
rect 5184 7002 5212 7686
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 4986 6352 5042 6361
rect 4986 6287 5042 6296
rect 5184 6254 5212 6938
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5368 6322 5396 6802
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 4622 5468 4918 5488
rect 4678 5466 4702 5468
rect 4758 5466 4782 5468
rect 4838 5466 4862 5468
rect 4700 5414 4702 5466
rect 4764 5414 4776 5466
rect 4838 5414 4840 5466
rect 4678 5412 4702 5414
rect 4758 5412 4782 5414
rect 4838 5412 4862 5414
rect 4622 5392 4918 5412
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4172 4593 4200 4626
rect 4158 4584 4214 4593
rect 4158 4519 4214 4528
rect 4356 4282 4384 4626
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4252 4140 4304 4146
rect 4304 4100 4384 4128
rect 4252 4082 4304 4088
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4080 3738 4108 4014
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3712 2650 3740 2926
rect 3976 2916 4028 2922
rect 4080 2904 4108 3130
rect 4264 3058 4292 3946
rect 4356 3602 4384 4100
rect 4540 4078 4568 4762
rect 5000 4690 5028 6122
rect 5184 5778 5212 6190
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5184 5352 5212 5714
rect 5264 5704 5316 5710
rect 5368 5692 5396 6258
rect 5460 5914 5488 7822
rect 5552 7041 5580 8928
rect 5828 8634 5856 9046
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5920 7478 5948 8026
rect 5908 7472 5960 7478
rect 5630 7440 5686 7449
rect 5908 7414 5960 7420
rect 5630 7375 5686 7384
rect 5644 7342 5672 7375
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5538 7032 5594 7041
rect 5538 6967 5594 6976
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5316 5664 5396 5692
rect 5264 5646 5316 5652
rect 5092 5324 5212 5352
rect 5092 5030 5120 5324
rect 5172 5228 5224 5234
rect 5276 5216 5304 5646
rect 5224 5188 5304 5216
rect 5172 5170 5224 5176
rect 5276 5030 5304 5188
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5276 4690 5304 4966
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 4622 4380 4918 4400
rect 4678 4378 4702 4380
rect 4758 4378 4782 4380
rect 4838 4378 4862 4380
rect 4700 4326 4702 4378
rect 4764 4326 4776 4378
rect 4838 4326 4840 4378
rect 4678 4324 4702 4326
rect 4758 4324 4782 4326
rect 4838 4324 4862 4326
rect 4622 4304 4918 4324
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4448 3398 4476 3946
rect 5000 3942 5028 4626
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4526 3768 4582 3777
rect 4526 3703 4582 3712
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4028 2876 4108 2904
rect 3976 2858 4028 2864
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3608 2576 3660 2582
rect 3608 2518 3660 2524
rect 3712 2378 3740 2586
rect 4540 2514 4568 3703
rect 5000 3584 5028 3878
rect 5092 3738 5120 4626
rect 5170 4584 5226 4593
rect 5170 4519 5226 4528
rect 5264 4548 5316 4554
rect 5184 4486 5212 4519
rect 5264 4490 5316 4496
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5184 4078 5212 4422
rect 5276 4214 5304 4490
rect 5460 4486 5488 5714
rect 5552 5710 5580 6967
rect 5920 6934 5948 7414
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5736 6458 5764 6802
rect 5920 6458 5948 6870
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6012 5234 6040 5510
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5276 3942 5304 4014
rect 5460 3942 5488 4150
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5080 3596 5132 3602
rect 5000 3556 5080 3584
rect 5080 3538 5132 3544
rect 4622 3292 4918 3312
rect 4678 3290 4702 3292
rect 4758 3290 4782 3292
rect 4838 3290 4862 3292
rect 4700 3238 4702 3290
rect 4764 3238 4776 3290
rect 4838 3238 4840 3290
rect 4678 3236 4702 3238
rect 4758 3236 4782 3238
rect 4838 3236 4862 3238
rect 4622 3216 4918 3236
rect 5092 3126 5120 3538
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 5092 2854 5120 3062
rect 5460 2990 5488 3878
rect 5552 3602 5580 4014
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 4724 2582 4752 2790
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 5092 2496 5120 2790
rect 5552 2514 5580 3538
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5644 2990 5672 3470
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5644 2582 5672 2926
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 5722 2544 5778 2553
rect 5172 2508 5224 2514
rect 5092 2468 5172 2496
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 4540 2106 4568 2314
rect 5092 2310 5120 2468
rect 5172 2450 5224 2456
rect 5540 2508 5592 2514
rect 5828 2514 5856 3878
rect 6012 2961 6040 5170
rect 5998 2952 6054 2961
rect 5998 2887 6054 2896
rect 5722 2479 5778 2488
rect 5816 2508 5868 2514
rect 5540 2450 5592 2456
rect 5356 2372 5408 2378
rect 5356 2314 5408 2320
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 4622 2204 4918 2224
rect 4678 2202 4702 2204
rect 4758 2202 4782 2204
rect 4838 2202 4862 2204
rect 4700 2150 4702 2202
rect 4764 2150 4776 2202
rect 4838 2150 4840 2202
rect 4678 2148 4702 2150
rect 4758 2148 4782 2150
rect 4838 2148 4862 2150
rect 4622 2128 4918 2148
rect 4528 2100 4580 2106
rect 4528 2042 4580 2048
rect 3054 2000 3110 2009
rect 3054 1935 3110 1944
rect 2594 82 2650 480
rect 2240 54 2650 82
rect 846 0 902 40
rect 2594 0 2650 54
rect 4434 82 4490 480
rect 4540 82 4568 2042
rect 5092 1737 5120 2246
rect 5368 2106 5396 2314
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 5552 2009 5580 2450
rect 5736 2446 5764 2479
rect 5816 2450 5868 2456
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5828 2378 5856 2450
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5538 2000 5594 2009
rect 5538 1935 5594 1944
rect 5078 1728 5134 1737
rect 5078 1663 5134 1672
rect 4434 54 4568 82
rect 6104 82 6132 9318
rect 6288 8498 6316 12940
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 9926 6408 11494
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9722 6408 9862
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6472 7342 6500 12854
rect 6564 11150 6592 13126
rect 6656 12714 6684 13670
rect 6644 12708 6696 12714
rect 6644 12650 6696 12656
rect 6656 12442 6684 12650
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6656 11898 6684 12378
rect 6748 12306 6776 18022
rect 6840 17542 6868 18158
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6840 13814 6868 17478
rect 6932 17202 6960 19110
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7576 17882 7604 18770
rect 7656 18148 7708 18154
rect 7656 18090 7708 18096
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7576 17610 7604 17818
rect 7564 17604 7616 17610
rect 7564 17546 7616 17552
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6932 16794 6960 17138
rect 7392 17066 7420 17478
rect 7668 17202 7696 18090
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7656 16720 7708 16726
rect 7656 16662 7708 16668
rect 7484 16250 7512 16662
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7392 15026 7420 15370
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7484 14890 7512 15302
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7208 14074 7236 14554
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 6840 13786 6960 13814
rect 7208 13802 7236 14010
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6840 12850 6868 13398
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6656 10810 6684 11222
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6656 8294 6684 9046
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7857 6684 8230
rect 6642 7848 6698 7857
rect 6642 7783 6698 7792
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6564 6769 6592 7142
rect 6656 6866 6684 7142
rect 6748 6934 6776 9454
rect 6840 9178 6868 11086
rect 6932 11082 6960 13786
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7300 12986 7328 13398
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7300 12442 7328 12922
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7208 11762 7236 12106
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7300 11626 7328 12378
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7300 11354 7328 11562
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6932 10169 6960 11018
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 6918 10160 6974 10169
rect 6918 10095 6974 10104
rect 6932 10062 6960 10095
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6932 9518 6960 9998
rect 7300 9926 7328 10610
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 7274 6960 8774
rect 7024 8090 7052 8910
rect 7300 8537 7328 9862
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7392 8634 7420 9454
rect 7668 9081 7696 16662
rect 7760 15570 7788 21542
rect 9770 21542 9904 21570
rect 9770 21520 9826 21542
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 7840 18828 7892 18834
rect 7840 18770 7892 18776
rect 7852 18426 7880 18770
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7852 18222 7880 18362
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 8128 17746 8156 18294
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 7944 16522 7972 17002
rect 8128 16998 8156 17682
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 8128 16726 8156 16934
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 7932 16516 7984 16522
rect 7932 16458 7984 16464
rect 7748 15564 7800 15570
rect 7748 15506 7800 15512
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 13938 7788 14214
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7852 11762 7880 15370
rect 7944 15094 7972 16458
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 8036 13938 8064 16526
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8128 14074 8156 14418
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 8036 13258 8064 13874
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8128 13326 8156 13806
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 8128 12986 8156 13262
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 8128 11898 8156 12310
rect 8220 12238 8248 19110
rect 8289 19068 8585 19088
rect 8345 19066 8369 19068
rect 8425 19066 8449 19068
rect 8505 19066 8529 19068
rect 8367 19014 8369 19066
rect 8431 19014 8443 19066
rect 8505 19014 8507 19066
rect 8345 19012 8369 19014
rect 8425 19012 8449 19014
rect 8505 19012 8529 19014
rect 8289 18992 8585 19012
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8289 17980 8585 18000
rect 8345 17978 8369 17980
rect 8425 17978 8449 17980
rect 8505 17978 8529 17980
rect 8367 17926 8369 17978
rect 8431 17926 8443 17978
rect 8505 17926 8507 17978
rect 8345 17924 8369 17926
rect 8425 17924 8449 17926
rect 8505 17924 8529 17926
rect 8289 17904 8585 17924
rect 8576 17740 8628 17746
rect 8680 17728 8708 18022
rect 8628 17700 8708 17728
rect 8576 17682 8628 17688
rect 8588 17134 8616 17682
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 8576 17128 8628 17134
rect 8628 17088 8708 17116
rect 8576 17070 8628 17076
rect 8289 16892 8585 16912
rect 8345 16890 8369 16892
rect 8425 16890 8449 16892
rect 8505 16890 8529 16892
rect 8367 16838 8369 16890
rect 8431 16838 8443 16890
rect 8505 16838 8507 16890
rect 8345 16836 8369 16838
rect 8425 16836 8449 16838
rect 8505 16836 8529 16838
rect 8289 16816 8585 16836
rect 8680 16794 8708 17088
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8772 16658 8800 17614
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8404 16250 8432 16526
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8289 15804 8585 15824
rect 8345 15802 8369 15804
rect 8425 15802 8449 15804
rect 8505 15802 8529 15804
rect 8367 15750 8369 15802
rect 8431 15750 8443 15802
rect 8505 15750 8507 15802
rect 8345 15748 8369 15750
rect 8425 15748 8449 15750
rect 8505 15748 8529 15750
rect 8289 15728 8585 15748
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 15162 8340 15506
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8289 14716 8585 14736
rect 8345 14714 8369 14716
rect 8425 14714 8449 14716
rect 8505 14714 8529 14716
rect 8367 14662 8369 14714
rect 8431 14662 8443 14714
rect 8505 14662 8507 14714
rect 8345 14660 8369 14662
rect 8425 14660 8449 14662
rect 8505 14660 8529 14662
rect 8289 14640 8585 14660
rect 8680 14346 8708 16390
rect 8956 15026 8984 18566
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 9048 16454 9076 17070
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 9048 15026 9076 15370
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8772 14618 8800 14826
rect 8956 14618 8984 14962
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8850 14376 8906 14385
rect 8668 14340 8720 14346
rect 8850 14311 8906 14320
rect 8668 14282 8720 14288
rect 8289 13628 8585 13648
rect 8345 13626 8369 13628
rect 8425 13626 8449 13628
rect 8505 13626 8529 13628
rect 8367 13574 8369 13626
rect 8431 13574 8443 13626
rect 8505 13574 8507 13626
rect 8345 13572 8369 13574
rect 8425 13572 8449 13574
rect 8505 13572 8529 13574
rect 8289 13552 8585 13572
rect 8289 12540 8585 12560
rect 8345 12538 8369 12540
rect 8425 12538 8449 12540
rect 8505 12538 8529 12540
rect 8367 12486 8369 12538
rect 8431 12486 8443 12538
rect 8505 12486 8507 12538
rect 8345 12484 8369 12486
rect 8425 12484 8449 12486
rect 8505 12484 8529 12486
rect 8289 12464 8585 12484
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 11898 8248 12174
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 11354 7880 11698
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 8128 11286 8156 11834
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 8128 10810 8156 11222
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7944 10198 7972 10406
rect 7932 10192 7984 10198
rect 7932 10134 7984 10140
rect 7944 9178 7972 10134
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8036 9586 8064 9998
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8036 9489 8064 9522
rect 8022 9480 8078 9489
rect 8022 9415 8078 9424
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7654 9072 7710 9081
rect 7654 9007 7710 9016
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7286 8528 7342 8537
rect 7286 8463 7342 8472
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 7024 6769 7052 7210
rect 7116 7177 7144 8230
rect 7208 7818 7236 8298
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7102 7168 7158 7177
rect 7102 7103 7158 7112
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 6550 6760 6606 6769
rect 6550 6695 6606 6704
rect 7010 6760 7066 6769
rect 7010 6695 7066 6704
rect 6564 6662 6592 6695
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6380 4758 6408 5510
rect 6472 5030 6500 5714
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 4865 6500 4966
rect 6458 4856 6514 4865
rect 6458 4791 6514 4800
rect 6368 4752 6420 4758
rect 6366 4720 6368 4729
rect 6420 4720 6422 4729
rect 6184 4684 6236 4690
rect 6366 4655 6422 4664
rect 6184 4626 6236 4632
rect 6380 4629 6408 4655
rect 6196 4486 6224 4626
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6196 3398 6224 4422
rect 6380 3942 6408 4490
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6472 3505 6500 4791
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6458 3496 6514 3505
rect 6276 3460 6328 3466
rect 6564 3466 6592 4626
rect 6656 4282 6684 6122
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6656 4078 6684 4218
rect 6644 4072 6696 4078
rect 6748 4049 6776 5510
rect 6840 5370 6868 6598
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6644 4014 6696 4020
rect 6734 4040 6790 4049
rect 6734 3975 6790 3984
rect 6840 3602 6868 5034
rect 6932 4622 6960 6598
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6932 4185 6960 4558
rect 6918 4176 6974 4185
rect 6918 4111 6974 4120
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6458 3431 6514 3440
rect 6552 3460 6604 3466
rect 6276 3402 6328 3408
rect 6552 3402 6604 3408
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6196 1601 6224 3334
rect 6288 2854 6316 3402
rect 6564 3097 6592 3402
rect 6656 3194 6684 3538
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6550 3088 6606 3097
rect 6550 3023 6552 3032
rect 6604 3023 6606 3032
rect 6552 2994 6604 3000
rect 6564 2963 6592 2994
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6182 1592 6238 1601
rect 6182 1527 6238 1536
rect 6472 1465 6500 2382
rect 6458 1456 6514 1465
rect 6458 1391 6514 1400
rect 6656 1329 6684 3130
rect 6840 2922 6868 3538
rect 7024 3058 7052 5510
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 6828 2916 6880 2922
rect 6828 2858 6880 2864
rect 7024 2446 7052 2994
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7116 2378 7144 6870
rect 7392 6322 7420 8570
rect 7576 7886 7604 8842
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7668 7886 7696 8434
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7576 7274 7604 7822
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7576 6730 7604 7210
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7470 6352 7526 6361
rect 7380 6316 7432 6322
rect 7470 6287 7526 6296
rect 7380 6258 7432 6264
rect 7196 6248 7248 6254
rect 7194 6216 7196 6225
rect 7248 6216 7250 6225
rect 7194 6151 7250 6160
rect 7208 3670 7236 6151
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7300 4146 7328 5102
rect 7484 4826 7512 6287
rect 7562 5400 7618 5409
rect 7562 5335 7618 5344
rect 7576 5302 7604 5335
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7484 4282 7512 4762
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7576 3738 7604 4218
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7576 2922 7604 3674
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7288 2508 7340 2514
rect 7564 2508 7616 2514
rect 7340 2468 7564 2496
rect 7288 2450 7340 2456
rect 7564 2450 7616 2456
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7668 2310 7696 7686
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7760 7002 7788 7210
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7852 6254 7880 7278
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7944 5846 7972 6802
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8036 6186 8064 6394
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8036 5846 8064 6122
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7852 4826 7880 5646
rect 7840 4820 7892 4826
rect 7760 4780 7840 4808
rect 7760 2990 7788 4780
rect 7840 4762 7892 4768
rect 7840 4684 7892 4690
rect 7944 4672 7972 5782
rect 8036 5370 8064 5782
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8036 5098 8064 5306
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8128 4758 8156 9658
rect 8220 8566 8248 11630
rect 8289 11452 8585 11472
rect 8345 11450 8369 11452
rect 8425 11450 8449 11452
rect 8505 11450 8529 11452
rect 8367 11398 8369 11450
rect 8431 11398 8443 11450
rect 8505 11398 8507 11450
rect 8345 11396 8369 11398
rect 8425 11396 8449 11398
rect 8505 11396 8529 11398
rect 8289 11376 8585 11396
rect 8289 10364 8585 10384
rect 8345 10362 8369 10364
rect 8425 10362 8449 10364
rect 8505 10362 8529 10364
rect 8367 10310 8369 10362
rect 8431 10310 8443 10362
rect 8505 10310 8507 10362
rect 8345 10308 8369 10310
rect 8425 10308 8449 10310
rect 8505 10308 8529 10310
rect 8289 10288 8585 10308
rect 8680 9722 8708 14282
rect 8864 13734 8892 14311
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8850 13288 8906 13297
rect 8760 13252 8812 13258
rect 8850 13223 8906 13232
rect 8760 13194 8812 13200
rect 8772 12374 8800 13194
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 8758 12200 8814 12209
rect 8758 12135 8814 12144
rect 8772 11150 8800 12135
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8864 10742 8892 13223
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8289 9276 8585 9296
rect 8345 9274 8369 9276
rect 8425 9274 8449 9276
rect 8505 9274 8529 9276
rect 8367 9222 8369 9274
rect 8431 9222 8443 9274
rect 8505 9222 8507 9274
rect 8345 9220 8369 9222
rect 8425 9220 8449 9222
rect 8505 9220 8529 9222
rect 8289 9200 8585 9220
rect 8680 9178 8708 9522
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8864 9042 8892 10678
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 9048 9926 9076 10542
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9625 9076 9862
rect 9034 9616 9090 9625
rect 9232 9586 9260 19110
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9416 17814 9444 18158
rect 9692 18086 9720 18770
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9416 17270 9444 17750
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 9312 17060 9364 17066
rect 9312 17002 9364 17008
rect 9324 15570 9352 17002
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9508 13938 9536 17818
rect 9692 16017 9720 18022
rect 9784 16114 9812 18090
rect 9876 16250 9904 21542
rect 11716 21542 12034 21570
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9968 16998 9996 17682
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9678 16008 9734 16017
rect 9588 15972 9640 15978
rect 9678 15943 9734 15952
rect 9588 15914 9640 15920
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9600 13814 9628 15914
rect 9692 15609 9720 15943
rect 9864 15904 9916 15910
rect 9968 15892 9996 16730
rect 10060 16522 10088 17546
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 9916 15864 9996 15892
rect 9864 15846 9916 15852
rect 9876 15706 9904 15846
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9678 15600 9734 15609
rect 9678 15535 9734 15544
rect 9876 15162 9904 15642
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 10060 14618 10088 15506
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10152 13870 10180 17546
rect 9508 13786 9628 13814
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 9680 13796 9732 13802
rect 9508 13734 9536 13786
rect 9680 13738 9732 13744
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9034 9551 9090 9560
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 8864 8634 8892 8978
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8289 8188 8585 8208
rect 8345 8186 8369 8188
rect 8425 8186 8449 8188
rect 8505 8186 8529 8188
rect 8367 8134 8369 8186
rect 8431 8134 8443 8186
rect 8505 8134 8507 8186
rect 8345 8132 8369 8134
rect 8425 8132 8449 8134
rect 8505 8132 8529 8134
rect 8289 8112 8585 8132
rect 8484 8016 8536 8022
rect 8680 7993 8708 8366
rect 8484 7958 8536 7964
rect 8666 7984 8722 7993
rect 8496 7750 8524 7958
rect 8666 7919 8722 7928
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8496 7274 8524 7686
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 8680 7177 8708 7278
rect 8666 7168 8722 7177
rect 8289 7100 8585 7120
rect 8666 7103 8722 7112
rect 8345 7098 8369 7100
rect 8425 7098 8449 7100
rect 8505 7098 8529 7100
rect 8367 7046 8369 7098
rect 8431 7046 8443 7098
rect 8505 7046 8507 7098
rect 8345 7044 8369 7046
rect 8425 7044 8449 7046
rect 8505 7044 8529 7046
rect 8289 7024 8585 7044
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8680 6254 8708 6598
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8772 6089 8800 6870
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8758 6080 8814 6089
rect 8289 6012 8585 6032
rect 8758 6015 8814 6024
rect 8345 6010 8369 6012
rect 8425 6010 8449 6012
rect 8505 6010 8529 6012
rect 8367 5958 8369 6010
rect 8431 5958 8443 6010
rect 8505 5958 8507 6010
rect 8345 5956 8369 5958
rect 8425 5956 8449 5958
rect 8505 5956 8529 5958
rect 8289 5936 8585 5956
rect 8289 4924 8585 4944
rect 8345 4922 8369 4924
rect 8425 4922 8449 4924
rect 8505 4922 8529 4924
rect 8367 4870 8369 4922
rect 8431 4870 8443 4922
rect 8505 4870 8507 4922
rect 8345 4868 8369 4870
rect 8425 4868 8449 4870
rect 8505 4868 8529 4870
rect 8289 4848 8585 4868
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8024 4684 8076 4690
rect 7944 4644 8024 4672
rect 7840 4626 7892 4632
rect 8024 4626 8076 4632
rect 7852 3534 7880 4626
rect 8220 4146 8248 4694
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8128 2990 8156 4014
rect 8289 3836 8585 3856
rect 8345 3834 8369 3836
rect 8425 3834 8449 3836
rect 8505 3834 8529 3836
rect 8367 3782 8369 3834
rect 8431 3782 8443 3834
rect 8505 3782 8507 3834
rect 8345 3780 8369 3782
rect 8425 3780 8449 3782
rect 8505 3780 8529 3782
rect 8289 3760 8585 3780
rect 8680 3738 8708 4558
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8220 3126 8248 3606
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8680 3058 8708 3674
rect 8772 3194 8800 3946
rect 8864 3466 8892 6598
rect 8956 5846 8984 8774
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9048 7546 9076 7686
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8956 4826 8984 5102
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 9048 3380 9076 7210
rect 9140 4706 9168 7754
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9232 7313 9260 7346
rect 9324 7342 9352 13466
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9416 12102 9444 12718
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9416 11529 9444 12038
rect 9508 11694 9536 13670
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9600 12918 9628 13330
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9692 12646 9720 13738
rect 10336 13161 10364 19110
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10612 17882 10640 18022
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10612 17202 10640 17818
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10600 17060 10652 17066
rect 10600 17002 10652 17008
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10416 16176 10468 16182
rect 10416 16118 10468 16124
rect 10322 13152 10378 13161
rect 10244 13110 10322 13138
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12374 9720 12582
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9692 11558 9720 12310
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9680 11552 9732 11558
rect 9402 11520 9458 11529
rect 9680 11494 9732 11500
rect 9402 11455 9458 11464
rect 9692 10538 9720 11494
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9692 10146 9720 10474
rect 9600 10130 9720 10146
rect 9588 10124 9720 10130
rect 9640 10118 9720 10124
rect 9588 10066 9640 10072
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9508 9042 9536 9998
rect 9692 9654 9720 10118
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9692 9450 9720 9590
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 9110 9628 9318
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9508 8945 9536 8978
rect 9494 8936 9550 8945
rect 9494 8871 9550 8880
rect 9600 8634 9628 9046
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9586 8392 9642 8401
rect 9692 8362 9720 9386
rect 9784 8974 9812 11834
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9876 10198 9904 10610
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9586 8327 9642 8336
rect 9680 8356 9732 8362
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9312 7336 9364 7342
rect 9218 7304 9274 7313
rect 9312 7278 9364 7284
rect 9218 7239 9274 7248
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9232 4826 9260 6734
rect 9312 6248 9364 6254
rect 9416 6225 9444 7142
rect 9508 7002 9536 7346
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9312 6190 9364 6196
rect 9402 6216 9458 6225
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9140 4678 9260 4706
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9140 3641 9168 4558
rect 9126 3632 9182 3641
rect 9126 3567 9182 3576
rect 9128 3392 9180 3398
rect 9048 3352 9128 3380
rect 9128 3334 9180 3340
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8772 2922 8800 3130
rect 9232 3058 9260 4678
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 8289 2748 8585 2768
rect 8345 2746 8369 2748
rect 8425 2746 8449 2748
rect 8505 2746 8529 2748
rect 8367 2694 8369 2746
rect 8431 2694 8443 2746
rect 8505 2694 8507 2746
rect 8345 2692 8369 2694
rect 8425 2692 8449 2694
rect 8505 2692 8529 2694
rect 8289 2672 8585 2692
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 8036 2038 8064 2246
rect 8024 2032 8076 2038
rect 8024 1974 8076 1980
rect 6642 1320 6698 1329
rect 6642 1255 6698 1264
rect 6274 82 6330 480
rect 6104 54 6330 82
rect 4434 0 4490 54
rect 6274 0 6330 54
rect 8114 82 8170 480
rect 8220 82 8248 2586
rect 8680 2417 8708 2790
rect 9232 2650 9260 2790
rect 9324 2650 9352 6190
rect 9402 6151 9458 6160
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9416 5914 9444 6054
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9416 4826 9444 5306
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9416 4282 9444 4762
rect 9600 4622 9628 8327
rect 9680 8298 9732 8304
rect 9692 7954 9720 8298
rect 9784 8022 9812 8910
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 7546 9720 7890
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9784 7478 9812 7822
rect 10244 7546 10272 13110
rect 10322 13087 10378 13096
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10336 11626 10364 12582
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10336 11354 10364 11562
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10336 10810 10364 11290
rect 10428 11286 10456 16118
rect 10520 14532 10548 16934
rect 10612 16794 10640 17002
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10612 15162 10640 15846
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10612 14822 10640 15098
rect 10704 15094 10732 18158
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10888 17066 10916 18022
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10876 17060 10928 17066
rect 10876 17002 10928 17008
rect 10888 15094 10916 17002
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10704 14634 10732 15030
rect 10704 14606 10916 14634
rect 10784 14544 10836 14550
rect 10520 14504 10640 14532
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10520 13297 10548 14214
rect 10506 13288 10562 13297
rect 10506 13223 10562 13232
rect 10508 11620 10560 11626
rect 10508 11562 10560 11568
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10428 10266 10456 11222
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10520 10033 10548 11562
rect 10612 11558 10640 14504
rect 10784 14486 10836 14492
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10704 14006 10732 14350
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10796 13938 10824 14486
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10888 13870 10916 14606
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10876 13456 10928 13462
rect 10876 13398 10928 13404
rect 10888 12986 10916 13398
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10888 12442 10916 12922
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10980 12170 11008 17478
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 11072 13326 11100 14486
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 10968 12164 11020 12170
rect 10968 12106 11020 12112
rect 11072 11762 11100 13262
rect 11164 12374 11192 19110
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11440 18086 11468 18770
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 11348 16998 11376 17682
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11256 16250 11284 16594
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11242 15600 11298 15609
rect 11348 15586 11376 16934
rect 11532 16590 11560 16934
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11532 15910 11560 16526
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11298 15558 11376 15586
rect 11242 15535 11298 15544
rect 11256 13734 11284 15535
rect 11532 14822 11560 15846
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11624 15026 11652 15302
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11256 12782 11284 13670
rect 11532 13530 11560 14758
rect 11624 13734 11652 14962
rect 11716 14278 11744 21542
rect 11978 21520 12034 21542
rect 14186 21570 14242 22000
rect 16394 21570 16450 22000
rect 18602 21570 18658 22000
rect 20810 21570 20866 22000
rect 14186 21542 14320 21570
rect 14186 21520 14242 21542
rect 11956 19612 12252 19632
rect 12012 19610 12036 19612
rect 12092 19610 12116 19612
rect 12172 19610 12196 19612
rect 12034 19558 12036 19610
rect 12098 19558 12110 19610
rect 12172 19558 12174 19610
rect 12012 19556 12036 19558
rect 12092 19556 12116 19558
rect 12172 19556 12196 19558
rect 11956 19536 12252 19556
rect 11956 18524 12252 18544
rect 12012 18522 12036 18524
rect 12092 18522 12116 18524
rect 12172 18522 12196 18524
rect 12034 18470 12036 18522
rect 12098 18470 12110 18522
rect 12172 18470 12174 18522
rect 12012 18468 12036 18470
rect 12092 18468 12116 18470
rect 12172 18468 12196 18470
rect 11956 18448 12252 18468
rect 14292 18426 14320 21542
rect 16040 21542 16450 21570
rect 15622 19068 15918 19088
rect 15678 19066 15702 19068
rect 15758 19066 15782 19068
rect 15838 19066 15862 19068
rect 15700 19014 15702 19066
rect 15764 19014 15776 19066
rect 15838 19014 15840 19066
rect 15678 19012 15702 19014
rect 15758 19012 15782 19014
rect 15838 19012 15862 19014
rect 15622 18992 15918 19012
rect 16040 18426 16068 21542
rect 16394 21520 16450 21542
rect 18340 21542 18658 21570
rect 17866 19000 17922 19009
rect 17866 18935 17922 18944
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 11956 17436 12252 17456
rect 12012 17434 12036 17436
rect 12092 17434 12116 17436
rect 12172 17434 12196 17436
rect 12034 17382 12036 17434
rect 12098 17382 12110 17434
rect 12172 17382 12174 17434
rect 12012 17380 12036 17382
rect 12092 17380 12116 17382
rect 12172 17380 12196 17382
rect 11956 17360 12252 17380
rect 12360 17338 12388 17682
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11808 16250 11836 16594
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 11956 16348 12252 16368
rect 12012 16346 12036 16348
rect 12092 16346 12116 16348
rect 12172 16346 12196 16348
rect 12034 16294 12036 16346
rect 12098 16294 12110 16346
rect 12172 16294 12174 16346
rect 12012 16292 12036 16294
rect 12092 16292 12116 16294
rect 12172 16292 12196 16294
rect 11956 16272 12252 16292
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11808 15162 11836 15642
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11900 14618 11928 15438
rect 11956 15260 12252 15280
rect 12012 15258 12036 15260
rect 12092 15258 12116 15260
rect 12172 15258 12196 15260
rect 12034 15206 12036 15258
rect 12098 15206 12110 15258
rect 12172 15206 12174 15258
rect 12012 15204 12036 15206
rect 12092 15204 12116 15206
rect 12172 15204 12196 15206
rect 11956 15184 12252 15204
rect 12360 15094 12388 15438
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 12360 14346 12388 14894
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 13841 11744 14214
rect 11956 14172 12252 14192
rect 12012 14170 12036 14172
rect 12092 14170 12116 14172
rect 12172 14170 12196 14172
rect 12034 14118 12036 14170
rect 12098 14118 12110 14170
rect 12172 14118 12174 14170
rect 12012 14116 12036 14118
rect 12092 14116 12116 14118
rect 12172 14116 12196 14118
rect 11956 14096 12252 14116
rect 11702 13832 11758 13841
rect 11702 13767 11758 13776
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 12452 13530 12480 16458
rect 12544 14618 12572 17478
rect 13464 17338 13492 17682
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12636 16794 12664 17070
rect 13452 17060 13504 17066
rect 13452 17002 13504 17008
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12636 16454 12664 16730
rect 13268 16720 13320 16726
rect 13268 16662 13320 16668
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 13188 15706 13216 16526
rect 13280 15978 13308 16662
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13280 15638 13308 15914
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13280 14890 13308 15574
rect 13372 15026 13400 15982
rect 13464 15570 13492 17002
rect 13648 16114 13676 18158
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 15622 17980 15918 18000
rect 15678 17978 15702 17980
rect 15758 17978 15782 17980
rect 15838 17978 15862 17980
rect 15700 17926 15702 17978
rect 15764 17926 15776 17978
rect 15838 17926 15840 17978
rect 15678 17924 15702 17926
rect 15758 17924 15782 17926
rect 15838 17924 15862 17926
rect 15622 17904 15918 17924
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14568 16794 14596 17002
rect 15304 16998 15332 17682
rect 15948 17338 15976 18022
rect 16868 17814 16896 18158
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13464 15162 13492 15506
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13268 14884 13320 14890
rect 13268 14826 13320 14832
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12544 13938 12572 14554
rect 13280 14550 13308 14826
rect 14108 14618 14136 15302
rect 14292 15162 14320 15846
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14292 14890 14320 15098
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 13268 14544 13320 14550
rect 13188 14504 13268 14532
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12728 13530 12756 14350
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12820 13734 12848 13874
rect 13188 13802 13216 14504
rect 13268 14486 13320 14492
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13176 13796 13228 13802
rect 13176 13738 13228 13744
rect 13648 13734 13676 14214
rect 14108 13938 14136 14554
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11440 12374 11468 13194
rect 11956 13084 12252 13104
rect 12012 13082 12036 13084
rect 12092 13082 12116 13084
rect 12172 13082 12196 13084
rect 12034 13030 12036 13082
rect 12098 13030 12110 13082
rect 12172 13030 12174 13082
rect 12012 13028 12036 13030
rect 12092 13028 12116 13030
rect 12172 13028 12196 13030
rect 11956 13008 12252 13028
rect 12452 12918 12480 13466
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11164 11830 11192 12310
rect 11900 12306 11928 12854
rect 12820 12850 12848 13670
rect 13740 13462 13768 13738
rect 14200 13705 14228 13738
rect 14186 13696 14242 13705
rect 14186 13631 14242 13640
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12912 12986 12940 13262
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12636 12442 12664 12650
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11256 11830 11284 12174
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11244 11824 11296 11830
rect 11900 11801 11928 12242
rect 11956 11996 12252 12016
rect 12012 11994 12036 11996
rect 12092 11994 12116 11996
rect 12172 11994 12196 11996
rect 12034 11942 12036 11994
rect 12098 11942 12110 11994
rect 12172 11942 12174 11994
rect 12012 11940 12036 11942
rect 12092 11940 12116 11942
rect 12172 11940 12196 11942
rect 11956 11920 12252 11940
rect 11244 11766 11296 11772
rect 11886 11792 11942 11801
rect 11060 11756 11112 11762
rect 11886 11727 11888 11736
rect 11060 11698 11112 11704
rect 11940 11727 11942 11736
rect 11888 11698 11940 11704
rect 11900 11667 11928 11698
rect 12348 11688 12400 11694
rect 11334 11656 11390 11665
rect 12348 11630 12400 11636
rect 11334 11591 11390 11600
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10784 10532 10836 10538
rect 10784 10474 10836 10480
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10796 10198 10824 10474
rect 10888 10266 10916 10474
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10506 10024 10562 10033
rect 10506 9959 10562 9968
rect 10796 9110 10824 10134
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10784 9104 10836 9110
rect 10888 9081 10916 9454
rect 11348 9110 11376 11591
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11520 11076 11572 11082
rect 11520 11018 11572 11024
rect 11532 10062 11560 11018
rect 11808 10810 11836 11222
rect 11956 10908 12252 10928
rect 12012 10906 12036 10908
rect 12092 10906 12116 10908
rect 12172 10906 12196 10908
rect 12034 10854 12036 10906
rect 12098 10854 12110 10906
rect 12172 10854 12174 10906
rect 12012 10852 12036 10854
rect 12092 10852 12116 10854
rect 12172 10852 12196 10854
rect 11956 10832 12252 10852
rect 11796 10804 11848 10810
rect 11716 10764 11796 10792
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11624 10198 11652 10406
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11532 9586 11560 9998
rect 11624 9722 11652 10134
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11716 9654 11744 10764
rect 11796 10746 11848 10752
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11808 10198 11836 10610
rect 12360 10577 12388 11630
rect 12820 11354 12848 12786
rect 13740 12646 13768 13398
rect 14292 13258 14320 13874
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 13832 12986 13860 13126
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 14108 12850 14136 13126
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14200 12714 14228 12922
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13464 12238 13492 12582
rect 13740 12374 13768 12582
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13740 12102 13768 12310
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 13280 11286 13308 11494
rect 13464 11354 13492 11630
rect 13740 11626 13768 12038
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 14384 11286 14412 11494
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12346 10568 12402 10577
rect 12346 10503 12402 10512
rect 12452 10266 12480 11086
rect 13280 10470 13308 11222
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13372 10674 13400 10950
rect 13464 10742 13492 11086
rect 14476 11082 14504 15846
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11808 10062 11836 10134
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 13464 9926 13492 10406
rect 14384 10198 14412 10950
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 14462 10160 14518 10169
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 11956 9820 12252 9840
rect 12012 9818 12036 9820
rect 12092 9818 12116 9820
rect 12172 9818 12196 9820
rect 12034 9766 12036 9818
rect 12098 9766 12110 9818
rect 12172 9766 12174 9818
rect 12012 9764 12036 9766
rect 12092 9764 12116 9766
rect 12172 9764 12196 9766
rect 11956 9744 12252 9764
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11520 9580 11572 9586
rect 11572 9540 11652 9568
rect 11520 9522 11572 9528
rect 11336 9104 11388 9110
rect 10784 9046 10836 9052
rect 10874 9072 10930 9081
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8344 10732 8774
rect 10796 8498 10824 9046
rect 11336 9046 11388 9052
rect 10874 9007 10930 9016
rect 10888 8974 10916 9007
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10784 8356 10836 8362
rect 10704 8316 10784 8344
rect 10784 8298 10836 8304
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 6798 9812 7142
rect 10060 7002 10088 7210
rect 10048 6996 10100 7002
rect 9968 6956 10048 6984
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9680 5908 9732 5914
rect 9784 5896 9812 6734
rect 9876 6118 9904 6870
rect 9968 6390 9996 6956
rect 10048 6938 10100 6944
rect 10612 6934 10640 7210
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9732 5868 9812 5896
rect 9680 5850 9732 5856
rect 9968 5846 9996 6326
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10060 5914 10088 6122
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 9968 5370 9996 5782
rect 10152 5710 10180 6258
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9876 4758 9904 4966
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9876 4282 9904 4694
rect 10152 4622 10180 5646
rect 10612 5302 10640 6870
rect 10796 6662 10824 8298
rect 10888 7818 10916 8298
rect 11348 8022 11376 9046
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11348 6934 11376 7754
rect 11440 7274 11468 7890
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11532 7410 11560 7686
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11428 7268 11480 7274
rect 11428 7210 11480 7216
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11426 6896 11482 6905
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 11348 6458 11376 6870
rect 11426 6831 11482 6840
rect 11440 6798 11468 6831
rect 11624 6798 11652 9540
rect 11716 9110 11744 9590
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11716 8634 11744 9046
rect 11956 8732 12252 8752
rect 12012 8730 12036 8732
rect 12092 8730 12116 8732
rect 12172 8730 12196 8732
rect 12034 8678 12036 8730
rect 12098 8678 12110 8730
rect 12172 8678 12174 8730
rect 12012 8676 12036 8678
rect 12092 8676 12116 8678
rect 12172 8676 12196 8678
rect 11956 8656 12252 8676
rect 12622 8664 12678 8673
rect 11704 8628 11756 8634
rect 12728 8634 12756 9386
rect 12912 9178 12940 9454
rect 13464 9450 13492 9862
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13556 9110 13584 9998
rect 13832 9722 13860 10134
rect 14462 10095 14518 10104
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 14384 9110 14412 9998
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 12622 8599 12678 8608
rect 12716 8628 12768 8634
rect 11704 8570 11756 8576
rect 11956 7644 12252 7664
rect 12012 7642 12036 7644
rect 12092 7642 12116 7644
rect 12172 7642 12196 7644
rect 12034 7590 12036 7642
rect 12098 7590 12110 7642
rect 12172 7590 12174 7642
rect 12012 7588 12036 7590
rect 12092 7588 12116 7590
rect 12172 7588 12196 7590
rect 11956 7568 12252 7588
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11242 5808 11298 5817
rect 11440 5778 11468 6734
rect 11956 6556 12252 6576
rect 12012 6554 12036 6556
rect 12092 6554 12116 6556
rect 12172 6554 12196 6556
rect 12034 6502 12036 6554
rect 12098 6502 12110 6554
rect 12172 6502 12174 6554
rect 12012 6500 12036 6502
rect 12092 6500 12116 6502
rect 12172 6500 12196 6502
rect 11956 6480 12252 6500
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12452 5914 12480 6190
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 11242 5743 11298 5752
rect 11428 5772 11480 5778
rect 11256 5642 11284 5743
rect 11428 5714 11480 5720
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10600 5296 10652 5302
rect 11072 5273 11100 5510
rect 11256 5370 11284 5578
rect 11956 5468 12252 5488
rect 12012 5466 12036 5468
rect 12092 5466 12116 5468
rect 12172 5466 12196 5468
rect 12034 5414 12036 5466
rect 12098 5414 12110 5466
rect 12172 5414 12174 5466
rect 12012 5412 12036 5414
rect 12092 5412 12116 5414
rect 12172 5412 12196 5414
rect 11956 5392 12252 5412
rect 12544 5370 12572 5646
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 10600 5238 10652 5244
rect 11058 5264 11114 5273
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9416 2689 9444 3470
rect 9402 2680 9458 2689
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9312 2644 9364 2650
rect 9402 2615 9458 2624
rect 9312 2586 9364 2592
rect 9508 2582 9536 3878
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9876 3194 9904 3606
rect 10152 3534 10180 4558
rect 10612 4214 10640 5238
rect 10692 5228 10744 5234
rect 11058 5199 11114 5208
rect 10692 5170 10744 5176
rect 10704 4826 10732 5170
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 11072 4282 11100 4490
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10244 3738 10272 3946
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10428 3466 10456 4082
rect 11256 4049 11284 4422
rect 11348 4214 11376 4694
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11716 4214 11744 4558
rect 11956 4380 12252 4400
rect 12012 4378 12036 4380
rect 12092 4378 12116 4380
rect 12172 4378 12196 4380
rect 12034 4326 12036 4378
rect 12098 4326 12110 4378
rect 12172 4326 12174 4378
rect 12012 4324 12036 4326
rect 12092 4324 12116 4326
rect 12172 4324 12196 4326
rect 11956 4304 12252 4324
rect 11336 4208 11388 4214
rect 11336 4150 11388 4156
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 12360 4146 12388 4626
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 11242 4040 11298 4049
rect 11242 3975 11298 3984
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10612 2990 10640 3334
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 11164 2650 11192 3470
rect 11956 3292 12252 3312
rect 12012 3290 12036 3292
rect 12092 3290 12116 3292
rect 12172 3290 12196 3292
rect 12034 3238 12036 3290
rect 12098 3238 12110 3290
rect 12172 3238 12174 3290
rect 12012 3236 12036 3238
rect 12092 3236 12116 3238
rect 12172 3236 12196 3238
rect 11956 3216 12252 3236
rect 12452 2650 12480 3674
rect 12636 3505 12664 8599
rect 12716 8570 12768 8576
rect 12728 8362 12756 8570
rect 13556 8566 13584 9046
rect 13832 8634 13860 9046
rect 14476 9042 14504 10095
rect 14568 9382 14596 14418
rect 14752 14278 14780 14962
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 13802 14780 14214
rect 14936 13870 14964 16594
rect 15304 15026 15332 16934
rect 15622 16892 15918 16912
rect 15678 16890 15702 16892
rect 15758 16890 15782 16892
rect 15838 16890 15862 16892
rect 15700 16838 15702 16890
rect 15764 16838 15776 16890
rect 15838 16838 15840 16890
rect 15678 16836 15702 16838
rect 15758 16836 15782 16838
rect 15838 16836 15862 16838
rect 15622 16816 15918 16836
rect 15948 15910 15976 17274
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16132 15910 16160 16594
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16302 16144 16358 16153
rect 16302 16079 16358 16088
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 15622 15804 15918 15824
rect 15678 15802 15702 15804
rect 15758 15802 15782 15804
rect 15838 15802 15862 15804
rect 15700 15750 15702 15802
rect 15764 15750 15776 15802
rect 15838 15750 15840 15802
rect 15678 15748 15702 15750
rect 15758 15748 15782 15750
rect 15838 15748 15862 15750
rect 15622 15728 15918 15748
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15396 15094 15424 15438
rect 15488 15162 15516 15574
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15672 15026 15700 15438
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 15028 14074 15056 14214
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14740 13796 14792 13802
rect 14792 13756 14872 13784
rect 14740 13738 14792 13744
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14660 13530 14688 13670
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14660 12238 14688 13262
rect 14844 12918 14872 13756
rect 14936 13734 14964 13806
rect 14924 13728 14976 13734
rect 15120 13705 15148 14486
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 14924 13670 14976 13676
rect 15106 13696 15162 13705
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14660 10169 14688 11494
rect 14844 10266 14872 12038
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14646 10160 14702 10169
rect 14936 10146 14964 13670
rect 15106 13631 15162 13640
rect 15120 13462 15148 13631
rect 15108 13456 15160 13462
rect 15108 13398 15160 13404
rect 15212 12209 15240 14214
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15198 12200 15254 12209
rect 15198 12135 15254 12144
rect 15198 11928 15254 11937
rect 15304 11898 15332 14010
rect 15488 13870 15516 14758
rect 15622 14716 15918 14736
rect 15678 14714 15702 14716
rect 15758 14714 15782 14716
rect 15838 14714 15862 14716
rect 15700 14662 15702 14714
rect 15764 14662 15776 14714
rect 15838 14662 15840 14714
rect 15678 14660 15702 14662
rect 15758 14660 15782 14662
rect 15838 14660 15862 14662
rect 15622 14640 15918 14660
rect 15476 13864 15528 13870
rect 15752 13864 15804 13870
rect 15528 13824 15752 13852
rect 15476 13806 15528 13812
rect 15752 13806 15804 13812
rect 15622 13628 15918 13648
rect 15678 13626 15702 13628
rect 15758 13626 15782 13628
rect 15838 13626 15862 13628
rect 15700 13574 15702 13626
rect 15764 13574 15776 13626
rect 15838 13574 15840 13626
rect 15678 13572 15702 13574
rect 15758 13572 15782 13574
rect 15838 13572 15862 13574
rect 15622 13552 15918 13572
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15488 12986 15516 13398
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15488 12374 15516 12582
rect 15622 12540 15918 12560
rect 15678 12538 15702 12540
rect 15758 12538 15782 12540
rect 15838 12538 15862 12540
rect 15700 12486 15702 12538
rect 15764 12486 15776 12538
rect 15838 12486 15840 12538
rect 15678 12484 15702 12486
rect 15758 12484 15782 12486
rect 15838 12484 15862 12486
rect 15622 12464 15918 12484
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15488 11898 15516 12310
rect 15198 11863 15254 11872
rect 15292 11892 15344 11898
rect 15212 11694 15240 11863
rect 15292 11834 15344 11840
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15108 11552 15160 11558
rect 15028 11529 15108 11540
rect 15014 11520 15108 11529
rect 15070 11512 15108 11520
rect 15108 11494 15160 11500
rect 15014 11455 15070 11464
rect 15016 11280 15068 11286
rect 15016 11222 15068 11228
rect 15028 10266 15056 11222
rect 15304 11082 15332 11698
rect 15396 11150 15424 11698
rect 15622 11452 15918 11472
rect 15678 11450 15702 11452
rect 15758 11450 15782 11452
rect 15838 11450 15862 11452
rect 15700 11398 15702 11450
rect 15764 11398 15776 11450
rect 15838 11398 15840 11450
rect 15678 11396 15702 11398
rect 15758 11396 15782 11398
rect 15838 11396 15862 11398
rect 15622 11376 15918 11396
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15212 10538 15240 10950
rect 15396 10810 15424 11086
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15108 10192 15160 10198
rect 14936 10118 15056 10146
rect 15108 10134 15160 10140
rect 14646 10095 14702 10104
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14752 9586 14780 9862
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14844 9450 14872 9658
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12728 8022 12756 8298
rect 13832 8090 13860 8570
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12728 7002 12756 7822
rect 13280 7546 13308 7958
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12728 6730 12756 6938
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 13280 6458 13308 7482
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13832 7002 13860 7346
rect 13924 7274 13952 7958
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13634 6624 13690 6633
rect 13634 6559 13690 6568
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12728 5846 12756 6054
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12728 5302 12756 5782
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 12716 5296 12768 5302
rect 12716 5238 12768 5244
rect 12728 4758 12756 5238
rect 13004 5098 13032 5714
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 12900 4752 12952 4758
rect 13004 4740 13032 5034
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12952 4712 13032 4740
rect 12900 4694 12952 4700
rect 12728 4282 12756 4694
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 13096 3738 13124 4762
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13556 4146 13584 4422
rect 13648 4154 13676 6559
rect 13740 6458 13768 6870
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13832 6390 13860 6734
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13832 5778 13860 6326
rect 14200 6118 14228 8230
rect 14292 7206 14320 8842
rect 14372 8288 14424 8294
rect 14476 8276 14504 8978
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 8634 14780 8774
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14936 8498 14964 9590
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14424 8248 14504 8276
rect 14556 8288 14608 8294
rect 14372 8230 14424 8236
rect 14556 8230 14608 8236
rect 14568 7954 14596 8230
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14660 7274 14688 8434
rect 14740 8356 14792 8362
rect 14740 8298 14792 8304
rect 14752 8090 14780 8298
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14936 7410 14964 8434
rect 15028 8378 15056 10118
rect 15120 9110 15148 10134
rect 15212 9654 15240 10474
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 15028 8350 15148 8378
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14830 7304 14886 7313
rect 14648 7268 14700 7274
rect 15028 7290 15056 7686
rect 14830 7239 14886 7248
rect 14936 7262 15056 7290
rect 14648 7210 14700 7216
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14292 6497 14320 7142
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14278 6488 14334 6497
rect 14278 6423 14334 6432
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14292 5778 14320 6258
rect 14384 6186 14412 6394
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13832 4826 13860 5034
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 14016 4622 14044 5306
rect 14476 5098 14504 6666
rect 14568 6361 14596 7142
rect 14844 6361 14872 7239
rect 14554 6352 14610 6361
rect 14554 6287 14610 6296
rect 14830 6352 14886 6361
rect 14830 6287 14886 6296
rect 14844 6118 14872 6287
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14384 4282 14412 4966
rect 14568 4282 14596 6054
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 13544 4140 13596 4146
rect 13648 4126 13768 4154
rect 13544 4082 13596 4088
rect 13740 4010 13768 4126
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13452 3528 13504 3534
rect 12622 3496 12678 3505
rect 13452 3470 13504 3476
rect 12622 3431 12678 3440
rect 12530 3088 12586 3097
rect 12530 3023 12586 3032
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 10152 2514 10180 2586
rect 12544 2553 12572 3023
rect 12636 2582 12664 3431
rect 13464 3194 13492 3470
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12728 2650 12756 2790
rect 13280 2650 13308 2926
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 12624 2576 12676 2582
rect 12530 2544 12586 2553
rect 10140 2508 10192 2514
rect 12624 2518 12676 2524
rect 12530 2479 12586 2488
rect 10140 2450 10192 2456
rect 13636 2440 13688 2446
rect 8666 2408 8722 2417
rect 13740 2428 13768 3946
rect 13924 3942 13952 4218
rect 14660 4214 14688 4762
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13924 3670 13952 3878
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 13924 2990 13952 3606
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 14200 2446 14228 2994
rect 14660 2922 14688 3334
rect 14648 2916 14700 2922
rect 14648 2858 14700 2864
rect 14660 2650 14688 2858
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 13688 2400 13768 2428
rect 13636 2382 13688 2388
rect 8666 2343 8722 2352
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 8114 54 8248 82
rect 9954 82 10010 480
rect 10060 82 10088 2314
rect 11956 2204 12252 2224
rect 12012 2202 12036 2204
rect 12092 2202 12116 2204
rect 12172 2202 12196 2204
rect 12034 2150 12036 2202
rect 12098 2150 12110 2202
rect 12172 2150 12174 2202
rect 12012 2148 12036 2150
rect 12092 2148 12116 2150
rect 12172 2148 12196 2150
rect 11956 2128 12252 2148
rect 12072 1964 12124 1970
rect 12072 1906 12124 1912
rect 9954 54 10088 82
rect 11794 82 11850 480
rect 12084 82 12112 1906
rect 11794 54 12112 82
rect 13634 82 13690 480
rect 13740 82 13768 2400
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14844 2310 14872 2450
rect 14936 2446 14964 7262
rect 15016 6860 15068 6866
rect 15120 6848 15148 8350
rect 15488 8072 15516 10406
rect 15622 10364 15918 10384
rect 15678 10362 15702 10364
rect 15758 10362 15782 10364
rect 15838 10362 15862 10364
rect 15700 10310 15702 10362
rect 15764 10310 15776 10362
rect 15838 10310 15840 10362
rect 15678 10308 15702 10310
rect 15758 10308 15782 10310
rect 15838 10308 15862 10310
rect 15622 10288 15918 10308
rect 15622 9276 15918 9296
rect 15678 9274 15702 9276
rect 15758 9274 15782 9276
rect 15838 9274 15862 9276
rect 15700 9222 15702 9274
rect 15764 9222 15776 9274
rect 15838 9222 15840 9274
rect 15678 9220 15702 9222
rect 15758 9220 15782 9222
rect 15838 9220 15862 9222
rect 15622 9200 15918 9220
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15672 8498 15700 8978
rect 15948 8906 15976 15846
rect 16028 15088 16080 15094
rect 16028 15030 16080 15036
rect 16040 14550 16068 15030
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 16040 13326 16068 14486
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16040 12374 16068 13262
rect 16132 12889 16160 15846
rect 16118 12880 16174 12889
rect 16118 12815 16174 12824
rect 16132 12714 16160 12815
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 16028 12368 16080 12374
rect 16028 12310 16080 12316
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 16040 11150 16068 11562
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16040 10538 16068 11086
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 16040 10198 16068 10474
rect 16132 10470 16160 11154
rect 16316 10792 16344 16079
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16408 12374 16436 12786
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16500 11218 16528 16186
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16316 10764 16436 10792
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16132 10198 16160 10406
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16132 9042 16160 9386
rect 16224 9042 16252 9454
rect 16316 9382 16344 10610
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15936 8492 15988 8498
rect 16212 8492 16264 8498
rect 15936 8434 15988 8440
rect 16132 8452 16212 8480
rect 15672 8401 15700 8434
rect 15658 8392 15714 8401
rect 15658 8327 15714 8336
rect 15622 8188 15918 8208
rect 15678 8186 15702 8188
rect 15758 8186 15782 8188
rect 15838 8186 15862 8188
rect 15700 8134 15702 8186
rect 15764 8134 15776 8186
rect 15838 8134 15840 8186
rect 15678 8132 15702 8134
rect 15758 8132 15782 8134
rect 15838 8132 15862 8134
rect 15622 8112 15918 8132
rect 15488 8044 15608 8072
rect 15200 7880 15252 7886
rect 15476 7880 15528 7886
rect 15396 7857 15476 7868
rect 15200 7822 15252 7828
rect 15382 7848 15476 7857
rect 15212 6934 15240 7822
rect 15292 7812 15344 7818
rect 15438 7840 15476 7848
rect 15476 7822 15528 7828
rect 15382 7783 15438 7792
rect 15292 7754 15344 7760
rect 15304 7177 15332 7754
rect 15580 7750 15608 8044
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15764 7342 15792 7686
rect 15948 7342 15976 8434
rect 16028 7472 16080 7478
rect 16028 7414 16080 7420
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15290 7168 15346 7177
rect 15290 7103 15346 7112
rect 15622 7100 15918 7120
rect 15678 7098 15702 7100
rect 15758 7098 15782 7100
rect 15838 7098 15862 7100
rect 15700 7046 15702 7098
rect 15764 7046 15776 7098
rect 15838 7046 15840 7098
rect 15678 7044 15702 7046
rect 15758 7044 15782 7046
rect 15838 7044 15862 7046
rect 15622 7024 15918 7044
rect 15200 6928 15252 6934
rect 15200 6870 15252 6876
rect 15948 6866 15976 7278
rect 15068 6820 15148 6848
rect 15016 6802 15068 6808
rect 15120 6254 15148 6820
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15948 6458 15976 6802
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15396 6276 15700 6304
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15120 5778 15148 6190
rect 15396 6089 15424 6276
rect 15672 6186 15700 6276
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15382 6080 15438 6089
rect 15382 6015 15438 6024
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15200 5636 15252 5642
rect 15200 5578 15252 5584
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 15028 3602 15056 3946
rect 15120 3942 15148 4694
rect 15212 4690 15240 5578
rect 15396 5370 15424 5782
rect 15488 5710 15516 6122
rect 16040 6118 16068 7414
rect 16132 6338 16160 8452
rect 16212 8434 16264 8440
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16224 7993 16252 8230
rect 16304 8016 16356 8022
rect 16210 7984 16266 7993
rect 16304 7958 16356 7964
rect 16210 7919 16266 7928
rect 16316 7546 16344 7958
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16408 7410 16436 10764
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16592 9217 16620 10406
rect 16684 10130 16712 16390
rect 16868 14958 16896 17750
rect 17590 16008 17646 16017
rect 17590 15943 17646 15952
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16960 14822 16988 15506
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 16960 14385 16988 14758
rect 16946 14376 17002 14385
rect 16946 14311 17002 14320
rect 17052 13190 17080 14758
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17144 14006 17172 14214
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 17144 12782 17172 13806
rect 17328 13734 17356 14418
rect 17408 13796 17460 13802
rect 17408 13738 17460 13744
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17236 12646 17264 13330
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 12306 17264 12582
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17144 11937 17172 12242
rect 17130 11928 17186 11937
rect 17130 11863 17186 11872
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 16960 10266 16988 10678
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16578 9208 16634 9217
rect 16578 9143 16634 9152
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16500 8480 16528 8910
rect 16580 8832 16632 8838
rect 16684 8820 16712 10066
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16632 8792 16712 8820
rect 16580 8774 16632 8780
rect 16500 8452 16620 8480
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16500 7750 16528 8298
rect 16592 7954 16620 8452
rect 16776 8022 16804 8978
rect 16960 8945 16988 9114
rect 16946 8936 17002 8945
rect 16946 8871 17002 8880
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16868 8090 16896 8774
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16764 8016 16816 8022
rect 16764 7958 16816 7964
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16408 6798 16436 7346
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16210 6352 16266 6361
rect 16132 6310 16210 6338
rect 16210 6287 16266 6296
rect 16224 6254 16252 6287
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 15622 6012 15918 6032
rect 15678 6010 15702 6012
rect 15758 6010 15782 6012
rect 15838 6010 15862 6012
rect 15700 5958 15702 6010
rect 15764 5958 15776 6010
rect 15838 5958 15840 6010
rect 15678 5956 15702 5958
rect 15758 5956 15782 5958
rect 15838 5956 15862 5958
rect 15622 5936 15918 5956
rect 16132 5846 16160 6190
rect 16120 5840 16172 5846
rect 16120 5782 16172 5788
rect 16304 5840 16356 5846
rect 16304 5782 16356 5788
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15488 5216 15516 5646
rect 15764 5302 15792 5646
rect 15752 5296 15804 5302
rect 15752 5238 15804 5244
rect 15304 5188 15516 5216
rect 15936 5228 15988 5234
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15304 3942 15332 5188
rect 15936 5170 15988 5176
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15488 4729 15516 4966
rect 15622 4924 15918 4944
rect 15678 4922 15702 4924
rect 15758 4922 15782 4924
rect 15838 4922 15862 4924
rect 15700 4870 15702 4922
rect 15764 4870 15776 4922
rect 15838 4870 15840 4922
rect 15678 4868 15702 4870
rect 15758 4868 15782 4870
rect 15838 4868 15862 4870
rect 15622 4848 15918 4868
rect 15474 4720 15530 4729
rect 15384 4684 15436 4690
rect 15474 4655 15530 4664
rect 15384 4626 15436 4632
rect 15396 4282 15424 4626
rect 15948 4593 15976 5170
rect 16120 5092 16172 5098
rect 16120 5034 16172 5040
rect 15934 4584 15990 4593
rect 15934 4519 15990 4528
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 16132 4010 16160 5034
rect 16316 4690 16344 5782
rect 16500 5778 16528 7686
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16592 6633 16620 7278
rect 16684 7206 16712 7890
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16672 7200 16724 7206
rect 16776 7177 16804 7210
rect 16856 7200 16908 7206
rect 16672 7142 16724 7148
rect 16762 7168 16818 7177
rect 16684 6769 16712 7142
rect 16856 7142 16908 7148
rect 16762 7103 16818 7112
rect 16868 7002 16896 7142
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16960 6882 16988 8434
rect 17052 8362 17080 11630
rect 17144 11626 17172 11863
rect 17236 11694 17264 12242
rect 17328 11801 17356 13670
rect 17420 13394 17448 13738
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17420 12850 17448 13330
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 12374 17448 12582
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17420 11830 17448 12174
rect 17408 11824 17460 11830
rect 17314 11792 17370 11801
rect 17408 11766 17460 11772
rect 17314 11727 17370 11736
rect 17224 11688 17276 11694
rect 17328 11676 17356 11727
rect 17328 11648 17448 11676
rect 17224 11630 17276 11636
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17328 10674 17356 11154
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17144 8673 17172 10542
rect 17328 10130 17356 10610
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 9722 17356 10066
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17328 9518 17356 9658
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 9042 17356 9318
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17130 8664 17186 8673
rect 17130 8599 17186 8608
rect 17040 8356 17092 8362
rect 17144 8344 17172 8599
rect 17328 8430 17356 8978
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17224 8356 17276 8362
rect 17144 8316 17224 8344
rect 17040 8298 17092 8304
rect 17224 8298 17276 8304
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 16868 6866 16988 6882
rect 17144 6866 17172 7142
rect 16856 6860 16988 6866
rect 16908 6854 16988 6860
rect 17132 6860 17184 6866
rect 16856 6802 16908 6808
rect 17132 6802 17184 6808
rect 16670 6760 16726 6769
rect 16670 6695 16726 6704
rect 16578 6624 16634 6633
rect 16578 6559 16634 6568
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16592 5234 16620 6559
rect 16868 6458 16896 6802
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16960 6458 16988 6734
rect 17040 6724 17092 6730
rect 17040 6666 17092 6672
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17052 6322 17080 6666
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17144 6186 17172 6802
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17144 5370 17172 5714
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16302 4176 16358 4185
rect 16592 4162 16620 4422
rect 16684 4282 16712 4626
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16592 4134 16712 4162
rect 17236 4154 17264 7958
rect 17316 6792 17368 6798
rect 17420 6780 17448 11648
rect 17512 6905 17540 13126
rect 17604 10033 17632 15943
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17788 13841 17816 14418
rect 17774 13832 17830 13841
rect 17774 13767 17776 13776
rect 17828 13767 17830 13776
rect 17776 13738 17828 13744
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17590 10024 17646 10033
rect 17590 9959 17646 9968
rect 17696 9042 17724 12718
rect 17880 11898 17908 18935
rect 18340 18426 18368 21542
rect 18602 21520 18658 21542
rect 20456 21542 20866 21570
rect 19289 19612 19585 19632
rect 19345 19610 19369 19612
rect 19425 19610 19449 19612
rect 19505 19610 19529 19612
rect 19367 19558 19369 19610
rect 19431 19558 19443 19610
rect 19505 19558 19507 19610
rect 19345 19556 19369 19558
rect 19425 19556 19449 19558
rect 19505 19556 19529 19558
rect 19289 19536 19585 19556
rect 19289 18524 19585 18544
rect 19345 18522 19369 18524
rect 19425 18522 19449 18524
rect 19505 18522 19529 18524
rect 19367 18470 19369 18522
rect 19431 18470 19443 18522
rect 19505 18470 19507 18522
rect 19345 18468 19369 18470
rect 19425 18468 19449 18470
rect 19505 18468 19529 18470
rect 19289 18448 19585 18468
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 20456 17882 20484 21542
rect 20810 21520 20866 21542
rect 21546 21176 21602 21185
rect 21546 21111 21602 21120
rect 21560 18970 21588 21111
rect 21548 18964 21600 18970
rect 21548 18906 21600 18912
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 19289 17436 19585 17456
rect 19345 17434 19369 17436
rect 19425 17434 19449 17436
rect 19505 17434 19529 17436
rect 19367 17382 19369 17434
rect 19431 17382 19443 17434
rect 19505 17382 19507 17434
rect 19345 17380 19369 17382
rect 19425 17380 19449 17382
rect 19505 17380 19529 17382
rect 19289 17360 19585 17380
rect 19246 17232 19302 17241
rect 19246 17167 19302 17176
rect 19260 16794 19288 17167
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 18142 16688 18198 16697
rect 18142 16623 18198 16632
rect 19064 16652 19116 16658
rect 18156 13530 18184 16623
rect 19064 16594 19116 16600
rect 19076 15910 19104 16594
rect 19289 16348 19585 16368
rect 19345 16346 19369 16348
rect 19425 16346 19449 16348
rect 19505 16346 19529 16348
rect 19367 16294 19369 16346
rect 19431 16294 19443 16346
rect 19505 16294 19507 16346
rect 19345 16292 19369 16294
rect 19425 16292 19449 16294
rect 19505 16292 19529 16294
rect 19289 16272 19585 16292
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17774 11248 17830 11257
rect 17774 11183 17830 11192
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17788 8498 17816 11183
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17880 9450 17908 10406
rect 17972 10062 18000 10542
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 18064 9518 18092 11494
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18156 9625 18184 10406
rect 18142 9616 18198 9625
rect 18142 9551 18198 9560
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 18064 9110 18092 9454
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18052 9104 18104 9110
rect 18156 9081 18184 9318
rect 18052 9046 18104 9052
rect 18142 9072 18198 9081
rect 18142 9007 18198 9016
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 18248 8090 18276 11562
rect 18432 11558 18460 12242
rect 18524 11694 18552 12650
rect 18616 12306 18644 12786
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18616 11898 18644 12242
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18432 9178 18460 10066
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18524 8537 18552 10202
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18510 8528 18566 8537
rect 18510 8463 18566 8472
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18432 7750 18460 8230
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 17774 7440 17830 7449
rect 17774 7375 17830 7384
rect 17788 7342 17816 7375
rect 18432 7342 18460 7686
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 17498 6896 17554 6905
rect 17498 6831 17554 6840
rect 17420 6752 17540 6780
rect 17316 6734 17368 6740
rect 17328 6225 17356 6734
rect 17314 6216 17370 6225
rect 17314 6151 17370 6160
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17328 5030 17356 5714
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17328 4690 17356 4966
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 16302 4111 16358 4120
rect 15476 4004 15528 4010
rect 15476 3946 15528 3952
rect 15844 4004 15896 4010
rect 16120 4004 16172 4010
rect 15896 3964 15976 3992
rect 15844 3946 15896 3952
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15120 2854 15148 3878
rect 15488 3738 15516 3946
rect 15622 3836 15918 3856
rect 15678 3834 15702 3836
rect 15758 3834 15782 3836
rect 15838 3834 15862 3836
rect 15700 3782 15702 3834
rect 15764 3782 15776 3834
rect 15838 3782 15840 3834
rect 15678 3780 15702 3782
rect 15758 3780 15782 3782
rect 15838 3780 15862 3782
rect 15622 3760 15918 3780
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 14844 1601 14872 2246
rect 15120 2009 15148 2246
rect 15106 2000 15162 2009
rect 15106 1935 15162 1944
rect 15212 1737 15240 2790
rect 15304 2514 15332 3470
rect 15580 3058 15608 3538
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15948 2990 15976 3964
rect 16120 3946 16172 3952
rect 16316 3738 16344 4111
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 15936 2984 15988 2990
rect 16132 2961 16160 2994
rect 16316 2990 16344 3674
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16304 2984 16356 2990
rect 15936 2926 15988 2932
rect 16118 2952 16174 2961
rect 16304 2926 16356 2932
rect 16118 2887 16174 2896
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 15936 2848 15988 2854
rect 16120 2848 16172 2854
rect 15988 2808 16120 2836
rect 15936 2790 15988 2796
rect 16120 2790 16172 2796
rect 15622 2748 15918 2768
rect 15678 2746 15702 2748
rect 15758 2746 15782 2748
rect 15838 2746 15862 2748
rect 15700 2694 15702 2746
rect 15764 2694 15776 2746
rect 15838 2694 15840 2746
rect 15678 2692 15702 2694
rect 15758 2692 15782 2694
rect 15838 2692 15862 2694
rect 15622 2672 15918 2692
rect 16500 2553 16528 2858
rect 16592 2650 16620 3470
rect 16684 2854 16712 4134
rect 17144 4126 17264 4154
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16486 2544 16542 2553
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15752 2508 15804 2514
rect 16776 2514 16804 4014
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16868 3126 16896 3878
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16960 3194 16988 3674
rect 17144 3602 17172 4126
rect 17328 3942 17356 4626
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17328 3602 17356 3878
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17144 3194 17172 3538
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 17328 2990 17356 3538
rect 17420 3466 17448 4966
rect 17512 4146 17540 6752
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17960 5160 18012 5166
rect 18064 5137 18092 6054
rect 17960 5102 18012 5108
rect 18050 5128 18106 5137
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17408 3460 17460 3466
rect 17408 3402 17460 3408
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17512 2650 17540 4082
rect 17972 3097 18000 5102
rect 18050 5063 18106 5072
rect 18328 4208 18380 4214
rect 18328 4150 18380 4156
rect 18052 4072 18104 4078
rect 18236 4072 18288 4078
rect 18104 4032 18236 4060
rect 18052 4014 18104 4020
rect 18236 4014 18288 4020
rect 17958 3088 18014 3097
rect 17958 3023 18014 3032
rect 17776 2984 17828 2990
rect 18248 2961 18276 4014
rect 18340 3233 18368 4150
rect 18326 3224 18382 3233
rect 18326 3159 18382 3168
rect 17776 2926 17828 2932
rect 18234 2952 18290 2961
rect 17788 2854 17816 2926
rect 18234 2887 18290 2896
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 16486 2479 16542 2488
rect 16764 2508 16816 2514
rect 15752 2450 15804 2456
rect 16764 2450 16816 2456
rect 15580 2417 15608 2450
rect 15566 2408 15622 2417
rect 15384 2372 15436 2378
rect 15566 2343 15622 2352
rect 15384 2314 15436 2320
rect 15198 1728 15254 1737
rect 15198 1663 15254 1672
rect 14830 1592 14886 1601
rect 14830 1527 14886 1536
rect 13634 54 13768 82
rect 15396 82 15424 2314
rect 15764 2310 15792 2450
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 15474 82 15530 480
rect 15396 54 15530 82
rect 17236 82 17264 2246
rect 17788 1329 17816 2790
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 18064 2310 18092 2450
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18064 1737 18092 2246
rect 18432 2038 18460 7278
rect 18512 5772 18564 5778
rect 18616 5760 18644 9454
rect 18708 7449 18736 12922
rect 18800 12646 18828 13330
rect 18984 12782 19012 14826
rect 19076 13870 19104 15846
rect 19289 15260 19585 15280
rect 19345 15258 19369 15260
rect 19425 15258 19449 15260
rect 19505 15258 19529 15260
rect 19367 15206 19369 15258
rect 19431 15206 19443 15258
rect 19505 15206 19507 15258
rect 19345 15204 19369 15206
rect 19425 15204 19449 15206
rect 19505 15204 19529 15206
rect 19289 15184 19585 15204
rect 21548 15088 21600 15094
rect 21548 15030 21600 15036
rect 21560 14385 21588 15030
rect 21546 14376 21602 14385
rect 21546 14311 21602 14320
rect 19289 14172 19585 14192
rect 19345 14170 19369 14172
rect 19425 14170 19449 14172
rect 19505 14170 19529 14172
rect 19367 14118 19369 14170
rect 19431 14118 19443 14170
rect 19505 14118 19507 14170
rect 19345 14116 19369 14118
rect 19425 14116 19449 14118
rect 19505 14116 19529 14118
rect 19289 14096 19585 14116
rect 19076 13864 19151 13870
rect 19076 13812 19099 13864
rect 19076 13806 19151 13812
rect 19076 13734 19104 13806
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18800 12102 18828 12582
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18984 11665 19012 12582
rect 18970 11656 19026 11665
rect 18970 11591 19026 11600
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18892 9450 18920 10066
rect 18880 9444 18932 9450
rect 18880 9386 18932 9392
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18892 8276 18920 8978
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18984 8566 19012 8774
rect 18972 8560 19024 8566
rect 19076 8537 19104 13670
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19289 13084 19585 13104
rect 19345 13082 19369 13084
rect 19425 13082 19449 13084
rect 19505 13082 19529 13084
rect 19367 13030 19369 13082
rect 19431 13030 19443 13082
rect 19505 13030 19507 13082
rect 19345 13028 19369 13030
rect 19425 13028 19449 13030
rect 19505 13028 19529 13030
rect 19289 13008 19585 13028
rect 19628 12986 19656 13330
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19289 11996 19585 12016
rect 19345 11994 19369 11996
rect 19425 11994 19449 11996
rect 19505 11994 19529 11996
rect 19367 11942 19369 11994
rect 19431 11942 19443 11994
rect 19505 11942 19507 11994
rect 19345 11940 19369 11942
rect 19425 11940 19449 11942
rect 19505 11940 19529 11942
rect 19289 11920 19585 11940
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 19168 10810 19196 11018
rect 19289 10908 19585 10928
rect 19345 10906 19369 10908
rect 19425 10906 19449 10908
rect 19505 10906 19529 10908
rect 19367 10854 19369 10906
rect 19431 10854 19443 10906
rect 19505 10854 19507 10906
rect 19345 10852 19369 10854
rect 19425 10852 19449 10854
rect 19505 10852 19529 10854
rect 19289 10832 19585 10852
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 19289 9820 19585 9840
rect 19345 9818 19369 9820
rect 19425 9818 19449 9820
rect 19505 9818 19529 9820
rect 19367 9766 19369 9818
rect 19431 9766 19443 9818
rect 19505 9766 19507 9818
rect 19345 9764 19369 9766
rect 19425 9764 19449 9766
rect 19505 9764 19529 9766
rect 19289 9744 19585 9764
rect 19628 9489 19656 10406
rect 19706 10024 19762 10033
rect 19706 9959 19762 9968
rect 19614 9480 19670 9489
rect 19614 9415 19670 9424
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 18972 8502 19024 8508
rect 19062 8528 19118 8537
rect 19062 8463 19118 8472
rect 19168 8362 19196 8978
rect 19289 8732 19585 8752
rect 19345 8730 19369 8732
rect 19425 8730 19449 8732
rect 19505 8730 19529 8732
rect 19367 8678 19369 8730
rect 19431 8678 19443 8730
rect 19505 8678 19507 8730
rect 19345 8676 19369 8678
rect 19425 8676 19449 8678
rect 19505 8676 19529 8678
rect 19289 8656 19585 8676
rect 19156 8356 19208 8362
rect 19076 8316 19156 8344
rect 18972 8288 19024 8294
rect 18892 8248 18972 8276
rect 18972 8230 19024 8236
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18694 7440 18750 7449
rect 18800 7410 18828 7686
rect 18694 7375 18750 7384
rect 18788 7404 18840 7410
rect 18708 6866 18736 7375
rect 18788 7346 18840 7352
rect 18800 7002 18828 7346
rect 18892 7206 18920 7822
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18708 6458 18736 6802
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18564 5732 18644 5760
rect 18512 5714 18564 5720
rect 18524 5030 18552 5714
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18420 2032 18472 2038
rect 18420 1974 18472 1980
rect 18524 1970 18552 4966
rect 18708 4690 18736 6394
rect 18800 5370 18828 6598
rect 18788 5364 18840 5370
rect 18788 5306 18840 5312
rect 18892 5250 18920 7142
rect 18984 5817 19012 8230
rect 18970 5808 19026 5817
rect 19076 5778 19104 8316
rect 19156 8298 19208 8304
rect 19156 7812 19208 7818
rect 19156 7754 19208 7760
rect 19168 7002 19196 7754
rect 19289 7644 19585 7664
rect 19345 7642 19369 7644
rect 19425 7642 19449 7644
rect 19505 7642 19529 7644
rect 19367 7590 19369 7642
rect 19431 7590 19443 7642
rect 19505 7590 19507 7642
rect 19345 7588 19369 7590
rect 19425 7588 19449 7590
rect 19505 7588 19529 7590
rect 19289 7568 19585 7588
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 19720 6866 19748 9959
rect 19812 8430 19840 10746
rect 19904 9518 19932 12582
rect 20074 12200 20130 12209
rect 20074 12135 20130 12144
rect 20088 11898 20116 12135
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20442 11248 20498 11257
rect 20442 11183 20498 11192
rect 20456 11014 20484 11183
rect 20444 11008 20496 11014
rect 20444 10950 20496 10956
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19289 6556 19585 6576
rect 19345 6554 19369 6556
rect 19425 6554 19449 6556
rect 19505 6554 19529 6556
rect 19367 6502 19369 6554
rect 19431 6502 19443 6554
rect 19505 6502 19507 6554
rect 19345 6500 19369 6502
rect 19425 6500 19449 6502
rect 19505 6500 19529 6502
rect 19289 6480 19585 6500
rect 19720 6458 19748 6802
rect 19812 6458 19840 8366
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19812 6254 19840 6394
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 18970 5743 19026 5752
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 19076 5302 19104 5714
rect 19289 5468 19585 5488
rect 19345 5466 19369 5468
rect 19425 5466 19449 5468
rect 19505 5466 19529 5468
rect 19367 5414 19369 5466
rect 19431 5414 19443 5466
rect 19505 5414 19507 5466
rect 19345 5412 19369 5414
rect 19425 5412 19449 5414
rect 19505 5412 19529 5414
rect 19289 5392 19585 5412
rect 18800 5222 18920 5250
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 18696 4684 18748 4690
rect 18696 4626 18748 4632
rect 18800 2650 18828 5222
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 18512 1964 18564 1970
rect 18512 1906 18564 1912
rect 18050 1728 18106 1737
rect 18050 1663 18106 1672
rect 17774 1320 17830 1329
rect 17774 1255 17830 1264
rect 17314 82 17370 480
rect 17236 54 17370 82
rect 18892 82 18920 4422
rect 19168 4282 19196 4626
rect 19289 4380 19585 4400
rect 19345 4378 19369 4380
rect 19425 4378 19449 4380
rect 19505 4378 19529 4380
rect 19367 4326 19369 4378
rect 19431 4326 19443 4378
rect 19505 4326 19507 4378
rect 19345 4324 19369 4326
rect 19425 4324 19449 4326
rect 19505 4324 19529 4326
rect 19289 4304 19585 4324
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 21638 4176 21694 4185
rect 21560 4146 21638 4154
rect 21548 4140 21638 4146
rect 21600 4126 21638 4140
rect 21638 4111 21694 4120
rect 21548 4082 21600 4088
rect 21088 4004 21140 4010
rect 21088 3946 21140 3952
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 19076 2854 19104 3538
rect 19289 3292 19585 3312
rect 19345 3290 19369 3292
rect 19425 3290 19449 3292
rect 19505 3290 19529 3292
rect 19367 3238 19369 3290
rect 19431 3238 19443 3290
rect 19505 3238 19507 3290
rect 19345 3236 19369 3238
rect 19425 3236 19449 3238
rect 19505 3236 19529 3238
rect 19289 3216 19585 3236
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 19076 1465 19104 2790
rect 19289 2204 19585 2224
rect 19345 2202 19369 2204
rect 19425 2202 19449 2204
rect 19505 2202 19529 2204
rect 19367 2150 19369 2202
rect 19431 2150 19443 2202
rect 19505 2150 19507 2202
rect 19345 2148 19369 2150
rect 19425 2148 19449 2150
rect 19505 2148 19529 2150
rect 19289 2128 19585 2148
rect 19062 1456 19118 1465
rect 19062 1391 19118 1400
rect 19154 82 19210 480
rect 18892 54 19210 82
rect 8114 0 8170 54
rect 9954 0 10010 54
rect 11794 0 11850 54
rect 13634 0 13690 54
rect 15474 0 15530 54
rect 17314 0 17370 54
rect 19154 0 19210 54
rect 20994 82 21050 480
rect 21100 82 21128 3946
rect 20994 54 21128 82
rect 20994 0 21050 54
<< via2 >>
rect 1030 21528 1086 21584
rect 18 20304 74 20360
rect 2962 20848 3018 20904
rect 110 19216 166 19272
rect 110 17176 166 17232
rect 110 9832 166 9888
rect 294 16632 350 16688
rect 18 8744 74 8800
rect 1214 17720 1270 17776
rect 1306 17584 1362 17640
rect 1398 14592 1454 14648
rect 1582 16360 1638 16416
rect 2042 15544 2098 15600
rect 4622 19610 4678 19612
rect 4702 19610 4758 19612
rect 4782 19610 4838 19612
rect 4862 19610 4918 19612
rect 4622 19558 4648 19610
rect 4648 19558 4678 19610
rect 4702 19558 4712 19610
rect 4712 19558 4758 19610
rect 4782 19558 4828 19610
rect 4828 19558 4838 19610
rect 4862 19558 4892 19610
rect 4892 19558 4918 19610
rect 4622 19556 4678 19558
rect 4702 19556 4758 19558
rect 4782 19556 4838 19558
rect 4862 19556 4918 19558
rect 1950 8880 2006 8936
rect 2318 8880 2374 8936
rect 1950 6160 2006 6216
rect 1582 5208 1638 5264
rect 2502 9016 2558 9072
rect 3146 10512 3202 10568
rect 2686 6160 2742 6216
rect 1674 4936 1730 4992
rect 1858 3984 1914 4040
rect 3422 9968 3478 10024
rect 3606 13232 3662 13288
rect 3422 6432 3478 6488
rect 4622 18522 4678 18524
rect 4702 18522 4758 18524
rect 4782 18522 4838 18524
rect 4862 18522 4918 18524
rect 4622 18470 4648 18522
rect 4648 18470 4678 18522
rect 4702 18470 4712 18522
rect 4712 18470 4758 18522
rect 4782 18470 4828 18522
rect 4828 18470 4838 18522
rect 4862 18470 4892 18522
rect 4892 18470 4918 18522
rect 4622 18468 4678 18470
rect 4702 18468 4758 18470
rect 4782 18468 4838 18470
rect 4862 18468 4918 18470
rect 4622 17434 4678 17436
rect 4702 17434 4758 17436
rect 4782 17434 4838 17436
rect 4862 17434 4918 17436
rect 4622 17382 4648 17434
rect 4648 17382 4678 17434
rect 4702 17382 4712 17434
rect 4712 17382 4758 17434
rect 4782 17382 4828 17434
rect 4828 17382 4838 17434
rect 4862 17382 4892 17434
rect 4892 17382 4918 17434
rect 4622 17380 4678 17382
rect 4702 17380 4758 17382
rect 4782 17380 4838 17382
rect 4862 17380 4918 17382
rect 4622 16346 4678 16348
rect 4702 16346 4758 16348
rect 4782 16346 4838 16348
rect 4862 16346 4918 16348
rect 4622 16294 4648 16346
rect 4648 16294 4678 16346
rect 4702 16294 4712 16346
rect 4712 16294 4758 16346
rect 4782 16294 4828 16346
rect 4828 16294 4838 16346
rect 4862 16294 4892 16346
rect 4892 16294 4918 16346
rect 4622 16292 4678 16294
rect 4702 16292 4758 16294
rect 4782 16292 4838 16294
rect 4862 16292 4918 16294
rect 4622 15258 4678 15260
rect 4702 15258 4758 15260
rect 4782 15258 4838 15260
rect 4862 15258 4918 15260
rect 4622 15206 4648 15258
rect 4648 15206 4678 15258
rect 4702 15206 4712 15258
rect 4712 15206 4758 15258
rect 4782 15206 4828 15258
rect 4828 15206 4838 15258
rect 4862 15206 4892 15258
rect 4892 15206 4918 15258
rect 4622 15204 4678 15206
rect 4702 15204 4758 15206
rect 4782 15204 4838 15206
rect 4862 15204 4918 15206
rect 5354 16088 5410 16144
rect 4622 14170 4678 14172
rect 4702 14170 4758 14172
rect 4782 14170 4838 14172
rect 4862 14170 4918 14172
rect 4622 14118 4648 14170
rect 4648 14118 4678 14170
rect 4702 14118 4712 14170
rect 4712 14118 4758 14170
rect 4782 14118 4828 14170
rect 4828 14118 4838 14170
rect 4862 14118 4892 14170
rect 4892 14118 4918 14170
rect 4622 14116 4678 14118
rect 4702 14116 4758 14118
rect 4782 14116 4838 14118
rect 4862 14116 4918 14118
rect 3790 11192 3846 11248
rect 4342 10376 4398 10432
rect 3698 7248 3754 7304
rect 3238 5208 3294 5264
rect 110 3576 166 3632
rect 110 2488 166 2544
rect 1674 992 1730 1048
rect 846 40 902 96
rect 2778 3576 2834 3632
rect 4622 13082 4678 13084
rect 4702 13082 4758 13084
rect 4782 13082 4838 13084
rect 4862 13082 4918 13084
rect 4622 13030 4648 13082
rect 4648 13030 4678 13082
rect 4702 13030 4712 13082
rect 4712 13030 4758 13082
rect 4782 13030 4828 13082
rect 4828 13030 4838 13082
rect 4862 13030 4892 13082
rect 4892 13030 4918 13082
rect 4622 13028 4678 13030
rect 4702 13028 4758 13030
rect 4782 13028 4838 13030
rect 4862 13028 4918 13030
rect 4622 11994 4678 11996
rect 4702 11994 4758 11996
rect 4782 11994 4838 11996
rect 4862 11994 4918 11996
rect 4622 11942 4648 11994
rect 4648 11942 4678 11994
rect 4702 11942 4712 11994
rect 4712 11942 4758 11994
rect 4782 11942 4828 11994
rect 4828 11942 4838 11994
rect 4862 11942 4892 11994
rect 4892 11942 4918 11994
rect 4622 11940 4678 11942
rect 4702 11940 4758 11942
rect 4782 11940 4838 11942
rect 4862 11940 4918 11942
rect 4622 10906 4678 10908
rect 4702 10906 4758 10908
rect 4782 10906 4838 10908
rect 4862 10906 4918 10908
rect 4622 10854 4648 10906
rect 4648 10854 4678 10906
rect 4702 10854 4712 10906
rect 4712 10854 4758 10906
rect 4782 10854 4828 10906
rect 4828 10854 4838 10906
rect 4862 10854 4892 10906
rect 4892 10854 4918 10906
rect 4622 10852 4678 10854
rect 4702 10852 4758 10854
rect 4782 10852 4838 10854
rect 4862 10852 4918 10854
rect 4622 9818 4678 9820
rect 4702 9818 4758 9820
rect 4782 9818 4838 9820
rect 4862 9818 4918 9820
rect 4622 9766 4648 9818
rect 4648 9766 4678 9818
rect 4702 9766 4712 9818
rect 4712 9766 4758 9818
rect 4782 9766 4828 9818
rect 4828 9766 4838 9818
rect 4862 9766 4892 9818
rect 4892 9766 4918 9818
rect 4622 9764 4678 9766
rect 4702 9764 4758 9766
rect 4782 9764 4838 9766
rect 4862 9764 4918 9766
rect 4622 8730 4678 8732
rect 4702 8730 4758 8732
rect 4782 8730 4838 8732
rect 4862 8730 4918 8732
rect 4622 8678 4648 8730
rect 4648 8678 4678 8730
rect 4702 8678 4712 8730
rect 4712 8678 4758 8730
rect 4782 8678 4828 8730
rect 4828 8678 4838 8730
rect 4862 8678 4892 8730
rect 4892 8678 4918 8730
rect 4622 8676 4678 8678
rect 4702 8676 4758 8678
rect 4782 8676 4838 8678
rect 4862 8676 4918 8678
rect 4622 7642 4678 7644
rect 4702 7642 4758 7644
rect 4782 7642 4838 7644
rect 4862 7642 4918 7644
rect 4622 7590 4648 7642
rect 4648 7590 4678 7642
rect 4702 7590 4712 7642
rect 4712 7590 4758 7642
rect 4782 7590 4828 7642
rect 4828 7590 4838 7642
rect 4862 7590 4892 7642
rect 4892 7590 4918 7642
rect 4622 7588 4678 7590
rect 4702 7588 4758 7590
rect 4782 7588 4838 7590
rect 4862 7588 4918 7590
rect 5722 17584 5778 17640
rect 5630 13776 5686 13832
rect 6458 13232 6514 13288
rect 6090 12824 6146 12880
rect 6090 12416 6146 12472
rect 5446 9152 5502 9208
rect 4622 6554 4678 6556
rect 4702 6554 4758 6556
rect 4782 6554 4838 6556
rect 4862 6554 4918 6556
rect 4622 6502 4648 6554
rect 4648 6502 4678 6554
rect 4702 6502 4712 6554
rect 4712 6502 4758 6554
rect 4782 6502 4828 6554
rect 4828 6502 4838 6554
rect 4862 6502 4892 6554
rect 4892 6502 4918 6554
rect 4622 6500 4678 6502
rect 4702 6500 4758 6502
rect 4782 6500 4838 6502
rect 4862 6500 4918 6502
rect 4986 6296 5042 6352
rect 4622 5466 4678 5468
rect 4702 5466 4758 5468
rect 4782 5466 4838 5468
rect 4862 5466 4918 5468
rect 4622 5414 4648 5466
rect 4648 5414 4678 5466
rect 4702 5414 4712 5466
rect 4712 5414 4758 5466
rect 4782 5414 4828 5466
rect 4828 5414 4838 5466
rect 4862 5414 4892 5466
rect 4892 5414 4918 5466
rect 4622 5412 4678 5414
rect 4702 5412 4758 5414
rect 4782 5412 4838 5414
rect 4862 5412 4918 5414
rect 4158 4528 4214 4584
rect 5630 7384 5686 7440
rect 5538 6976 5594 7032
rect 4622 4378 4678 4380
rect 4702 4378 4758 4380
rect 4782 4378 4838 4380
rect 4862 4378 4918 4380
rect 4622 4326 4648 4378
rect 4648 4326 4678 4378
rect 4702 4326 4712 4378
rect 4712 4326 4758 4378
rect 4782 4326 4828 4378
rect 4828 4326 4838 4378
rect 4862 4326 4892 4378
rect 4892 4326 4918 4378
rect 4622 4324 4678 4326
rect 4702 4324 4758 4326
rect 4782 4324 4838 4326
rect 4862 4324 4918 4326
rect 4526 3712 4582 3768
rect 5170 4528 5226 4584
rect 4622 3290 4678 3292
rect 4702 3290 4758 3292
rect 4782 3290 4838 3292
rect 4862 3290 4918 3292
rect 4622 3238 4648 3290
rect 4648 3238 4678 3290
rect 4702 3238 4712 3290
rect 4712 3238 4758 3290
rect 4782 3238 4828 3290
rect 4828 3238 4838 3290
rect 4862 3238 4892 3290
rect 4892 3238 4918 3290
rect 4622 3236 4678 3238
rect 4702 3236 4758 3238
rect 4782 3236 4838 3238
rect 4862 3236 4918 3238
rect 5722 2488 5778 2544
rect 5998 2896 6054 2952
rect 4622 2202 4678 2204
rect 4702 2202 4758 2204
rect 4782 2202 4838 2204
rect 4862 2202 4918 2204
rect 4622 2150 4648 2202
rect 4648 2150 4678 2202
rect 4702 2150 4712 2202
rect 4712 2150 4758 2202
rect 4782 2150 4828 2202
rect 4828 2150 4838 2202
rect 4862 2150 4892 2202
rect 4892 2150 4918 2202
rect 4622 2148 4678 2150
rect 4702 2148 4758 2150
rect 4782 2148 4838 2150
rect 4862 2148 4918 2150
rect 3054 1944 3110 2000
rect 5538 1944 5594 2000
rect 5078 1672 5134 1728
rect 6642 7792 6698 7848
rect 6918 10104 6974 10160
rect 8289 19066 8345 19068
rect 8369 19066 8425 19068
rect 8449 19066 8505 19068
rect 8529 19066 8585 19068
rect 8289 19014 8315 19066
rect 8315 19014 8345 19066
rect 8369 19014 8379 19066
rect 8379 19014 8425 19066
rect 8449 19014 8495 19066
rect 8495 19014 8505 19066
rect 8529 19014 8559 19066
rect 8559 19014 8585 19066
rect 8289 19012 8345 19014
rect 8369 19012 8425 19014
rect 8449 19012 8505 19014
rect 8529 19012 8585 19014
rect 8289 17978 8345 17980
rect 8369 17978 8425 17980
rect 8449 17978 8505 17980
rect 8529 17978 8585 17980
rect 8289 17926 8315 17978
rect 8315 17926 8345 17978
rect 8369 17926 8379 17978
rect 8379 17926 8425 17978
rect 8449 17926 8495 17978
rect 8495 17926 8505 17978
rect 8529 17926 8559 17978
rect 8559 17926 8585 17978
rect 8289 17924 8345 17926
rect 8369 17924 8425 17926
rect 8449 17924 8505 17926
rect 8529 17924 8585 17926
rect 8289 16890 8345 16892
rect 8369 16890 8425 16892
rect 8449 16890 8505 16892
rect 8529 16890 8585 16892
rect 8289 16838 8315 16890
rect 8315 16838 8345 16890
rect 8369 16838 8379 16890
rect 8379 16838 8425 16890
rect 8449 16838 8495 16890
rect 8495 16838 8505 16890
rect 8529 16838 8559 16890
rect 8559 16838 8585 16890
rect 8289 16836 8345 16838
rect 8369 16836 8425 16838
rect 8449 16836 8505 16838
rect 8529 16836 8585 16838
rect 8289 15802 8345 15804
rect 8369 15802 8425 15804
rect 8449 15802 8505 15804
rect 8529 15802 8585 15804
rect 8289 15750 8315 15802
rect 8315 15750 8345 15802
rect 8369 15750 8379 15802
rect 8379 15750 8425 15802
rect 8449 15750 8495 15802
rect 8495 15750 8505 15802
rect 8529 15750 8559 15802
rect 8559 15750 8585 15802
rect 8289 15748 8345 15750
rect 8369 15748 8425 15750
rect 8449 15748 8505 15750
rect 8529 15748 8585 15750
rect 8289 14714 8345 14716
rect 8369 14714 8425 14716
rect 8449 14714 8505 14716
rect 8529 14714 8585 14716
rect 8289 14662 8315 14714
rect 8315 14662 8345 14714
rect 8369 14662 8379 14714
rect 8379 14662 8425 14714
rect 8449 14662 8495 14714
rect 8495 14662 8505 14714
rect 8529 14662 8559 14714
rect 8559 14662 8585 14714
rect 8289 14660 8345 14662
rect 8369 14660 8425 14662
rect 8449 14660 8505 14662
rect 8529 14660 8585 14662
rect 8850 14320 8906 14376
rect 8289 13626 8345 13628
rect 8369 13626 8425 13628
rect 8449 13626 8505 13628
rect 8529 13626 8585 13628
rect 8289 13574 8315 13626
rect 8315 13574 8345 13626
rect 8369 13574 8379 13626
rect 8379 13574 8425 13626
rect 8449 13574 8495 13626
rect 8495 13574 8505 13626
rect 8529 13574 8559 13626
rect 8559 13574 8585 13626
rect 8289 13572 8345 13574
rect 8369 13572 8425 13574
rect 8449 13572 8505 13574
rect 8529 13572 8585 13574
rect 8289 12538 8345 12540
rect 8369 12538 8425 12540
rect 8449 12538 8505 12540
rect 8529 12538 8585 12540
rect 8289 12486 8315 12538
rect 8315 12486 8345 12538
rect 8369 12486 8379 12538
rect 8379 12486 8425 12538
rect 8449 12486 8495 12538
rect 8495 12486 8505 12538
rect 8529 12486 8559 12538
rect 8559 12486 8585 12538
rect 8289 12484 8345 12486
rect 8369 12484 8425 12486
rect 8449 12484 8505 12486
rect 8529 12484 8585 12486
rect 8022 9424 8078 9480
rect 7654 9016 7710 9072
rect 7286 8472 7342 8528
rect 7102 7112 7158 7168
rect 6550 6704 6606 6760
rect 7010 6704 7066 6760
rect 6458 4800 6514 4856
rect 6366 4700 6368 4720
rect 6368 4700 6420 4720
rect 6420 4700 6422 4720
rect 6366 4664 6422 4700
rect 6458 3440 6514 3496
rect 6734 3984 6790 4040
rect 6918 4120 6974 4176
rect 6550 3052 6606 3088
rect 6550 3032 6552 3052
rect 6552 3032 6604 3052
rect 6604 3032 6606 3052
rect 6182 1536 6238 1592
rect 6458 1400 6514 1456
rect 7470 6296 7526 6352
rect 7194 6196 7196 6216
rect 7196 6196 7248 6216
rect 7248 6196 7250 6216
rect 7194 6160 7250 6196
rect 7562 5344 7618 5400
rect 8289 11450 8345 11452
rect 8369 11450 8425 11452
rect 8449 11450 8505 11452
rect 8529 11450 8585 11452
rect 8289 11398 8315 11450
rect 8315 11398 8345 11450
rect 8369 11398 8379 11450
rect 8379 11398 8425 11450
rect 8449 11398 8495 11450
rect 8495 11398 8505 11450
rect 8529 11398 8559 11450
rect 8559 11398 8585 11450
rect 8289 11396 8345 11398
rect 8369 11396 8425 11398
rect 8449 11396 8505 11398
rect 8529 11396 8585 11398
rect 8289 10362 8345 10364
rect 8369 10362 8425 10364
rect 8449 10362 8505 10364
rect 8529 10362 8585 10364
rect 8289 10310 8315 10362
rect 8315 10310 8345 10362
rect 8369 10310 8379 10362
rect 8379 10310 8425 10362
rect 8449 10310 8495 10362
rect 8495 10310 8505 10362
rect 8529 10310 8559 10362
rect 8559 10310 8585 10362
rect 8289 10308 8345 10310
rect 8369 10308 8425 10310
rect 8449 10308 8505 10310
rect 8529 10308 8585 10310
rect 8850 13232 8906 13288
rect 8758 12144 8814 12200
rect 8289 9274 8345 9276
rect 8369 9274 8425 9276
rect 8449 9274 8505 9276
rect 8529 9274 8585 9276
rect 8289 9222 8315 9274
rect 8315 9222 8345 9274
rect 8369 9222 8379 9274
rect 8379 9222 8425 9274
rect 8449 9222 8495 9274
rect 8495 9222 8505 9274
rect 8529 9222 8559 9274
rect 8559 9222 8585 9274
rect 8289 9220 8345 9222
rect 8369 9220 8425 9222
rect 8449 9220 8505 9222
rect 8529 9220 8585 9222
rect 9034 9560 9090 9616
rect 9678 15952 9734 16008
rect 9678 15544 9734 15600
rect 8289 8186 8345 8188
rect 8369 8186 8425 8188
rect 8449 8186 8505 8188
rect 8529 8186 8585 8188
rect 8289 8134 8315 8186
rect 8315 8134 8345 8186
rect 8369 8134 8379 8186
rect 8379 8134 8425 8186
rect 8449 8134 8495 8186
rect 8495 8134 8505 8186
rect 8529 8134 8559 8186
rect 8559 8134 8585 8186
rect 8289 8132 8345 8134
rect 8369 8132 8425 8134
rect 8449 8132 8505 8134
rect 8529 8132 8585 8134
rect 8666 7928 8722 7984
rect 8666 7112 8722 7168
rect 8289 7098 8345 7100
rect 8369 7098 8425 7100
rect 8449 7098 8505 7100
rect 8529 7098 8585 7100
rect 8289 7046 8315 7098
rect 8315 7046 8345 7098
rect 8369 7046 8379 7098
rect 8379 7046 8425 7098
rect 8449 7046 8495 7098
rect 8495 7046 8505 7098
rect 8529 7046 8559 7098
rect 8559 7046 8585 7098
rect 8289 7044 8345 7046
rect 8369 7044 8425 7046
rect 8449 7044 8505 7046
rect 8529 7044 8585 7046
rect 8758 6024 8814 6080
rect 8289 6010 8345 6012
rect 8369 6010 8425 6012
rect 8449 6010 8505 6012
rect 8529 6010 8585 6012
rect 8289 5958 8315 6010
rect 8315 5958 8345 6010
rect 8369 5958 8379 6010
rect 8379 5958 8425 6010
rect 8449 5958 8495 6010
rect 8495 5958 8505 6010
rect 8529 5958 8559 6010
rect 8559 5958 8585 6010
rect 8289 5956 8345 5958
rect 8369 5956 8425 5958
rect 8449 5956 8505 5958
rect 8529 5956 8585 5958
rect 8289 4922 8345 4924
rect 8369 4922 8425 4924
rect 8449 4922 8505 4924
rect 8529 4922 8585 4924
rect 8289 4870 8315 4922
rect 8315 4870 8345 4922
rect 8369 4870 8379 4922
rect 8379 4870 8425 4922
rect 8449 4870 8495 4922
rect 8495 4870 8505 4922
rect 8529 4870 8559 4922
rect 8559 4870 8585 4922
rect 8289 4868 8345 4870
rect 8369 4868 8425 4870
rect 8449 4868 8505 4870
rect 8529 4868 8585 4870
rect 8289 3834 8345 3836
rect 8369 3834 8425 3836
rect 8449 3834 8505 3836
rect 8529 3834 8585 3836
rect 8289 3782 8315 3834
rect 8315 3782 8345 3834
rect 8369 3782 8379 3834
rect 8379 3782 8425 3834
rect 8449 3782 8495 3834
rect 8495 3782 8505 3834
rect 8529 3782 8559 3834
rect 8559 3782 8585 3834
rect 8289 3780 8345 3782
rect 8369 3780 8425 3782
rect 8449 3780 8505 3782
rect 8529 3780 8585 3782
rect 9402 11464 9458 11520
rect 9494 8880 9550 8936
rect 9586 8336 9642 8392
rect 9218 7248 9274 7304
rect 9126 3576 9182 3632
rect 8289 2746 8345 2748
rect 8369 2746 8425 2748
rect 8449 2746 8505 2748
rect 8529 2746 8585 2748
rect 8289 2694 8315 2746
rect 8315 2694 8345 2746
rect 8369 2694 8379 2746
rect 8379 2694 8425 2746
rect 8449 2694 8495 2746
rect 8495 2694 8505 2746
rect 8529 2694 8559 2746
rect 8559 2694 8585 2746
rect 8289 2692 8345 2694
rect 8369 2692 8425 2694
rect 8449 2692 8505 2694
rect 8529 2692 8585 2694
rect 6642 1264 6698 1320
rect 9402 6160 9458 6216
rect 10322 13096 10378 13152
rect 10506 13232 10562 13288
rect 11242 15544 11298 15600
rect 11956 19610 12012 19612
rect 12036 19610 12092 19612
rect 12116 19610 12172 19612
rect 12196 19610 12252 19612
rect 11956 19558 11982 19610
rect 11982 19558 12012 19610
rect 12036 19558 12046 19610
rect 12046 19558 12092 19610
rect 12116 19558 12162 19610
rect 12162 19558 12172 19610
rect 12196 19558 12226 19610
rect 12226 19558 12252 19610
rect 11956 19556 12012 19558
rect 12036 19556 12092 19558
rect 12116 19556 12172 19558
rect 12196 19556 12252 19558
rect 11956 18522 12012 18524
rect 12036 18522 12092 18524
rect 12116 18522 12172 18524
rect 12196 18522 12252 18524
rect 11956 18470 11982 18522
rect 11982 18470 12012 18522
rect 12036 18470 12046 18522
rect 12046 18470 12092 18522
rect 12116 18470 12162 18522
rect 12162 18470 12172 18522
rect 12196 18470 12226 18522
rect 12226 18470 12252 18522
rect 11956 18468 12012 18470
rect 12036 18468 12092 18470
rect 12116 18468 12172 18470
rect 12196 18468 12252 18470
rect 15622 19066 15678 19068
rect 15702 19066 15758 19068
rect 15782 19066 15838 19068
rect 15862 19066 15918 19068
rect 15622 19014 15648 19066
rect 15648 19014 15678 19066
rect 15702 19014 15712 19066
rect 15712 19014 15758 19066
rect 15782 19014 15828 19066
rect 15828 19014 15838 19066
rect 15862 19014 15892 19066
rect 15892 19014 15918 19066
rect 15622 19012 15678 19014
rect 15702 19012 15758 19014
rect 15782 19012 15838 19014
rect 15862 19012 15918 19014
rect 17866 18944 17922 19000
rect 11956 17434 12012 17436
rect 12036 17434 12092 17436
rect 12116 17434 12172 17436
rect 12196 17434 12252 17436
rect 11956 17382 11982 17434
rect 11982 17382 12012 17434
rect 12036 17382 12046 17434
rect 12046 17382 12092 17434
rect 12116 17382 12162 17434
rect 12162 17382 12172 17434
rect 12196 17382 12226 17434
rect 12226 17382 12252 17434
rect 11956 17380 12012 17382
rect 12036 17380 12092 17382
rect 12116 17380 12172 17382
rect 12196 17380 12252 17382
rect 11956 16346 12012 16348
rect 12036 16346 12092 16348
rect 12116 16346 12172 16348
rect 12196 16346 12252 16348
rect 11956 16294 11982 16346
rect 11982 16294 12012 16346
rect 12036 16294 12046 16346
rect 12046 16294 12092 16346
rect 12116 16294 12162 16346
rect 12162 16294 12172 16346
rect 12196 16294 12226 16346
rect 12226 16294 12252 16346
rect 11956 16292 12012 16294
rect 12036 16292 12092 16294
rect 12116 16292 12172 16294
rect 12196 16292 12252 16294
rect 11956 15258 12012 15260
rect 12036 15258 12092 15260
rect 12116 15258 12172 15260
rect 12196 15258 12252 15260
rect 11956 15206 11982 15258
rect 11982 15206 12012 15258
rect 12036 15206 12046 15258
rect 12046 15206 12092 15258
rect 12116 15206 12162 15258
rect 12162 15206 12172 15258
rect 12196 15206 12226 15258
rect 12226 15206 12252 15258
rect 11956 15204 12012 15206
rect 12036 15204 12092 15206
rect 12116 15204 12172 15206
rect 12196 15204 12252 15206
rect 11956 14170 12012 14172
rect 12036 14170 12092 14172
rect 12116 14170 12172 14172
rect 12196 14170 12252 14172
rect 11956 14118 11982 14170
rect 11982 14118 12012 14170
rect 12036 14118 12046 14170
rect 12046 14118 12092 14170
rect 12116 14118 12162 14170
rect 12162 14118 12172 14170
rect 12196 14118 12226 14170
rect 12226 14118 12252 14170
rect 11956 14116 12012 14118
rect 12036 14116 12092 14118
rect 12116 14116 12172 14118
rect 12196 14116 12252 14118
rect 11702 13776 11758 13832
rect 15622 17978 15678 17980
rect 15702 17978 15758 17980
rect 15782 17978 15838 17980
rect 15862 17978 15918 17980
rect 15622 17926 15648 17978
rect 15648 17926 15678 17978
rect 15702 17926 15712 17978
rect 15712 17926 15758 17978
rect 15782 17926 15828 17978
rect 15828 17926 15838 17978
rect 15862 17926 15892 17978
rect 15892 17926 15918 17978
rect 15622 17924 15678 17926
rect 15702 17924 15758 17926
rect 15782 17924 15838 17926
rect 15862 17924 15918 17926
rect 11956 13082 12012 13084
rect 12036 13082 12092 13084
rect 12116 13082 12172 13084
rect 12196 13082 12252 13084
rect 11956 13030 11982 13082
rect 11982 13030 12012 13082
rect 12036 13030 12046 13082
rect 12046 13030 12092 13082
rect 12116 13030 12162 13082
rect 12162 13030 12172 13082
rect 12196 13030 12226 13082
rect 12226 13030 12252 13082
rect 11956 13028 12012 13030
rect 12036 13028 12092 13030
rect 12116 13028 12172 13030
rect 12196 13028 12252 13030
rect 14186 13640 14242 13696
rect 11956 11994 12012 11996
rect 12036 11994 12092 11996
rect 12116 11994 12172 11996
rect 12196 11994 12252 11996
rect 11956 11942 11982 11994
rect 11982 11942 12012 11994
rect 12036 11942 12046 11994
rect 12046 11942 12092 11994
rect 12116 11942 12162 11994
rect 12162 11942 12172 11994
rect 12196 11942 12226 11994
rect 12226 11942 12252 11994
rect 11956 11940 12012 11942
rect 12036 11940 12092 11942
rect 12116 11940 12172 11942
rect 12196 11940 12252 11942
rect 11886 11756 11942 11792
rect 11886 11736 11888 11756
rect 11888 11736 11940 11756
rect 11940 11736 11942 11756
rect 11334 11600 11390 11656
rect 10506 9968 10562 10024
rect 11956 10906 12012 10908
rect 12036 10906 12092 10908
rect 12116 10906 12172 10908
rect 12196 10906 12252 10908
rect 11956 10854 11982 10906
rect 11982 10854 12012 10906
rect 12036 10854 12046 10906
rect 12046 10854 12092 10906
rect 12116 10854 12162 10906
rect 12162 10854 12172 10906
rect 12196 10854 12226 10906
rect 12226 10854 12252 10906
rect 11956 10852 12012 10854
rect 12036 10852 12092 10854
rect 12116 10852 12172 10854
rect 12196 10852 12252 10854
rect 12346 10512 12402 10568
rect 11956 9818 12012 9820
rect 12036 9818 12092 9820
rect 12116 9818 12172 9820
rect 12196 9818 12252 9820
rect 11956 9766 11982 9818
rect 11982 9766 12012 9818
rect 12036 9766 12046 9818
rect 12046 9766 12092 9818
rect 12116 9766 12162 9818
rect 12162 9766 12172 9818
rect 12196 9766 12226 9818
rect 12226 9766 12252 9818
rect 11956 9764 12012 9766
rect 12036 9764 12092 9766
rect 12116 9764 12172 9766
rect 12196 9764 12252 9766
rect 10874 9016 10930 9072
rect 11426 6840 11482 6896
rect 11956 8730 12012 8732
rect 12036 8730 12092 8732
rect 12116 8730 12172 8732
rect 12196 8730 12252 8732
rect 11956 8678 11982 8730
rect 11982 8678 12012 8730
rect 12036 8678 12046 8730
rect 12046 8678 12092 8730
rect 12116 8678 12162 8730
rect 12162 8678 12172 8730
rect 12196 8678 12226 8730
rect 12226 8678 12252 8730
rect 11956 8676 12012 8678
rect 12036 8676 12092 8678
rect 12116 8676 12172 8678
rect 12196 8676 12252 8678
rect 12622 8608 12678 8664
rect 14462 10104 14518 10160
rect 11956 7642 12012 7644
rect 12036 7642 12092 7644
rect 12116 7642 12172 7644
rect 12196 7642 12252 7644
rect 11956 7590 11982 7642
rect 11982 7590 12012 7642
rect 12036 7590 12046 7642
rect 12046 7590 12092 7642
rect 12116 7590 12162 7642
rect 12162 7590 12172 7642
rect 12196 7590 12226 7642
rect 12226 7590 12252 7642
rect 11956 7588 12012 7590
rect 12036 7588 12092 7590
rect 12116 7588 12172 7590
rect 12196 7588 12252 7590
rect 11242 5752 11298 5808
rect 11956 6554 12012 6556
rect 12036 6554 12092 6556
rect 12116 6554 12172 6556
rect 12196 6554 12252 6556
rect 11956 6502 11982 6554
rect 11982 6502 12012 6554
rect 12036 6502 12046 6554
rect 12046 6502 12092 6554
rect 12116 6502 12162 6554
rect 12162 6502 12172 6554
rect 12196 6502 12226 6554
rect 12226 6502 12252 6554
rect 11956 6500 12012 6502
rect 12036 6500 12092 6502
rect 12116 6500 12172 6502
rect 12196 6500 12252 6502
rect 11956 5466 12012 5468
rect 12036 5466 12092 5468
rect 12116 5466 12172 5468
rect 12196 5466 12252 5468
rect 11956 5414 11982 5466
rect 11982 5414 12012 5466
rect 12036 5414 12046 5466
rect 12046 5414 12092 5466
rect 12116 5414 12162 5466
rect 12162 5414 12172 5466
rect 12196 5414 12226 5466
rect 12226 5414 12252 5466
rect 11956 5412 12012 5414
rect 12036 5412 12092 5414
rect 12116 5412 12172 5414
rect 12196 5412 12252 5414
rect 9402 2624 9458 2680
rect 11058 5208 11114 5264
rect 11956 4378 12012 4380
rect 12036 4378 12092 4380
rect 12116 4378 12172 4380
rect 12196 4378 12252 4380
rect 11956 4326 11982 4378
rect 11982 4326 12012 4378
rect 12036 4326 12046 4378
rect 12046 4326 12092 4378
rect 12116 4326 12162 4378
rect 12162 4326 12172 4378
rect 12196 4326 12226 4378
rect 12226 4326 12252 4378
rect 11956 4324 12012 4326
rect 12036 4324 12092 4326
rect 12116 4324 12172 4326
rect 12196 4324 12252 4326
rect 11242 3984 11298 4040
rect 11956 3290 12012 3292
rect 12036 3290 12092 3292
rect 12116 3290 12172 3292
rect 12196 3290 12252 3292
rect 11956 3238 11982 3290
rect 11982 3238 12012 3290
rect 12036 3238 12046 3290
rect 12046 3238 12092 3290
rect 12116 3238 12162 3290
rect 12162 3238 12172 3290
rect 12196 3238 12226 3290
rect 12226 3238 12252 3290
rect 11956 3236 12012 3238
rect 12036 3236 12092 3238
rect 12116 3236 12172 3238
rect 12196 3236 12252 3238
rect 15622 16890 15678 16892
rect 15702 16890 15758 16892
rect 15782 16890 15838 16892
rect 15862 16890 15918 16892
rect 15622 16838 15648 16890
rect 15648 16838 15678 16890
rect 15702 16838 15712 16890
rect 15712 16838 15758 16890
rect 15782 16838 15828 16890
rect 15828 16838 15838 16890
rect 15862 16838 15892 16890
rect 15892 16838 15918 16890
rect 15622 16836 15678 16838
rect 15702 16836 15758 16838
rect 15782 16836 15838 16838
rect 15862 16836 15918 16838
rect 16302 16088 16358 16144
rect 15622 15802 15678 15804
rect 15702 15802 15758 15804
rect 15782 15802 15838 15804
rect 15862 15802 15918 15804
rect 15622 15750 15648 15802
rect 15648 15750 15678 15802
rect 15702 15750 15712 15802
rect 15712 15750 15758 15802
rect 15782 15750 15828 15802
rect 15828 15750 15838 15802
rect 15862 15750 15892 15802
rect 15892 15750 15918 15802
rect 15622 15748 15678 15750
rect 15702 15748 15758 15750
rect 15782 15748 15838 15750
rect 15862 15748 15918 15750
rect 14646 10104 14702 10160
rect 15106 13640 15162 13696
rect 15198 12144 15254 12200
rect 15198 11872 15254 11928
rect 15622 14714 15678 14716
rect 15702 14714 15758 14716
rect 15782 14714 15838 14716
rect 15862 14714 15918 14716
rect 15622 14662 15648 14714
rect 15648 14662 15678 14714
rect 15702 14662 15712 14714
rect 15712 14662 15758 14714
rect 15782 14662 15828 14714
rect 15828 14662 15838 14714
rect 15862 14662 15892 14714
rect 15892 14662 15918 14714
rect 15622 14660 15678 14662
rect 15702 14660 15758 14662
rect 15782 14660 15838 14662
rect 15862 14660 15918 14662
rect 15622 13626 15678 13628
rect 15702 13626 15758 13628
rect 15782 13626 15838 13628
rect 15862 13626 15918 13628
rect 15622 13574 15648 13626
rect 15648 13574 15678 13626
rect 15702 13574 15712 13626
rect 15712 13574 15758 13626
rect 15782 13574 15828 13626
rect 15828 13574 15838 13626
rect 15862 13574 15892 13626
rect 15892 13574 15918 13626
rect 15622 13572 15678 13574
rect 15702 13572 15758 13574
rect 15782 13572 15838 13574
rect 15862 13572 15918 13574
rect 15622 12538 15678 12540
rect 15702 12538 15758 12540
rect 15782 12538 15838 12540
rect 15862 12538 15918 12540
rect 15622 12486 15648 12538
rect 15648 12486 15678 12538
rect 15702 12486 15712 12538
rect 15712 12486 15758 12538
rect 15782 12486 15828 12538
rect 15828 12486 15838 12538
rect 15862 12486 15892 12538
rect 15892 12486 15918 12538
rect 15622 12484 15678 12486
rect 15702 12484 15758 12486
rect 15782 12484 15838 12486
rect 15862 12484 15918 12486
rect 15014 11464 15070 11520
rect 15622 11450 15678 11452
rect 15702 11450 15758 11452
rect 15782 11450 15838 11452
rect 15862 11450 15918 11452
rect 15622 11398 15648 11450
rect 15648 11398 15678 11450
rect 15702 11398 15712 11450
rect 15712 11398 15758 11450
rect 15782 11398 15828 11450
rect 15828 11398 15838 11450
rect 15862 11398 15892 11450
rect 15892 11398 15918 11450
rect 15622 11396 15678 11398
rect 15702 11396 15758 11398
rect 15782 11396 15838 11398
rect 15862 11396 15918 11398
rect 13634 6568 13690 6624
rect 14830 7248 14886 7304
rect 14278 6432 14334 6488
rect 14554 6296 14610 6352
rect 14830 6296 14886 6352
rect 12622 3440 12678 3496
rect 12530 3032 12586 3088
rect 12530 2488 12586 2544
rect 8666 2352 8722 2408
rect 11956 2202 12012 2204
rect 12036 2202 12092 2204
rect 12116 2202 12172 2204
rect 12196 2202 12252 2204
rect 11956 2150 11982 2202
rect 11982 2150 12012 2202
rect 12036 2150 12046 2202
rect 12046 2150 12092 2202
rect 12116 2150 12162 2202
rect 12162 2150 12172 2202
rect 12196 2150 12226 2202
rect 12226 2150 12252 2202
rect 11956 2148 12012 2150
rect 12036 2148 12092 2150
rect 12116 2148 12172 2150
rect 12196 2148 12252 2150
rect 15622 10362 15678 10364
rect 15702 10362 15758 10364
rect 15782 10362 15838 10364
rect 15862 10362 15918 10364
rect 15622 10310 15648 10362
rect 15648 10310 15678 10362
rect 15702 10310 15712 10362
rect 15712 10310 15758 10362
rect 15782 10310 15828 10362
rect 15828 10310 15838 10362
rect 15862 10310 15892 10362
rect 15892 10310 15918 10362
rect 15622 10308 15678 10310
rect 15702 10308 15758 10310
rect 15782 10308 15838 10310
rect 15862 10308 15918 10310
rect 15622 9274 15678 9276
rect 15702 9274 15758 9276
rect 15782 9274 15838 9276
rect 15862 9274 15918 9276
rect 15622 9222 15648 9274
rect 15648 9222 15678 9274
rect 15702 9222 15712 9274
rect 15712 9222 15758 9274
rect 15782 9222 15828 9274
rect 15828 9222 15838 9274
rect 15862 9222 15892 9274
rect 15892 9222 15918 9274
rect 15622 9220 15678 9222
rect 15702 9220 15758 9222
rect 15782 9220 15838 9222
rect 15862 9220 15918 9222
rect 16118 12824 16174 12880
rect 15658 8336 15714 8392
rect 15622 8186 15678 8188
rect 15702 8186 15758 8188
rect 15782 8186 15838 8188
rect 15862 8186 15918 8188
rect 15622 8134 15648 8186
rect 15648 8134 15678 8186
rect 15702 8134 15712 8186
rect 15712 8134 15758 8186
rect 15782 8134 15828 8186
rect 15828 8134 15838 8186
rect 15862 8134 15892 8186
rect 15892 8134 15918 8186
rect 15622 8132 15678 8134
rect 15702 8132 15758 8134
rect 15782 8132 15838 8134
rect 15862 8132 15918 8134
rect 15382 7792 15438 7848
rect 15290 7112 15346 7168
rect 15622 7098 15678 7100
rect 15702 7098 15758 7100
rect 15782 7098 15838 7100
rect 15862 7098 15918 7100
rect 15622 7046 15648 7098
rect 15648 7046 15678 7098
rect 15702 7046 15712 7098
rect 15712 7046 15758 7098
rect 15782 7046 15828 7098
rect 15828 7046 15838 7098
rect 15862 7046 15892 7098
rect 15892 7046 15918 7098
rect 15622 7044 15678 7046
rect 15702 7044 15758 7046
rect 15782 7044 15838 7046
rect 15862 7044 15918 7046
rect 15382 6024 15438 6080
rect 16210 7928 16266 7984
rect 17590 15952 17646 16008
rect 16946 14320 17002 14376
rect 17130 11872 17186 11928
rect 16578 9152 16634 9208
rect 16946 8880 17002 8936
rect 16210 6296 16266 6352
rect 15622 6010 15678 6012
rect 15702 6010 15758 6012
rect 15782 6010 15838 6012
rect 15862 6010 15918 6012
rect 15622 5958 15648 6010
rect 15648 5958 15678 6010
rect 15702 5958 15712 6010
rect 15712 5958 15758 6010
rect 15782 5958 15828 6010
rect 15828 5958 15838 6010
rect 15862 5958 15892 6010
rect 15892 5958 15918 6010
rect 15622 5956 15678 5958
rect 15702 5956 15758 5958
rect 15782 5956 15838 5958
rect 15862 5956 15918 5958
rect 15622 4922 15678 4924
rect 15702 4922 15758 4924
rect 15782 4922 15838 4924
rect 15862 4922 15918 4924
rect 15622 4870 15648 4922
rect 15648 4870 15678 4922
rect 15702 4870 15712 4922
rect 15712 4870 15758 4922
rect 15782 4870 15828 4922
rect 15828 4870 15838 4922
rect 15862 4870 15892 4922
rect 15892 4870 15918 4922
rect 15622 4868 15678 4870
rect 15702 4868 15758 4870
rect 15782 4868 15838 4870
rect 15862 4868 15918 4870
rect 15474 4664 15530 4720
rect 15934 4528 15990 4584
rect 16762 7112 16818 7168
rect 17314 11736 17370 11792
rect 17130 8608 17186 8664
rect 16670 6704 16726 6760
rect 16578 6568 16634 6624
rect 16302 4120 16358 4176
rect 17774 13796 17830 13832
rect 17774 13776 17776 13796
rect 17776 13776 17828 13796
rect 17828 13776 17830 13796
rect 17590 9968 17646 10024
rect 19289 19610 19345 19612
rect 19369 19610 19425 19612
rect 19449 19610 19505 19612
rect 19529 19610 19585 19612
rect 19289 19558 19315 19610
rect 19315 19558 19345 19610
rect 19369 19558 19379 19610
rect 19379 19558 19425 19610
rect 19449 19558 19495 19610
rect 19495 19558 19505 19610
rect 19529 19558 19559 19610
rect 19559 19558 19585 19610
rect 19289 19556 19345 19558
rect 19369 19556 19425 19558
rect 19449 19556 19505 19558
rect 19529 19556 19585 19558
rect 19289 18522 19345 18524
rect 19369 18522 19425 18524
rect 19449 18522 19505 18524
rect 19529 18522 19585 18524
rect 19289 18470 19315 18522
rect 19315 18470 19345 18522
rect 19369 18470 19379 18522
rect 19379 18470 19425 18522
rect 19449 18470 19495 18522
rect 19495 18470 19505 18522
rect 19529 18470 19559 18522
rect 19559 18470 19585 18522
rect 19289 18468 19345 18470
rect 19369 18468 19425 18470
rect 19449 18468 19505 18470
rect 19529 18468 19585 18470
rect 21546 21120 21602 21176
rect 19289 17434 19345 17436
rect 19369 17434 19425 17436
rect 19449 17434 19505 17436
rect 19529 17434 19585 17436
rect 19289 17382 19315 17434
rect 19315 17382 19345 17434
rect 19369 17382 19379 17434
rect 19379 17382 19425 17434
rect 19449 17382 19495 17434
rect 19495 17382 19505 17434
rect 19529 17382 19559 17434
rect 19559 17382 19585 17434
rect 19289 17380 19345 17382
rect 19369 17380 19425 17382
rect 19449 17380 19505 17382
rect 19529 17380 19585 17382
rect 19246 17176 19302 17232
rect 18142 16632 18198 16688
rect 19289 16346 19345 16348
rect 19369 16346 19425 16348
rect 19449 16346 19505 16348
rect 19529 16346 19585 16348
rect 19289 16294 19315 16346
rect 19315 16294 19345 16346
rect 19369 16294 19379 16346
rect 19379 16294 19425 16346
rect 19449 16294 19495 16346
rect 19495 16294 19505 16346
rect 19529 16294 19559 16346
rect 19559 16294 19585 16346
rect 19289 16292 19345 16294
rect 19369 16292 19425 16294
rect 19449 16292 19505 16294
rect 19529 16292 19585 16294
rect 17774 11192 17830 11248
rect 18142 9560 18198 9616
rect 18142 9016 18198 9072
rect 18510 8472 18566 8528
rect 17774 7384 17830 7440
rect 17498 6840 17554 6896
rect 17314 6160 17370 6216
rect 15622 3834 15678 3836
rect 15702 3834 15758 3836
rect 15782 3834 15838 3836
rect 15862 3834 15918 3836
rect 15622 3782 15648 3834
rect 15648 3782 15678 3834
rect 15702 3782 15712 3834
rect 15712 3782 15758 3834
rect 15782 3782 15828 3834
rect 15828 3782 15838 3834
rect 15862 3782 15892 3834
rect 15892 3782 15918 3834
rect 15622 3780 15678 3782
rect 15702 3780 15758 3782
rect 15782 3780 15838 3782
rect 15862 3780 15918 3782
rect 15106 1944 15162 2000
rect 16118 2896 16174 2952
rect 15622 2746 15678 2748
rect 15702 2746 15758 2748
rect 15782 2746 15838 2748
rect 15862 2746 15918 2748
rect 15622 2694 15648 2746
rect 15648 2694 15678 2746
rect 15702 2694 15712 2746
rect 15712 2694 15758 2746
rect 15782 2694 15828 2746
rect 15828 2694 15838 2746
rect 15862 2694 15892 2746
rect 15892 2694 15918 2746
rect 15622 2692 15678 2694
rect 15702 2692 15758 2694
rect 15782 2692 15838 2694
rect 15862 2692 15918 2694
rect 16486 2488 16542 2544
rect 18050 5072 18106 5128
rect 17958 3032 18014 3088
rect 18326 3168 18382 3224
rect 18234 2896 18290 2952
rect 15566 2352 15622 2408
rect 15198 1672 15254 1728
rect 14830 1536 14886 1592
rect 19289 15258 19345 15260
rect 19369 15258 19425 15260
rect 19449 15258 19505 15260
rect 19529 15258 19585 15260
rect 19289 15206 19315 15258
rect 19315 15206 19345 15258
rect 19369 15206 19379 15258
rect 19379 15206 19425 15258
rect 19449 15206 19495 15258
rect 19495 15206 19505 15258
rect 19529 15206 19559 15258
rect 19559 15206 19585 15258
rect 19289 15204 19345 15206
rect 19369 15204 19425 15206
rect 19449 15204 19505 15206
rect 19529 15204 19585 15206
rect 21546 14320 21602 14376
rect 19289 14170 19345 14172
rect 19369 14170 19425 14172
rect 19449 14170 19505 14172
rect 19529 14170 19585 14172
rect 19289 14118 19315 14170
rect 19315 14118 19345 14170
rect 19369 14118 19379 14170
rect 19379 14118 19425 14170
rect 19449 14118 19495 14170
rect 19495 14118 19505 14170
rect 19529 14118 19559 14170
rect 19559 14118 19585 14170
rect 19289 14116 19345 14118
rect 19369 14116 19425 14118
rect 19449 14116 19505 14118
rect 19529 14116 19585 14118
rect 18970 11600 19026 11656
rect 19289 13082 19345 13084
rect 19369 13082 19425 13084
rect 19449 13082 19505 13084
rect 19529 13082 19585 13084
rect 19289 13030 19315 13082
rect 19315 13030 19345 13082
rect 19369 13030 19379 13082
rect 19379 13030 19425 13082
rect 19449 13030 19495 13082
rect 19495 13030 19505 13082
rect 19529 13030 19559 13082
rect 19559 13030 19585 13082
rect 19289 13028 19345 13030
rect 19369 13028 19425 13030
rect 19449 13028 19505 13030
rect 19529 13028 19585 13030
rect 19289 11994 19345 11996
rect 19369 11994 19425 11996
rect 19449 11994 19505 11996
rect 19529 11994 19585 11996
rect 19289 11942 19315 11994
rect 19315 11942 19345 11994
rect 19369 11942 19379 11994
rect 19379 11942 19425 11994
rect 19449 11942 19495 11994
rect 19495 11942 19505 11994
rect 19529 11942 19559 11994
rect 19559 11942 19585 11994
rect 19289 11940 19345 11942
rect 19369 11940 19425 11942
rect 19449 11940 19505 11942
rect 19529 11940 19585 11942
rect 19289 10906 19345 10908
rect 19369 10906 19425 10908
rect 19449 10906 19505 10908
rect 19529 10906 19585 10908
rect 19289 10854 19315 10906
rect 19315 10854 19345 10906
rect 19369 10854 19379 10906
rect 19379 10854 19425 10906
rect 19449 10854 19495 10906
rect 19495 10854 19505 10906
rect 19529 10854 19559 10906
rect 19559 10854 19585 10906
rect 19289 10852 19345 10854
rect 19369 10852 19425 10854
rect 19449 10852 19505 10854
rect 19529 10852 19585 10854
rect 19289 9818 19345 9820
rect 19369 9818 19425 9820
rect 19449 9818 19505 9820
rect 19529 9818 19585 9820
rect 19289 9766 19315 9818
rect 19315 9766 19345 9818
rect 19369 9766 19379 9818
rect 19379 9766 19425 9818
rect 19449 9766 19495 9818
rect 19495 9766 19505 9818
rect 19529 9766 19559 9818
rect 19559 9766 19585 9818
rect 19289 9764 19345 9766
rect 19369 9764 19425 9766
rect 19449 9764 19505 9766
rect 19529 9764 19585 9766
rect 19706 9968 19762 10024
rect 19614 9424 19670 9480
rect 19062 8472 19118 8528
rect 19289 8730 19345 8732
rect 19369 8730 19425 8732
rect 19449 8730 19505 8732
rect 19529 8730 19585 8732
rect 19289 8678 19315 8730
rect 19315 8678 19345 8730
rect 19369 8678 19379 8730
rect 19379 8678 19425 8730
rect 19449 8678 19495 8730
rect 19495 8678 19505 8730
rect 19529 8678 19559 8730
rect 19559 8678 19585 8730
rect 19289 8676 19345 8678
rect 19369 8676 19425 8678
rect 19449 8676 19505 8678
rect 19529 8676 19585 8678
rect 18694 7384 18750 7440
rect 18970 5752 19026 5808
rect 19289 7642 19345 7644
rect 19369 7642 19425 7644
rect 19449 7642 19505 7644
rect 19529 7642 19585 7644
rect 19289 7590 19315 7642
rect 19315 7590 19345 7642
rect 19369 7590 19379 7642
rect 19379 7590 19425 7642
rect 19449 7590 19495 7642
rect 19495 7590 19505 7642
rect 19529 7590 19559 7642
rect 19559 7590 19585 7642
rect 19289 7588 19345 7590
rect 19369 7588 19425 7590
rect 19449 7588 19505 7590
rect 19529 7588 19585 7590
rect 20074 12144 20130 12200
rect 20442 11192 20498 11248
rect 19289 6554 19345 6556
rect 19369 6554 19425 6556
rect 19449 6554 19505 6556
rect 19529 6554 19585 6556
rect 19289 6502 19315 6554
rect 19315 6502 19345 6554
rect 19369 6502 19379 6554
rect 19379 6502 19425 6554
rect 19449 6502 19495 6554
rect 19495 6502 19505 6554
rect 19529 6502 19559 6554
rect 19559 6502 19585 6554
rect 19289 6500 19345 6502
rect 19369 6500 19425 6502
rect 19449 6500 19505 6502
rect 19529 6500 19585 6502
rect 19289 5466 19345 5468
rect 19369 5466 19425 5468
rect 19449 5466 19505 5468
rect 19529 5466 19585 5468
rect 19289 5414 19315 5466
rect 19315 5414 19345 5466
rect 19369 5414 19379 5466
rect 19379 5414 19425 5466
rect 19449 5414 19495 5466
rect 19495 5414 19505 5466
rect 19529 5414 19559 5466
rect 19559 5414 19585 5466
rect 19289 5412 19345 5414
rect 19369 5412 19425 5414
rect 19449 5412 19505 5414
rect 19529 5412 19585 5414
rect 18050 1672 18106 1728
rect 17774 1264 17830 1320
rect 19289 4378 19345 4380
rect 19369 4378 19425 4380
rect 19449 4378 19505 4380
rect 19529 4378 19585 4380
rect 19289 4326 19315 4378
rect 19315 4326 19345 4378
rect 19369 4326 19379 4378
rect 19379 4326 19425 4378
rect 19449 4326 19495 4378
rect 19495 4326 19505 4378
rect 19529 4326 19559 4378
rect 19559 4326 19585 4378
rect 19289 4324 19345 4326
rect 19369 4324 19425 4326
rect 19449 4324 19505 4326
rect 19529 4324 19585 4326
rect 21638 4120 21694 4176
rect 19289 3290 19345 3292
rect 19369 3290 19425 3292
rect 19449 3290 19505 3292
rect 19529 3290 19585 3292
rect 19289 3238 19315 3290
rect 19315 3238 19345 3290
rect 19369 3238 19379 3290
rect 19379 3238 19425 3290
rect 19449 3238 19495 3290
rect 19495 3238 19505 3290
rect 19529 3238 19559 3290
rect 19559 3238 19585 3290
rect 19289 3236 19345 3238
rect 19369 3236 19425 3238
rect 19449 3236 19505 3238
rect 19529 3236 19585 3238
rect 19289 2202 19345 2204
rect 19369 2202 19425 2204
rect 19449 2202 19505 2204
rect 19529 2202 19585 2204
rect 19289 2150 19315 2202
rect 19315 2150 19345 2202
rect 19369 2150 19379 2202
rect 19379 2150 19425 2202
rect 19449 2150 19495 2202
rect 19495 2150 19505 2202
rect 19529 2150 19559 2202
rect 19559 2150 19585 2202
rect 19289 2148 19345 2150
rect 19369 2148 19425 2150
rect 19449 2148 19505 2150
rect 19529 2148 19585 2150
rect 19062 1400 19118 1456
<< metal3 >>
rect 1025 21586 1091 21589
rect 2630 21586 2636 21588
rect 1025 21584 2636 21586
rect 1025 21528 1030 21584
rect 1086 21528 2636 21584
rect 1025 21526 2636 21528
rect 1025 21523 1091 21526
rect 2630 21524 2636 21526
rect 2700 21524 2706 21588
rect 0 21360 480 21480
rect 62 20906 122 21360
rect 21520 21178 22000 21208
rect 21460 21176 22000 21178
rect 21460 21120 21546 21176
rect 21602 21120 22000 21176
rect 21460 21118 22000 21120
rect 21520 21088 22000 21118
rect 2957 20906 3023 20909
rect 62 20904 3023 20906
rect 62 20848 2962 20904
rect 3018 20848 3023 20904
rect 62 20846 3023 20848
rect 2957 20843 3023 20846
rect 0 20360 480 20392
rect 0 20304 18 20360
rect 74 20304 480 20360
rect 0 20272 480 20304
rect 4610 19616 4930 19617
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4930 19616
rect 4610 19551 4930 19552
rect 11944 19616 12264 19617
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 19551 12264 19552
rect 19277 19616 19597 19617
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 19551 19597 19552
rect 21520 19456 22000 19576
rect 0 19272 480 19304
rect 0 19216 110 19272
rect 166 19216 480 19272
rect 0 19184 480 19216
rect 8277 19072 8597 19073
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 19007 8597 19008
rect 15610 19072 15930 19073
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 19007 15930 19008
rect 17861 19002 17927 19005
rect 21590 19002 21650 19456
rect 17861 19000 21650 19002
rect 17861 18944 17866 19000
rect 17922 18944 21650 19000
rect 17861 18942 21650 18944
rect 17861 18939 17927 18942
rect 4610 18528 4930 18529
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4930 18528
rect 4610 18463 4930 18464
rect 11944 18528 12264 18529
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 18463 12264 18464
rect 19277 18528 19597 18529
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 19277 18463 19597 18464
rect 0 18232 480 18352
rect 62 17778 122 18232
rect 8277 17984 8597 17985
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 8277 17919 8597 17920
rect 15610 17984 15930 17985
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 15610 17919 15930 17920
rect 1209 17778 1275 17781
rect 62 17776 1275 17778
rect 62 17720 1214 17776
rect 1270 17720 1275 17776
rect 62 17718 1275 17720
rect 1209 17715 1275 17718
rect 21520 17688 22000 17808
rect 1301 17642 1367 17645
rect 5717 17642 5783 17645
rect 1301 17640 5783 17642
rect 1301 17584 1306 17640
rect 1362 17584 5722 17640
rect 5778 17584 5783 17640
rect 1301 17582 5783 17584
rect 1301 17579 1367 17582
rect 5717 17579 5783 17582
rect 4610 17440 4930 17441
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4930 17440
rect 4610 17375 4930 17376
rect 11944 17440 12264 17441
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 11944 17375 12264 17376
rect 19277 17440 19597 17441
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 17375 19597 17376
rect 0 17232 480 17264
rect 0 17176 110 17232
rect 166 17176 480 17232
rect 0 17144 480 17176
rect 19241 17234 19307 17237
rect 21590 17234 21650 17688
rect 19241 17232 21650 17234
rect 19241 17176 19246 17232
rect 19302 17176 21650 17232
rect 19241 17174 21650 17176
rect 19241 17171 19307 17174
rect 8277 16896 8597 16897
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 8277 16831 8597 16832
rect 15610 16896 15930 16897
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 15610 16831 15930 16832
rect 289 16690 355 16693
rect 18137 16690 18203 16693
rect 289 16688 18203 16690
rect 289 16632 294 16688
rect 350 16632 18142 16688
rect 18198 16632 18203 16688
rect 289 16630 18203 16632
rect 289 16627 355 16630
rect 18137 16627 18203 16630
rect 54 16356 60 16420
rect 124 16418 130 16420
rect 1577 16418 1643 16421
rect 124 16416 1643 16418
rect 124 16360 1582 16416
rect 1638 16360 1643 16416
rect 124 16358 1643 16360
rect 124 16356 130 16358
rect 1577 16355 1643 16358
rect 4610 16352 4930 16353
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4930 16352
rect 4610 16287 4930 16288
rect 11944 16352 12264 16353
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11944 16287 12264 16288
rect 19277 16352 19597 16353
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 16287 19597 16288
rect 0 16148 480 16176
rect 0 16084 60 16148
rect 124 16084 480 16148
rect 0 16056 480 16084
rect 5349 16146 5415 16149
rect 16297 16146 16363 16149
rect 5349 16144 16363 16146
rect 5349 16088 5354 16144
rect 5410 16088 16302 16144
rect 16358 16088 16363 16144
rect 5349 16086 16363 16088
rect 5349 16083 5415 16086
rect 16297 16083 16363 16086
rect 21520 16056 22000 16176
rect 9673 16010 9739 16013
rect 17585 16010 17651 16013
rect 9673 16008 17651 16010
rect 9673 15952 9678 16008
rect 9734 15952 17590 16008
rect 17646 15952 17651 16008
rect 9673 15950 17651 15952
rect 9673 15947 9739 15950
rect 17585 15947 17651 15950
rect 8277 15808 8597 15809
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 8277 15743 8597 15744
rect 15610 15808 15930 15809
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 15743 15930 15744
rect 2037 15602 2103 15605
rect 9673 15602 9739 15605
rect 2037 15600 9739 15602
rect 2037 15544 2042 15600
rect 2098 15544 9678 15600
rect 9734 15544 9739 15600
rect 2037 15542 9739 15544
rect 2037 15539 2103 15542
rect 9673 15539 9739 15542
rect 11237 15602 11303 15605
rect 21590 15602 21650 16056
rect 11237 15600 21650 15602
rect 11237 15544 11242 15600
rect 11298 15544 21650 15600
rect 11237 15542 21650 15544
rect 11237 15539 11303 15542
rect 4610 15264 4930 15265
rect 0 15104 480 15224
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4930 15264
rect 4610 15199 4930 15200
rect 11944 15264 12264 15265
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11944 15199 12264 15200
rect 19277 15264 19597 15265
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 19277 15199 19597 15200
rect 62 14650 122 15104
rect 8277 14720 8597 14721
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 8277 14655 8597 14656
rect 15610 14720 15930 14721
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 15610 14655 15930 14656
rect 1393 14650 1459 14653
rect 62 14648 1459 14650
rect 62 14592 1398 14648
rect 1454 14592 1459 14648
rect 62 14590 1459 14592
rect 1393 14587 1459 14590
rect 8845 14378 8911 14381
rect 16941 14378 17007 14381
rect 21520 14378 22000 14408
rect 8845 14376 17007 14378
rect 8845 14320 8850 14376
rect 8906 14320 16946 14376
rect 17002 14320 17007 14376
rect 8845 14318 17007 14320
rect 21460 14376 22000 14378
rect 21460 14320 21546 14376
rect 21602 14320 22000 14376
rect 21460 14318 22000 14320
rect 8845 14315 8911 14318
rect 16941 14315 17007 14318
rect 21520 14288 22000 14318
rect 4610 14176 4930 14177
rect 0 14108 480 14136
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4930 14176
rect 4610 14111 4930 14112
rect 11944 14176 12264 14177
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11944 14111 12264 14112
rect 19277 14176 19597 14177
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 14111 19597 14112
rect 0 14044 60 14108
rect 124 14044 480 14108
rect 0 14016 480 14044
rect 54 13772 60 13836
rect 124 13834 130 13836
rect 5625 13834 5691 13837
rect 124 13832 5691 13834
rect 124 13776 5630 13832
rect 5686 13776 5691 13832
rect 124 13774 5691 13776
rect 124 13772 130 13774
rect 5625 13771 5691 13774
rect 11697 13834 11763 13837
rect 17769 13834 17835 13837
rect 11697 13832 17835 13834
rect 11697 13776 11702 13832
rect 11758 13776 17774 13832
rect 17830 13776 17835 13832
rect 11697 13774 17835 13776
rect 11697 13771 11763 13774
rect 17769 13771 17835 13774
rect 14181 13698 14247 13701
rect 15101 13698 15167 13701
rect 14181 13696 15167 13698
rect 14181 13640 14186 13696
rect 14242 13640 15106 13696
rect 15162 13640 15167 13696
rect 14181 13638 15167 13640
rect 14181 13635 14247 13638
rect 15101 13635 15167 13638
rect 8277 13632 8597 13633
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 8277 13567 8597 13568
rect 15610 13632 15930 13633
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 15610 13567 15930 13568
rect 3601 13290 3667 13293
rect 6453 13290 6519 13293
rect 8845 13290 8911 13293
rect 10501 13290 10567 13293
rect 62 13288 6378 13290
rect 62 13232 3606 13288
rect 3662 13232 6378 13288
rect 62 13230 6378 13232
rect 62 13048 122 13230
rect 3601 13227 3667 13230
rect 6318 13154 6378 13230
rect 6453 13288 10567 13290
rect 6453 13232 6458 13288
rect 6514 13232 8850 13288
rect 8906 13232 10506 13288
rect 10562 13232 10567 13288
rect 6453 13230 10567 13232
rect 6453 13227 6519 13230
rect 8845 13227 8911 13230
rect 10501 13227 10567 13230
rect 10317 13154 10383 13157
rect 6318 13152 10383 13154
rect 6318 13096 10322 13152
rect 10378 13096 10383 13152
rect 6318 13094 10383 13096
rect 10317 13091 10383 13094
rect 4610 13088 4930 13089
rect 0 12928 480 13048
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4930 13088
rect 4610 13023 4930 13024
rect 11944 13088 12264 13089
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 13023 12264 13024
rect 19277 13088 19597 13089
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 19277 13023 19597 13024
rect 6085 12882 6151 12885
rect 16113 12882 16179 12885
rect 6085 12880 16179 12882
rect 6085 12824 6090 12880
rect 6146 12824 16118 12880
rect 16174 12824 16179 12880
rect 6085 12822 16179 12824
rect 6085 12819 6151 12822
rect 16113 12819 16179 12822
rect 21520 12656 22000 12776
rect 8277 12544 8597 12545
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 12479 8597 12480
rect 15610 12544 15930 12545
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 12479 15930 12480
rect 6085 12474 6151 12477
rect 62 12472 6151 12474
rect 62 12416 6090 12472
rect 6146 12416 6151 12472
rect 62 12414 6151 12416
rect 62 11960 122 12414
rect 6085 12411 6151 12414
rect 8753 12202 8819 12205
rect 15193 12202 15259 12205
rect 8753 12200 15259 12202
rect 8753 12144 8758 12200
rect 8814 12144 15198 12200
rect 15254 12144 15259 12200
rect 8753 12142 15259 12144
rect 8753 12139 8819 12142
rect 15193 12139 15259 12142
rect 20069 12202 20135 12205
rect 21590 12202 21650 12656
rect 20069 12200 21650 12202
rect 20069 12144 20074 12200
rect 20130 12144 21650 12200
rect 20069 12142 21650 12144
rect 20069 12139 20135 12142
rect 4610 12000 4930 12001
rect 0 11840 480 11960
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4930 12000
rect 4610 11935 4930 11936
rect 11944 12000 12264 12001
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 11935 12264 11936
rect 19277 12000 19597 12001
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 11935 19597 11936
rect 15193 11930 15259 11933
rect 17125 11930 17191 11933
rect 15193 11928 17191 11930
rect 15193 11872 15198 11928
rect 15254 11872 17130 11928
rect 17186 11872 17191 11928
rect 15193 11870 17191 11872
rect 15193 11867 15259 11870
rect 17125 11867 17191 11870
rect 11881 11794 11947 11797
rect 17309 11794 17375 11797
rect 11881 11792 17375 11794
rect 11881 11736 11886 11792
rect 11942 11736 17314 11792
rect 17370 11736 17375 11792
rect 11881 11734 17375 11736
rect 11881 11731 11947 11734
rect 17309 11731 17375 11734
rect 11329 11658 11395 11661
rect 18965 11658 19031 11661
rect 11329 11656 19031 11658
rect 11329 11600 11334 11656
rect 11390 11600 18970 11656
rect 19026 11600 19031 11656
rect 11329 11598 19031 11600
rect 11329 11595 11395 11598
rect 18965 11595 19031 11598
rect 9397 11522 9463 11525
rect 15009 11522 15075 11525
rect 9397 11520 15075 11522
rect 9397 11464 9402 11520
rect 9458 11464 15014 11520
rect 15070 11464 15075 11520
rect 9397 11462 15075 11464
rect 9397 11459 9463 11462
rect 15009 11459 15075 11462
rect 8277 11456 8597 11457
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 11391 8597 11392
rect 15610 11456 15930 11457
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 15610 11391 15930 11392
rect 2630 11188 2636 11252
rect 2700 11250 2706 11252
rect 3785 11250 3851 11253
rect 2700 11248 3851 11250
rect 2700 11192 3790 11248
rect 3846 11192 3851 11248
rect 2700 11190 3851 11192
rect 2700 11188 2706 11190
rect 3785 11187 3851 11190
rect 4102 11188 4108 11252
rect 4172 11250 4178 11252
rect 17769 11250 17835 11253
rect 4172 11248 17835 11250
rect 4172 11192 17774 11248
rect 17830 11192 17835 11248
rect 4172 11190 17835 11192
rect 4172 11188 4178 11190
rect 17769 11187 17835 11190
rect 20437 11250 20503 11253
rect 21582 11250 21588 11252
rect 20437 11248 21588 11250
rect 20437 11192 20442 11248
rect 20498 11192 21588 11248
rect 20437 11190 21588 11192
rect 20437 11187 20503 11190
rect 21582 11188 21588 11190
rect 21652 11188 21658 11252
rect 0 10888 480 11008
rect 21520 10980 22000 11008
rect 21520 10978 21588 10980
rect 21460 10918 21588 10978
rect 21520 10916 21588 10918
rect 21652 10916 22000 10980
rect 4610 10912 4930 10913
rect 62 10570 122 10888
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4930 10912
rect 4610 10847 4930 10848
rect 11944 10912 12264 10913
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11944 10847 12264 10848
rect 19277 10912 19597 10913
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 21520 10888 22000 10916
rect 19277 10847 19597 10848
rect 3141 10570 3207 10573
rect 12341 10570 12407 10573
rect 62 10568 12407 10570
rect 62 10512 3146 10568
rect 3202 10512 12346 10568
rect 12402 10512 12407 10568
rect 62 10510 12407 10512
rect 3141 10507 3207 10510
rect 12341 10507 12407 10510
rect 4337 10434 4403 10437
rect 4470 10434 4476 10436
rect 4337 10432 4476 10434
rect 4337 10376 4342 10432
rect 4398 10376 4476 10432
rect 4337 10374 4476 10376
rect 4337 10371 4403 10374
rect 4470 10372 4476 10374
rect 4540 10372 4546 10436
rect 8277 10368 8597 10369
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 10303 8597 10304
rect 15610 10368 15930 10369
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 10303 15930 10304
rect 6913 10162 6979 10165
rect 14457 10162 14523 10165
rect 14641 10162 14707 10165
rect 6913 10160 14707 10162
rect 6913 10104 6918 10160
rect 6974 10104 14462 10160
rect 14518 10104 14646 10160
rect 14702 10104 14707 10160
rect 6913 10102 14707 10104
rect 6913 10099 6979 10102
rect 14457 10099 14523 10102
rect 14641 10099 14707 10102
rect 3417 10026 3483 10029
rect 10501 10026 10567 10029
rect 3417 10024 10567 10026
rect 3417 9968 3422 10024
rect 3478 9968 10506 10024
rect 10562 9968 10567 10024
rect 3417 9966 10567 9968
rect 3417 9963 3483 9966
rect 10501 9963 10567 9966
rect 17585 10026 17651 10029
rect 19701 10026 19767 10029
rect 17585 10024 21650 10026
rect 17585 9968 17590 10024
rect 17646 9968 19706 10024
rect 19762 9968 21650 10024
rect 17585 9966 21650 9968
rect 17585 9963 17651 9966
rect 19701 9963 19767 9966
rect 0 9888 480 9920
rect 0 9832 110 9888
rect 166 9832 480 9888
rect 0 9800 480 9832
rect 4610 9824 4930 9825
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4930 9824
rect 4610 9759 4930 9760
rect 11944 9824 12264 9825
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 11944 9759 12264 9760
rect 19277 9824 19597 9825
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 19277 9759 19597 9760
rect 9029 9618 9095 9621
rect 18137 9618 18203 9621
rect 9029 9616 18203 9618
rect 9029 9560 9034 9616
rect 9090 9560 18142 9616
rect 18198 9560 18203 9616
rect 9029 9558 18203 9560
rect 9029 9555 9095 9558
rect 18137 9555 18203 9558
rect 8017 9482 8083 9485
rect 19609 9482 19675 9485
rect 8017 9480 19675 9482
rect 8017 9424 8022 9480
rect 8078 9424 19614 9480
rect 19670 9424 19675 9480
rect 8017 9422 19675 9424
rect 8017 9419 8083 9422
rect 19609 9419 19675 9422
rect 21590 9376 21650 9966
rect 8277 9280 8597 9281
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 8277 9215 8597 9216
rect 15610 9280 15930 9281
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 21520 9256 22000 9376
rect 15610 9215 15930 9216
rect 5441 9210 5507 9213
rect 5574 9210 5580 9212
rect 5441 9208 5580 9210
rect 5441 9152 5446 9208
rect 5502 9152 5580 9208
rect 5441 9150 5580 9152
rect 5441 9147 5507 9150
rect 5574 9148 5580 9150
rect 5644 9148 5650 9212
rect 16246 9148 16252 9212
rect 16316 9210 16322 9212
rect 16573 9210 16639 9213
rect 16316 9208 16639 9210
rect 16316 9152 16578 9208
rect 16634 9152 16639 9208
rect 16316 9150 16639 9152
rect 16316 9148 16322 9150
rect 16573 9147 16639 9150
rect 2497 9074 2563 9077
rect 7649 9074 7715 9077
rect 2497 9072 7715 9074
rect 2497 9016 2502 9072
rect 2558 9016 7654 9072
rect 7710 9016 7715 9072
rect 2497 9014 7715 9016
rect 2497 9011 2563 9014
rect 7649 9011 7715 9014
rect 10869 9074 10935 9077
rect 18137 9074 18203 9077
rect 10869 9072 18203 9074
rect 10869 9016 10874 9072
rect 10930 9016 18142 9072
rect 18198 9016 18203 9072
rect 10869 9014 18203 9016
rect 10869 9011 10935 9014
rect 18137 9011 18203 9014
rect 1945 8938 2011 8941
rect 2313 8938 2379 8941
rect 4102 8938 4108 8940
rect 1945 8936 4108 8938
rect 1945 8880 1950 8936
rect 2006 8880 2318 8936
rect 2374 8880 4108 8936
rect 1945 8878 4108 8880
rect 1945 8875 2011 8878
rect 2313 8875 2379 8878
rect 4102 8876 4108 8878
rect 4172 8876 4178 8940
rect 9489 8938 9555 8941
rect 16941 8938 17007 8941
rect 9489 8936 17007 8938
rect 9489 8880 9494 8936
rect 9550 8880 16946 8936
rect 17002 8880 17007 8936
rect 9489 8878 17007 8880
rect 9489 8875 9555 8878
rect 16941 8875 17007 8878
rect 0 8800 480 8832
rect 0 8744 18 8800
rect 74 8744 480 8800
rect 0 8712 480 8744
rect 4610 8736 4930 8737
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4930 8736
rect 4610 8671 4930 8672
rect 11944 8736 12264 8737
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 11944 8671 12264 8672
rect 19277 8736 19597 8737
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 19277 8671 19597 8672
rect 12617 8666 12683 8669
rect 17125 8666 17191 8669
rect 12617 8664 17191 8666
rect 12617 8608 12622 8664
rect 12678 8608 17130 8664
rect 17186 8608 17191 8664
rect 12617 8606 17191 8608
rect 12617 8603 12683 8606
rect 17125 8603 17191 8606
rect 7281 8530 7347 8533
rect 18505 8530 18571 8533
rect 7281 8528 18571 8530
rect 7281 8472 7286 8528
rect 7342 8472 18510 8528
rect 18566 8472 18571 8528
rect 7281 8470 18571 8472
rect 7281 8467 7347 8470
rect 18505 8467 18571 8470
rect 18638 8468 18644 8532
rect 18708 8530 18714 8532
rect 19057 8530 19123 8533
rect 18708 8528 19123 8530
rect 18708 8472 19062 8528
rect 19118 8472 19123 8528
rect 18708 8470 19123 8472
rect 18708 8468 18714 8470
rect 19057 8467 19123 8470
rect 9581 8394 9647 8397
rect 15653 8394 15719 8397
rect 9581 8392 15719 8394
rect 9581 8336 9586 8392
rect 9642 8336 15658 8392
rect 15714 8336 15719 8392
rect 9581 8334 15719 8336
rect 9581 8331 9647 8334
rect 15653 8331 15719 8334
rect 8277 8192 8597 8193
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 8127 8597 8128
rect 15610 8192 15930 8193
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 15610 8127 15930 8128
rect 8661 7986 8727 7989
rect 16205 7986 16271 7989
rect 8661 7984 16271 7986
rect 8661 7928 8666 7984
rect 8722 7928 16210 7984
rect 16266 7928 16271 7984
rect 8661 7926 16271 7928
rect 8661 7923 8727 7926
rect 16205 7923 16271 7926
rect 0 7760 480 7880
rect 6637 7850 6703 7853
rect 15377 7850 15443 7853
rect 6637 7848 15443 7850
rect 6637 7792 6642 7848
rect 6698 7792 15382 7848
rect 15438 7792 15443 7848
rect 6637 7790 15443 7792
rect 6637 7787 6703 7790
rect 15377 7787 15443 7790
rect 62 7306 122 7760
rect 4610 7648 4930 7649
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4930 7648
rect 4610 7583 4930 7584
rect 11944 7648 12264 7649
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 7583 12264 7584
rect 19277 7648 19597 7649
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 19277 7583 19597 7584
rect 21520 7580 22000 7608
rect 21520 7578 21588 7580
rect 21460 7518 21588 7578
rect 21520 7516 21588 7518
rect 21652 7516 22000 7580
rect 21520 7488 22000 7516
rect 5625 7442 5691 7445
rect 17769 7442 17835 7445
rect 5625 7440 17835 7442
rect 5625 7384 5630 7440
rect 5686 7384 17774 7440
rect 17830 7384 17835 7440
rect 5625 7382 17835 7384
rect 5625 7379 5691 7382
rect 17769 7379 17835 7382
rect 18689 7442 18755 7445
rect 18689 7440 19350 7442
rect 18689 7384 18694 7440
rect 18750 7384 19350 7440
rect 18689 7382 19350 7384
rect 18689 7379 18755 7382
rect 3693 7306 3759 7309
rect 62 7304 3759 7306
rect 62 7248 3698 7304
rect 3754 7248 3759 7304
rect 62 7246 3759 7248
rect 3693 7243 3759 7246
rect 9213 7306 9279 7309
rect 14825 7306 14891 7309
rect 9213 7304 14891 7306
rect 9213 7248 9218 7304
rect 9274 7248 14830 7304
rect 14886 7248 14891 7304
rect 9213 7246 14891 7248
rect 19290 7306 19350 7382
rect 21582 7306 21588 7308
rect 19290 7246 21588 7306
rect 9213 7243 9279 7246
rect 14825 7243 14891 7246
rect 21582 7244 21588 7246
rect 21652 7244 21658 7308
rect 7097 7170 7163 7173
rect 7966 7170 7972 7172
rect 7097 7168 7972 7170
rect 7097 7112 7102 7168
rect 7158 7112 7972 7168
rect 7097 7110 7972 7112
rect 7097 7107 7163 7110
rect 7966 7108 7972 7110
rect 8036 7108 8042 7172
rect 8661 7170 8727 7173
rect 15285 7170 15351 7173
rect 8661 7168 15351 7170
rect 8661 7112 8666 7168
rect 8722 7112 15290 7168
rect 15346 7112 15351 7168
rect 8661 7110 15351 7112
rect 8661 7107 8727 7110
rect 15285 7107 15351 7110
rect 16614 7108 16620 7172
rect 16684 7170 16690 7172
rect 16757 7170 16823 7173
rect 16684 7168 16823 7170
rect 16684 7112 16762 7168
rect 16818 7112 16823 7168
rect 16684 7110 16823 7112
rect 16684 7108 16690 7110
rect 16757 7107 16823 7110
rect 8277 7104 8597 7105
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 8277 7039 8597 7040
rect 15610 7104 15930 7105
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 15610 7039 15930 7040
rect 54 6972 60 7036
rect 124 7034 130 7036
rect 5533 7034 5599 7037
rect 124 7032 5599 7034
rect 124 6976 5538 7032
rect 5594 6976 5599 7032
rect 124 6974 5599 6976
rect 124 6972 130 6974
rect 5533 6971 5599 6974
rect 11421 6898 11487 6901
rect 17493 6898 17559 6901
rect 11421 6896 17559 6898
rect 11421 6840 11426 6896
rect 11482 6840 17498 6896
rect 17554 6840 17559 6896
rect 11421 6838 17559 6840
rect 11421 6835 11487 6838
rect 17493 6835 17559 6838
rect 0 6764 480 6792
rect 0 6700 60 6764
rect 124 6700 480 6764
rect 0 6672 480 6700
rect 6545 6762 6611 6765
rect 7005 6762 7071 6765
rect 16665 6762 16731 6765
rect 6545 6760 16731 6762
rect 6545 6704 6550 6760
rect 6606 6704 7010 6760
rect 7066 6704 16670 6760
rect 16726 6704 16731 6760
rect 6545 6702 16731 6704
rect 6545 6699 6611 6702
rect 7005 6699 7071 6702
rect 16665 6699 16731 6702
rect 13629 6626 13695 6629
rect 16573 6626 16639 6629
rect 13629 6624 16639 6626
rect 13629 6568 13634 6624
rect 13690 6568 16578 6624
rect 16634 6568 16639 6624
rect 13629 6566 16639 6568
rect 13629 6563 13695 6566
rect 16573 6563 16639 6566
rect 4610 6560 4930 6561
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4930 6560
rect 4610 6495 4930 6496
rect 11944 6560 12264 6561
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 6495 12264 6496
rect 19277 6560 19597 6561
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 6495 19597 6496
rect 3417 6490 3483 6493
rect 3550 6490 3556 6492
rect 3417 6488 3556 6490
rect 3417 6432 3422 6488
rect 3478 6432 3556 6488
rect 3417 6430 3556 6432
rect 3417 6427 3483 6430
rect 3550 6428 3556 6430
rect 3620 6428 3626 6492
rect 14273 6490 14339 6493
rect 14273 6488 16452 6490
rect 14273 6432 14278 6488
rect 14334 6432 16452 6488
rect 14273 6430 16452 6432
rect 14273 6427 14339 6430
rect 4981 6354 5047 6357
rect 7465 6354 7531 6357
rect 14549 6354 14615 6357
rect 4981 6352 14615 6354
rect 4981 6296 4986 6352
rect 5042 6296 7470 6352
rect 7526 6296 14554 6352
rect 14610 6296 14615 6352
rect 4981 6294 14615 6296
rect 4981 6291 5047 6294
rect 7465 6291 7531 6294
rect 14549 6291 14615 6294
rect 14825 6354 14891 6357
rect 16205 6354 16271 6357
rect 14825 6352 16271 6354
rect 14825 6296 14830 6352
rect 14886 6296 16210 6352
rect 16266 6296 16271 6352
rect 14825 6294 16271 6296
rect 16392 6354 16452 6430
rect 16392 6294 21650 6354
rect 14825 6291 14891 6294
rect 16205 6291 16271 6294
rect 1945 6218 2011 6221
rect 62 6216 2011 6218
rect 62 6160 1950 6216
rect 2006 6160 2011 6216
rect 62 6158 2011 6160
rect 62 5704 122 6158
rect 1945 6155 2011 6158
rect 2681 6218 2747 6221
rect 7189 6218 7255 6221
rect 2681 6216 7255 6218
rect 2681 6160 2686 6216
rect 2742 6160 7194 6216
rect 7250 6160 7255 6216
rect 2681 6158 7255 6160
rect 2681 6155 2747 6158
rect 7189 6155 7255 6158
rect 9397 6218 9463 6221
rect 17309 6218 17375 6221
rect 9397 6216 17375 6218
rect 9397 6160 9402 6216
rect 9458 6160 17314 6216
rect 17370 6160 17375 6216
rect 9397 6158 17375 6160
rect 9397 6155 9463 6158
rect 17309 6155 17375 6158
rect 8753 6082 8819 6085
rect 15377 6082 15443 6085
rect 8753 6080 15443 6082
rect 8753 6024 8758 6080
rect 8814 6024 15382 6080
rect 15438 6024 15443 6080
rect 8753 6022 15443 6024
rect 8753 6019 8819 6022
rect 15377 6019 15443 6022
rect 8277 6016 8597 6017
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 8277 5951 8597 5952
rect 15610 6016 15930 6017
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 21590 5976 21650 6294
rect 15610 5951 15930 5952
rect 21520 5856 22000 5976
rect 11237 5810 11303 5813
rect 18965 5810 19031 5813
rect 11237 5808 19031 5810
rect 11237 5752 11242 5808
rect 11298 5752 18970 5808
rect 19026 5752 19031 5808
rect 11237 5750 19031 5752
rect 11237 5747 11303 5750
rect 18965 5747 19031 5750
rect 0 5584 480 5704
rect 4610 5472 4930 5473
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4930 5472
rect 4610 5407 4930 5408
rect 11944 5472 12264 5473
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 11944 5407 12264 5408
rect 19277 5472 19597 5473
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 19277 5407 19597 5408
rect 7414 5340 7420 5404
rect 7484 5402 7490 5404
rect 7557 5402 7623 5405
rect 7484 5400 7623 5402
rect 7484 5344 7562 5400
rect 7618 5344 7623 5400
rect 7484 5342 7623 5344
rect 7484 5340 7490 5342
rect 7557 5339 7623 5342
rect 1577 5266 1643 5269
rect 3233 5266 3299 5269
rect 11053 5266 11119 5269
rect 1577 5264 11119 5266
rect 1577 5208 1582 5264
rect 1638 5208 3238 5264
rect 3294 5208 11058 5264
rect 11114 5208 11119 5264
rect 1577 5206 11119 5208
rect 1577 5203 1643 5206
rect 3233 5203 3299 5206
rect 11053 5203 11119 5206
rect 4102 5068 4108 5132
rect 4172 5130 4178 5132
rect 18045 5130 18111 5133
rect 4172 5128 18111 5130
rect 4172 5072 18050 5128
rect 18106 5072 18111 5128
rect 4172 5070 18111 5072
rect 4172 5068 4178 5070
rect 18045 5067 18111 5070
rect 1669 4994 1735 4997
rect 1894 4994 1900 4996
rect 1669 4992 1900 4994
rect 1669 4936 1674 4992
rect 1730 4936 1900 4992
rect 1669 4934 1900 4936
rect 1669 4931 1735 4934
rect 1894 4932 1900 4934
rect 1964 4932 1970 4996
rect 8277 4928 8597 4929
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 8277 4863 8597 4864
rect 15610 4928 15930 4929
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 15610 4863 15930 4864
rect 6453 4858 6519 4861
rect 62 4856 6519 4858
rect 62 4800 6458 4856
rect 6514 4800 6519 4856
rect 62 4798 6519 4800
rect 62 4616 122 4798
rect 6453 4795 6519 4798
rect 6361 4722 6427 4725
rect 15469 4722 15535 4725
rect 6361 4720 15535 4722
rect 6361 4664 6366 4720
rect 6422 4664 15474 4720
rect 15530 4664 15535 4720
rect 6361 4662 15535 4664
rect 6361 4659 6427 4662
rect 15469 4659 15535 4662
rect 0 4496 480 4616
rect 4153 4586 4219 4589
rect 5165 4586 5231 4589
rect 4153 4584 5231 4586
rect 4153 4528 4158 4584
rect 4214 4528 5170 4584
rect 5226 4528 5231 4584
rect 4153 4526 5231 4528
rect 4153 4523 4219 4526
rect 5165 4523 5231 4526
rect 9622 4524 9628 4588
rect 9692 4586 9698 4588
rect 15929 4586 15995 4589
rect 9692 4584 15995 4586
rect 9692 4528 15934 4584
rect 15990 4528 15995 4584
rect 9692 4526 15995 4528
rect 9692 4524 9698 4526
rect 15929 4523 15995 4526
rect 4610 4384 4930 4385
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4930 4384
rect 4610 4319 4930 4320
rect 11944 4384 12264 4385
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 11944 4319 12264 4320
rect 19277 4384 19597 4385
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 19277 4319 19597 4320
rect 6913 4178 6979 4181
rect 16297 4178 16363 4181
rect 6913 4176 16363 4178
rect 6913 4120 6918 4176
rect 6974 4120 16302 4176
rect 16358 4120 16363 4176
rect 6913 4118 16363 4120
rect 6913 4115 6979 4118
rect 16297 4115 16363 4118
rect 21520 4176 22000 4208
rect 21520 4120 21638 4176
rect 21694 4120 22000 4176
rect 21520 4088 22000 4120
rect 1853 4042 1919 4045
rect 6729 4042 6795 4045
rect 11237 4042 11303 4045
rect 1853 4040 11303 4042
rect 1853 3984 1858 4040
rect 1914 3984 6734 4040
rect 6790 3984 11242 4040
rect 11298 3984 11303 4040
rect 1853 3982 11303 3984
rect 1853 3979 1919 3982
rect 6729 3979 6795 3982
rect 11237 3979 11303 3982
rect 8277 3840 8597 3841
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 8277 3775 8597 3776
rect 15610 3840 15930 3841
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 15610 3775 15930 3776
rect 4286 3708 4292 3772
rect 4356 3770 4362 3772
rect 4521 3770 4587 3773
rect 4356 3768 4587 3770
rect 4356 3712 4526 3768
rect 4582 3712 4587 3768
rect 4356 3710 4587 3712
rect 4356 3708 4362 3710
rect 4521 3707 4587 3710
rect 0 3632 480 3664
rect 0 3576 110 3632
rect 166 3576 480 3632
rect 0 3544 480 3576
rect 2773 3634 2839 3637
rect 9121 3634 9187 3637
rect 2773 3632 9187 3634
rect 2773 3576 2778 3632
rect 2834 3576 9126 3632
rect 9182 3576 9187 3632
rect 2773 3574 9187 3576
rect 2773 3571 2839 3574
rect 9121 3571 9187 3574
rect 6453 3498 6519 3501
rect 12617 3498 12683 3501
rect 6453 3496 12683 3498
rect 6453 3440 6458 3496
rect 6514 3440 12622 3496
rect 12678 3440 12683 3496
rect 6453 3438 12683 3440
rect 6453 3435 6519 3438
rect 12617 3435 12683 3438
rect 4610 3296 4930 3297
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4930 3296
rect 4610 3231 4930 3232
rect 11944 3296 12264 3297
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 3231 12264 3232
rect 19277 3296 19597 3297
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 19277 3231 19597 3232
rect 18321 3226 18387 3229
rect 12390 3224 18387 3226
rect 12390 3168 18326 3224
rect 18382 3168 18387 3224
rect 12390 3166 18387 3168
rect 6545 3090 6611 3093
rect 12390 3090 12450 3166
rect 18321 3163 18387 3166
rect 6545 3088 12450 3090
rect 6545 3032 6550 3088
rect 6606 3032 12450 3088
rect 6545 3030 12450 3032
rect 12525 3090 12591 3093
rect 17953 3090 18019 3093
rect 12525 3088 18019 3090
rect 12525 3032 12530 3088
rect 12586 3032 17958 3088
rect 18014 3032 18019 3088
rect 12525 3030 18019 3032
rect 6545 3027 6611 3030
rect 12525 3027 12591 3030
rect 17953 3027 18019 3030
rect 5993 2954 6059 2957
rect 16113 2954 16179 2957
rect 5993 2952 16179 2954
rect 5993 2896 5998 2952
rect 6054 2896 16118 2952
rect 16174 2896 16179 2952
rect 5993 2894 16179 2896
rect 5993 2891 6059 2894
rect 16113 2891 16179 2894
rect 18229 2954 18295 2957
rect 18229 2952 21650 2954
rect 18229 2896 18234 2952
rect 18290 2896 21650 2952
rect 18229 2894 21650 2896
rect 18229 2891 18295 2894
rect 8277 2752 8597 2753
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2687 8597 2688
rect 15610 2752 15930 2753
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 15610 2687 15930 2688
rect 9397 2682 9463 2685
rect 9397 2680 12818 2682
rect 9397 2624 9402 2680
rect 9458 2624 12818 2680
rect 9397 2622 12818 2624
rect 9397 2619 9463 2622
rect 0 2544 480 2576
rect 0 2488 110 2544
rect 166 2488 480 2544
rect 0 2456 480 2488
rect 5717 2546 5783 2549
rect 12525 2546 12591 2549
rect 5717 2544 12591 2546
rect 5717 2488 5722 2544
rect 5778 2488 12530 2544
rect 12586 2488 12591 2544
rect 5717 2486 12591 2488
rect 12758 2546 12818 2622
rect 21590 2576 21650 2894
rect 16481 2546 16547 2549
rect 12758 2544 16547 2546
rect 12758 2488 16486 2544
rect 16542 2488 16547 2544
rect 12758 2486 16547 2488
rect 5717 2483 5783 2486
rect 12525 2483 12591 2486
rect 16481 2483 16547 2486
rect 21520 2456 22000 2576
rect 8661 2410 8727 2413
rect 15561 2410 15627 2413
rect 8661 2408 15627 2410
rect 8661 2352 8666 2408
rect 8722 2352 15566 2408
rect 15622 2352 15627 2408
rect 8661 2350 15627 2352
rect 8661 2347 8727 2350
rect 15561 2347 15627 2350
rect 4610 2208 4930 2209
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4930 2208
rect 4610 2143 4930 2144
rect 11944 2208 12264 2209
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2143 12264 2144
rect 19277 2208 19597 2209
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2143 19597 2144
rect 3049 2002 3115 2005
rect 62 2000 3115 2002
rect 62 1944 3054 2000
rect 3110 1944 3115 2000
rect 62 1942 3115 1944
rect 62 1488 122 1942
rect 3049 1939 3115 1942
rect 5533 2002 5599 2005
rect 15101 2002 15167 2005
rect 5533 2000 15167 2002
rect 5533 1944 5538 2000
rect 5594 1944 15106 2000
rect 15162 1944 15167 2000
rect 5533 1942 15167 1944
rect 5533 1939 5599 1942
rect 15101 1939 15167 1942
rect 5073 1730 5139 1733
rect 15193 1730 15259 1733
rect 5073 1728 16498 1730
rect 5073 1672 5078 1728
rect 5134 1672 15198 1728
rect 15254 1672 16498 1728
rect 5073 1670 16498 1672
rect 5073 1667 5139 1670
rect 15193 1667 15259 1670
rect 6177 1594 6243 1597
rect 14825 1594 14891 1597
rect 6177 1592 14891 1594
rect 6177 1536 6182 1592
rect 6238 1536 14830 1592
rect 14886 1536 14891 1592
rect 6177 1534 14891 1536
rect 16438 1594 16498 1670
rect 17902 1668 17908 1732
rect 17972 1730 17978 1732
rect 18045 1730 18111 1733
rect 17972 1728 18111 1730
rect 17972 1672 18050 1728
rect 18106 1672 18111 1728
rect 17972 1670 18111 1672
rect 17972 1668 17978 1670
rect 18045 1667 18111 1670
rect 16438 1534 21650 1594
rect 6177 1531 6243 1534
rect 14825 1531 14891 1534
rect 0 1368 480 1488
rect 6453 1458 6519 1461
rect 19057 1458 19123 1461
rect 6453 1456 19123 1458
rect 6453 1400 6458 1456
rect 6514 1400 19062 1456
rect 19118 1400 19123 1456
rect 6453 1398 19123 1400
rect 6453 1395 6519 1398
rect 19057 1395 19123 1398
rect 6637 1322 6703 1325
rect 17769 1322 17835 1325
rect 6637 1320 17835 1322
rect 6637 1264 6642 1320
rect 6698 1264 17774 1320
rect 17830 1264 17835 1320
rect 6637 1262 17835 1264
rect 6637 1259 6703 1262
rect 17769 1259 17835 1262
rect 1669 1050 1735 1053
rect 62 1048 1735 1050
rect 62 992 1674 1048
rect 1730 992 1735 1048
rect 62 990 1735 992
rect 62 536 122 990
rect 1669 987 1735 990
rect 21590 944 21650 1534
rect 21520 824 22000 944
rect 0 416 480 536
rect 841 98 907 101
rect 4102 98 4108 100
rect 841 96 4108 98
rect 841 40 846 96
rect 902 40 4108 96
rect 841 38 4108 40
rect 841 35 907 38
rect 4102 36 4108 38
rect 4172 36 4178 100
<< via3 >>
rect 2636 21524 2700 21588
rect 4618 19612 4682 19616
rect 4618 19556 4622 19612
rect 4622 19556 4678 19612
rect 4678 19556 4682 19612
rect 4618 19552 4682 19556
rect 4698 19612 4762 19616
rect 4698 19556 4702 19612
rect 4702 19556 4758 19612
rect 4758 19556 4762 19612
rect 4698 19552 4762 19556
rect 4778 19612 4842 19616
rect 4778 19556 4782 19612
rect 4782 19556 4838 19612
rect 4838 19556 4842 19612
rect 4778 19552 4842 19556
rect 4858 19612 4922 19616
rect 4858 19556 4862 19612
rect 4862 19556 4918 19612
rect 4918 19556 4922 19612
rect 4858 19552 4922 19556
rect 11952 19612 12016 19616
rect 11952 19556 11956 19612
rect 11956 19556 12012 19612
rect 12012 19556 12016 19612
rect 11952 19552 12016 19556
rect 12032 19612 12096 19616
rect 12032 19556 12036 19612
rect 12036 19556 12092 19612
rect 12092 19556 12096 19612
rect 12032 19552 12096 19556
rect 12112 19612 12176 19616
rect 12112 19556 12116 19612
rect 12116 19556 12172 19612
rect 12172 19556 12176 19612
rect 12112 19552 12176 19556
rect 12192 19612 12256 19616
rect 12192 19556 12196 19612
rect 12196 19556 12252 19612
rect 12252 19556 12256 19612
rect 12192 19552 12256 19556
rect 19285 19612 19349 19616
rect 19285 19556 19289 19612
rect 19289 19556 19345 19612
rect 19345 19556 19349 19612
rect 19285 19552 19349 19556
rect 19365 19612 19429 19616
rect 19365 19556 19369 19612
rect 19369 19556 19425 19612
rect 19425 19556 19429 19612
rect 19365 19552 19429 19556
rect 19445 19612 19509 19616
rect 19445 19556 19449 19612
rect 19449 19556 19505 19612
rect 19505 19556 19509 19612
rect 19445 19552 19509 19556
rect 19525 19612 19589 19616
rect 19525 19556 19529 19612
rect 19529 19556 19585 19612
rect 19585 19556 19589 19612
rect 19525 19552 19589 19556
rect 8285 19068 8349 19072
rect 8285 19012 8289 19068
rect 8289 19012 8345 19068
rect 8345 19012 8349 19068
rect 8285 19008 8349 19012
rect 8365 19068 8429 19072
rect 8365 19012 8369 19068
rect 8369 19012 8425 19068
rect 8425 19012 8429 19068
rect 8365 19008 8429 19012
rect 8445 19068 8509 19072
rect 8445 19012 8449 19068
rect 8449 19012 8505 19068
rect 8505 19012 8509 19068
rect 8445 19008 8509 19012
rect 8525 19068 8589 19072
rect 8525 19012 8529 19068
rect 8529 19012 8585 19068
rect 8585 19012 8589 19068
rect 8525 19008 8589 19012
rect 15618 19068 15682 19072
rect 15618 19012 15622 19068
rect 15622 19012 15678 19068
rect 15678 19012 15682 19068
rect 15618 19008 15682 19012
rect 15698 19068 15762 19072
rect 15698 19012 15702 19068
rect 15702 19012 15758 19068
rect 15758 19012 15762 19068
rect 15698 19008 15762 19012
rect 15778 19068 15842 19072
rect 15778 19012 15782 19068
rect 15782 19012 15838 19068
rect 15838 19012 15842 19068
rect 15778 19008 15842 19012
rect 15858 19068 15922 19072
rect 15858 19012 15862 19068
rect 15862 19012 15918 19068
rect 15918 19012 15922 19068
rect 15858 19008 15922 19012
rect 4618 18524 4682 18528
rect 4618 18468 4622 18524
rect 4622 18468 4678 18524
rect 4678 18468 4682 18524
rect 4618 18464 4682 18468
rect 4698 18524 4762 18528
rect 4698 18468 4702 18524
rect 4702 18468 4758 18524
rect 4758 18468 4762 18524
rect 4698 18464 4762 18468
rect 4778 18524 4842 18528
rect 4778 18468 4782 18524
rect 4782 18468 4838 18524
rect 4838 18468 4842 18524
rect 4778 18464 4842 18468
rect 4858 18524 4922 18528
rect 4858 18468 4862 18524
rect 4862 18468 4918 18524
rect 4918 18468 4922 18524
rect 4858 18464 4922 18468
rect 11952 18524 12016 18528
rect 11952 18468 11956 18524
rect 11956 18468 12012 18524
rect 12012 18468 12016 18524
rect 11952 18464 12016 18468
rect 12032 18524 12096 18528
rect 12032 18468 12036 18524
rect 12036 18468 12092 18524
rect 12092 18468 12096 18524
rect 12032 18464 12096 18468
rect 12112 18524 12176 18528
rect 12112 18468 12116 18524
rect 12116 18468 12172 18524
rect 12172 18468 12176 18524
rect 12112 18464 12176 18468
rect 12192 18524 12256 18528
rect 12192 18468 12196 18524
rect 12196 18468 12252 18524
rect 12252 18468 12256 18524
rect 12192 18464 12256 18468
rect 19285 18524 19349 18528
rect 19285 18468 19289 18524
rect 19289 18468 19345 18524
rect 19345 18468 19349 18524
rect 19285 18464 19349 18468
rect 19365 18524 19429 18528
rect 19365 18468 19369 18524
rect 19369 18468 19425 18524
rect 19425 18468 19429 18524
rect 19365 18464 19429 18468
rect 19445 18524 19509 18528
rect 19445 18468 19449 18524
rect 19449 18468 19505 18524
rect 19505 18468 19509 18524
rect 19445 18464 19509 18468
rect 19525 18524 19589 18528
rect 19525 18468 19529 18524
rect 19529 18468 19585 18524
rect 19585 18468 19589 18524
rect 19525 18464 19589 18468
rect 8285 17980 8349 17984
rect 8285 17924 8289 17980
rect 8289 17924 8345 17980
rect 8345 17924 8349 17980
rect 8285 17920 8349 17924
rect 8365 17980 8429 17984
rect 8365 17924 8369 17980
rect 8369 17924 8425 17980
rect 8425 17924 8429 17980
rect 8365 17920 8429 17924
rect 8445 17980 8509 17984
rect 8445 17924 8449 17980
rect 8449 17924 8505 17980
rect 8505 17924 8509 17980
rect 8445 17920 8509 17924
rect 8525 17980 8589 17984
rect 8525 17924 8529 17980
rect 8529 17924 8585 17980
rect 8585 17924 8589 17980
rect 8525 17920 8589 17924
rect 15618 17980 15682 17984
rect 15618 17924 15622 17980
rect 15622 17924 15678 17980
rect 15678 17924 15682 17980
rect 15618 17920 15682 17924
rect 15698 17980 15762 17984
rect 15698 17924 15702 17980
rect 15702 17924 15758 17980
rect 15758 17924 15762 17980
rect 15698 17920 15762 17924
rect 15778 17980 15842 17984
rect 15778 17924 15782 17980
rect 15782 17924 15838 17980
rect 15838 17924 15842 17980
rect 15778 17920 15842 17924
rect 15858 17980 15922 17984
rect 15858 17924 15862 17980
rect 15862 17924 15918 17980
rect 15918 17924 15922 17980
rect 15858 17920 15922 17924
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 4698 17436 4762 17440
rect 4698 17380 4702 17436
rect 4702 17380 4758 17436
rect 4758 17380 4762 17436
rect 4698 17376 4762 17380
rect 4778 17436 4842 17440
rect 4778 17380 4782 17436
rect 4782 17380 4838 17436
rect 4838 17380 4842 17436
rect 4778 17376 4842 17380
rect 4858 17436 4922 17440
rect 4858 17380 4862 17436
rect 4862 17380 4918 17436
rect 4918 17380 4922 17436
rect 4858 17376 4922 17380
rect 11952 17436 12016 17440
rect 11952 17380 11956 17436
rect 11956 17380 12012 17436
rect 12012 17380 12016 17436
rect 11952 17376 12016 17380
rect 12032 17436 12096 17440
rect 12032 17380 12036 17436
rect 12036 17380 12092 17436
rect 12092 17380 12096 17436
rect 12032 17376 12096 17380
rect 12112 17436 12176 17440
rect 12112 17380 12116 17436
rect 12116 17380 12172 17436
rect 12172 17380 12176 17436
rect 12112 17376 12176 17380
rect 12192 17436 12256 17440
rect 12192 17380 12196 17436
rect 12196 17380 12252 17436
rect 12252 17380 12256 17436
rect 12192 17376 12256 17380
rect 19285 17436 19349 17440
rect 19285 17380 19289 17436
rect 19289 17380 19345 17436
rect 19345 17380 19349 17436
rect 19285 17376 19349 17380
rect 19365 17436 19429 17440
rect 19365 17380 19369 17436
rect 19369 17380 19425 17436
rect 19425 17380 19429 17436
rect 19365 17376 19429 17380
rect 19445 17436 19509 17440
rect 19445 17380 19449 17436
rect 19449 17380 19505 17436
rect 19505 17380 19509 17436
rect 19445 17376 19509 17380
rect 19525 17436 19589 17440
rect 19525 17380 19529 17436
rect 19529 17380 19585 17436
rect 19585 17380 19589 17436
rect 19525 17376 19589 17380
rect 8285 16892 8349 16896
rect 8285 16836 8289 16892
rect 8289 16836 8345 16892
rect 8345 16836 8349 16892
rect 8285 16832 8349 16836
rect 8365 16892 8429 16896
rect 8365 16836 8369 16892
rect 8369 16836 8425 16892
rect 8425 16836 8429 16892
rect 8365 16832 8429 16836
rect 8445 16892 8509 16896
rect 8445 16836 8449 16892
rect 8449 16836 8505 16892
rect 8505 16836 8509 16892
rect 8445 16832 8509 16836
rect 8525 16892 8589 16896
rect 8525 16836 8529 16892
rect 8529 16836 8585 16892
rect 8585 16836 8589 16892
rect 8525 16832 8589 16836
rect 15618 16892 15682 16896
rect 15618 16836 15622 16892
rect 15622 16836 15678 16892
rect 15678 16836 15682 16892
rect 15618 16832 15682 16836
rect 15698 16892 15762 16896
rect 15698 16836 15702 16892
rect 15702 16836 15758 16892
rect 15758 16836 15762 16892
rect 15698 16832 15762 16836
rect 15778 16892 15842 16896
rect 15778 16836 15782 16892
rect 15782 16836 15838 16892
rect 15838 16836 15842 16892
rect 15778 16832 15842 16836
rect 15858 16892 15922 16896
rect 15858 16836 15862 16892
rect 15862 16836 15918 16892
rect 15918 16836 15922 16892
rect 15858 16832 15922 16836
rect 60 16356 124 16420
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 4698 16348 4762 16352
rect 4698 16292 4702 16348
rect 4702 16292 4758 16348
rect 4758 16292 4762 16348
rect 4698 16288 4762 16292
rect 4778 16348 4842 16352
rect 4778 16292 4782 16348
rect 4782 16292 4838 16348
rect 4838 16292 4842 16348
rect 4778 16288 4842 16292
rect 4858 16348 4922 16352
rect 4858 16292 4862 16348
rect 4862 16292 4918 16348
rect 4918 16292 4922 16348
rect 4858 16288 4922 16292
rect 11952 16348 12016 16352
rect 11952 16292 11956 16348
rect 11956 16292 12012 16348
rect 12012 16292 12016 16348
rect 11952 16288 12016 16292
rect 12032 16348 12096 16352
rect 12032 16292 12036 16348
rect 12036 16292 12092 16348
rect 12092 16292 12096 16348
rect 12032 16288 12096 16292
rect 12112 16348 12176 16352
rect 12112 16292 12116 16348
rect 12116 16292 12172 16348
rect 12172 16292 12176 16348
rect 12112 16288 12176 16292
rect 12192 16348 12256 16352
rect 12192 16292 12196 16348
rect 12196 16292 12252 16348
rect 12252 16292 12256 16348
rect 12192 16288 12256 16292
rect 19285 16348 19349 16352
rect 19285 16292 19289 16348
rect 19289 16292 19345 16348
rect 19345 16292 19349 16348
rect 19285 16288 19349 16292
rect 19365 16348 19429 16352
rect 19365 16292 19369 16348
rect 19369 16292 19425 16348
rect 19425 16292 19429 16348
rect 19365 16288 19429 16292
rect 19445 16348 19509 16352
rect 19445 16292 19449 16348
rect 19449 16292 19505 16348
rect 19505 16292 19509 16348
rect 19445 16288 19509 16292
rect 19525 16348 19589 16352
rect 19525 16292 19529 16348
rect 19529 16292 19585 16348
rect 19585 16292 19589 16348
rect 19525 16288 19589 16292
rect 60 16084 124 16148
rect 8285 15804 8349 15808
rect 8285 15748 8289 15804
rect 8289 15748 8345 15804
rect 8345 15748 8349 15804
rect 8285 15744 8349 15748
rect 8365 15804 8429 15808
rect 8365 15748 8369 15804
rect 8369 15748 8425 15804
rect 8425 15748 8429 15804
rect 8365 15744 8429 15748
rect 8445 15804 8509 15808
rect 8445 15748 8449 15804
rect 8449 15748 8505 15804
rect 8505 15748 8509 15804
rect 8445 15744 8509 15748
rect 8525 15804 8589 15808
rect 8525 15748 8529 15804
rect 8529 15748 8585 15804
rect 8585 15748 8589 15804
rect 8525 15744 8589 15748
rect 15618 15804 15682 15808
rect 15618 15748 15622 15804
rect 15622 15748 15678 15804
rect 15678 15748 15682 15804
rect 15618 15744 15682 15748
rect 15698 15804 15762 15808
rect 15698 15748 15702 15804
rect 15702 15748 15758 15804
rect 15758 15748 15762 15804
rect 15698 15744 15762 15748
rect 15778 15804 15842 15808
rect 15778 15748 15782 15804
rect 15782 15748 15838 15804
rect 15838 15748 15842 15804
rect 15778 15744 15842 15748
rect 15858 15804 15922 15808
rect 15858 15748 15862 15804
rect 15862 15748 15918 15804
rect 15918 15748 15922 15804
rect 15858 15744 15922 15748
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 4698 15260 4762 15264
rect 4698 15204 4702 15260
rect 4702 15204 4758 15260
rect 4758 15204 4762 15260
rect 4698 15200 4762 15204
rect 4778 15260 4842 15264
rect 4778 15204 4782 15260
rect 4782 15204 4838 15260
rect 4838 15204 4842 15260
rect 4778 15200 4842 15204
rect 4858 15260 4922 15264
rect 4858 15204 4862 15260
rect 4862 15204 4918 15260
rect 4918 15204 4922 15260
rect 4858 15200 4922 15204
rect 11952 15260 12016 15264
rect 11952 15204 11956 15260
rect 11956 15204 12012 15260
rect 12012 15204 12016 15260
rect 11952 15200 12016 15204
rect 12032 15260 12096 15264
rect 12032 15204 12036 15260
rect 12036 15204 12092 15260
rect 12092 15204 12096 15260
rect 12032 15200 12096 15204
rect 12112 15260 12176 15264
rect 12112 15204 12116 15260
rect 12116 15204 12172 15260
rect 12172 15204 12176 15260
rect 12112 15200 12176 15204
rect 12192 15260 12256 15264
rect 12192 15204 12196 15260
rect 12196 15204 12252 15260
rect 12252 15204 12256 15260
rect 12192 15200 12256 15204
rect 19285 15260 19349 15264
rect 19285 15204 19289 15260
rect 19289 15204 19345 15260
rect 19345 15204 19349 15260
rect 19285 15200 19349 15204
rect 19365 15260 19429 15264
rect 19365 15204 19369 15260
rect 19369 15204 19425 15260
rect 19425 15204 19429 15260
rect 19365 15200 19429 15204
rect 19445 15260 19509 15264
rect 19445 15204 19449 15260
rect 19449 15204 19505 15260
rect 19505 15204 19509 15260
rect 19445 15200 19509 15204
rect 19525 15260 19589 15264
rect 19525 15204 19529 15260
rect 19529 15204 19585 15260
rect 19585 15204 19589 15260
rect 19525 15200 19589 15204
rect 8285 14716 8349 14720
rect 8285 14660 8289 14716
rect 8289 14660 8345 14716
rect 8345 14660 8349 14716
rect 8285 14656 8349 14660
rect 8365 14716 8429 14720
rect 8365 14660 8369 14716
rect 8369 14660 8425 14716
rect 8425 14660 8429 14716
rect 8365 14656 8429 14660
rect 8445 14716 8509 14720
rect 8445 14660 8449 14716
rect 8449 14660 8505 14716
rect 8505 14660 8509 14716
rect 8445 14656 8509 14660
rect 8525 14716 8589 14720
rect 8525 14660 8529 14716
rect 8529 14660 8585 14716
rect 8585 14660 8589 14716
rect 8525 14656 8589 14660
rect 15618 14716 15682 14720
rect 15618 14660 15622 14716
rect 15622 14660 15678 14716
rect 15678 14660 15682 14716
rect 15618 14656 15682 14660
rect 15698 14716 15762 14720
rect 15698 14660 15702 14716
rect 15702 14660 15758 14716
rect 15758 14660 15762 14716
rect 15698 14656 15762 14660
rect 15778 14716 15842 14720
rect 15778 14660 15782 14716
rect 15782 14660 15838 14716
rect 15838 14660 15842 14716
rect 15778 14656 15842 14660
rect 15858 14716 15922 14720
rect 15858 14660 15862 14716
rect 15862 14660 15918 14716
rect 15918 14660 15922 14716
rect 15858 14656 15922 14660
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 4698 14172 4762 14176
rect 4698 14116 4702 14172
rect 4702 14116 4758 14172
rect 4758 14116 4762 14172
rect 4698 14112 4762 14116
rect 4778 14172 4842 14176
rect 4778 14116 4782 14172
rect 4782 14116 4838 14172
rect 4838 14116 4842 14172
rect 4778 14112 4842 14116
rect 4858 14172 4922 14176
rect 4858 14116 4862 14172
rect 4862 14116 4918 14172
rect 4918 14116 4922 14172
rect 4858 14112 4922 14116
rect 11952 14172 12016 14176
rect 11952 14116 11956 14172
rect 11956 14116 12012 14172
rect 12012 14116 12016 14172
rect 11952 14112 12016 14116
rect 12032 14172 12096 14176
rect 12032 14116 12036 14172
rect 12036 14116 12092 14172
rect 12092 14116 12096 14172
rect 12032 14112 12096 14116
rect 12112 14172 12176 14176
rect 12112 14116 12116 14172
rect 12116 14116 12172 14172
rect 12172 14116 12176 14172
rect 12112 14112 12176 14116
rect 12192 14172 12256 14176
rect 12192 14116 12196 14172
rect 12196 14116 12252 14172
rect 12252 14116 12256 14172
rect 12192 14112 12256 14116
rect 19285 14172 19349 14176
rect 19285 14116 19289 14172
rect 19289 14116 19345 14172
rect 19345 14116 19349 14172
rect 19285 14112 19349 14116
rect 19365 14172 19429 14176
rect 19365 14116 19369 14172
rect 19369 14116 19425 14172
rect 19425 14116 19429 14172
rect 19365 14112 19429 14116
rect 19445 14172 19509 14176
rect 19445 14116 19449 14172
rect 19449 14116 19505 14172
rect 19505 14116 19509 14172
rect 19445 14112 19509 14116
rect 19525 14172 19589 14176
rect 19525 14116 19529 14172
rect 19529 14116 19585 14172
rect 19585 14116 19589 14172
rect 19525 14112 19589 14116
rect 60 14044 124 14108
rect 60 13772 124 13836
rect 8285 13628 8349 13632
rect 8285 13572 8289 13628
rect 8289 13572 8345 13628
rect 8345 13572 8349 13628
rect 8285 13568 8349 13572
rect 8365 13628 8429 13632
rect 8365 13572 8369 13628
rect 8369 13572 8425 13628
rect 8425 13572 8429 13628
rect 8365 13568 8429 13572
rect 8445 13628 8509 13632
rect 8445 13572 8449 13628
rect 8449 13572 8505 13628
rect 8505 13572 8509 13628
rect 8445 13568 8509 13572
rect 8525 13628 8589 13632
rect 8525 13572 8529 13628
rect 8529 13572 8585 13628
rect 8585 13572 8589 13628
rect 8525 13568 8589 13572
rect 15618 13628 15682 13632
rect 15618 13572 15622 13628
rect 15622 13572 15678 13628
rect 15678 13572 15682 13628
rect 15618 13568 15682 13572
rect 15698 13628 15762 13632
rect 15698 13572 15702 13628
rect 15702 13572 15758 13628
rect 15758 13572 15762 13628
rect 15698 13568 15762 13572
rect 15778 13628 15842 13632
rect 15778 13572 15782 13628
rect 15782 13572 15838 13628
rect 15838 13572 15842 13628
rect 15778 13568 15842 13572
rect 15858 13628 15922 13632
rect 15858 13572 15862 13628
rect 15862 13572 15918 13628
rect 15918 13572 15922 13628
rect 15858 13568 15922 13572
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 4698 13084 4762 13088
rect 4698 13028 4702 13084
rect 4702 13028 4758 13084
rect 4758 13028 4762 13084
rect 4698 13024 4762 13028
rect 4778 13084 4842 13088
rect 4778 13028 4782 13084
rect 4782 13028 4838 13084
rect 4838 13028 4842 13084
rect 4778 13024 4842 13028
rect 4858 13084 4922 13088
rect 4858 13028 4862 13084
rect 4862 13028 4918 13084
rect 4918 13028 4922 13084
rect 4858 13024 4922 13028
rect 11952 13084 12016 13088
rect 11952 13028 11956 13084
rect 11956 13028 12012 13084
rect 12012 13028 12016 13084
rect 11952 13024 12016 13028
rect 12032 13084 12096 13088
rect 12032 13028 12036 13084
rect 12036 13028 12092 13084
rect 12092 13028 12096 13084
rect 12032 13024 12096 13028
rect 12112 13084 12176 13088
rect 12112 13028 12116 13084
rect 12116 13028 12172 13084
rect 12172 13028 12176 13084
rect 12112 13024 12176 13028
rect 12192 13084 12256 13088
rect 12192 13028 12196 13084
rect 12196 13028 12252 13084
rect 12252 13028 12256 13084
rect 12192 13024 12256 13028
rect 19285 13084 19349 13088
rect 19285 13028 19289 13084
rect 19289 13028 19345 13084
rect 19345 13028 19349 13084
rect 19285 13024 19349 13028
rect 19365 13084 19429 13088
rect 19365 13028 19369 13084
rect 19369 13028 19425 13084
rect 19425 13028 19429 13084
rect 19365 13024 19429 13028
rect 19445 13084 19509 13088
rect 19445 13028 19449 13084
rect 19449 13028 19505 13084
rect 19505 13028 19509 13084
rect 19445 13024 19509 13028
rect 19525 13084 19589 13088
rect 19525 13028 19529 13084
rect 19529 13028 19585 13084
rect 19585 13028 19589 13084
rect 19525 13024 19589 13028
rect 8285 12540 8349 12544
rect 8285 12484 8289 12540
rect 8289 12484 8345 12540
rect 8345 12484 8349 12540
rect 8285 12480 8349 12484
rect 8365 12540 8429 12544
rect 8365 12484 8369 12540
rect 8369 12484 8425 12540
rect 8425 12484 8429 12540
rect 8365 12480 8429 12484
rect 8445 12540 8509 12544
rect 8445 12484 8449 12540
rect 8449 12484 8505 12540
rect 8505 12484 8509 12540
rect 8445 12480 8509 12484
rect 8525 12540 8589 12544
rect 8525 12484 8529 12540
rect 8529 12484 8585 12540
rect 8585 12484 8589 12540
rect 8525 12480 8589 12484
rect 15618 12540 15682 12544
rect 15618 12484 15622 12540
rect 15622 12484 15678 12540
rect 15678 12484 15682 12540
rect 15618 12480 15682 12484
rect 15698 12540 15762 12544
rect 15698 12484 15702 12540
rect 15702 12484 15758 12540
rect 15758 12484 15762 12540
rect 15698 12480 15762 12484
rect 15778 12540 15842 12544
rect 15778 12484 15782 12540
rect 15782 12484 15838 12540
rect 15838 12484 15842 12540
rect 15778 12480 15842 12484
rect 15858 12540 15922 12544
rect 15858 12484 15862 12540
rect 15862 12484 15918 12540
rect 15918 12484 15922 12540
rect 15858 12480 15922 12484
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 4698 11996 4762 12000
rect 4698 11940 4702 11996
rect 4702 11940 4758 11996
rect 4758 11940 4762 11996
rect 4698 11936 4762 11940
rect 4778 11996 4842 12000
rect 4778 11940 4782 11996
rect 4782 11940 4838 11996
rect 4838 11940 4842 11996
rect 4778 11936 4842 11940
rect 4858 11996 4922 12000
rect 4858 11940 4862 11996
rect 4862 11940 4918 11996
rect 4918 11940 4922 11996
rect 4858 11936 4922 11940
rect 11952 11996 12016 12000
rect 11952 11940 11956 11996
rect 11956 11940 12012 11996
rect 12012 11940 12016 11996
rect 11952 11936 12016 11940
rect 12032 11996 12096 12000
rect 12032 11940 12036 11996
rect 12036 11940 12092 11996
rect 12092 11940 12096 11996
rect 12032 11936 12096 11940
rect 12112 11996 12176 12000
rect 12112 11940 12116 11996
rect 12116 11940 12172 11996
rect 12172 11940 12176 11996
rect 12112 11936 12176 11940
rect 12192 11996 12256 12000
rect 12192 11940 12196 11996
rect 12196 11940 12252 11996
rect 12252 11940 12256 11996
rect 12192 11936 12256 11940
rect 19285 11996 19349 12000
rect 19285 11940 19289 11996
rect 19289 11940 19345 11996
rect 19345 11940 19349 11996
rect 19285 11936 19349 11940
rect 19365 11996 19429 12000
rect 19365 11940 19369 11996
rect 19369 11940 19425 11996
rect 19425 11940 19429 11996
rect 19365 11936 19429 11940
rect 19445 11996 19509 12000
rect 19445 11940 19449 11996
rect 19449 11940 19505 11996
rect 19505 11940 19509 11996
rect 19445 11936 19509 11940
rect 19525 11996 19589 12000
rect 19525 11940 19529 11996
rect 19529 11940 19585 11996
rect 19585 11940 19589 11996
rect 19525 11936 19589 11940
rect 8285 11452 8349 11456
rect 8285 11396 8289 11452
rect 8289 11396 8345 11452
rect 8345 11396 8349 11452
rect 8285 11392 8349 11396
rect 8365 11452 8429 11456
rect 8365 11396 8369 11452
rect 8369 11396 8425 11452
rect 8425 11396 8429 11452
rect 8365 11392 8429 11396
rect 8445 11452 8509 11456
rect 8445 11396 8449 11452
rect 8449 11396 8505 11452
rect 8505 11396 8509 11452
rect 8445 11392 8509 11396
rect 8525 11452 8589 11456
rect 8525 11396 8529 11452
rect 8529 11396 8585 11452
rect 8585 11396 8589 11452
rect 8525 11392 8589 11396
rect 15618 11452 15682 11456
rect 15618 11396 15622 11452
rect 15622 11396 15678 11452
rect 15678 11396 15682 11452
rect 15618 11392 15682 11396
rect 15698 11452 15762 11456
rect 15698 11396 15702 11452
rect 15702 11396 15758 11452
rect 15758 11396 15762 11452
rect 15698 11392 15762 11396
rect 15778 11452 15842 11456
rect 15778 11396 15782 11452
rect 15782 11396 15838 11452
rect 15838 11396 15842 11452
rect 15778 11392 15842 11396
rect 15858 11452 15922 11456
rect 15858 11396 15862 11452
rect 15862 11396 15918 11452
rect 15918 11396 15922 11452
rect 15858 11392 15922 11396
rect 2636 11188 2700 11252
rect 4108 11188 4172 11252
rect 21588 11188 21652 11252
rect 21588 10916 21652 10980
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 4698 10908 4762 10912
rect 4698 10852 4702 10908
rect 4702 10852 4758 10908
rect 4758 10852 4762 10908
rect 4698 10848 4762 10852
rect 4778 10908 4842 10912
rect 4778 10852 4782 10908
rect 4782 10852 4838 10908
rect 4838 10852 4842 10908
rect 4778 10848 4842 10852
rect 4858 10908 4922 10912
rect 4858 10852 4862 10908
rect 4862 10852 4918 10908
rect 4918 10852 4922 10908
rect 4858 10848 4922 10852
rect 11952 10908 12016 10912
rect 11952 10852 11956 10908
rect 11956 10852 12012 10908
rect 12012 10852 12016 10908
rect 11952 10848 12016 10852
rect 12032 10908 12096 10912
rect 12032 10852 12036 10908
rect 12036 10852 12092 10908
rect 12092 10852 12096 10908
rect 12032 10848 12096 10852
rect 12112 10908 12176 10912
rect 12112 10852 12116 10908
rect 12116 10852 12172 10908
rect 12172 10852 12176 10908
rect 12112 10848 12176 10852
rect 12192 10908 12256 10912
rect 12192 10852 12196 10908
rect 12196 10852 12252 10908
rect 12252 10852 12256 10908
rect 12192 10848 12256 10852
rect 19285 10908 19349 10912
rect 19285 10852 19289 10908
rect 19289 10852 19345 10908
rect 19345 10852 19349 10908
rect 19285 10848 19349 10852
rect 19365 10908 19429 10912
rect 19365 10852 19369 10908
rect 19369 10852 19425 10908
rect 19425 10852 19429 10908
rect 19365 10848 19429 10852
rect 19445 10908 19509 10912
rect 19445 10852 19449 10908
rect 19449 10852 19505 10908
rect 19505 10852 19509 10908
rect 19445 10848 19509 10852
rect 19525 10908 19589 10912
rect 19525 10852 19529 10908
rect 19529 10852 19585 10908
rect 19585 10852 19589 10908
rect 19525 10848 19589 10852
rect 4476 10372 4540 10436
rect 8285 10364 8349 10368
rect 8285 10308 8289 10364
rect 8289 10308 8345 10364
rect 8345 10308 8349 10364
rect 8285 10304 8349 10308
rect 8365 10364 8429 10368
rect 8365 10308 8369 10364
rect 8369 10308 8425 10364
rect 8425 10308 8429 10364
rect 8365 10304 8429 10308
rect 8445 10364 8509 10368
rect 8445 10308 8449 10364
rect 8449 10308 8505 10364
rect 8505 10308 8509 10364
rect 8445 10304 8509 10308
rect 8525 10364 8589 10368
rect 8525 10308 8529 10364
rect 8529 10308 8585 10364
rect 8585 10308 8589 10364
rect 8525 10304 8589 10308
rect 15618 10364 15682 10368
rect 15618 10308 15622 10364
rect 15622 10308 15678 10364
rect 15678 10308 15682 10364
rect 15618 10304 15682 10308
rect 15698 10364 15762 10368
rect 15698 10308 15702 10364
rect 15702 10308 15758 10364
rect 15758 10308 15762 10364
rect 15698 10304 15762 10308
rect 15778 10364 15842 10368
rect 15778 10308 15782 10364
rect 15782 10308 15838 10364
rect 15838 10308 15842 10364
rect 15778 10304 15842 10308
rect 15858 10364 15922 10368
rect 15858 10308 15862 10364
rect 15862 10308 15918 10364
rect 15918 10308 15922 10364
rect 15858 10304 15922 10308
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 4698 9820 4762 9824
rect 4698 9764 4702 9820
rect 4702 9764 4758 9820
rect 4758 9764 4762 9820
rect 4698 9760 4762 9764
rect 4778 9820 4842 9824
rect 4778 9764 4782 9820
rect 4782 9764 4838 9820
rect 4838 9764 4842 9820
rect 4778 9760 4842 9764
rect 4858 9820 4922 9824
rect 4858 9764 4862 9820
rect 4862 9764 4918 9820
rect 4918 9764 4922 9820
rect 4858 9760 4922 9764
rect 11952 9820 12016 9824
rect 11952 9764 11956 9820
rect 11956 9764 12012 9820
rect 12012 9764 12016 9820
rect 11952 9760 12016 9764
rect 12032 9820 12096 9824
rect 12032 9764 12036 9820
rect 12036 9764 12092 9820
rect 12092 9764 12096 9820
rect 12032 9760 12096 9764
rect 12112 9820 12176 9824
rect 12112 9764 12116 9820
rect 12116 9764 12172 9820
rect 12172 9764 12176 9820
rect 12112 9760 12176 9764
rect 12192 9820 12256 9824
rect 12192 9764 12196 9820
rect 12196 9764 12252 9820
rect 12252 9764 12256 9820
rect 12192 9760 12256 9764
rect 19285 9820 19349 9824
rect 19285 9764 19289 9820
rect 19289 9764 19345 9820
rect 19345 9764 19349 9820
rect 19285 9760 19349 9764
rect 19365 9820 19429 9824
rect 19365 9764 19369 9820
rect 19369 9764 19425 9820
rect 19425 9764 19429 9820
rect 19365 9760 19429 9764
rect 19445 9820 19509 9824
rect 19445 9764 19449 9820
rect 19449 9764 19505 9820
rect 19505 9764 19509 9820
rect 19445 9760 19509 9764
rect 19525 9820 19589 9824
rect 19525 9764 19529 9820
rect 19529 9764 19585 9820
rect 19585 9764 19589 9820
rect 19525 9760 19589 9764
rect 8285 9276 8349 9280
rect 8285 9220 8289 9276
rect 8289 9220 8345 9276
rect 8345 9220 8349 9276
rect 8285 9216 8349 9220
rect 8365 9276 8429 9280
rect 8365 9220 8369 9276
rect 8369 9220 8425 9276
rect 8425 9220 8429 9276
rect 8365 9216 8429 9220
rect 8445 9276 8509 9280
rect 8445 9220 8449 9276
rect 8449 9220 8505 9276
rect 8505 9220 8509 9276
rect 8445 9216 8509 9220
rect 8525 9276 8589 9280
rect 8525 9220 8529 9276
rect 8529 9220 8585 9276
rect 8585 9220 8589 9276
rect 8525 9216 8589 9220
rect 15618 9276 15682 9280
rect 15618 9220 15622 9276
rect 15622 9220 15678 9276
rect 15678 9220 15682 9276
rect 15618 9216 15682 9220
rect 15698 9276 15762 9280
rect 15698 9220 15702 9276
rect 15702 9220 15758 9276
rect 15758 9220 15762 9276
rect 15698 9216 15762 9220
rect 15778 9276 15842 9280
rect 15778 9220 15782 9276
rect 15782 9220 15838 9276
rect 15838 9220 15842 9276
rect 15778 9216 15842 9220
rect 15858 9276 15922 9280
rect 15858 9220 15862 9276
rect 15862 9220 15918 9276
rect 15918 9220 15922 9276
rect 15858 9216 15922 9220
rect 5580 9148 5644 9212
rect 16252 9148 16316 9212
rect 4108 8876 4172 8940
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 4698 8732 4762 8736
rect 4698 8676 4702 8732
rect 4702 8676 4758 8732
rect 4758 8676 4762 8732
rect 4698 8672 4762 8676
rect 4778 8732 4842 8736
rect 4778 8676 4782 8732
rect 4782 8676 4838 8732
rect 4838 8676 4842 8732
rect 4778 8672 4842 8676
rect 4858 8732 4922 8736
rect 4858 8676 4862 8732
rect 4862 8676 4918 8732
rect 4918 8676 4922 8732
rect 4858 8672 4922 8676
rect 11952 8732 12016 8736
rect 11952 8676 11956 8732
rect 11956 8676 12012 8732
rect 12012 8676 12016 8732
rect 11952 8672 12016 8676
rect 12032 8732 12096 8736
rect 12032 8676 12036 8732
rect 12036 8676 12092 8732
rect 12092 8676 12096 8732
rect 12032 8672 12096 8676
rect 12112 8732 12176 8736
rect 12112 8676 12116 8732
rect 12116 8676 12172 8732
rect 12172 8676 12176 8732
rect 12112 8672 12176 8676
rect 12192 8732 12256 8736
rect 12192 8676 12196 8732
rect 12196 8676 12252 8732
rect 12252 8676 12256 8732
rect 12192 8672 12256 8676
rect 19285 8732 19349 8736
rect 19285 8676 19289 8732
rect 19289 8676 19345 8732
rect 19345 8676 19349 8732
rect 19285 8672 19349 8676
rect 19365 8732 19429 8736
rect 19365 8676 19369 8732
rect 19369 8676 19425 8732
rect 19425 8676 19429 8732
rect 19365 8672 19429 8676
rect 19445 8732 19509 8736
rect 19445 8676 19449 8732
rect 19449 8676 19505 8732
rect 19505 8676 19509 8732
rect 19445 8672 19509 8676
rect 19525 8732 19589 8736
rect 19525 8676 19529 8732
rect 19529 8676 19585 8732
rect 19585 8676 19589 8732
rect 19525 8672 19589 8676
rect 18644 8468 18708 8532
rect 8285 8188 8349 8192
rect 8285 8132 8289 8188
rect 8289 8132 8345 8188
rect 8345 8132 8349 8188
rect 8285 8128 8349 8132
rect 8365 8188 8429 8192
rect 8365 8132 8369 8188
rect 8369 8132 8425 8188
rect 8425 8132 8429 8188
rect 8365 8128 8429 8132
rect 8445 8188 8509 8192
rect 8445 8132 8449 8188
rect 8449 8132 8505 8188
rect 8505 8132 8509 8188
rect 8445 8128 8509 8132
rect 8525 8188 8589 8192
rect 8525 8132 8529 8188
rect 8529 8132 8585 8188
rect 8585 8132 8589 8188
rect 8525 8128 8589 8132
rect 15618 8188 15682 8192
rect 15618 8132 15622 8188
rect 15622 8132 15678 8188
rect 15678 8132 15682 8188
rect 15618 8128 15682 8132
rect 15698 8188 15762 8192
rect 15698 8132 15702 8188
rect 15702 8132 15758 8188
rect 15758 8132 15762 8188
rect 15698 8128 15762 8132
rect 15778 8188 15842 8192
rect 15778 8132 15782 8188
rect 15782 8132 15838 8188
rect 15838 8132 15842 8188
rect 15778 8128 15842 8132
rect 15858 8188 15922 8192
rect 15858 8132 15862 8188
rect 15862 8132 15918 8188
rect 15918 8132 15922 8188
rect 15858 8128 15922 8132
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 4698 7644 4762 7648
rect 4698 7588 4702 7644
rect 4702 7588 4758 7644
rect 4758 7588 4762 7644
rect 4698 7584 4762 7588
rect 4778 7644 4842 7648
rect 4778 7588 4782 7644
rect 4782 7588 4838 7644
rect 4838 7588 4842 7644
rect 4778 7584 4842 7588
rect 4858 7644 4922 7648
rect 4858 7588 4862 7644
rect 4862 7588 4918 7644
rect 4918 7588 4922 7644
rect 4858 7584 4922 7588
rect 11952 7644 12016 7648
rect 11952 7588 11956 7644
rect 11956 7588 12012 7644
rect 12012 7588 12016 7644
rect 11952 7584 12016 7588
rect 12032 7644 12096 7648
rect 12032 7588 12036 7644
rect 12036 7588 12092 7644
rect 12092 7588 12096 7644
rect 12032 7584 12096 7588
rect 12112 7644 12176 7648
rect 12112 7588 12116 7644
rect 12116 7588 12172 7644
rect 12172 7588 12176 7644
rect 12112 7584 12176 7588
rect 12192 7644 12256 7648
rect 12192 7588 12196 7644
rect 12196 7588 12252 7644
rect 12252 7588 12256 7644
rect 12192 7584 12256 7588
rect 19285 7644 19349 7648
rect 19285 7588 19289 7644
rect 19289 7588 19345 7644
rect 19345 7588 19349 7644
rect 19285 7584 19349 7588
rect 19365 7644 19429 7648
rect 19365 7588 19369 7644
rect 19369 7588 19425 7644
rect 19425 7588 19429 7644
rect 19365 7584 19429 7588
rect 19445 7644 19509 7648
rect 19445 7588 19449 7644
rect 19449 7588 19505 7644
rect 19505 7588 19509 7644
rect 19445 7584 19509 7588
rect 19525 7644 19589 7648
rect 19525 7588 19529 7644
rect 19529 7588 19585 7644
rect 19585 7588 19589 7644
rect 19525 7584 19589 7588
rect 21588 7516 21652 7580
rect 21588 7244 21652 7308
rect 7972 7108 8036 7172
rect 16620 7108 16684 7172
rect 8285 7100 8349 7104
rect 8285 7044 8289 7100
rect 8289 7044 8345 7100
rect 8345 7044 8349 7100
rect 8285 7040 8349 7044
rect 8365 7100 8429 7104
rect 8365 7044 8369 7100
rect 8369 7044 8425 7100
rect 8425 7044 8429 7100
rect 8365 7040 8429 7044
rect 8445 7100 8509 7104
rect 8445 7044 8449 7100
rect 8449 7044 8505 7100
rect 8505 7044 8509 7100
rect 8445 7040 8509 7044
rect 8525 7100 8589 7104
rect 8525 7044 8529 7100
rect 8529 7044 8585 7100
rect 8585 7044 8589 7100
rect 8525 7040 8589 7044
rect 15618 7100 15682 7104
rect 15618 7044 15622 7100
rect 15622 7044 15678 7100
rect 15678 7044 15682 7100
rect 15618 7040 15682 7044
rect 15698 7100 15762 7104
rect 15698 7044 15702 7100
rect 15702 7044 15758 7100
rect 15758 7044 15762 7100
rect 15698 7040 15762 7044
rect 15778 7100 15842 7104
rect 15778 7044 15782 7100
rect 15782 7044 15838 7100
rect 15838 7044 15842 7100
rect 15778 7040 15842 7044
rect 15858 7100 15922 7104
rect 15858 7044 15862 7100
rect 15862 7044 15918 7100
rect 15918 7044 15922 7100
rect 15858 7040 15922 7044
rect 60 6972 124 7036
rect 60 6700 124 6764
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 4698 6556 4762 6560
rect 4698 6500 4702 6556
rect 4702 6500 4758 6556
rect 4758 6500 4762 6556
rect 4698 6496 4762 6500
rect 4778 6556 4842 6560
rect 4778 6500 4782 6556
rect 4782 6500 4838 6556
rect 4838 6500 4842 6556
rect 4778 6496 4842 6500
rect 4858 6556 4922 6560
rect 4858 6500 4862 6556
rect 4862 6500 4918 6556
rect 4918 6500 4922 6556
rect 4858 6496 4922 6500
rect 11952 6556 12016 6560
rect 11952 6500 11956 6556
rect 11956 6500 12012 6556
rect 12012 6500 12016 6556
rect 11952 6496 12016 6500
rect 12032 6556 12096 6560
rect 12032 6500 12036 6556
rect 12036 6500 12092 6556
rect 12092 6500 12096 6556
rect 12032 6496 12096 6500
rect 12112 6556 12176 6560
rect 12112 6500 12116 6556
rect 12116 6500 12172 6556
rect 12172 6500 12176 6556
rect 12112 6496 12176 6500
rect 12192 6556 12256 6560
rect 12192 6500 12196 6556
rect 12196 6500 12252 6556
rect 12252 6500 12256 6556
rect 12192 6496 12256 6500
rect 19285 6556 19349 6560
rect 19285 6500 19289 6556
rect 19289 6500 19345 6556
rect 19345 6500 19349 6556
rect 19285 6496 19349 6500
rect 19365 6556 19429 6560
rect 19365 6500 19369 6556
rect 19369 6500 19425 6556
rect 19425 6500 19429 6556
rect 19365 6496 19429 6500
rect 19445 6556 19509 6560
rect 19445 6500 19449 6556
rect 19449 6500 19505 6556
rect 19505 6500 19509 6556
rect 19445 6496 19509 6500
rect 19525 6556 19589 6560
rect 19525 6500 19529 6556
rect 19529 6500 19585 6556
rect 19585 6500 19589 6556
rect 19525 6496 19589 6500
rect 3556 6428 3620 6492
rect 8285 6012 8349 6016
rect 8285 5956 8289 6012
rect 8289 5956 8345 6012
rect 8345 5956 8349 6012
rect 8285 5952 8349 5956
rect 8365 6012 8429 6016
rect 8365 5956 8369 6012
rect 8369 5956 8425 6012
rect 8425 5956 8429 6012
rect 8365 5952 8429 5956
rect 8445 6012 8509 6016
rect 8445 5956 8449 6012
rect 8449 5956 8505 6012
rect 8505 5956 8509 6012
rect 8445 5952 8509 5956
rect 8525 6012 8589 6016
rect 8525 5956 8529 6012
rect 8529 5956 8585 6012
rect 8585 5956 8589 6012
rect 8525 5952 8589 5956
rect 15618 6012 15682 6016
rect 15618 5956 15622 6012
rect 15622 5956 15678 6012
rect 15678 5956 15682 6012
rect 15618 5952 15682 5956
rect 15698 6012 15762 6016
rect 15698 5956 15702 6012
rect 15702 5956 15758 6012
rect 15758 5956 15762 6012
rect 15698 5952 15762 5956
rect 15778 6012 15842 6016
rect 15778 5956 15782 6012
rect 15782 5956 15838 6012
rect 15838 5956 15842 6012
rect 15778 5952 15842 5956
rect 15858 6012 15922 6016
rect 15858 5956 15862 6012
rect 15862 5956 15918 6012
rect 15918 5956 15922 6012
rect 15858 5952 15922 5956
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 4698 5468 4762 5472
rect 4698 5412 4702 5468
rect 4702 5412 4758 5468
rect 4758 5412 4762 5468
rect 4698 5408 4762 5412
rect 4778 5468 4842 5472
rect 4778 5412 4782 5468
rect 4782 5412 4838 5468
rect 4838 5412 4842 5468
rect 4778 5408 4842 5412
rect 4858 5468 4922 5472
rect 4858 5412 4862 5468
rect 4862 5412 4918 5468
rect 4918 5412 4922 5468
rect 4858 5408 4922 5412
rect 11952 5468 12016 5472
rect 11952 5412 11956 5468
rect 11956 5412 12012 5468
rect 12012 5412 12016 5468
rect 11952 5408 12016 5412
rect 12032 5468 12096 5472
rect 12032 5412 12036 5468
rect 12036 5412 12092 5468
rect 12092 5412 12096 5468
rect 12032 5408 12096 5412
rect 12112 5468 12176 5472
rect 12112 5412 12116 5468
rect 12116 5412 12172 5468
rect 12172 5412 12176 5468
rect 12112 5408 12176 5412
rect 12192 5468 12256 5472
rect 12192 5412 12196 5468
rect 12196 5412 12252 5468
rect 12252 5412 12256 5468
rect 12192 5408 12256 5412
rect 19285 5468 19349 5472
rect 19285 5412 19289 5468
rect 19289 5412 19345 5468
rect 19345 5412 19349 5468
rect 19285 5408 19349 5412
rect 19365 5468 19429 5472
rect 19365 5412 19369 5468
rect 19369 5412 19425 5468
rect 19425 5412 19429 5468
rect 19365 5408 19429 5412
rect 19445 5468 19509 5472
rect 19445 5412 19449 5468
rect 19449 5412 19505 5468
rect 19505 5412 19509 5468
rect 19445 5408 19509 5412
rect 19525 5468 19589 5472
rect 19525 5412 19529 5468
rect 19529 5412 19585 5468
rect 19585 5412 19589 5468
rect 19525 5408 19589 5412
rect 7420 5340 7484 5404
rect 4108 5068 4172 5132
rect 1900 4932 1964 4996
rect 8285 4924 8349 4928
rect 8285 4868 8289 4924
rect 8289 4868 8345 4924
rect 8345 4868 8349 4924
rect 8285 4864 8349 4868
rect 8365 4924 8429 4928
rect 8365 4868 8369 4924
rect 8369 4868 8425 4924
rect 8425 4868 8429 4924
rect 8365 4864 8429 4868
rect 8445 4924 8509 4928
rect 8445 4868 8449 4924
rect 8449 4868 8505 4924
rect 8505 4868 8509 4924
rect 8445 4864 8509 4868
rect 8525 4924 8589 4928
rect 8525 4868 8529 4924
rect 8529 4868 8585 4924
rect 8585 4868 8589 4924
rect 8525 4864 8589 4868
rect 15618 4924 15682 4928
rect 15618 4868 15622 4924
rect 15622 4868 15678 4924
rect 15678 4868 15682 4924
rect 15618 4864 15682 4868
rect 15698 4924 15762 4928
rect 15698 4868 15702 4924
rect 15702 4868 15758 4924
rect 15758 4868 15762 4924
rect 15698 4864 15762 4868
rect 15778 4924 15842 4928
rect 15778 4868 15782 4924
rect 15782 4868 15838 4924
rect 15838 4868 15842 4924
rect 15778 4864 15842 4868
rect 15858 4924 15922 4928
rect 15858 4868 15862 4924
rect 15862 4868 15918 4924
rect 15918 4868 15922 4924
rect 15858 4864 15922 4868
rect 9628 4524 9692 4588
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 4698 4380 4762 4384
rect 4698 4324 4702 4380
rect 4702 4324 4758 4380
rect 4758 4324 4762 4380
rect 4698 4320 4762 4324
rect 4778 4380 4842 4384
rect 4778 4324 4782 4380
rect 4782 4324 4838 4380
rect 4838 4324 4842 4380
rect 4778 4320 4842 4324
rect 4858 4380 4922 4384
rect 4858 4324 4862 4380
rect 4862 4324 4918 4380
rect 4918 4324 4922 4380
rect 4858 4320 4922 4324
rect 11952 4380 12016 4384
rect 11952 4324 11956 4380
rect 11956 4324 12012 4380
rect 12012 4324 12016 4380
rect 11952 4320 12016 4324
rect 12032 4380 12096 4384
rect 12032 4324 12036 4380
rect 12036 4324 12092 4380
rect 12092 4324 12096 4380
rect 12032 4320 12096 4324
rect 12112 4380 12176 4384
rect 12112 4324 12116 4380
rect 12116 4324 12172 4380
rect 12172 4324 12176 4380
rect 12112 4320 12176 4324
rect 12192 4380 12256 4384
rect 12192 4324 12196 4380
rect 12196 4324 12252 4380
rect 12252 4324 12256 4380
rect 12192 4320 12256 4324
rect 19285 4380 19349 4384
rect 19285 4324 19289 4380
rect 19289 4324 19345 4380
rect 19345 4324 19349 4380
rect 19285 4320 19349 4324
rect 19365 4380 19429 4384
rect 19365 4324 19369 4380
rect 19369 4324 19425 4380
rect 19425 4324 19429 4380
rect 19365 4320 19429 4324
rect 19445 4380 19509 4384
rect 19445 4324 19449 4380
rect 19449 4324 19505 4380
rect 19505 4324 19509 4380
rect 19445 4320 19509 4324
rect 19525 4380 19589 4384
rect 19525 4324 19529 4380
rect 19529 4324 19585 4380
rect 19585 4324 19589 4380
rect 19525 4320 19589 4324
rect 8285 3836 8349 3840
rect 8285 3780 8289 3836
rect 8289 3780 8345 3836
rect 8345 3780 8349 3836
rect 8285 3776 8349 3780
rect 8365 3836 8429 3840
rect 8365 3780 8369 3836
rect 8369 3780 8425 3836
rect 8425 3780 8429 3836
rect 8365 3776 8429 3780
rect 8445 3836 8509 3840
rect 8445 3780 8449 3836
rect 8449 3780 8505 3836
rect 8505 3780 8509 3836
rect 8445 3776 8509 3780
rect 8525 3836 8589 3840
rect 8525 3780 8529 3836
rect 8529 3780 8585 3836
rect 8585 3780 8589 3836
rect 8525 3776 8589 3780
rect 15618 3836 15682 3840
rect 15618 3780 15622 3836
rect 15622 3780 15678 3836
rect 15678 3780 15682 3836
rect 15618 3776 15682 3780
rect 15698 3836 15762 3840
rect 15698 3780 15702 3836
rect 15702 3780 15758 3836
rect 15758 3780 15762 3836
rect 15698 3776 15762 3780
rect 15778 3836 15842 3840
rect 15778 3780 15782 3836
rect 15782 3780 15838 3836
rect 15838 3780 15842 3836
rect 15778 3776 15842 3780
rect 15858 3836 15922 3840
rect 15858 3780 15862 3836
rect 15862 3780 15918 3836
rect 15918 3780 15922 3836
rect 15858 3776 15922 3780
rect 4292 3708 4356 3772
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 4698 3292 4762 3296
rect 4698 3236 4702 3292
rect 4702 3236 4758 3292
rect 4758 3236 4762 3292
rect 4698 3232 4762 3236
rect 4778 3292 4842 3296
rect 4778 3236 4782 3292
rect 4782 3236 4838 3292
rect 4838 3236 4842 3292
rect 4778 3232 4842 3236
rect 4858 3292 4922 3296
rect 4858 3236 4862 3292
rect 4862 3236 4918 3292
rect 4918 3236 4922 3292
rect 4858 3232 4922 3236
rect 11952 3292 12016 3296
rect 11952 3236 11956 3292
rect 11956 3236 12012 3292
rect 12012 3236 12016 3292
rect 11952 3232 12016 3236
rect 12032 3292 12096 3296
rect 12032 3236 12036 3292
rect 12036 3236 12092 3292
rect 12092 3236 12096 3292
rect 12032 3232 12096 3236
rect 12112 3292 12176 3296
rect 12112 3236 12116 3292
rect 12116 3236 12172 3292
rect 12172 3236 12176 3292
rect 12112 3232 12176 3236
rect 12192 3292 12256 3296
rect 12192 3236 12196 3292
rect 12196 3236 12252 3292
rect 12252 3236 12256 3292
rect 12192 3232 12256 3236
rect 19285 3292 19349 3296
rect 19285 3236 19289 3292
rect 19289 3236 19345 3292
rect 19345 3236 19349 3292
rect 19285 3232 19349 3236
rect 19365 3292 19429 3296
rect 19365 3236 19369 3292
rect 19369 3236 19425 3292
rect 19425 3236 19429 3292
rect 19365 3232 19429 3236
rect 19445 3292 19509 3296
rect 19445 3236 19449 3292
rect 19449 3236 19505 3292
rect 19505 3236 19509 3292
rect 19445 3232 19509 3236
rect 19525 3292 19589 3296
rect 19525 3236 19529 3292
rect 19529 3236 19585 3292
rect 19585 3236 19589 3292
rect 19525 3232 19589 3236
rect 8285 2748 8349 2752
rect 8285 2692 8289 2748
rect 8289 2692 8345 2748
rect 8345 2692 8349 2748
rect 8285 2688 8349 2692
rect 8365 2748 8429 2752
rect 8365 2692 8369 2748
rect 8369 2692 8425 2748
rect 8425 2692 8429 2748
rect 8365 2688 8429 2692
rect 8445 2748 8509 2752
rect 8445 2692 8449 2748
rect 8449 2692 8505 2748
rect 8505 2692 8509 2748
rect 8445 2688 8509 2692
rect 8525 2748 8589 2752
rect 8525 2692 8529 2748
rect 8529 2692 8585 2748
rect 8585 2692 8589 2748
rect 8525 2688 8589 2692
rect 15618 2748 15682 2752
rect 15618 2692 15622 2748
rect 15622 2692 15678 2748
rect 15678 2692 15682 2748
rect 15618 2688 15682 2692
rect 15698 2748 15762 2752
rect 15698 2692 15702 2748
rect 15702 2692 15758 2748
rect 15758 2692 15762 2748
rect 15698 2688 15762 2692
rect 15778 2748 15842 2752
rect 15778 2692 15782 2748
rect 15782 2692 15838 2748
rect 15838 2692 15842 2748
rect 15778 2688 15842 2692
rect 15858 2748 15922 2752
rect 15858 2692 15862 2748
rect 15862 2692 15918 2748
rect 15918 2692 15922 2748
rect 15858 2688 15922 2692
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 4698 2204 4762 2208
rect 4698 2148 4702 2204
rect 4702 2148 4758 2204
rect 4758 2148 4762 2204
rect 4698 2144 4762 2148
rect 4778 2204 4842 2208
rect 4778 2148 4782 2204
rect 4782 2148 4838 2204
rect 4838 2148 4842 2204
rect 4778 2144 4842 2148
rect 4858 2204 4922 2208
rect 4858 2148 4862 2204
rect 4862 2148 4918 2204
rect 4918 2148 4922 2204
rect 4858 2144 4922 2148
rect 11952 2204 12016 2208
rect 11952 2148 11956 2204
rect 11956 2148 12012 2204
rect 12012 2148 12016 2204
rect 11952 2144 12016 2148
rect 12032 2204 12096 2208
rect 12032 2148 12036 2204
rect 12036 2148 12092 2204
rect 12092 2148 12096 2204
rect 12032 2144 12096 2148
rect 12112 2204 12176 2208
rect 12112 2148 12116 2204
rect 12116 2148 12172 2204
rect 12172 2148 12176 2204
rect 12112 2144 12176 2148
rect 12192 2204 12256 2208
rect 12192 2148 12196 2204
rect 12196 2148 12252 2204
rect 12252 2148 12256 2204
rect 12192 2144 12256 2148
rect 19285 2204 19349 2208
rect 19285 2148 19289 2204
rect 19289 2148 19345 2204
rect 19345 2148 19349 2204
rect 19285 2144 19349 2148
rect 19365 2204 19429 2208
rect 19365 2148 19369 2204
rect 19369 2148 19425 2204
rect 19425 2148 19429 2204
rect 19365 2144 19429 2148
rect 19445 2204 19509 2208
rect 19445 2148 19449 2204
rect 19449 2148 19505 2204
rect 19505 2148 19509 2204
rect 19445 2144 19509 2148
rect 19525 2204 19589 2208
rect 19525 2148 19529 2204
rect 19529 2148 19585 2204
rect 19585 2148 19589 2204
rect 19525 2144 19589 2148
rect 17908 1668 17972 1732
rect 4108 36 4172 100
<< metal4 >>
rect 2635 21588 2701 21589
rect 2635 21524 2636 21588
rect 2700 21524 2701 21588
rect 2635 21523 2701 21524
rect 59 16420 125 16421
rect 59 16356 60 16420
rect 124 16356 125 16420
rect 59 16355 125 16356
rect 62 16149 122 16355
rect 59 16148 125 16149
rect 59 16084 60 16148
rect 124 16084 125 16148
rect 59 16083 125 16084
rect 59 14108 125 14109
rect 59 14044 60 14108
rect 124 14044 125 14108
rect 59 14043 125 14044
rect 62 13837 122 14043
rect 59 13836 125 13837
rect 59 13772 60 13836
rect 124 13772 125 13836
rect 59 13771 125 13772
rect 2638 11338 2698 21523
rect 4610 19616 4931 19632
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4931 19616
rect 4610 18528 4931 19552
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4931 18528
rect 4610 17440 4931 18464
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4931 17440
rect 4610 16352 4931 17376
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4931 16352
rect 4610 15264 4931 16288
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4931 15264
rect 4610 14176 4931 15200
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4931 14176
rect 4610 13088 4931 14112
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4931 13088
rect 4610 12000 4931 13024
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4931 12000
rect 2638 11060 2698 11102
rect 4610 10912 4931 11936
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4931 10912
rect 4475 10436 4541 10437
rect 4475 10372 4476 10436
rect 4540 10372 4541 10436
rect 4475 10371 4541 10372
rect 4107 8940 4173 8941
rect 4107 8876 4108 8940
rect 4172 8876 4173 8940
rect 4107 8875 4173 8876
rect 4110 8618 4170 8875
rect 59 7036 125 7037
rect 59 6972 60 7036
rect 124 6972 125 7036
rect 59 6971 125 6972
rect 62 6765 122 6971
rect 59 6764 125 6765
rect 59 6700 60 6764
rect 124 6700 125 6764
rect 59 6699 125 6700
rect 3555 6492 3621 6493
rect 3555 6428 3556 6492
rect 3620 6428 3621 6492
rect 3555 6427 3621 6428
rect 3558 5218 3618 6427
rect 1899 4996 1965 4997
rect 1899 4932 1900 4996
rect 1964 4932 1965 4996
rect 1899 4931 1965 4932
rect 1902 3858 1962 4931
rect 4478 4170 4538 10371
rect 4294 4110 4538 4170
rect 4610 9824 4931 10848
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4931 9824
rect 4610 8736 4931 9760
rect 8277 19072 8597 19632
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 17984 8597 19008
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 8277 16896 8597 17920
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 8277 15808 8597 16832
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 8277 14720 8597 15744
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 8277 13632 8597 14656
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 8277 12544 8597 13568
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 11456 8597 12480
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 10368 8597 11392
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 9280 8597 10304
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4931 8736
rect 4610 7648 4931 8672
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4931 7648
rect 4610 6560 4931 7584
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4931 6560
rect 4610 5472 4931 6496
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4931 5472
rect 4610 4384 4931 5408
rect 7422 5405 7482 8382
rect 8277 8192 8597 9216
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 7104 8597 8128
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 8277 6016 8597 7040
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 7419 5404 7485 5405
rect 7419 5340 7420 5404
rect 7484 5340 7485 5404
rect 7419 5339 7485 5340
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4931 4384
rect 4294 3773 4354 4110
rect 4291 3772 4357 3773
rect 4291 3708 4292 3772
rect 4356 3708 4357 3772
rect 4291 3707 4357 3708
rect 4610 3296 4931 4320
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4931 3296
rect 4610 2208 4931 3232
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4931 2208
rect 4610 2128 4931 2144
rect 8277 4928 8597 5952
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 8277 3840 8597 4864
rect 11944 19616 12264 19632
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 18528 12264 19552
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 17440 12264 18464
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 11944 16352 12264 17376
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11944 15264 12264 16288
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11944 14176 12264 15200
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11944 13088 12264 14112
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 12000 12264 13024
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 10912 12264 11936
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11944 9824 12264 10848
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 11944 8736 12264 9760
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 11944 7648 12264 8672
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 6560 12264 7584
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 5472 12264 6496
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 9627 4588 9693 4589
rect 9627 4524 9628 4588
rect 9692 4524 9693 4588
rect 9627 4523 9693 4524
rect 9630 3858 9690 4523
rect 11944 4384 12264 5408
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 8277 2752 8597 3776
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2128 8597 2688
rect 11944 3296 12264 4320
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 2208 12264 3232
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2128 12264 2144
rect 15610 19072 15930 19632
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 17984 15930 19008
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 15610 16896 15930 17920
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 15610 15808 15930 16832
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 14720 15930 15744
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 15610 13632 15930 14656
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 15610 12544 15930 13568
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 11456 15930 12480
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 15610 10368 15930 11392
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 9280 15930 10304
rect 19277 19616 19597 19632
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 18528 19597 19552
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 19277 17440 19597 18464
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 16352 19597 17376
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 15264 19597 16288
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 19277 14176 19597 15200
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 13088 19597 14112
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 19277 12000 19597 13024
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 10912 19597 11936
rect 21587 11252 21653 11253
rect 21587 11188 21588 11252
rect 21652 11188 21653 11252
rect 21587 11187 21653 11188
rect 21590 10981 21650 11187
rect 21587 10980 21653 10981
rect 21587 10916 21588 10980
rect 21652 10916 21653 10980
rect 21587 10915 21653 10916
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 19277 9824 19597 10848
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 15610 8192 15930 9216
rect 19277 8736 19597 9760
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 15610 7104 15930 8128
rect 19277 7648 19597 8672
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 15610 6016 15930 7040
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 15610 4928 15930 5952
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 15610 3840 15930 4864
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 15610 2752 15930 3776
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 15610 2128 15930 2688
rect 19277 6560 19597 7584
rect 21587 7580 21653 7581
rect 21587 7516 21588 7580
rect 21652 7516 21653 7580
rect 21587 7515 21653 7516
rect 21590 7309 21650 7515
rect 21587 7308 21653 7309
rect 21587 7244 21588 7308
rect 21652 7244 21653 7308
rect 21587 7243 21653 7244
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 5472 19597 6496
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 19277 4384 19597 5408
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 19277 3296 19597 4320
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 19277 2208 19597 3232
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2128 19597 2144
rect 4110 101 4170 1582
rect 4107 100 4173 101
rect 4107 36 4108 100
rect 4172 36 4173 100
rect 4107 35 4173 36
<< via4 >>
rect 2550 11252 2786 11338
rect 2550 11188 2636 11252
rect 2636 11188 2700 11252
rect 2700 11188 2786 11252
rect 2550 11102 2786 11188
rect 4022 11252 4258 11338
rect 4022 11188 4108 11252
rect 4108 11188 4172 11252
rect 4172 11188 4258 11252
rect 4022 11102 4258 11188
rect 4022 8382 4258 8618
rect 3470 4982 3706 5218
rect 4022 5132 4258 5218
rect 4022 5068 4108 5132
rect 4108 5068 4172 5132
rect 4172 5068 4258 5132
rect 4022 4982 4258 5068
rect 5494 9212 5730 9298
rect 5494 9148 5580 9212
rect 5580 9148 5644 9212
rect 5644 9148 5730 9212
rect 5494 9062 5730 9148
rect 7334 8382 7570 8618
rect 7886 7172 8122 7258
rect 7886 7108 7972 7172
rect 7972 7108 8036 7172
rect 8036 7108 8122 7172
rect 7886 7022 8122 7108
rect 1814 3622 2050 3858
rect 9542 3622 9778 3858
rect 16166 9212 16402 9298
rect 16166 9148 16252 9212
rect 16252 9148 16316 9212
rect 16316 9148 16402 9212
rect 16166 9062 16402 9148
rect 18558 8532 18794 8618
rect 18558 8468 18644 8532
rect 18644 8468 18708 8532
rect 18708 8468 18794 8532
rect 18558 8382 18794 8468
rect 16534 7172 16770 7258
rect 16534 7108 16620 7172
rect 16620 7108 16684 7172
rect 16684 7108 16770 7172
rect 16534 7022 16770 7108
rect 4022 1582 4258 1818
rect 17822 1732 18058 1818
rect 17822 1668 17908 1732
rect 17908 1668 17972 1732
rect 17972 1668 18058 1732
rect 17822 1582 18058 1668
<< metal5 >>
rect 2508 11338 4300 11380
rect 2508 11102 2550 11338
rect 2786 11102 4022 11338
rect 4258 11102 4300 11338
rect 2508 11060 4300 11102
rect 5452 9298 16444 9340
rect 5452 9062 5494 9298
rect 5730 9062 16166 9298
rect 16402 9062 16444 9298
rect 5452 9020 16444 9062
rect 3980 8618 18836 8660
rect 3980 8382 4022 8618
rect 4258 8382 7334 8618
rect 7570 8382 18558 8618
rect 18794 8382 18836 8618
rect 3980 8340 18836 8382
rect 7844 7258 16812 7300
rect 7844 7022 7886 7258
rect 8122 7022 16534 7258
rect 16770 7022 16812 7258
rect 7844 6980 16812 7022
rect 3428 5218 4300 5260
rect 3428 4982 3470 5218
rect 3706 4982 4022 5218
rect 4258 4982 4300 5218
rect 3428 4940 4300 4982
rect 1772 3858 9820 3900
rect 1772 3622 1814 3858
rect 2050 3622 9542 3858
rect 9778 3622 9820 3858
rect 1772 3580 9820 3622
rect 3980 1818 18100 1860
rect 3980 1582 4022 1818
rect 4258 1582 17822 1818
rect 18058 1582 18100 1818
rect 3980 1540 18100 1582
use scs8hd_decap_4  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__B tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_8 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_or4_4  _110_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 866 592
use scs8hd_or3_4  _075_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _061_
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__061__C
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__B
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_21
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_25
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_19
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_29
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_64 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _145_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_or3_4  _065_
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _104_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__065__C
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__C
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__B
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 1050 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_79
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_80
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _142_
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 1050 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_94
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _045_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_115
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_111
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_111
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _159_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_nor2_4  _077_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__053__C
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_144
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_148
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_140
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_or3_4  _053_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__053__B
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _158_
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_177
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _049_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _050_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_181
timestamp 1586364061
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _139_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_196 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_204 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 20884 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 20884 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 406 592
use scs8hd_nand2_4  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_12
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_22
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_26
timestamp 1586364061
transform 1 0 3496 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 4508 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_29
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_35
timestamp 1586364061
transform 1 0 4324 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_39
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 222 592
use scs8hd_or3_4  _057_
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__059__C
timestamp 1586364061
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_52
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 222 592
use scs8hd_or2_4  _054_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_110
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_114
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _042_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_4  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_8  _048_
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_180
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_197
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_14
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_18
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__C
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _063_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_or2_4  _076_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_69
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8280 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_89
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_93
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_106
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_126
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_130
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_146
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_150
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_163
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _136_
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_167
timestamp 1586364061
transform 1 0 16468 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_174
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 314 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 20884 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_16
timestamp 1586364061
transform 1 0 2576 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_20
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_4_26
timestamp 1586364061
transform 1 0 3496 0 -1 4896
box -38 -48 314 592
use scs8hd_nor3_4  _107_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__C
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_or3_4  _059_
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__C
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_45
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_49
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_62
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_66
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_70
timestamp 1586364061
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_87
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_138
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_142
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_146
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_150
timestamp 1586364061
transform 1 0 14904 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use scs8hd_buf_2  _155_
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_8  FILLER_4_192
timestamp 1586364061
transform 1 0 18768 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_203
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_211
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_13
timestamp 1586364061
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use scs8hd_nor3_4  _106_
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_17
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_21
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_37
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_41
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_or2_4  _098_
timestamp 1586364061
transform 1 0 5244 0 1 4896
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_52
timestamp 1586364061
transform 1 0 5888 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_56
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_68
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_72
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_87
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_91
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_104
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_108
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_140
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _044_
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_157
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_182
timestamp 1586364061
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_187
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_198
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_202
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_206 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20056 0 1 4896
box -38 -48 590 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 20884 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 1050 592
use scs8hd_buf_2  _147_
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_20
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_26
timestamp 1586364061
transform 1 0 3496 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_18
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_22
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_30
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__D
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_36
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__C
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_nor3_4  _109_
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 1234 592
use scs8hd_nor3_4  _108_
timestamp 1586364061
transform 1 0 4508 0 -1 5984
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_50
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_54
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_61
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_69
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_or2_4  _117_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 682 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_73
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_109
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_113
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_135
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_139
timestamp 1586364061
transform 1 0 13892 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_150
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_155
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_168
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_173
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _140_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_180
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_181
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_187
timestamp 1586364061
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_191
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_198
timestamp 1586364061
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_202
timestamp 1586364061
transform 1 0 19688 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_206
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 590 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 20884 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 20884 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_14
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_18
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_22
timestamp 1586364061
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_26
timestamp 1586364061
transform 1 0 3496 0 -1 7072
box -38 -48 314 592
use scs8hd_or4_4  _099_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__D
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_60
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_128
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_134
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_148
timestamp 1586364061
transform 1 0 14720 0 -1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__055__B
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_180
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_191
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__055__D
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_195
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _043_
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 406 592
use scs8hd_or4_4  _068_
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_28
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_41
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_45
timestamp 1586364061
transform 1 0 5244 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_or2_4  _124_
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_104
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_108
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_126
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_146
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_150
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_163
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_167
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use scs8hd_inv_8  _051_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _141_
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__C
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_204
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 20884 0 1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_12
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_or2_4  _084_
timestamp 1586364061
transform 1 0 4140 0 -1 8160
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_40
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_59
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9752 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_109
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_112
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_116
timestamp 1586364061
transform 1 0 11776 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_148
timestamp 1586364061
transform 1 0 14720 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _046_
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_or4_4  _055_
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_180
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_197
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_209
timestamp 1586364061
transform 1 0 20332 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_46
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_50
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_54
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_117
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _073_
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_172
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_176
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 406 592
use scs8hd_inv_8  _052_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_204
timestamp 1586364061
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 20884 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_12
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_16
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_38
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_42
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_76
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_130
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_167
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_180
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_191
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_195
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_2  _151_
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_17
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_21
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_33
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_58
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_107
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_115
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_111
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_119
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_139
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_160
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_177
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _069_
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_180
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_197
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 20884 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_2  _143_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_25
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_29
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_79
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_102
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13340 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_129
timestamp 1586364061
transform 1 0 12972 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_148
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_161
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_165
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_172
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_176
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _071_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_180
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _135_
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 406 592
use scs8hd_decap_8  FILLER_15_204
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 20884 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_21
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_25
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4692 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_29
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_50
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_54
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_67
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_4  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_97
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_109
timestamp 1586364061
transform 1 0 11132 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_126
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_130
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_12  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_16_192
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_2  _150_
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _144_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_28
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_45
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_49
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_54
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_58
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_78
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_85
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_89
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_107
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_111
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 590 592
use scs8hd_decap_3  FILLER_17_119
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_149
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _066_
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_166
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_173
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_177
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _131_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_187
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_191
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _148_
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_199
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_203
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 20884 0 1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_17_211
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1472 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 2668 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_19
timestamp 1586364061
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_45
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_53
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_71
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9752 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_109
timestamp 1586364061
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_120
timestamp 1586364061
transform 1 0 12144 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_124
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_139
timestamp 1586364061
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_143
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_180
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_197
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_209
timestamp 1586364061
transform 1 0 20332 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_8
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_17
timestamp 1586364061
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_21
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_25
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_41
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_29
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_45
timestamp 1586364061
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_52
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_47
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_55
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_60
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_73
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_74
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_85
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_86
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_8  FILLER_20_96
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_100
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_104
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_108
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_124
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_113
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_149
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_139
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_143
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_153
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_166
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_170
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_187
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_191
timestamp 1586364061
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_191
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_198
timestamp 1586364061
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_202
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_206
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 590 592
use scs8hd_decap_8  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 20884 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_6
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_10
timestamp 1586364061
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_23
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_42
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_46
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_76
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_84
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_87
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_102
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_106
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_149
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_166
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_170
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_173
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_187
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_191
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_198
timestamp 1586364061
transform 1 0 19320 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_202
timestamp 1586364061
transform 1 0 19688 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 20884 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_210
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2116 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_8
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_22
timestamp 1586364061
transform 1 0 3128 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_26
timestamp 1586364061
transform 1 0 3496 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_43
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_22_55
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_22_69
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_73
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_86
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_4  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_99
timestamp 1586364061
transform 1 0 10212 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_112
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_137
timestamp 1586364061
transform 1 0 13708 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_147
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_174
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_185
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_197
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_209
timestamp 1586364061
transform 1 0 20332 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 1656 0 1 14688
box -38 -48 1050 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_17
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_21
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_26
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_41
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_45
timestamp 1586364061
transform 1 0 5244 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_52
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_76
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_80
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_140
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 314 592
use scs8hd_buf_2  _146_
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_166
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_170
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_174
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_182
timestamp 1586364061
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_187
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_191
timestamp 1586364061
transform 1 0 18676 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_203
timestamp 1586364061
transform 1 0 19780 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 20884 0 1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_23_211
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_8
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_47
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_55
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_74
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_4  FILLER_24_112
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_133
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_174
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_186
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_198
timestamp 1586364061
transform 1 0 19320 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_2  _154_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_28
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_32
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_36
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_47
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_buf_2  _149_
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_73
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_89
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_104
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_108
timestamp 1586364061
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_116
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_120
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13340 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_129
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_144
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_148
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_155
timestamp 1586364061
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_166
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_170
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_25_192
timestamp 1586364061
transform 1 0 18768 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 20884 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_209
timestamp 1586364061
transform 1 0 20332 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1564 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_16
timestamp 1586364061
transform 1 0 2576 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_20
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_24
timestamp 1586364061
transform 1 0 3312 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_21
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_25
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_28
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_38
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_37
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__D
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_42
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_46
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _058_
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 8280 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_76
timestamp 1586364061
transform 1 0 8096 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_71
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_27_90
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_95
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_108
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_27_107
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 11592 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_123
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_112
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_127
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_142
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_146
timestamp 1586364061
transform 1 0 14536 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_152
timestamp 1586364061
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use scs8hd_conb_1  _133_
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_157
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_164
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_169
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_176
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_181
timestamp 1586364061
transform 1 0 17756 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_26_193
timestamp 1586364061
transform 1 0 18860 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_182
timestamp 1586364061
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_2  _152_
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_199
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 20884 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 406 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_12
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_16
timestamp 1586364061
transform 1 0 2576 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_or4_4  _091_
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_41
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_45
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_49
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_59
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _056_
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_73
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _062_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__060__B
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_113
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_124
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_147
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_158
timestamp 1586364061
transform 1 0 15640 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_170
timestamp 1586364061
transform 1 0 16744 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_182
timestamp 1586364061
transform 1 0 17848 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_194
timestamp 1586364061
transform 1 0 18952 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_29
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_48
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_52
timestamp 1586364061
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_56
timestamp 1586364061
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_75
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _060_
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _134_
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_99
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 406 592
use scs8hd_decap_6  FILLER_29_106
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use scs8hd_decap_6  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 590 592
use scs8hd_buf_2  _157_
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_129
timestamp 1586364061
transform 1 0 12972 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_134
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_138
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_29_150
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 590 592
use scs8hd_buf_2  _156_
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_160
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_164
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 590 592
use scs8hd_buf_2  _153_
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 20884 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_22
timestamp 1586364061
transform 1 0 3128 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_38
timestamp 1586364061
transform 1 0 4600 0 -1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 5704 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_42
timestamp 1586364061
transform 1 0 4968 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_47
timestamp 1586364061
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_59
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_76
timestamp 1586364061
transform 1 0 8096 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_96
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_108
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_115
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_127
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_139
timestamp 1586364061
transform 1 0 13892 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_151
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_210
timestamp 1586364061
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use scs8hd_conb_1  _132_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_6
timestamp 1586364061
transform 1 0 1656 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_10
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_17
timestamp 1586364061
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_21
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 774 592
use scs8hd_conb_1  _138_
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_29
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_35
timestamp 1586364061
transform 1 0 4324 0 1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 5244 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_54
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 774 592
use scs8hd_conb_1  _137_
timestamp 1586364061
transform 1 0 6900 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_66
timestamp 1586364061
transform 1 0 7176 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_77
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_81
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_108
timestamp 1586364061
transform 1 0 11040 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_112
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_125
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_137
timestamp 1586364061
transform 1 0 13708 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_168
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_180
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_187
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_199
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 20884 0 1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_31_211
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 130 592
<< labels >>
rlabel metal3 s 21520 824 22000 944 6 address[0]
port 0 nsew default input
rlabel metal3 s 21520 2456 22000 2576 6 address[1]
port 1 nsew default input
rlabel metal2 s 4434 0 4490 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 1030 21520 1086 22000 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 416 480 536 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 1368 480 1488 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 2456 480 2576 6 address[6]
port 6 nsew default input
rlabel metal3 s 0 3544 480 3664 6 bottom_grid_pin_0_
port 7 nsew default tristate
rlabel metal2 s 3146 21520 3202 22000 6 bottom_grid_pin_4_
port 8 nsew default tristate
rlabel metal2 s 5354 21520 5410 22000 6 bottom_grid_pin_8_
port 9 nsew default tristate
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 21520 4088 22000 4208 6 chanx_left_in[1]
port 11 nsew default input
rlabel metal2 s 7562 21520 7618 22000 6 chanx_left_in[2]
port 12 nsew default input
rlabel metal3 s 21520 5856 22000 5976 6 chanx_left_in[3]
port 13 nsew default input
rlabel metal3 s 21520 7488 22000 7608 6 chanx_left_in[4]
port 14 nsew default input
rlabel metal3 s 21520 9256 22000 9376 6 chanx_left_in[5]
port 15 nsew default input
rlabel metal2 s 6274 0 6330 480 6 chanx_left_in[6]
port 16 nsew default input
rlabel metal3 s 0 5584 480 5704 6 chanx_left_in[7]
port 17 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[8]
port 18 nsew default input
rlabel metal3 s 21520 10888 22000 11008 6 chanx_left_out[0]
port 19 nsew default tristate
rlabel metal2 s 9770 21520 9826 22000 6 chanx_left_out[1]
port 20 nsew default tristate
rlabel metal3 s 21520 12656 22000 12776 6 chanx_left_out[2]
port 21 nsew default tristate
rlabel metal3 s 0 7760 480 7880 6 chanx_left_out[3]
port 22 nsew default tristate
rlabel metal3 s 21520 14288 22000 14408 6 chanx_left_out[4]
port 23 nsew default tristate
rlabel metal2 s 8114 0 8170 480 6 chanx_left_out[5]
port 24 nsew default tristate
rlabel metal3 s 0 8712 480 8832 6 chanx_left_out[6]
port 25 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[7]
port 26 nsew default tristate
rlabel metal2 s 9954 0 10010 480 6 chanx_left_out[8]
port 27 nsew default tristate
rlabel metal3 s 0 10888 480 11008 6 chanx_right_in[0]
port 28 nsew default input
rlabel metal3 s 21520 16056 22000 16176 6 chanx_right_in[1]
port 29 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_right_in[2]
port 30 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_right_in[3]
port 31 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chanx_right_in[4]
port 32 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_right_in[5]
port 33 nsew default input
rlabel metal3 s 0 15104 480 15224 6 chanx_right_in[6]
port 34 nsew default input
rlabel metal2 s 11978 21520 12034 22000 6 chanx_right_in[7]
port 35 nsew default input
rlabel metal2 s 13634 0 13690 480 6 chanx_right_in[8]
port 36 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chanx_right_out[0]
port 37 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chanx_right_out[1]
port 38 nsew default tristate
rlabel metal2 s 14186 21520 14242 22000 6 chanx_right_out[2]
port 39 nsew default tristate
rlabel metal2 s 16394 21520 16450 22000 6 chanx_right_out[3]
port 40 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chanx_right_out[4]
port 41 nsew default tristate
rlabel metal3 s 0 16056 480 16176 6 chanx_right_out[5]
port 42 nsew default tristate
rlabel metal2 s 18602 21520 18658 22000 6 chanx_right_out[6]
port 43 nsew default tristate
rlabel metal3 s 21520 17688 22000 17808 6 chanx_right_out[7]
port 44 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chanx_right_out[8]
port 45 nsew default tristate
rlabel metal2 s 2594 0 2650 480 6 data_in
port 46 nsew default input
rlabel metal2 s 846 0 902 480 6 enable
port 47 nsew default input
rlabel metal3 s 21520 19456 22000 19576 6 top_grid_pin_0_
port 48 nsew default tristate
rlabel metal2 s 20994 0 21050 480 6 top_grid_pin_10_
port 49 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 top_grid_pin_12_
port 50 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 top_grid_pin_14_
port 51 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 top_grid_pin_2_
port 52 nsew default tristate
rlabel metal2 s 20810 21520 20866 22000 6 top_grid_pin_4_
port 53 nsew default tristate
rlabel metal3 s 21520 21088 22000 21208 6 top_grid_pin_6_
port 54 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 top_grid_pin_8_
port 55 nsew default tristate
rlabel metal4 s 4611 2128 4931 19632 6 vpwr
port 56 nsew default input
rlabel metal4 s 8277 2128 8597 19632 6 vgnd
port 57 nsew default input
<< end >>
