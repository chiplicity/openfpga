VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__2_
  CLASS BLOCK ;
  FOREIGN sb_0__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 115.000 BY 115.000 ;
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 111.000 28.890 115.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END SC_OUT_BOT
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END bottom_left_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 111.000 86.390 115.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 19.080 115.000 19.680 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 41.520 115.000 42.120 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 44.240 115.000 44.840 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 46.280 115.000 46.880 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 48.320 115.000 48.920 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 51.040 115.000 51.640 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 53.080 115.000 53.680 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 55.800 115.000 56.400 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 57.840 115.000 58.440 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 59.880 115.000 60.480 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 62.600 115.000 63.200 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 21.120 115.000 21.720 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 23.160 115.000 23.760 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 25.880 115.000 26.480 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 27.920 115.000 28.520 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 29.960 115.000 30.560 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 32.680 115.000 33.280 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 34.720 115.000 35.320 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 37.440 115.000 38.040 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 39.480 115.000 40.080 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 64.640 115.000 65.240 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 87.760 115.000 88.360 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 89.800 115.000 90.400 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 92.520 115.000 93.120 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 94.560 115.000 95.160 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 96.600 115.000 97.200 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 99.320 115.000 99.920 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 101.360 115.000 101.960 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 104.080 115.000 104.680 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 106.120 115.000 106.720 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 108.160 115.000 108.760 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 67.360 115.000 67.960 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 69.400 115.000 70.000 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 71.440 115.000 72.040 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 74.160 115.000 74.760 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 76.200 115.000 76.800 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 78.240 115.000 78.840 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 80.960 115.000 81.560 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 83.000 115.000 83.600 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 85.720 115.000 86.320 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END chany_bottom_out[9]
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 110.880 115.000 111.480 ;
    END
  END prog_clk_0_E_in
  PIN right_bottom_grid_pin_34_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 0.720 115.000 1.320 ;
    END
  END right_bottom_grid_pin_34_
  PIN right_bottom_grid_pin_35_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 2.760 115.000 3.360 ;
    END
  END right_bottom_grid_pin_35_
  PIN right_bottom_grid_pin_36_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 4.800 115.000 5.400 ;
    END
  END right_bottom_grid_pin_36_
  PIN right_bottom_grid_pin_37_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 7.520 115.000 8.120 ;
    END
  END right_bottom_grid_pin_37_
  PIN right_bottom_grid_pin_38_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 9.560 115.000 10.160 ;
    END
  END right_bottom_grid_pin_38_
  PIN right_bottom_grid_pin_39_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 11.600 115.000 12.200 ;
    END
  END right_bottom_grid_pin_39_
  PIN right_bottom_grid_pin_40_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 14.320 115.000 14.920 ;
    END
  END right_bottom_grid_pin_40_
  PIN right_bottom_grid_pin_41_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 16.360 115.000 16.960 ;
    END
  END right_bottom_grid_pin_41_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 112.920 115.000 113.520 ;
    END
  END right_top_grid_pin_1_
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 91.355 10.640 92.955 103.600 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 56.700 10.640 58.300 103.600 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.045 10.640 23.645 103.600 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.025 10.640 75.625 103.600 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.375 10.640 40.975 103.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 110.255 103.445 ;
      LAYER met1 ;
        RECT 3.290 6.840 110.790 103.600 ;
      LAYER met2 ;
        RECT 1.010 110.720 28.330 113.405 ;
        RECT 29.170 110.720 85.830 113.405 ;
        RECT 86.670 110.720 113.530 113.405 ;
        RECT 1.010 4.280 113.530 110.720 ;
        RECT 1.570 0.835 3.030 4.280 ;
        RECT 3.870 0.835 5.790 4.280 ;
        RECT 6.630 0.835 8.550 4.280 ;
        RECT 9.390 0.835 11.310 4.280 ;
        RECT 12.150 0.835 14.070 4.280 ;
        RECT 14.910 0.835 16.830 4.280 ;
        RECT 17.670 0.835 19.590 4.280 ;
        RECT 20.430 0.835 22.350 4.280 ;
        RECT 23.190 0.835 25.110 4.280 ;
        RECT 25.950 0.835 27.870 4.280 ;
        RECT 28.710 0.835 30.630 4.280 ;
        RECT 31.470 0.835 33.390 4.280 ;
        RECT 34.230 0.835 36.150 4.280 ;
        RECT 36.990 0.835 38.910 4.280 ;
        RECT 39.750 0.835 41.670 4.280 ;
        RECT 42.510 0.835 44.430 4.280 ;
        RECT 45.270 0.835 47.190 4.280 ;
        RECT 48.030 0.835 49.950 4.280 ;
        RECT 50.790 0.835 52.710 4.280 ;
        RECT 53.550 0.835 55.470 4.280 ;
        RECT 56.310 0.835 58.230 4.280 ;
        RECT 59.070 0.835 60.530 4.280 ;
        RECT 61.370 0.835 63.290 4.280 ;
        RECT 64.130 0.835 66.050 4.280 ;
        RECT 66.890 0.835 68.810 4.280 ;
        RECT 69.650 0.835 71.570 4.280 ;
        RECT 72.410 0.835 74.330 4.280 ;
        RECT 75.170 0.835 77.090 4.280 ;
        RECT 77.930 0.835 79.850 4.280 ;
        RECT 80.690 0.835 82.610 4.280 ;
        RECT 83.450 0.835 85.370 4.280 ;
        RECT 86.210 0.835 88.130 4.280 ;
        RECT 88.970 0.835 90.890 4.280 ;
        RECT 91.730 0.835 93.650 4.280 ;
        RECT 94.490 0.835 96.410 4.280 ;
        RECT 97.250 0.835 99.170 4.280 ;
        RECT 100.010 0.835 101.930 4.280 ;
        RECT 102.770 0.835 104.690 4.280 ;
        RECT 105.530 0.835 107.450 4.280 ;
        RECT 108.290 0.835 110.210 4.280 ;
        RECT 111.050 0.835 112.970 4.280 ;
      LAYER met3 ;
        RECT 0.985 112.520 110.600 113.385 ;
        RECT 0.985 111.880 113.555 112.520 ;
        RECT 0.985 110.480 110.600 111.880 ;
        RECT 0.985 109.160 113.555 110.480 ;
        RECT 0.985 107.760 110.600 109.160 ;
        RECT 0.985 107.120 113.555 107.760 ;
        RECT 0.985 105.720 110.600 107.120 ;
        RECT 0.985 105.080 113.555 105.720 ;
        RECT 0.985 103.680 110.600 105.080 ;
        RECT 0.985 102.360 113.555 103.680 ;
        RECT 0.985 100.960 110.600 102.360 ;
        RECT 0.985 100.320 113.555 100.960 ;
        RECT 0.985 98.920 110.600 100.320 ;
        RECT 0.985 97.600 113.555 98.920 ;
        RECT 0.985 96.200 110.600 97.600 ;
        RECT 0.985 95.560 113.555 96.200 ;
        RECT 0.985 94.160 110.600 95.560 ;
        RECT 0.985 93.520 113.555 94.160 ;
        RECT 0.985 92.120 110.600 93.520 ;
        RECT 0.985 90.800 113.555 92.120 ;
        RECT 0.985 89.400 110.600 90.800 ;
        RECT 0.985 88.760 113.555 89.400 ;
        RECT 0.985 87.360 110.600 88.760 ;
        RECT 0.985 86.720 113.555 87.360 ;
        RECT 0.985 85.320 110.600 86.720 ;
        RECT 0.985 84.000 113.555 85.320 ;
        RECT 0.985 82.600 110.600 84.000 ;
        RECT 0.985 81.960 113.555 82.600 ;
        RECT 0.985 80.560 110.600 81.960 ;
        RECT 0.985 79.240 113.555 80.560 ;
        RECT 0.985 77.840 110.600 79.240 ;
        RECT 0.985 77.200 113.555 77.840 ;
        RECT 0.985 75.800 110.600 77.200 ;
        RECT 0.985 75.160 113.555 75.800 ;
        RECT 0.985 73.760 110.600 75.160 ;
        RECT 0.985 72.440 113.555 73.760 ;
        RECT 0.985 71.040 110.600 72.440 ;
        RECT 0.985 70.400 113.555 71.040 ;
        RECT 0.985 69.000 110.600 70.400 ;
        RECT 0.985 68.360 113.555 69.000 ;
        RECT 0.985 66.960 110.600 68.360 ;
        RECT 0.985 65.640 113.555 66.960 ;
        RECT 0.985 64.240 110.600 65.640 ;
        RECT 0.985 63.600 113.555 64.240 ;
        RECT 0.985 62.200 110.600 63.600 ;
        RECT 0.985 60.880 113.555 62.200 ;
        RECT 0.985 59.480 110.600 60.880 ;
        RECT 0.985 58.840 113.555 59.480 ;
        RECT 0.985 58.160 110.600 58.840 ;
        RECT 4.400 57.440 110.600 58.160 ;
        RECT 4.400 56.800 113.555 57.440 ;
        RECT 4.400 56.760 110.600 56.800 ;
        RECT 0.985 55.400 110.600 56.760 ;
        RECT 0.985 54.080 113.555 55.400 ;
        RECT 0.985 52.680 110.600 54.080 ;
        RECT 0.985 52.040 113.555 52.680 ;
        RECT 0.985 50.640 110.600 52.040 ;
        RECT 0.985 49.320 113.555 50.640 ;
        RECT 0.985 47.920 110.600 49.320 ;
        RECT 0.985 47.280 113.555 47.920 ;
        RECT 0.985 45.880 110.600 47.280 ;
        RECT 0.985 45.240 113.555 45.880 ;
        RECT 0.985 43.840 110.600 45.240 ;
        RECT 0.985 42.520 113.555 43.840 ;
        RECT 0.985 41.120 110.600 42.520 ;
        RECT 0.985 40.480 113.555 41.120 ;
        RECT 0.985 39.080 110.600 40.480 ;
        RECT 0.985 38.440 113.555 39.080 ;
        RECT 0.985 37.040 110.600 38.440 ;
        RECT 0.985 35.720 113.555 37.040 ;
        RECT 0.985 34.320 110.600 35.720 ;
        RECT 0.985 33.680 113.555 34.320 ;
        RECT 0.985 32.280 110.600 33.680 ;
        RECT 0.985 30.960 113.555 32.280 ;
        RECT 0.985 29.560 110.600 30.960 ;
        RECT 0.985 28.920 113.555 29.560 ;
        RECT 0.985 27.520 110.600 28.920 ;
        RECT 0.985 26.880 113.555 27.520 ;
        RECT 0.985 25.480 110.600 26.880 ;
        RECT 0.985 24.160 113.555 25.480 ;
        RECT 0.985 22.760 110.600 24.160 ;
        RECT 0.985 22.120 113.555 22.760 ;
        RECT 0.985 20.720 110.600 22.120 ;
        RECT 0.985 20.080 113.555 20.720 ;
        RECT 0.985 18.680 110.600 20.080 ;
        RECT 0.985 17.360 113.555 18.680 ;
        RECT 0.985 15.960 110.600 17.360 ;
        RECT 0.985 15.320 113.555 15.960 ;
        RECT 0.985 13.920 110.600 15.320 ;
        RECT 0.985 12.600 113.555 13.920 ;
        RECT 0.985 11.200 110.600 12.600 ;
        RECT 0.985 10.560 113.555 11.200 ;
        RECT 0.985 9.160 110.600 10.560 ;
        RECT 0.985 8.520 113.555 9.160 ;
        RECT 0.985 7.120 110.600 8.520 ;
        RECT 0.985 5.800 113.555 7.120 ;
        RECT 0.985 4.400 110.600 5.800 ;
        RECT 0.985 3.760 113.555 4.400 ;
        RECT 0.985 2.360 110.600 3.760 ;
        RECT 0.985 1.720 113.555 2.360 ;
        RECT 0.985 0.855 110.600 1.720 ;
      LAYER met4 ;
        RECT 41.375 10.640 56.300 103.600 ;
        RECT 58.700 10.640 73.625 103.600 ;
        RECT 76.025 10.640 90.955 103.600 ;
  END
END sb_0__2_
END LIBRARY

