* NGSPICE file created from sb_1__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt sb_1__0_ SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] left_bottom_grid_pin_11_ left_bottom_grid_pin_1_ left_bottom_grid_pin_3_
+ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_ prog_clk
+ right_bottom_grid_pin_11_ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_
+ right_bottom_grid_pin_7_ right_bottom_grid_pin_9_ top_left_grid_pin_42_ top_left_grid_pin_43_
+ top_left_grid_pin_44_ top_left_grid_pin_45_ top_left_grid_pin_46_ top_left_grid_pin_47_
+ top_left_grid_pin_48_ top_left_grid_pin_49_ VPWR VGND
XFILLER_39_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_0.mux_l3_in_0_/S mux_right_track_2.mux_l1_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_42_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_9.mux_l3_in_0_/S mux_left_track_17.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A1 mux_left_track_25.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 top_left_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_062_ _062_/A chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_10.mux_l3_in_0_ mux_top_track_10.mux_l2_in_1_/X mux_top_track_10.mux_l2_in_0_/X
+ mux_top_track_10.mux_l3_in_0_/S mux_top_track_10.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_6.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_114_ _114_/A chany_top_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_045_ _045_/HI _045_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l2_in_1__A1 left_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__S mux_left_track_17.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_10.mux_l2_in_1_ _030_/HI chanx_left_in[9] mux_top_track_10.mux_l2_in_0_/S
+ mux_top_track_10.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_9.mux_l1_in_3__A0 _049_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__S mux_right_track_16.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_028_ _028_/HI _028_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 right_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l2_in_1__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l3_in_0__A1 mux_left_track_33.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_6.mux_l1_in_2__S mux_top_track_6.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A mux_left_track_1.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_061_ chanx_right_in[16] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_10.mux_l2_in_0_/S mux_top_track_10.mux_l3_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_4.mux_l4_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l3_in_0_/X _074_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_left_track_1.mux_l2_in_2__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_113_ _113_/A chany_top_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_24.mux_l1_in_0__S mux_top_track_24.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_044_ _044_/HI _044_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_4.mux_l2_in_2__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l3_in_0__S mux_left_track_5.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l3_in_0__S mux_right_track_8.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_10.mux_l2_in_0_ chanx_right_in[19] mux_top_track_10.mux_l1_in_0_/X
+ mux_top_track_10.mux_l2_in_0_/S mux_top_track_10.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_3__A1 left_bottom_grid_pin_9_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A mux_top_track_20.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l3_in_0_/X _066_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_track_0.mux_l2_in_3_ _029_/HI chanx_left_in[2] mux_top_track_0.mux_l2_in_3_/S
+ mux_top_track_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_1__S mux_left_track_33.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l2_in_1__S mux_right_track_32.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_10.mux_l2_in_0__A0 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_3__A0 right_bottom_grid_pin_9_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_10.mux_l1_in_0_/S mux_top_track_10.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_060_ chanx_right_in[17] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S mux_top_track_0.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l2_in_0__S mux_top_track_16.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_track_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_2__A0 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__061__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_112_ _112_/A chany_top_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_043_ _043_/HI _043_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_0_/S mux_top_track_0.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__056__A SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l3_in_1__A0 mux_right_track_4.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l2_in_1__S mux_left_track_25.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_2_ chanx_left_in[0] chanx_right_in[2] mux_top_track_0.mux_l2_in_3_/S
+ mux_top_track_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_10.mux_l1_in_0_ chanx_right_in[9] top_left_grid_pin_43_ mux_top_track_10.mux_l1_in_0_/S
+ mux_top_track_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 top_left_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l4_in_0__A0 mux_right_track_4.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_22.mux_l2_in_0_ mux_top_track_22.mux_l1_in_1_/X mux_top_track_22.mux_l1_in_0_/X
+ mux_top_track_22.mux_l2_in_0_/S mux_top_track_22.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_10.mux_l2_in_0__A1 mux_top_track_10.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_3.mux_l1_in_0__S mux_left_track_3.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A mux_top_track_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__064__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l1_in_3_ _028_/HI chanx_left_in[16] mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_3__A1 right_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l1_in_2__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0__A0 mux_top_track_2.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__059__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_22.mux_l1_in_1_ _037_/HI chanx_left_in[17] mux_top_track_22.mux_l1_in_0_/S
+ mux_top_track_22.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_8.mux_l3_in_0_/S mux_top_track_10.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_6.mux_l2_in_0__S mux_top_track_6.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_2__A1 right_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_2__A0 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_111_ _111_/A chany_top_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_042_ _042_/HI _042_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S mux_top_track_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__072__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_4.mux_l3_in_1__A1 mux_right_track_4.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_16.mux_l1_in_1_/S mux_top_track_16.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_0.mux_l3_in_1__A0 mux_top_track_0.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_20.mux_l1_in_0__S mux_top_track_20.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l1_in_3__S mux_left_track_3.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__S mux_left_track_1.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__067__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_8.mux_l2_in_1_ mux_right_track_8.mux_l1_in_3_/X mux_right_track_8.mux_l1_in_2_/X
+ mux_right_track_8.mux_l2_in_1_/S mux_right_track_8.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ chanx_right_in[1] top_left_grid_pin_48_ mux_top_track_0.mux_l2_in_3_/S
+ mux_top_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A1 top_left_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l4_in_0__A1 mux_right_track_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l4_in_0__A0 mux_top_track_0.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_22.sky130_fd_sc_hd__buf_4_0_ mux_top_track_22.mux_l2_in_0_/X _107_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__080__A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l1_in_2_ chanx_left_in[6] right_bottom_grid_pin_9_ mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l2_in_0__A1 mux_top_track_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_14.mux_l1_in_0__A0 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A0 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l2_in_0_/X _110_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_track_22.mux_l1_in_0_ chanx_right_in[17] top_left_grid_pin_49_ mux_top_track_22.mux_l1_in_0_/S
+ mux_top_track_22.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__075__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_22.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_2__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_110_ _110_/A chany_top_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A mux_top_track_6.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_041_ _041_/HI _041_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_12.mux_l2_in_0__S mux_top_track_12.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_8.mux_l1_in_2__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_18.mux_l1_in_1__S mux_top_track_18.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_14.mux_l2_in_0_/S mux_top_track_16.mux_l1_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l3_in_1__A1 mux_top_track_0.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__083__A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l4_in_0_/X _118_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l2_in_0_ mux_right_track_8.mux_l1_in_1_/X mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_1_/S mux_right_track_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 mux_right_track_8.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ top_left_grid_pin_46_ mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_3_/S mux_top_track_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__078__A _078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l4_in_0__A1 mux_top_track_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_22.mux_l1_in_0__A0 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.mux_l1_in_1_ right_bottom_grid_pin_1_ chany_top_in[16] mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l3_in_0__A0 mux_right_track_8.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0__A1 top_left_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A1 mux_left_track_1.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__091__A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0__A0 top_left_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__086__A _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_38.sky130_fd_sc_hd__buf_4_0_ mux_top_track_38.mux_l2_in_0_/X _099_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_3_3_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_040_ _040_/HI _040_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_2.mux_l2_in_0__S mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_2__A1 right_bottom_grid_pin_9_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A0 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_24.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 mux_right_track_8.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_4.mux_l2_in_1__A0 mux_top_track_4.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A0 right_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__094__A _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_22.mux_l1_in_0__A1 top_left_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_3.mux_l2_in_1__S mux_left_track_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l1_in_0_ chany_top_in[9] chany_top_in[2] mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l3_in_0__A1 mux_right_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_38.mux_l1_in_0__S mux_top_track_38.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__089__A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A0 mux_top_track_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_44_ top_left_grid_pin_42_ mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2__S mux_left_track_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l4_in_0__S mux_top_track_0.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 mux_right_track_16.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l3_in_0_/X _094_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_6.mux_l1_in_0__A1 top_left_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_099_ _099_/A chany_top_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_2__A0 left_bottom_grid_pin_7_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A mux_right_track_0.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__097__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A0 right_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A mux_top_track_12.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l3_in_0_/X _082_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_15_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_24.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l1_in_1__S mux_top_track_14.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l2_in_1__A1 mux_top_track_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 _033_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_1__A0 mux_left_track_3.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_42_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 mux_right_track_24.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l2_in_3__A0 _043_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l3_in_0__A1 mux_top_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A0 mux_top_track_16.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A0 mux_left_track_3.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l4_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l3_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_098_ _098_/A chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.mux_l1_in_1__A0 right_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_2__A1 left_bottom_grid_pin_3_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_28_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_24.mux_l1_in_1__A0 _038_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_14.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_4.mux_l1_in_1__S mux_top_track_4.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l2_in_0__A0 mux_right_track_32.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 mux_left_track_3.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l4_in_0_/X _076_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 mux_top_track_24.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l2_in_3__A1 left_bottom_grid_pin_9_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_37_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A1 mux_left_track_3.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A1 mux_top_track_16.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A mux_top_track_18.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l3_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_3__A0 _041_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A mux_right_track_32.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_5.mux_l1_in_2__S mux_left_track_5.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l1_in_3_ _046_/HI left_bottom_grid_pin_11_ mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_2__S mux_right_track_8.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l2_in_3_ _055_/HI chanx_left_in[14] mux_right_track_4.mux_l2_in_1_/S
+ mux_right_track_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_097_ _097_/A chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.mux_l1_in_1__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_4.mux_l2_in_0_/S mux_top_track_4.mux_l3_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_17.mux_l1_in_1__A0 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l2_in_0__A1 mux_right_track_32.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_24.mux_l2_in_0__A1 mux_top_track_24.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_0_/S mux_right_track_4.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_17.mux_l2_in_0__A0 mux_left_track_17.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_1.mux_l1_in_0_/S mux_left_track_1.mux_l2_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_1_ mux_left_track_3.mux_l1_in_3_/X mux_left_track_3.mux_l1_in_2_/X
+ mux_left_track_3.mux_l2_in_0_/S mux_left_track_3.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_3.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_3__A0 left_bottom_grid_pin_5_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_3__A1 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_0__A1 mux_top_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A mux_left_track_33.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__100__A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_2.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l4_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l1_in_2_ left_bottom_grid_pin_7_ left_bottom_grid_pin_3_ mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_2_ chanx_left_in[5] right_bottom_grid_pin_11_ mux_right_track_4.mux_l2_in_1_/S
+ mux_right_track_4.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l2_in_2__A0 left_bottom_grid_pin_9_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_096_ _096_/A chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_4.mux_l1_in_0_/S mux_top_track_4.mux_l2_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_079_ chanx_left_in[18] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_3_ _051_/HI chanx_left_in[17] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_3_ right_bottom_grid_pin_9_ right_bottom_grid_pin_7_
+ mux_right_track_4.mux_l1_in_1_/S mux_right_track_4.mux_l1_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l3_in_1__A0 mux_left_track_5.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0__S mux_left_track_17.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A0 mux_left_track_25.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_1_ _033_/HI chanx_left_in[13] mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_20.mux_l1_in_0_/S mux_top_track_20.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_33.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_17.mux_l2_in_0__A1 mux_left_track_17.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__103__A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l4_in_0__A0 mux_left_track_5.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_32.mux_l3_in_0_/S mux_left_track_1.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_0_/S mux_left_track_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S mux_right_track_16.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_3__A1 left_bottom_grid_pin_3_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l1_in_1__A0 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__D mux_left_track_17.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l3_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l1_in_1_ chanx_right_in[13] chanx_right_in[4] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_1_ mux_right_track_16.mux_l1_in_3_/X mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_0_/S mux_right_track_16.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_3__S mux_left_track_17.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_095_ chanx_left_in[2] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_5.mux_l2_in_2__A1 left_bottom_grid_pin_7_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__111__A _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_2.mux_l3_in_0_/S mux_top_track_4.mux_l1_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_33.mux_l2_in_0__A0 mux_left_track_33.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_2__S mux_right_track_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_078_ _078_/A chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_0.mux_l1_in_3__A0 _050_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__106__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_12.sky130_fd_sc_hd__buf_4_0_ mux_top_track_12.mux_l2_in_0_/X _112_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_left_track_5.mux_l2_in_0__S mux_left_track_5.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_2_ chanx_left_in[8] right_bottom_grid_pin_11_ mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_2_ right_bottom_grid_pin_5_ right_bottom_grid_pin_3_
+ mux_right_track_4.mux_l1_in_1_/S mux_right_track_4.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l3_in_1__A1 mux_left_track_5.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l2_in_0__A1 mux_left_track_25.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l1_in_0_ chanx_right_in[13] top_left_grid_pin_46_ mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_18.mux_l2_in_0_/S mux_top_track_20.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_8.mux_l3_in_0__S mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l4_in_0__A1 mux_left_track_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l1_in_3_ _041_/HI chanx_left_in[6] mux_top_track_6.mux_l1_in_0_/S
+ mux_top_track_6.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__114__A _114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_32.mux_l1_in_1__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l1_in_1__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_22.mux_l2_in_0__S mux_top_track_22.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__109__A _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_4.mux_l1_in_1_/S mux_right_track_4.mux_l2_in_1_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_5.mux_l2_in_3__S mux_left_track_5.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[6] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__D mux_left_track_3.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_0_/S mux_right_track_16.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0__S mux_top_track_16.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l3_in_0_ mux_top_track_6.mux_l2_in_1_/X mux_top_track_6.mux_l2_in_0_/X
+ mux_top_track_6.mux_l3_in_0_/S mux_top_track_6.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_094_ _094_/A chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_17.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l2_in_0__A1 mux_left_track_33.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_3__A1 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2__A0 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_077_ _077_/A chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_1_ right_bottom_grid_pin_3_ chany_top_in[17] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_1_ chany_top_in[15] mux_right_track_4.mux_l1_in_1_/S
+ mux_right_track_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_6.mux_l2_in_1_ mux_top_track_6.mux_l1_in_3_/X mux_top_track_6.mux_l1_in_2_/X
+ mux_top_track_6.mux_l2_in_0_/S mux_top_track_6.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__117__A _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 mux_left_track_9.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_25.mux_l1_in_1__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_24.mux_l2_in_1__S mux_right_track_24.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__D mux_left_track_5.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l1_in_2_ chanx_right_in[11] chanx_right_in[6] mux_top_track_6.mux_l1_in_0_/S
+ mux_top_track_6.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l3_in_0__A0 mux_left_track_9.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_2.mux_l4_in_0_/S mux_right_track_4.mux_l1_in_1_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_6.mux_l1_in_0__S mux_top_track_6.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_093_ chanx_left_in[4] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l1_in_2__A1 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_076_ _076_/A chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l1_in_0_ chany_top_in[10] chany_top_in[3] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_0_ chany_top_in[8] chany_top_in[1] mux_right_track_4.mux_l1_in_1_/S
+ mux_right_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_10.mux_l1_in_0__A0 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l2_in_0_ mux_top_track_6.mux_l1_in_1_/X mux_top_track_6.mux_l1_in_0_/X
+ mux_top_track_6.mux_l2_in_0_/S mux_top_track_6.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l4_in_0_/X _096_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_left_track_17.mux_l2_in_1__S mux_left_track_17.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_059_ chanx_right_in[18] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_0.mux_l1_in_2__S mux_right_track_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 mux_left_track_9.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_6.sky130_fd_sc_hd__buf_4_0_ mux_top_track_6.mux_l3_in_0_/X _115_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_35_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_2__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l1_in_1_ top_left_grid_pin_49_ top_left_grid_pin_47_ mux_top_track_6.mux_l1_in_0_/S
+ mux_top_track_6.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 right_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_3__S mux_top_track_6.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_4.mux_l3_in_0__S mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l3_in_0__A1 mux_left_track_9.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A mux_right_track_24.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 mux_right_track_4.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_092_ chanx_left_in[5] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A mux_left_track_3.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_3__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_3__A0 _052_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_24.mux_l1_in_1__S mux_top_track_24.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_075_ chanx_right_in[2] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_20.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_3__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0__S mux_top_track_12.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l4_in_0__S mux_right_track_2.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l3_in_1__S mux_left_track_5.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l3_in_0_/X _090_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_10.mux_l1_in_0__A1 top_left_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_38.mux_l2_in_0__A0 _039_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ _058_/A SC_OUT_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 top_left_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_6.mux_l1_in_0_ top_left_grid_pin_45_ top_left_grid_pin_43_ mux_top_track_6.mux_l1_in_0_/S
+ mux_top_track_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 right_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_38.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A mux_left_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A mux_top_track_22.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 mux_right_track_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_10.mux_l3_in_0__S mux_top_track_10.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l4_in_0_/X _078_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_091_ chanx_left_in[6] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_3__A1 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__062__A _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_074_ _074_/A chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l3_in_0__A0 mux_top_track_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_12.mux_l1_in_0_/S mux_top_track_12.mux_l2_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_38.mux_l2_in_0__A1 mux_top_track_38.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_057_ _057_/A SC_OUT_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 top_left_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A mux_left_track_9.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_109_ _109_/A chany_top_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__070__A _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_1__S mux_left_track_3.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__065__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l1_in_3__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_0.mux_l3_in_0__S mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_0.mux_l2_in_1__A1 top_left_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.mux_l1_in_1__A0 _031_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_6.mux_l2_in_1__S mux_top_track_6.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_090_ _090_/A chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A mux_top_track_2.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_1__A0 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_073_ chanx_right_in[4] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_0.mux_l3_in_0__A1 mux_top_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_12.mux_l2_in_0__A0 mux_top_track_12.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_10.mux_l3_in_0_/S mux_top_track_12.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__073__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 mux_right_track_8.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_056_ SC_IN_BOT SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_38_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_20.mux_l1_in_1__S mux_top_track_20.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__068__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l3_in_1__S mux_left_track_1.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l3_in_1__S mux_right_track_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_108_ _108_/A chany_top_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l1_in_3_ _044_/HI left_bottom_grid_pin_11_ mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_039_ _039_/HI _039_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_18.mux_l1_in_1_/S mux_top_track_18.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_20.mux_l1_in_1__A0 _036_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_12.mux_l2_in_0_ mux_top_track_12.mux_l1_in_1_/X mux_top_track_12.mux_l1_in_0_/X
+ mux_top_track_12.mux_l2_in_0_/S mux_top_track_12.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__081__A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X _062_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_left_track_9.mux_l1_in_3_ _049_/HI left_bottom_grid_pin_9_ mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_12.mux_l1_in_1__A1 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_3_ _050_/HI chanx_left_in[12] mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__076__A _076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S mux_left_track_17.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_33.mux_l2_in_0__S mux_left_track_33.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_20.mux_l2_in_0__A0 mux_top_track_20.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_12.mux_l1_in_1_ _031_/HI chanx_left_in[10] mux_top_track_12.mux_l1_in_0_/S
+ mux_top_track_12.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_1__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l3_in_0__S mux_right_track_32.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_1__A0 top_left_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_072_ chanx_right_in[5] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_12.mux_l2_in_0__A1 mux_top_track_12.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l2_in_1_ mux_left_track_17.mux_l1_in_3_/X mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_3__A0 _035_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_055_ _055_/HI _055_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_4.mux_l2_in_0__A0 mux_top_track_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A mux_top_track_8.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__084__A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_038_ _038_/HI _038_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_2_ left_bottom_grid_pin_3_ chanx_right_in[17] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_107_ _107_/A chany_top_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l2_in_1_ mux_left_track_9.mux_l1_in_3_/X mux_left_track_9.mux_l1_in_2_/X
+ mux_left_track_9.mux_l2_in_0_/S mux_left_track_9.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_16.mux_l2_in_0_/S mux_top_track_18.mux_l1_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__079__A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.mux_l2_in_1_ mux_right_track_0.mux_l1_in_3_/X mux_right_track_0.mux_l1_in_2_/X
+ mux_right_track_0.mux_l2_in_1_/S mux_right_track_0.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_20.mux_l1_in_1__A1 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__S mux_left_track_25.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_9.mux_l1_in_2_ left_bottom_grid_pin_1_ chanx_right_in[16] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_2_ chanx_left_in[2] right_bottom_grid_pin_9_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__092__A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_20.mux_l2_in_0__A1 mux_top_track_20.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_12.mux_l1_in_0_ chanx_right_in[10] top_left_grid_pin_44_ mux_top_track_12.mux_l1_in_0_/S
+ mux_top_track_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S mux_top_track_24.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A1 top_left_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__087__A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_071_ chanx_right_in[6] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_2.mux_l2_in_1__S mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0__S mux_left_track_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l1_in_3_ _035_/HI chanx_left_in[4] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l1_in_3__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_054_ _054_/HI _054_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_track_24.mux_l1_in_1_ _038_/HI chanx_left_in[18] mux_top_track_24.mux_l1_in_1_/S
+ mux_top_track_24.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_0__A0 mux_left_track_3.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0__A1 mux_top_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_037_ _037_/HI _037_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_1_ chanx_right_in[8] chany_top_in[17] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_106_ _106_/A chany_top_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_0_/S mux_left_track_9.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l2_in_2__A0 left_bottom_grid_pin_5_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A mux_right_track_16.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__095__A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_1_/S mux_right_track_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S mux_top_track_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l1_in_1_ chanx_right_in[6] chany_top_in[18] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l3_in_1__A0 mux_left_track_1.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_3__S mux_left_track_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_5_ right_bottom_grid_pin_1_
+ mux_right_track_0.mux_l1_in_1_/S mux_right_track_0.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l2_in_1_ mux_top_track_2.mux_l1_in_3_/X mux_top_track_2.mux_l1_in_2_/X
+ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l2_in_1_ _053_/HI mux_right_track_24.mux_l1_in_2_/X mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l4_in_0__A0 mux_left_track_1.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_070_ _070_/A chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_track_0.mux_l3_in_0_/S mux_top_track_0.mux_l4_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l2_in_0_/X _106_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l1_in_2_ chanx_right_in[4] chanx_right_in[3] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_2_ chanx_left_in[18] chanx_left_in[9] mux_right_track_24.mux_l1_in_2_/S
+ mux_right_track_24.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_22.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__098__A _098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_053_ _053_/HI _053_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 top_left_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[18] top_left_grid_pin_42_ mux_top_track_24.mux_l1_in_1_/S
+ mux_top_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l2_in_0__A1 mux_left_track_3.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_32.mux_l2_in_1_/S
+ mux_right_track_32.mux_l3_in_0_/S clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_18.sky130_fd_sc_hd__buf_4_0_ mux_top_track_18.mux_l2_in_0_/X _109_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_105_ top_left_grid_pin_43_ chany_top_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A mux_right_track_2.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_036_ _036_/HI _036_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_0_ chany_top_in[10] chany_top_in[3] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_1.mux_l2_in_2__A1 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A mux_left_track_17.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_18.mux_l2_in_0__S mux_top_track_18.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A mux_top_track_14.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_6.mux_l1_in_2__A0 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l3_in_0_/X _098_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_38_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l3_in_1__A1 mux_left_track_1.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l1_in_0_ chany_top_in[11] chany_top_in[4] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_0_ chany_top_in[13] chany_top_in[6] mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X _117_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_8.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l2_in_1__A0 mux_top_track_6.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l4_in_0__A1 mux_left_track_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_0.mux_l2_in_3_/S mux_top_track_0.mux_l3_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 top_left_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_3__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l1_in_1_ top_left_grid_pin_49_ top_left_grid_pin_47_ mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_1_ right_bottom_grid_pin_5_ chany_top_in[18] mux_right_track_24.mux_l1_in_2_/S
+ mux_right_track_24.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_6.mux_l3_in_0__A0 mux_top_track_6.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_3__A0 _051_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_052_ _052_/HI _052_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l2_in_1_/S clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__S mux_left_track_5.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_2__S mux_top_track_4.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_035_ _035_/HI _035_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_104_ chanx_left_in[19] chany_top_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_34_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0__S mux_top_track_8.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_2__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A0 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A mux_right_track_8.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l2_in_1__A1 mux_top_track_6.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l1_in_1__A0 _034_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A0 mux_left_track_5.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_22.mux_l1_in_0__S mux_top_track_22.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_3.mux_l2_in_0_/S mux_left_track_3.mux_l3_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_2.mux_l2_in_2__S mux_right_track_2.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_3__S mux_left_track_5.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__S mux_left_track_3.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_0.mux_l1_in_0_/S mux_top_track_0.mux_l2_in_3_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_8.mux_l1_in_3__S mux_right_track_8.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D mux_left_track_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l2_in_1__S mux_left_track_9.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_45_ top_left_grid_pin_43_ mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l1_in_0_ chany_top_in[11] chany_top_in[4] mux_right_track_24.mux_l1_in_2_/S
+ mux_right_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_18.mux_l2_in_0__A0 mux_top_track_18.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l3_in_0__A1 mux_top_track_6.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A0 mux_left_track_5.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_3__A1 chanx_left_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_051_ _051_/HI _051_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_24.mux_l3_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_034_ _034_/HI _034_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_103_ chanx_left_in[15] chany_top_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_6.mux_l2_in_0_/S mux_top_track_6.mux_l3_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l1_in_1__S mux_right_track_24.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0__S mux_top_track_14.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__D mux_left_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_0.mux_l2_in_1_/S mux_right_track_0.mux_l3_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A1 mux_left_track_5.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l1_in_1__A1 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__101__A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_3.mux_l1_in_0_/S mux_left_track_3.mux_l2_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_top_track_0.mux_l1_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_3_ _048_/HI left_bottom_grid_pin_11_ mux_left_track_5.mux_l2_in_1_/S
+ mux_left_track_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_18.mux_l2_in_0__A1 mux_top_track_18.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A1 mux_left_track_5.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_050_ _050_/HI _050_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_9.mux_l2_in_0_/S mux_left_track_9.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_28_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 mux_right_track_0.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1__S mux_left_track_17.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_033_ _033_/HI _033_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_102_ chanx_left_in[11] chany_top_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_6.mux_l1_in_0_/S mux_top_track_6.mux_l2_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_16.mux_l2_in_1__S mux_right_track_16.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S mux_left_track_5.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__104__A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_22.mux_l1_in_0_/S mux_top_track_22.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0__S mux_top_track_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A1 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_0.mux_l1_in_1_/S mux_right_track_0.mux_l2_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_1.mux_l4_in_0_/S mux_left_track_3.mux_l1_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_17.mux_l1_in_3__A0 _044_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1__A0 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_2__A1 right_bottom_grid_pin_9_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__112__A _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_2_ left_bottom_grid_pin_9_ left_bottom_grid_pin_7_ mux_left_track_5.mux_l2_in_1_/S
+ mux_left_track_5.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_3__S mux_right_track_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__107__A _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l2_in_1__S mux_left_track_5.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 mux_left_track_9.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 mux_right_track_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_1__S mux_right_track_8.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_101_ chanx_left_in[7] chany_top_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_032_ _032_/HI _032_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_4.mux_l3_in_0_/S mux_top_track_6.mux_l1_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_3_ left_bottom_grid_pin_5_ left_bottom_grid_pin_3_ mux_left_track_5.mux_l1_in_1_/S
+ mux_left_track_5.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_38.sky130_fd_sc_hd__buf_4_0__A mux_top_track_38.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_20.mux_l2_in_0_/S mux_top_track_22.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l3_in_0_/X _070_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_28_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__115__A _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_38.mux_l2_in_0_/S mux_right_track_0.mux_l1_in_1_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_10.mux_l2_in_0__S mux_top_track_10.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_5.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l1_in_3__A1 left_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_16.mux_l1_in_1__S mux_top_track_16.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_9.mux_l1_in_1__A1 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l3_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_5.mux_l4_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_9.mux_l2_in_0__A1 mux_left_track_9.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_100_ chanx_left_in[3] chany_top_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_031_ _031_/HI _031_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_19_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__118__A _118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_2_ left_bottom_grid_pin_1_ chanx_right_in[14] mux_left_track_5.mux_l1_in_1_/S
+ mux_left_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_18.mux_l2_in_0_ mux_top_track_18.mux_l1_in_1_/X mux_top_track_18.mux_l1_in_0_/X
+ mux_top_track_18.mux_l2_in_0_/S mux_top_track_18.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l1_in_2__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_33.mux_l2_in_0_/S ccff_tail
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_20.mux_l2_in_0_ mux_top_track_20.mux_l1_in_1_/X mux_top_track_20.mux_l1_in_0_/X
+ mux_top_track_20.mux_l2_in_0_/S mux_top_track_20.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 mux_right_track_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_18.mux_l1_in_1_ _034_/HI chanx_left_in[14] mux_top_track_18.mux_l1_in_1_/S
+ mux_top_track_18.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S mux_left_track_25.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_20.mux_l1_in_1_ _036_/HI chanx_left_in[16] mux_top_track_20.mux_l1_in_0_/S
+ mux_top_track_20.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_38.mux_l1_in_0__A0 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_2__A0 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_1__S mux_top_track_6.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_24.mux_l1_in_2_/S
+ mux_right_track_24.mux_l2_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l2_in_1_ _045_/HI mux_left_track_25.mux_l1_in_2_/X mux_left_track_25.mux_l2_in_0_/S
+ mux_left_track_25.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_2.mux_l3_in_1__A0 mux_right_track_2.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_030_ _030_/HI _030_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_22_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_1_ chanx_right_in[5] chany_top_in[19] mux_left_track_5.mux_l1_in_1_/S
+ mux_left_track_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_2_ left_bottom_grid_pin_5_ chanx_right_in[18] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_0.mux_l1_in_3__S mux_right_track_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_1__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_20.sky130_fd_sc_hd__buf_4_0_ mux_top_track_20.mux_l2_in_0_/X _108_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_33.mux_l1_in_0_/S mux_left_track_33.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_2.mux_l4_in_0__A0 mux_right_track_2.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_3__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_14.sky130_fd_sc_hd__buf_4_0_ mux_top_track_14.mux_l2_in_0_/X _111_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_0.mux_l2_in_0__A0 top_left_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_18.mux_l1_in_0_ chanx_right_in[14] top_left_grid_pin_47_ mux_top_track_18.mux_l1_in_1_/S
+ mux_top_track_18.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_20.mux_l1_in_0_ chanx_right_in[16] top_left_grid_pin_48_ mux_top_track_20.mux_l1_in_0_/S
+ mux_top_track_20.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_38.mux_l1_in_0__A1 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_2__A1 right_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_0__S mux_left_track_33.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_16.mux_l3_in_0_/S
+ mux_right_track_24.mux_l1_in_2_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_32.mux_l2_in_0__S mux_right_track_32.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l3_in_1__A1 mux_right_track_2.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_12.mux_l1_in_1__S mux_top_track_12.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A mux_left_track_5.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_0_ chany_top_in[12] chany_top_in[5] mux_left_track_5.mux_l1_in_1_/S
+ mux_left_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_1_ chanx_right_in[9] chany_top_in[16] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_089_ chanx_left_in[8] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S mux_top_track_8.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__060__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_25.mux_l3_in_0_/S mux_left_track_33.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l4_in_0__A1 mux_right_track_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S mux_right_track_32.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_10.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l2_in_1_ _042_/HI chanx_left_in[8] mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_0.mux_l2_in_0__A1 mux_top_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0__A0 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l2_in_0__S mux_left_track_25.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_32.mux_l2_in_1_ _054_/HI chanx_left_in[10] mux_right_track_32.mux_l2_in_1_/S
+ mux_right_track_32.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l3_in_0__S mux_right_track_24.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A mux_top_track_24.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__063__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l1_in_1__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_10.mux_l2_in_1__A0 _030_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_25.mux_l1_in_0_ chany_top_in[9] chany_top_in[2] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_088_ chanx_left_in[9] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_14.mux_l1_in_0_/S mux_top_track_14.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_10.mux_l3_in_0__A0 mux_top_track_10.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_20.mux_l1_in_0__A0 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__A0 _055_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__071__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l3_in_0__S mux_left_track_17.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_6_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l2_in_0_ chanx_right_in[15] mux_top_track_8.mux_l1_in_0_/X mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0__A1 top_left_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_2__S mux_left_track_3.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__066__A _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_1_/S mux_right_track_32.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l3_in_1__S mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 top_left_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l3_in_0_/X _114_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l1_in_1_ right_bottom_grid_pin_7_ chany_top_in[19] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A mux_top_track_4.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_10.mux_l2_in_1__A1 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__074__A _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_087_ chanx_left_in[10] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A0 mux_top_track_2.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_20.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__069__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_12.mux_l2_in_0_/S mux_top_track_14.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_10.mux_l3_in_0__A1 mux_top_track_10.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l2_in_0__S mux_top_track_24.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X _086_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_30_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_20.mux_l1_in_0__A1 top_left_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l4_in_0__S mux_left_track_5.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__A1 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_3__A0 _029_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_18.mux_l1_in_0__S mux_top_track_18.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l3_in_0__A0 mux_top_track_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l2_in_3_ _043_/HI left_bottom_grid_pin_9_ mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__082__A _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_41_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_16.mux_l2_in_0_/S
+ mux_right_track_16.mux_l3_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__077__A _077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[8] top_left_grid_pin_42_ mux_top_track_8.mux_l1_in_0_/S
+ mux_top_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l2_in_1__S mux_left_track_33.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__D mux_left_track_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l1_in_0_ chany_top_in[12] chany_top_in[5] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l1_in_2__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S mux_left_track_1.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__090__A _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_086_ _086_/A chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 mux_top_track_2.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_1__A0 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_14.mux_l1_in_1__A0 _032_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l3_in_0_/X _077_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__085__A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_069_ chanx_right_in[8] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l2_in_3__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0__S mux_top_track_8.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0__A0 mux_top_track_14.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l3_in_0__A1 mux_top_track_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A0 mux_left_track_1.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_3__A0 _028_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_2_ left_bottom_grid_pin_5_ left_bottom_grid_pin_1_ mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l2_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__093__A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_3.mux_l2_in_0__S mux_left_track_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l2_in_3_ _052_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_2_/S
+ mux_right_track_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__088__A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_22.mux_l1_in_1__A0 _037_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1__S mux_left_track_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_32.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l3_in_0__S mux_top_track_6.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_25.mux_l1_in_0_/S mux_left_track_25.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_085_ chanx_left_in[12] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l1_in_1__A1 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_22.mux_l2_in_0__A0 mux_top_track_22.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_38.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A mux_top_track_10.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S mux_right_track_2.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_068_ chanx_right_in[9] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_6.mux_l1_in_1__A0 top_left_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__096__A _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l2_in_0__A1 mux_top_track_14.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A1 mux_left_track_1.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_20.mux_l2_in_0__S mux_top_track_20.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_3__A1 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ chanx_right_in[12] chanx_right_in[2] mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_4.mux_l1_in_3__A0 _040_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l4_in_0__S mux_left_track_1.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_6.mux_l2_in_0__A0 mux_top_track_6.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0__S mux_top_track_14.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_16.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l4_in_0__S mux_right_track_4.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_8.mux_l3_in_0_/S mux_right_track_16.mux_l1_in_3_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__D mux_left_track_1.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_2_ chanx_left_in[4] right_bottom_grid_pin_11_ mux_right_track_2.mux_l2_in_2_/S
+ mux_right_track_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_14.mux_l2_in_0_ mux_top_track_14.mux_l1_in_1_/X mux_top_track_14.mux_l1_in_0_/X
+ mux_top_track_14.mux_l2_in_0_/S mux_top_track_14.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_22.mux_l1_in_1__A1 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__099__A _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_24.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_17.mux_l3_in_0_/S mux_left_track_25.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_084_ chanx_left_in[13] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.mux_l2_in_1__A0 mux_right_track_16.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_14.mux_l1_in_1_ _032_/HI chanx_left_in[12] mux_top_track_14.mux_l1_in_0_/S
+ mux_top_track_14.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_22.mux_l2_in_0__A1 mux_top_track_22.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_38.mux_l1_in_0_/S mux_top_track_38.mux_l2_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_067_ chanx_right_in[10] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_16.mux_l1_in_1__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_1__A1 top_left_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l3_in_0__A0 mux_right_track_16.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l2_in_0_ chany_top_in[14] mux_left_track_1.mux_l1_in_0_/X mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_3__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A mux_right_track_4.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_3__A0 _046_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_6.mux_l2_in_0__A1 mux_top_track_6.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l1_in_0__A0 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A0 mux_left_track_5.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A mux_top_track_16.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_41_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ right_bottom_grid_pin_7_ right_bottom_grid_pin_3_
+ mux_right_track_2.mux_l2_in_2_/S mux_right_track_2.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2__A1 right_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l2_in_1__A0 _053_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_10.sky130_fd_sc_hd__buf_4_0_ mux_top_track_10.mux_l3_in_0_/X _113_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_083_ chanx_left_in[14] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l3_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A1 mux_right_track_16.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__S mux_left_track_5.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_14.mux_l1_in_0_ chanx_right_in[12] top_left_grid_pin_45_ mux_top_track_14.mux_l1_in_0_/S
+ mux_top_track_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l3_in_0__A0 mux_right_track_24.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1__S mux_right_track_8.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_3__S mux_top_track_4.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l3_in_0__S mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_24.mux_l2_in_0_/S mux_top_track_38.mux_l1_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_066_ _066_/A chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_8.mux_l2_in_1__S mux_top_track_8.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l3_in_0__A1 mux_right_track_16.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l1_in_3_ _040_/HI chanx_left_in[5] mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_118_ _118_/A chany_top_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_049_ _049_/HI _049_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l1_in_3__A1 left_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail mux_left_track_33.mux_l3_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_18.mux_l1_in_0__A1 top_left_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_5.mux_l2_in_0__A1 mux_left_track_5.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_24.mux_l1_in_2__A1 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_32.mux_l2_in_1__A0 _054_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 right_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l1_in_0_ chany_top_in[7] chany_top_in[0] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_22.mux_l1_in_1__S mux_top_track_22.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_3__S mux_right_track_2.mux_l2_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_10.mux_l1_in_0__S mux_top_track_10.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l2_in_0_ chany_top_in[14] mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_2_/S mux_right_track_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l2_in_1_ _047_/HI left_bottom_grid_pin_7_ mux_left_track_33.mux_l2_in_0_/S
+ mux_left_track_33.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_38.mux_l2_in_0__S mux_top_track_38.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l4_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_24.mux_l2_in_1__A1 mux_right_track_24.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l3_in_0__A0 mux_right_track_32.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 mux_right_track_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l3_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_082_ _082_/A chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_37_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_2.mux_l1_in_1_/S mux_top_track_2.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l1_in_3_/X mux_top_track_4.mux_l1_in_2_/X
+ mux_top_track_4.mux_l2_in_0_/S mux_top_track_4.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l3_in_0__A1 mux_right_track_24.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l2_in_1__A0 _042_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_065_ chanx_right_in[12] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_4.mux_l1_in_2_ chanx_right_in[7] chanx_right_in[5] mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_117_ _117_/A chany_top_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_048_ _048_/HI _048_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_24.mux_l1_in_2__S mux_right_track_24.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l3_in_0__A0 mux_top_track_8.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_8.mux_l2_in_1_/S mux_top_track_8.mux_l3_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_38.mux_l2_in_0_ _039_/HI mux_top_track_38.mux_l1_in_0_/X mux_top_track_38.mux_l2_in_0_/S
+ mux_top_track_38.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_17.mux_l1_in_2__A0 left_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l2_in_1__A1 chanx_left_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__102__A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__S mux_top_track_0.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_0_/S mux_left_track_33.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_2.mux_l2_in_2_/S mux_right_track_2.mux_l3_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_17.mux_l2_in_1__A0 mux_left_track_17.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_32.mux_l3_in_0__A1 mux_right_track_32.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l4_in_0_/X _097_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_5.mux_l1_in_1_/S mux_left_track_5.mux_l2_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_081_ chanx_left_in[16] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_6.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_2_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_2.mux_l1_in_0_ chany_top_in[7] chany_top_in[0] mux_right_track_2.mux_l1_in_0_/S
+ mux_right_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_0.mux_l4_in_0_/S mux_top_track_2.mux_l1_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_33.mux_l1_in_1_ chanx_right_in[10] chany_top_in[15] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_0_/S mux_top_track_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l3_in_0__A0 mux_left_track_17.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2__S mux_left_track_17.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X _116_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_8.mux_l2_in_1__A1 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_064_ chanx_right_in[13] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__110__A _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_4.mux_l1_in_1_ top_left_grid_pin_48_ top_left_grid_pin_46_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_116_ _116_/A chany_top_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_4.mux_l1_in_1__S mux_right_track_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_3__A0 _048_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__105__A top_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_047_ _047_/HI _047_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_25.mux_l1_in_2__A0 left_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l3_in_0__A1 mux_top_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_8.mux_l1_in_0_/S mux_top_track_8.mux_l2_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l2_in_1__S mux_top_track_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2__A1 chanx_right_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_24.mux_l1_in_1_/S mux_top_track_24.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_3_7_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l2_in_1__A0 _045_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_25.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_38.mux_l1_in_0_ chanx_left_in[1] chanx_right_in[0] mux_top_track_38.mux_l1_in_0_/S
+ mux_top_track_38.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_2.mux_l1_in_0_/S mux_right_track_2.mux_l2_in_2_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__113__A _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A1 mux_left_track_17.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_17.mux_l1_in_0_/S mux_left_track_17.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_32.mux_l1_in_0__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A0 mux_left_track_25.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_3.mux_l3_in_0_/S mux_left_track_5.mux_l1_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_080_ chanx_left_in[17] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l1_in_0_ chany_top_in[8] chany_top_in[1] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__108__A _108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l3_in_1__S mux_right_track_2.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_5.mux_l2_in_2__S mux_left_track_5.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l3_in_0__A1 mux_left_track_17.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_063_ chanx_right_in[14] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l3_in_0__S mux_left_track_9.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_8.mux_l2_in_1_/S mux_right_track_8.mux_l3_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__D mux_left_track_9.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_44_ top_left_grid_pin_42_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_115_ _115_/A chany_top_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_5.mux_l2_in_3__A1 left_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_046_ _046_/HI _046_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_2__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_6.mux_l3_in_0_/S mux_top_track_8.mux_l1_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l2_in_1__A0 _047_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__116__A _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_029_ _029_/HI _029_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 right_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_8.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_0__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l2_in_1__A1 mux_left_track_25.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_22.mux_l2_in_0_/S mux_top_track_24.mux_l1_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l3_in_0__A0 mux_left_track_33.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_10.mux_l2_in_1__S mux_top_track_10.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

