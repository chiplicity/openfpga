* NGSPICE file created from sb_0__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

.subckt sb_0__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4]
+ chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_out[0]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] data_in enable right_bottom_grid_pin_11_ right_bottom_grid_pin_13_
+ right_bottom_grid_pin_15_ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_
+ right_bottom_grid_pin_7_ right_bottom_grid_pin_9_ right_top_grid_pin_10_ top_left_grid_pin_11_
+ top_left_grid_pin_13_ top_left_grid_pin_15_ top_left_grid_pin_1_ top_left_grid_pin_3_
+ top_left_grid_pin_5_ top_left_grid_pin_7_ top_left_grid_pin_9_ top_right_grid_pin_11_
+ vpwr vgnd
Xmem_right_track_12.LATCH_1_.latch data_in _115_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_199 vgnd vpwr scs8hd_decap_12
XFILLER_7_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_144 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_9_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_181 vgnd vpwr scs8hd_decap_3
XFILLER_27_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _115_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__124__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ _200_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__209__A _209_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_20 vpwr vgnd scs8hd_fill_2
X_131_ _131_/A _131_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_42 vgnd vpwr scs8hd_decap_4
XFILLER_23_97 vpwr vgnd scs8hd_fill_2
XFILLER_2_154 vgnd vpwr scs8hd_decap_3
XFILLER_2_121 vpwr vgnd scs8hd_fill_2
XFILLER_9_33 vgnd vpwr scs8hd_decap_4
XFILLER_9_77 vgnd vpwr scs8hd_decap_4
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_64 vpwr vgnd scs8hd_fill_2
XFILLER_7_202 vgnd vpwr scs8hd_decap_3
XFILLER_7_224 vgnd vpwr scs8hd_decap_8
X_114_ _114_/A _114_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__121__B address[5] vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _182_/HI _119_/Y mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _187_/HI _086_/Y mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_45 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _146_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_4
Xmem_right_track_8.LATCH_1_.latch data_in _111_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_164 vgnd vpwr scs8hd_decap_12
XFILLER_31_31 vgnd vpwr scs8hd_decap_12
XFILLER_15_87 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _110_/A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_16_120 vgnd vpwr scs8hd_decap_3
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _114_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_134 vgnd vpwr scs8hd_decap_8
XFILLER_22_145 vgnd vpwr scs8hd_decap_4
Xmem_top_track_4.LATCH_0_.latch data_in _090_/A _132_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_101 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_6
XFILLER_9_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_119 vgnd vpwr scs8hd_decap_4
XFILLER_12_99 vgnd vpwr scs8hd_fill_1
XFILLER_33_218 vgnd vpwr scs8hd_decap_4
XFILLER_33_229 vgnd vpwr scs8hd_decap_4
XFILLER_5_174 vgnd vpwr scs8hd_decap_6
XANTENNA__124__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_6.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_7_ mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_15_229 vgnd vpwr scs8hd_decap_4
X_130_ address[3] _155_/B _139_/C _155_/D _131_/B vgnd vpwr scs8hd_or4_4
XFILLER_2_144 vgnd vpwr scs8hd_decap_8
XFILLER_2_133 vgnd vpwr scs8hd_decap_8
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_43 vpwr vgnd scs8hd_fill_2
X_113_ _113_/A _113_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_232 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _116_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_6.tap_buf4_0_.scs8hd_inv_1 mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _210_/A vgnd vpwr scs8hd_inv_1
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _118_/A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_118 vgnd vpwr scs8hd_decap_4
XFILLER_4_206 vgnd vpwr scs8hd_decap_8
XFILLER_20_22 vgnd vpwr scs8hd_decap_4
XFILLER_20_88 vgnd vpwr scs8hd_decap_4
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XFILLER_28_151 vpwr vgnd scs8hd_fill_2
XFILLER_6_24 vgnd vpwr scs8hd_fill_1
XFILLER_6_68 vgnd vpwr scs8hd_decap_3
XANTENNA__132__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_121 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_140 vgnd vpwr scs8hd_fill_1
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _102_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_176 vgnd vpwr scs8hd_decap_6
XFILLER_15_22 vpwr vgnd scs8hd_fill_2
XFILLER_31_43 vgnd vpwr scs8hd_decap_12
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_146 vpwr vgnd scs8hd_fill_2
XFILLER_31_135 vgnd vpwr scs8hd_decap_6
XFILLER_31_113 vpwr vgnd scs8hd_fill_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_102 vgnd vpwr scs8hd_decap_8
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _105_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _088_/Y mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_26_54 vgnd vpwr scs8hd_decap_8
XFILLER_3_69 vgnd vpwr scs8hd_decap_8
XANTENNA__138__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_33_208 vgnd vpwr scs8hd_decap_3
XFILLER_5_142 vpwr vgnd scs8hd_fill_2
XANTENNA__140__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XANTENNA__135__B _134_/B vgnd vpwr scs8hd_diode_2
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__151__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _088_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_88 vpwr vgnd scs8hd_fill_2
X_112_ _112_/A _112_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_222 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_5_ mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _107_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_10 vpwr vgnd scs8hd_fill_2
XFILLER_20_67 vgnd vpwr scs8hd_decap_4
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _105_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_87 vgnd vpwr scs8hd_decap_12
XFILLER_29_65 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_34_133 vgnd vpwr scs8hd_decap_12
XFILLER_19_196 vgnd vpwr scs8hd_decap_8
XFILLER_31_55 vgnd vpwr scs8hd_decap_6
XFILLER_0_221 vpwr vgnd scs8hd_fill_2
XFILLER_16_100 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _139_/C vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _143_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.LATCH_1_.latch data_in _107_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_66 vgnd vpwr scs8hd_decap_3
XFILLER_26_44 vgnd vpwr scs8hd_fill_1
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _185_/HI _109_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_26 vpwr vgnd scs8hd_fill_2
XANTENNA__138__B _137_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_151 vpwr vgnd scs8hd_fill_2
XFILLER_8_162 vpwr vgnd scs8hd_fill_2
XFILLER_8_173 vgnd vpwr scs8hd_decap_8
XANTENNA__154__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _090_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_217 vgnd vpwr scs8hd_decap_12
XFILLER_10_139 vgnd vpwr scs8hd_fill_1
XFILLER_5_7 vgnd vpwr scs8hd_fill_1
XFILLER_12_46 vpwr vgnd scs8hd_fill_2
XFILLER_12_57 vgnd vpwr scs8hd_decap_8
XFILLER_12_68 vgnd vpwr scs8hd_decap_4
XFILLER_18_206 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _195_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_198 vgnd vpwr scs8hd_decap_6
Xmem_top_track_0.LATCH_0_.latch data_in _085_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_23_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_179 vgnd vpwr scs8hd_decap_12
XFILLER_2_168 vpwr vgnd scs8hd_fill_2
XFILLER_0_38 vgnd vpwr scs8hd_decap_4
XFILLER_9_14 vpwr vgnd scs8hd_fill_2
XFILLER_9_69 vpwr vgnd scs8hd_fill_2
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__151__B _151_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_190 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _113_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_212 vpwr vgnd scs8hd_fill_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
X_111_ _111_/A _111_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__146__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_46 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _186_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_48 vpwr vgnd scs8hd_fill_2
XFILLER_6_59 vgnd vpwr scs8hd_decap_3
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XFILLER_34_145 vgnd vpwr scs8hd_decap_8
XANTENNA__157__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_3_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _181_/HI _117_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_123 vgnd vpwr scs8hd_fill_1
XFILLER_15_35 vpwr vgnd scs8hd_fill_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_68 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_145 vgnd vpwr scs8hd_decap_8
XFILLER_16_189 vgnd vpwr scs8hd_decap_12
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__D _139_/D vgnd vpwr scs8hd_diode_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_80 vgnd vpwr scs8hd_decap_3
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_13_159 vpwr vgnd scs8hd_fill_2
XFILLER_3_16 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _108_/A mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__154__B _154_/B vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_229 vgnd vpwr scs8hd_decap_4
XFILLER_10_107 vgnd vpwr scs8hd_decap_12
XFILLER_12_36 vpwr vgnd scs8hd_fill_2
XANTENNA__080__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA__149__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_232 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_24 vgnd vpwr scs8hd_decap_3
XFILLER_23_46 vgnd vpwr scs8hd_fill_1
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_2_125 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_37 vgnd vpwr scs8hd_fill_1
XFILLER_14_232 vgnd vpwr scs8hd_fill_1
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _112_/Y mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _110_/A _110_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _113_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__162__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_14 vpwr vgnd scs8hd_fill_2
XFILLER_28_143 vgnd vpwr scs8hd_decap_8
XFILLER_6_16 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XFILLER_19_132 vpwr vgnd scs8hd_fill_2
XFILLER_19_154 vpwr vgnd scs8hd_fill_2
XANTENNA__157__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA__173__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_25_135 vpwr vgnd scs8hd_fill_2
XANTENNA__083__A enable vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _116_/A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_212 vgnd vpwr scs8hd_decap_4
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_190 vgnd vpwr scs8hd_decap_12
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _131_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_1_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_8_186 vpwr vgnd scs8hd_fill_2
XANTENNA__170__B _155_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_230 vgnd vpwr scs8hd_decap_3
XFILLER_10_119 vgnd vpwr scs8hd_decap_4
XFILLER_26_230 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_7_ mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_0.LATCH_1_.latch data_in _103_/A _153_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_123 vpwr vgnd scs8hd_fill_2
XFILLER_5_101 vpwr vgnd scs8hd_fill_2
Xmem_top_track_8.LATCH_1_.latch data_in _093_/A _137_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _120_/Y mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _115_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _085_/Y mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__149__C _155_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_60 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_104 vpwr vgnd scs8hd_fill_2
X_186_ _186_/HI _186_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _108_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_170 vgnd vpwr scs8hd_decap_12
XANTENNA__176__A _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _101_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_14 vgnd vpwr scs8hd_decap_3
XFILLER_18_47 vpwr vgnd scs8hd_fill_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_7_207 vpwr vgnd scs8hd_fill_2
XFILLER_11_214 vgnd vpwr scs8hd_fill_1
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
X_169_ address[0] _167_/X _169_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_26 vgnd vpwr scs8hd_fill_1
XFILLER_29_57 vgnd vpwr scs8hd_decap_4
XFILLER_28_133 vgnd vpwr scs8hd_fill_1
XFILLER_3_221 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__173__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_25_103 vpwr vgnd scs8hd_fill_2
XFILLER_31_117 vgnd vpwr scs8hd_decap_4
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vgnd vpwr scs8hd_decap_3
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _103_/A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_150 vgnd vpwr scs8hd_decap_3
XFILLER_15_180 vgnd vpwr scs8hd_decap_3
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_14.LATCH_0_.latch data_in _100_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_154 vgnd vpwr scs8hd_decap_8
XFILLER_12_150 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _110_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__170__C _155_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _087_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _198_/A vgnd vpwr scs8hd_inv_1
XANTENNA__089__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_146 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _206_/A vgnd vpwr scs8hd_inv_1
XANTENNA__149__D _155_/D vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _184_/HI _107_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_83 vgnd vpwr scs8hd_decap_3
X_185_ _185_/HI _185_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_5_ mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_6 vpwr vgnd scs8hd_fill_2
XFILLER_1_182 vgnd vpwr scs8hd_fill_1
XANTENNA__176__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_204 vgnd vpwr scs8hd_decap_8
XFILLER_11_226 vgnd vpwr scs8hd_decap_6
XFILLER_6_230 vgnd vpwr scs8hd_decap_3
X_168_ _131_/A _167_/X _168_/Y vgnd vpwr scs8hd_nor2_4
X_099_ _099_/A _099_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_73 vgnd vpwr scs8hd_decap_4
XFILLER_29_69 vpwr vgnd scs8hd_fill_2
XFILLER_29_14 vgnd vpwr scs8hd_decap_12
XFILLER_28_123 vgnd vpwr scs8hd_decap_8
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_200 vgnd vpwr scs8hd_fill_1
XFILLER_10_82 vgnd vpwr scs8hd_fill_1
XFILLER_13_9 vpwr vgnd scs8hd_fill_2
XFILLER_19_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _089_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__173__C address[4] vgnd vpwr scs8hd_diode_2
XFILLER_25_115 vgnd vpwr scs8hd_fill_1
XFILLER_0_225 vgnd vpwr scs8hd_decap_8
XFILLER_16_104 vgnd vpwr scs8hd_decap_3
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_7_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _201_/A vgnd vpwr scs8hd_inv_1
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_21_162 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _180_/HI _115_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XFILLER_16_70 vpwr vgnd scs8hd_fill_2
XFILLER_12_140 vpwr vgnd scs8hd_fill_2
XFILLER_12_184 vpwr vgnd scs8hd_fill_2
XFILLER_8_199 vgnd vpwr scs8hd_decap_12
XANTENNA__170__D _139_/D vgnd vpwr scs8hd_diode_2
XFILLER_12_17 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_158 vgnd vpwr scs8hd_fill_1
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_210 vgnd vpwr scs8hd_decap_3
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_27_91 vgnd vpwr scs8hd_fill_1
XFILLER_17_232 vgnd vpwr scs8hd_fill_1
XFILLER_4_73 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _106_/A mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_23_16 vpwr vgnd scs8hd_fill_2
XFILLER_23_49 vgnd vpwr scs8hd_decap_6
XFILLER_9_18 vpwr vgnd scs8hd_fill_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
XFILLER_14_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_184_ _184_/HI _184_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_194 vgnd vpwr scs8hd_decap_12
Xmem_top_track_4.LATCH_1_.latch data_in _089_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__176__C _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vpwr vgnd scs8hd_fill_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_167_ _139_/A _155_/B _155_/C _155_/D _167_/X vgnd vpwr scs8hd_or4_4
X_098_ _098_/A _098_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_3_ mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_26 vgnd vpwr scs8hd_decap_12
XFILLER_28_157 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _110_/Y mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_212 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_61 vpwr vgnd scs8hd_fill_2
XFILLER_34_105 vgnd vpwr scs8hd_fill_1
XFILLER_19_179 vgnd vpwr scs8hd_decap_4
XANTENNA__173__D _148_/B vgnd vpwr scs8hd_diode_2
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_39 vgnd vpwr scs8hd_decap_3
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_116 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_60 vgnd vpwr scs8hd_fill_1
XFILLER_21_71 vgnd vpwr scs8hd_decap_12
XFILLER_11_7 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_160 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vgnd vpwr scs8hd_fill_1
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _116_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
XFILLER_32_81 vgnd vpwr scs8hd_decap_8
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _114_/A mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_35_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_70 vpwr vgnd scs8hd_fill_2
XFILLER_17_222 vpwr vgnd scs8hd_fill_2
Xmem_top_track_10.LATCH_0_.latch data_in _096_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _212_/A vgnd vpwr scs8hd_inv_1
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_184 vgnd vpwr scs8hd_decap_3
XFILLER_1_140 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _118_/Y mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_6 vpwr vgnd scs8hd_fill_2
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
X_166_ address[0] _164_/X _166_/Y vgnd vpwr scs8hd_nor2_4
X_097_ _097_/A _097_/Y vgnd vpwr scs8hd_inv_8
XFILLER_20_18 vpwr vgnd scs8hd_fill_2
XFILLER_20_29 vpwr vgnd scs8hd_fill_2
XFILLER_29_38 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _118_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_169 vgnd vpwr scs8hd_decap_12
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_136 vgnd vpwr scs8hd_decap_4
XFILLER_27_180 vgnd vpwr scs8hd_decap_3
XFILLER_19_158 vgnd vpwr scs8hd_decap_6
X_149_ address[3] address[2] _155_/C _155_/D _151_/B vgnd vpwr scs8hd_or4_4
XFILLER_25_139 vpwr vgnd scs8hd_fill_2
XFILLER_15_18 vpwr vgnd scs8hd_fill_2
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_1_ mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_83 vgnd vpwr scs8hd_fill_1
XFILLER_30_142 vgnd vpwr scs8hd_decap_8
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_172 vpwr vgnd scs8hd_fill_2
XFILLER_21_175 vgnd vpwr scs8hd_decap_8
XFILLER_8_102 vgnd vpwr scs8hd_decap_3
XFILLER_12_120 vgnd vpwr scs8hd_decap_8
XFILLER_16_61 vgnd vpwr scs8hd_decap_3
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _107_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_7_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_190 vpwr vgnd scs8hd_fill_2
XFILLER_5_127 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_29 vpwr vgnd scs8hd_fill_2
XFILLER_2_108 vgnd vpwr scs8hd_decap_4
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_73 vgnd vpwr scs8hd_decap_4
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_218 vgnd vpwr scs8hd_decap_12
XFILLER_11_218 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _183_/HI _105_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _090_/Y vgnd vpwr
+ scs8hd_diode_2
X_165_ _131_/A _164_/X _165_/Y vgnd vpwr scs8hd_nor2_4
X_096_ _096_/A _096_/Y vgnd vpwr scs8hd_inv_8
XFILLER_27_6 vpwr vgnd scs8hd_fill_2
XFILLER_1_10 vpwr vgnd scs8hd_fill_2
XFILLER_1_21 vgnd vpwr scs8hd_decap_8
XFILLER_1_43 vpwr vgnd scs8hd_fill_2
XFILLER_1_98 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_1_.latch data_in _086_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_85 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _109_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_83 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_148_ address[4] _148_/B _155_/C vgnd vpwr scs8hd_nand2_4
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_25_107 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_33_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_40 vpwr vgnd scs8hd_fill_2
XFILLER_21_95 vpwr vgnd scs8hd_fill_2
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XFILLER_7_42 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _096_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_125 vpwr vgnd scs8hd_fill_2
XFILLER_12_154 vgnd vpwr scs8hd_decap_3
XFILLER_12_176 vgnd vpwr scs8hd_decap_8
XFILLER_16_84 vgnd vpwr scs8hd_decap_6
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_26_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _092_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_6
XFILLER_27_94 vpwr vgnd scs8hd_fill_2
XFILLER_27_83 vpwr vgnd scs8hd_fill_2
XFILLER_17_202 vgnd vpwr scs8hd_decap_8
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _179_/HI _113_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_43 vgnd vpwr scs8hd_decap_8
XFILLER_4_21 vgnd vpwr scs8hd_decap_8
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_30 vpwr vgnd scs8hd_fill_2
Xmem_right_track_14.LATCH_0_.latch data_in _118_/A _175_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_153 vpwr vgnd scs8hd_fill_2
XFILLER_9_231 vpwr vgnd scs8hd_fill_2
XFILLER_18_19 vgnd vpwr scs8hd_decap_8
XFILLER_11_208 vgnd vpwr scs8hd_decap_6
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _104_/A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_6_201 vgnd vpwr scs8hd_decap_4
X_164_ _139_/A address[2] _155_/C _139_/D _164_/X vgnd vpwr scs8hd_or4_4
XFILLER_10_230 vgnd vpwr scs8hd_decap_3
X_095_ _095_/A _095_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_73 vgnd vpwr scs8hd_decap_8
XFILLER_24_84 vgnd vpwr scs8hd_decap_8
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_20 vgnd vpwr scs8hd_decap_3
XFILLER_10_53 vgnd vpwr scs8hd_decap_8
XFILLER_19_40 vpwr vgnd scs8hd_fill_2
XFILLER_19_73 vpwr vgnd scs8hd_fill_2
XFILLER_35_94 vgnd vpwr scs8hd_decap_12
X_147_ address[0] _147_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _179_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_3 vpwr vgnd scs8hd_fill_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XFILLER_31_19 vgnd vpwr scs8hd_decap_12
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_52 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _101_/A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_30_100 vgnd vpwr scs8hd_decap_4
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _108_/Y mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_196 vgnd vpwr scs8hd_decap_6
XFILLER_7_76 vpwr vgnd scs8hd_fill_2
XFILLER_7_98 vpwr vgnd scs8hd_fill_2
Xmux_top_track_12.INVTX1_1_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_144 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_41 vgnd vpwr scs8hd_decap_3
XFILLER_12_144 vgnd vpwr scs8hd_decap_4
XFILLER_12_188 vgnd vpwr scs8hd_decap_12
XFILLER_16_74 vgnd vpwr scs8hd_fill_1
XFILLER_16_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_151 vpwr vgnd scs8hd_fill_2
XFILLER_4_88 vgnd vpwr scs8hd_decap_4
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_53 vgnd vpwr scs8hd_decap_6
X_180_ _180_/HI _180_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XFILLER_1_143 vgnd vpwr scs8hd_decap_3
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_41 vgnd vpwr scs8hd_decap_6
X_094_ _094_/A _094_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_213 vgnd vpwr scs8hd_fill_1
X_163_ address[0] _163_/B _163_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_28_106 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _115_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _116_/Y mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__212__A _212_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_76 vgnd vpwr scs8hd_decap_6
XFILLER_34_109 vgnd vpwr scs8hd_decap_12
XANTENNA__122__A address[1] vgnd vpwr scs8hd_diode_2
X_146_ _131_/A _147_/B _146_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_6 vgnd vpwr scs8hd_decap_12
XFILLER_33_131 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_208 vpwr vgnd scs8hd_fill_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_153 vgnd vpwr scs8hd_fill_1
XFILLER_15_164 vgnd vpwr scs8hd_decap_8
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XFILLER_7_11 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
X_129_ address[0] _129_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_20 vgnd vpwr scs8hd_decap_8
XFILLER_32_30 vgnd vpwr scs8hd_fill_1
Xmux_top_track_10.INVTX1_1_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_226 vgnd vpwr scs8hd_decap_6
XANTENNA__130__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _117_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_207 vgnd vpwr scs8hd_decap_6
XFILLER_13_65 vpwr vgnd scs8hd_fill_2
XFILLER_1_166 vpwr vgnd scs8hd_fill_2
XFILLER_1_111 vpwr vgnd scs8hd_fill_2
XFILLER_8_3 vpwr vgnd scs8hd_fill_2
Xmem_top_track_14.LATCH_1_.latch data_in _099_/A _146_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _110_/Y vgnd vpwr
+ scs8hd_diode_2
X_162_ _131_/A _163_/B _162_/Y vgnd vpwr scs8hd_nor2_4
X_093_ _093_/A _093_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_79 vgnd vpwr scs8hd_decap_4
Xmem_right_track_10.LATCH_0_.latch data_in _114_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _188_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_217 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_63 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_27_140 vpwr vgnd scs8hd_fill_2
XFILLER_19_97 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _178_/HI _103_/Y mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_145_ _139_/A _155_/B _139_/C _139_/D _147_/B vgnd vpwr scs8hd_or4_4
XANTENNA__122__B _083_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_143 vgnd vpwr scs8hd_decap_12
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_173 vgnd vpwr scs8hd_decap_12
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_21 vpwr vgnd scs8hd_fill_2
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vpwr vgnd scs8hd_fill_2
XFILLER_15_176 vpwr vgnd scs8hd_fill_2
X_128_ _131_/A _129_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__133__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.tap_buf4_0_.scs8hd_inv_1 mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _208_/A vgnd vpwr scs8hd_inv_1
XFILLER_8_139 vgnd vpwr scs8hd_decap_12
XFILLER_12_168 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_161 vgnd vpwr scs8hd_decap_3
XFILLER_7_194 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _112_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _089_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XFILLER_4_186 vgnd vpwr scs8hd_decap_12
XFILLER_4_68 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__130__B _155_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_22 vpwr vgnd scs8hd_fill_2
XFILLER_13_88 vgnd vpwr scs8hd_decap_3
XFILLER_9_201 vgnd vpwr scs8hd_decap_3
Xmem_right_track_6.LATCH_0_.latch data_in _110_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A address[0] vgnd vpwr scs8hd_diode_2
X_161_ _139_/A address[2] _155_/C _155_/D _163_/B vgnd vpwr scs8hd_or4_4
XFILLER_24_10 vgnd vpwr scs8hd_decap_4
XFILLER_24_32 vgnd vpwr scs8hd_decap_6
X_092_ _092_/A _092_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_47 vgnd vpwr scs8hd_decap_12
XFILLER_1_69 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A _139_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _095_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_65 vpwr vgnd scs8hd_fill_2
XFILLER_35_75 vgnd vpwr scs8hd_decap_12
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_27_152 vpwr vgnd scs8hd_fill_2
X_213_ _213_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_144_ address[0] _143_/B _144_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
XFILLER_18_185 vpwr vgnd scs8hd_fill_2
XFILLER_33_177 vgnd vpwr scs8hd_decap_6
XFILLER_33_155 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _091_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_166 vgnd vpwr scs8hd_decap_12
XFILLER_21_44 vpwr vgnd scs8hd_fill_2
XFILLER_21_99 vgnd vpwr scs8hd_decap_12
XFILLER_15_100 vgnd vpwr scs8hd_decap_3
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_7_24 vpwr vgnd scs8hd_fill_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
X_127_ address[3] address[2] _139_/C _139_/D _129_/B vgnd vpwr scs8hd_or4_4
XANTENNA__133__B _155_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_21_136 vgnd vpwr scs8hd_decap_8
XFILLER_21_158 vpwr vgnd scs8hd_fill_2
XFILLER_29_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_107 vgnd vpwr scs8hd_decap_3
XFILLER_16_66 vpwr vgnd scs8hd_fill_2
XFILLER_32_76 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_8_129 vgnd vpwr scs8hd_fill_1
XFILLER_20_180 vgnd vpwr scs8hd_decap_12
XANTENNA__128__B _129_/B vgnd vpwr scs8hd_diode_2
XANTENNA__144__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_173 vpwr vgnd scs8hd_fill_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_4
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _099_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _106_/Y mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_27_98 vpwr vgnd scs8hd_fill_2
XFILLER_27_87 vgnd vpwr scs8hd_decap_4
XFILLER_27_65 vgnd vpwr scs8hd_decap_3
XFILLER_27_10 vpwr vgnd scs8hd_fill_2
XFILLER_4_198 vgnd vpwr scs8hd_decap_4
XFILLER_4_165 vpwr vgnd scs8hd_fill_2
XFILLER_4_143 vgnd vpwr scs8hd_decap_8
XANTENNA__130__C _139_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__141__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_091_ _091_/A _091_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_205 vgnd vpwr scs8hd_fill_1
X_160_ address[0] _160_/B _160_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__136__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__152__A address[3] vgnd vpwr scs8hd_diode_2
Xmem_top_track_10.LATCH_1_.latch data_in _095_/A _140_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_35 vpwr vgnd scs8hd_fill_2
XFILLER_19_22 vgnd vpwr scs8hd_decap_3
XFILLER_19_77 vgnd vpwr scs8hd_decap_6
XFILLER_35_87 vgnd vpwr scs8hd_decap_6
XFILLER_35_32 vgnd vpwr scs8hd_decap_12
X_212_ _212_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
X_143_ _131_/A _143_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_131 vgnd vpwr scs8hd_decap_4
XFILLER_33_167 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _180_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__147__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_8
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_178 vgnd vpwr scs8hd_decap_12
XFILLER_21_56 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _114_/Y mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_30_104 vgnd vpwr scs8hd_fill_1
XFILLER_15_156 vgnd vpwr scs8hd_fill_1
X_126_ address[1] enable _139_/D vgnd vpwr scs8hd_nand2_4
XANTENNA__133__C _139_/C vgnd vpwr scs8hd_diode_2
XFILLER_30_6 vgnd vpwr scs8hd_decap_12
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_119 vgnd vpwr scs8hd_decap_4
XFILLER_20_192 vgnd vpwr scs8hd_decap_12
XFILLER_35_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _118_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_170 vgnd vpwr scs8hd_decap_12
XANTENNA__144__B _143_/B vgnd vpwr scs8hd_diode_2
XANTENNA__160__A address[0] vgnd vpwr scs8hd_diode_2
X_109_ _109_/A _109_/Y vgnd vpwr scs8hd_inv_8
XFILLER_26_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_33 vgnd vpwr scs8hd_decap_4
XFILLER_17_218 vpwr vgnd scs8hd_fill_2
XANTENNA__130__D _155_/D vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_fill_1
XANTENNA__139__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__155__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_1_136 vgnd vpwr scs8hd_decap_4
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
XFILLER_24_56 vgnd vpwr scs8hd_decap_6
X_090_ _090_/A _090_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
XFILLER_6_3 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _102_/A mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__136__C _139_/C vgnd vpwr scs8hd_diode_2
XANTENNA__152__B address[2] vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_0_.latch data_in _106_/A _157_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_25 vgnd vpwr scs8hd_decap_4
XFILLER_35_44 vgnd vpwr scs8hd_decap_12
X_211_ _211_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
X_142_ _139_/A _155_/B _139_/C _155_/D _143_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _120_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__147__B _147_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_4
XANTENNA__163__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_3_ vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_135 vgnd vpwr scs8hd_decap_12
XFILLER_7_37 vgnd vpwr scs8hd_decap_3
X_125_ address[0] _125_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__133__D _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA__158__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_16_46 vgnd vpwr scs8hd_decap_4
XFILLER_32_89 vgnd vpwr scs8hd_decap_3
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
X_108_ _108_/A _108_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_142 vgnd vpwr scs8hd_decap_6
XFILLER_11_182 vgnd vpwr scs8hd_fill_1
XANTENNA__160__B _160_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _109_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _209_/A vgnd vpwr scs8hd_inv_1
XANTENNA__139__C _139_/C vgnd vpwr scs8hd_diode_2
XANTENNA__155__B _155_/B vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_211 vgnd vpwr scs8hd_decap_3
XFILLER_13_69 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_115 vgnd vpwr scs8hd_decap_4
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_9_215 vpwr vgnd scs8hd_fill_2
XANTENNA__166__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _096_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_17 vpwr vgnd scs8hd_fill_2
XANTENNA__136__D _155_/D vgnd vpwr scs8hd_diode_2
XANTENNA__152__C _155_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _092_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_56 vgnd vpwr scs8hd_decap_6
XFILLER_27_144 vgnd vpwr scs8hd_decap_8
XFILLER_27_111 vgnd vpwr scs8hd_decap_3
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
X_210_ _210_/A chany_top_out[3] vgnd vpwr scs8hd_buf_2
X_141_ address[0] _140_/B _141_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _093_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__163__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _111_/A vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _117_/A _174_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_147 vgnd vpwr scs8hd_decap_6
XFILLER_21_25 vpwr vgnd scs8hd_fill_2
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
X_124_ _131_/A _125_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__158__B _155_/B vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _155_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_217 vgnd vpwr scs8hd_decap_12
XFILLER_32_68 vgnd vpwr scs8hd_decap_8
XANTENNA__084__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_128 vgnd vpwr scs8hd_decap_3
X_107_ _107_/A _107_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_90 vpwr vgnd scs8hd_fill_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _098_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__169__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vgnd vpwr scs8hd_decap_4
XFILLER_4_113 vpwr vgnd scs8hd_fill_2
XFILLER_4_102 vgnd vpwr scs8hd_decap_3
XANTENNA__139__D _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _094_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__155__C _155_/C vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _172_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_149 vpwr vgnd scs8hd_fill_2
Xmux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _097_/A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _104_/Y mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_13_223 vpwr vgnd scs8hd_fill_2
XFILLER_0_160 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_82 vpwr vgnd scs8hd_fill_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_208 vgnd vpwr scs8hd_decap_3
XANTENNA__092__A _092_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_1_29 vgnd vpwr scs8hd_decap_3
XANTENNA__152__D _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA__177__A _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_14 vpwr vgnd scs8hd_fill_2
XFILLER_19_36 vpwr vgnd scs8hd_fill_2
XFILLER_19_69 vpwr vgnd scs8hd_fill_2
XFILLER_27_156 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vgnd vpwr scs8hd_decap_6
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
X_140_ _131_/A _140_/B _140_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _101_/Y mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_145 vgnd vpwr scs8hd_decap_8
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_189 vgnd vpwr scs8hd_decap_8
XFILLER_2_61 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_48 vpwr vgnd scs8hd_fill_2
Xmem_top_track_6.LATCH_0_.latch data_in _092_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_129 vgnd vpwr scs8hd_decap_4
XFILLER_30_107 vgnd vpwr scs8hd_fill_1
X_123_ address[3] address[2] _139_/C _155_/D _125_/B vgnd vpwr scs8hd_or4_4
XANTENNA__158__C _155_/C vgnd vpwr scs8hd_diode_2
XANTENNA__174__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XFILLER_29_229 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_111 vpwr vgnd scs8hd_fill_2
XFILLER_7_166 vpwr vgnd scs8hd_fill_2
XFILLER_7_177 vgnd vpwr scs8hd_decap_6
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
X_106_ _106_/A _106_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__169__B _167_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_25 vpwr vgnd scs8hd_fill_2
XFILLER_27_14 vpwr vgnd scs8hd_fill_2
XANTENNA__095__A _095_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_169 vgnd vpwr scs8hd_decap_8
XFILLER_4_125 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_91 vpwr vgnd scs8hd_fill_2
XANTENNA__155__D _155_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_49 vpwr vgnd scs8hd_fill_2
XFILLER_28_90 vpwr vgnd scs8hd_fill_2
XFILLER_0_172 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_50 vpwr vgnd scs8hd_fill_2
XFILLER_5_231 vpwr vgnd scs8hd_fill_2
XFILLER_14_81 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XANTENNA__177__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_39 vgnd vpwr scs8hd_decap_3
XFILLER_27_168 vgnd vpwr scs8hd_decap_12
XFILLER_4_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _117_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_127 vpwr vgnd scs8hd_fill_2
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
XFILLER_18_135 vgnd vpwr scs8hd_fill_1
XFILLER_26_190 vgnd vpwr scs8hd_decap_12
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _199_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _100_/A mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _181_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_105 vpwr vgnd scs8hd_fill_2
XANTENNA__098__A _098_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_149 vgnd vpwr scs8hd_decap_4
X_122_ address[1] _083_/Y _155_/D vgnd vpwr scs8hd_or2_4
XANTENNA__158__D _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__174__C _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_208 vgnd vpwr scs8hd_decap_6
XFILLER_16_16 vpwr vgnd scs8hd_fill_2
Xmem_right_track_10.LATCH_1_.latch data_in _113_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_163 vgnd vpwr scs8hd_decap_3
XFILLER_28_230 vgnd vpwr scs8hd_decap_3
XFILLER_7_123 vpwr vgnd scs8hd_fill_2
XFILLER_11_152 vgnd vpwr scs8hd_decap_3
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
X_105_ _105_/A _105_/Y vgnd vpwr scs8hd_inv_8
XFILLER_19_230 vgnd vpwr scs8hd_decap_3
XFILLER_27_37 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _119_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_184 vpwr vgnd scs8hd_fill_2
XFILLER_5_95 vgnd vpwr scs8hd_decap_4
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_24_38 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _112_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__177__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_180 vgnd vpwr scs8hd_decap_6
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XFILLER_33_106 vpwr vgnd scs8hd_fill_2
XFILLER_18_169 vpwr vgnd scs8hd_fill_2
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_81 vgnd vpwr scs8hd_decap_4
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
XFILLER_32_150 vgnd vpwr scs8hd_decap_3
Xmem_right_track_6.LATCH_1_.latch data_in _109_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_17 vpwr vgnd scs8hd_fill_2
XFILLER_7_19 vgnd vpwr scs8hd_decap_3
X_121_ address[4] address[5] _139_/C vgnd vpwr scs8hd_or2_4
XFILLER_11_83 vpwr vgnd scs8hd_fill_2
XFILLER_14_172 vpwr vgnd scs8hd_fill_2
XFILLER_14_183 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _091_/A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_28 vgnd vpwr scs8hd_fill_1
XFILLER_12_109 vgnd vpwr scs8hd_decap_8
XFILLER_20_142 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_2.LATCH_0_.latch data_in _088_/A _129_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_71 vgnd vpwr scs8hd_decap_12
X_104_ _104_/A _104_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _095_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_62 vgnd vpwr scs8hd_fill_1
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
XFILLER_16_201 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _091_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_171 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_1_119 vgnd vpwr scs8hd_fill_1
XFILLER_9_219 vgnd vpwr scs8hd_decap_12
XFILLER_10_218 vgnd vpwr scs8hd_decap_12
XFILLER_30_93 vgnd vpwr scs8hd_decap_4
Xmux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _095_/A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _197_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _104_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _197_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _097_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_75 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _205_/A vgnd vpwr scs8hd_inv_1
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _120_/A _120_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
XFILLER_11_40 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vgnd vpwr scs8hd_decap_8
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _093_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_195 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _099_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_121 vpwr vgnd scs8hd_fill_2
X_103_ _103_/A _103_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_50 vgnd vpwr scs8hd_decap_8
XFILLER_22_83 vgnd vpwr scs8hd_decap_4
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_8_30 vgnd vpwr scs8hd_fill_1
XFILLER_8_41 vgnd vpwr scs8hd_decap_3
XFILLER_4_139 vpwr vgnd scs8hd_fill_2
XFILLER_4_117 vgnd vpwr scs8hd_decap_6
XFILLER_16_213 vgnd vpwr scs8hd_fill_1
XFILLER_22_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_205 vgnd vpwr scs8hd_decap_3
XFILLER_13_227 vgnd vpwr scs8hd_decap_6
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _094_/A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_164 vgnd vpwr scs8hd_decap_4
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_4
XFILLER_28_82 vgnd vpwr scs8hd_decap_8
XFILLER_5_75 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _200_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_62 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_18 vpwr vgnd scs8hd_fill_2
XFILLER_27_116 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_127 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_25_50 vpwr vgnd scs8hd_fill_2
X_196_ _196_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vpwr vgnd scs8hd_fill_2
XFILLER_24_108 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_152 vgnd vpwr scs8hd_decap_4
XFILLER_23_163 vgnd vpwr scs8hd_decap_12
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
X_179_ _179_/HI _179_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_18 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _098_/A mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_1_.latch data_in _105_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_100 vpwr vgnd scs8hd_fill_2
XFILLER_11_111 vgnd vpwr scs8hd_decap_6
XFILLER_11_133 vpwr vgnd scs8hd_fill_2
XFILLER_11_144 vpwr vgnd scs8hd_fill_2
X_102_ _102_/A _102_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_115 vpwr vgnd scs8hd_fill_2
XFILLER_11_166 vpwr vgnd scs8hd_fill_2
XFILLER_22_40 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_222 vgnd vpwr scs8hd_decap_8
XFILLER_8_20 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_29 vpwr vgnd scs8hd_fill_2
XFILLER_25_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _120_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_129 vgnd vpwr scs8hd_fill_1
XFILLER_4_107 vgnd vpwr scs8hd_decap_3
XFILLER_17_40 vpwr vgnd scs8hd_fill_2
XFILLER_17_62 vpwr vgnd scs8hd_fill_2
XFILLER_17_95 vpwr vgnd scs8hd_fill_2
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _102_/Y mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_0_176 vgnd vpwr scs8hd_decap_8
XFILLER_5_21 vgnd vpwr scs8hd_decap_3
XFILLER_8_232 vgnd vpwr scs8hd_fill_1
XFILLER_5_54 vgnd vpwr scs8hd_decap_4
XFILLER_5_43 vpwr vgnd scs8hd_fill_2
XFILLER_10_209 vgnd vpwr scs8hd_decap_4
XFILLER_14_85 vgnd vpwr scs8hd_decap_4
XFILLER_30_62 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_6
XFILLER_2_205 vgnd vpwr scs8hd_decap_8
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_106 vpwr vgnd scs8hd_fill_2
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_150 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_73 vpwr vgnd scs8hd_fill_2
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/HI _195_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_11 vgnd vpwr scs8hd_fill_1
XANTENNA__112__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XFILLER_17_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _182_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in _102_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_109 vpwr vgnd scs8hd_fill_2
XFILLER_23_175 vgnd vpwr scs8hd_decap_8
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.tap_buf4_0_.scs8hd_inv_1 mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _211_/A vgnd vpwr scs8hd_inv_1
XANTENNA__107__A _107_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_164 vgnd vpwr scs8hd_decap_8
X_178_ _178_/HI _178_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_15_ mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_145 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
X_101_ _101_/A _101_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_127 vpwr vgnd scs8hd_fill_2
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
XFILLER_11_123 vgnd vpwr scs8hd_fill_1
XFILLER_14_9 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_65 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _089_/A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__210__A _210_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _111_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_196 vgnd vpwr scs8hd_decap_4
XANTENNA__120__A _120_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_111 vgnd vpwr scs8hd_fill_1
XFILLER_0_199 vgnd vpwr scs8hd_decap_6
XFILLER_8_211 vgnd vpwr scs8hd_decap_3
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _178_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _098_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _195_/HI _093_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_9_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _094_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_25_30 vpwr vgnd scs8hd_fill_2
XPHY_63 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_85 vgnd vpwr scs8hd_fill_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
X_194_ _194_/HI _194_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_67 vgnd vpwr scs8hd_decap_8
XFILLER_2_45 vgnd vpwr scs8hd_decap_12
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_17_184 vgnd vpwr scs8hd_decap_3
XFILLER_23_132 vgnd vpwr scs8hd_decap_12
XANTENNA__213__A _213_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_87 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_fill_1
X_177_ _139_/D _175_/B address[0] _177_/Y vgnd vpwr scs8hd_nor3_4
Xmux_top_track_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__123__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_102 vgnd vpwr scs8hd_decap_3
XFILLER_9_180 vgnd vpwr scs8hd_fill_1
XFILLER_20_168 vgnd vpwr scs8hd_decap_3
XFILLER_28_213 vgnd vpwr scs8hd_fill_1
X_100_ _100_/A _100_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__208__A _208_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_6
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_88 vgnd vpwr scs8hd_decap_4
Xmux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _189_/HI _097_/Y mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _100_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_12.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XFILLER_16_227 vgnd vpwr scs8hd_decap_6
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
Xmem_top_track_6.LATCH_1_.latch data_in _091_/A _134_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XFILLER_3_153 vgnd vpwr scs8hd_fill_1
XFILLER_3_131 vpwr vgnd scs8hd_fill_2
XFILLER_12_7 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_230 vgnd vpwr scs8hd_decap_3
XFILLER_13_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _103_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
XFILLER_0_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_230 vgnd vpwr scs8hd_decap_3
XANTENNA__131__A _131_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_15_ mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XFILLER_14_43 vpwr vgnd scs8hd_fill_2
XFILLER_14_54 vpwr vgnd scs8hd_fill_2
XFILLER_30_75 vgnd vpwr scs8hd_decap_3
XFILLER_5_215 vpwr vgnd scs8hd_fill_2
XFILLER_29_171 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _092_/A mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_18_119 vgnd vpwr scs8hd_decap_8
XPHY_42 vgnd vpwr scs8hd_decap_3
X_193_ _193_/HI _193_/LO vgnd vpwr scs8hd_conb_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_57 vgnd vpwr scs8hd_decap_4
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _085_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_111 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_11 vpwr vgnd scs8hd_fill_2
XFILLER_14_133 vgnd vpwr scs8hd_decap_3
X_176_ _139_/D _175_/B _131_/A _176_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__123__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_8
XFILLER_22_87 vgnd vpwr scs8hd_fill_1
Xmem_top_track_12.LATCH_0_.latch data_in _098_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_159_ _131_/A _160_/B _159_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_217 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_10 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_53 vgnd vpwr scs8hd_decap_8
XFILLER_33_31 vgnd vpwr scs8hd_decap_12
XFILLER_17_87 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _096_/A mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_121 vgnd vpwr scs8hd_fill_1
XANTENNA__129__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_224 vgnd vpwr scs8hd_decap_8
XFILLER_5_79 vgnd vpwr scs8hd_fill_1
XANTENNA__131__B _131_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_10.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_11_ mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_77 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XANTENNA__126__B enable vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _100_/Y mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _139_/A vgnd vpwr scs8hd_diode_2
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_54 vgnd vpwr scs8hd_decap_4
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
X_192_ _192_/HI _192_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_13_ mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_14 vgnd vpwr scs8hd_fill_1
XFILLER_1_230 vgnd vpwr scs8hd_decap_3
XFILLER_17_120 vpwr vgnd scs8hd_fill_2
XFILLER_17_131 vpwr vgnd scs8hd_fill_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _119_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_101 vpwr vgnd scs8hd_fill_2
XFILLER_2_7 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_34 vgnd vpwr scs8hd_decap_4
XFILLER_14_145 vpwr vgnd scs8hd_fill_2
X_175_ _155_/D _175_/B address[0] _175_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__123__C _139_/C vgnd vpwr scs8hd_diode_2
XFILLER_28_6 vgnd vpwr scs8hd_decap_8
XFILLER_9_193 vgnd vpwr scs8hd_decap_8
XFILLER_3_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_104 vgnd vpwr scs8hd_decap_4
XFILLER_7_119 vgnd vpwr scs8hd_decap_3
XFILLER_11_148 vpwr vgnd scs8hd_fill_2
XFILLER_19_204 vgnd vpwr scs8hd_decap_3
XFILLER_8_24 vgnd vpwr scs8hd_decap_4
XFILLER_8_46 vgnd vpwr scs8hd_decap_3
X_089_ _089_/A _089_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
X_158_ address[3] _155_/B _155_/C _139_/D _160_/B vgnd vpwr scs8hd_or4_4
XANTENNA__134__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA__150__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_229 vgnd vpwr scs8hd_decap_4
XFILLER_17_77 vgnd vpwr scs8hd_decap_8
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vpwr vgnd scs8hd_fill_2
XFILLER_33_43 vgnd vpwr scs8hd_decap_3
XANTENNA__129__B _129_/B vgnd vpwr scs8hd_diode_2
XANTENNA__145__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_fill_1
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _087_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_5_58 vgnd vpwr scs8hd_fill_1
Xmem_top_track_2.LATCH_1_.latch data_in _087_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_89 vgnd vpwr scs8hd_fill_1
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _155_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_187 vgnd vpwr scs8hd_decap_12
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_88 vpwr vgnd scs8hd_fill_2
XFILLER_25_77 vpwr vgnd scs8hd_fill_2
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_25_11 vpwr vgnd scs8hd_fill_2
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XFILLER_17_165 vpwr vgnd scs8hd_fill_2
XANTENNA__137__B _137_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_198 vpwr vgnd scs8hd_fill_2
Xmux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _194_/HI _091_/Y mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__153__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vgnd vpwr scs8hd_decap_4
XFILLER_14_102 vgnd vpwr scs8hd_decap_3
X_174_ _155_/D _175_/B _131_/A _174_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__123__D _155_/D vgnd vpwr scs8hd_diode_2
XANTENNA__148__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_11_ mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_138 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_205 vgnd vpwr scs8hd_decap_8
XFILLER_11_127 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _192_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_58 vgnd vpwr scs8hd_decap_4
XFILLER_8_69 vgnd vpwr scs8hd_decap_4
X_157_ address[0] _157_/B _157_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__B _151_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_175 vgnd vpwr scs8hd_decap_12
X_088_ _088_/A _088_/Y vgnd vpwr scs8hd_inv_8
XFILLER_25_208 vgnd vpwr scs8hd_decap_6
XFILLER_19_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _104_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _097_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_34 vgnd vpwr scs8hd_decap_4
XFILLER_33_11 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.LATCH_0_.latch data_in _120_/A _177_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_156 vgnd vpwr scs8hd_decap_4
XFILLER_3_123 vgnd vpwr scs8hd_decap_3
X_209_ _209_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__145__B _155_/B vgnd vpwr scs8hd_diode_2
XANTENNA__161__A _139_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _093_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_200 vgnd vpwr scs8hd_decap_8
XFILLER_5_26 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _188_/HI _095_/Y mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_7 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _199_/A vgnd vpwr scs8hd_inv_1
XANTENNA__156__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_24 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_6
XFILLER_30_67 vgnd vpwr scs8hd_decap_8
Xmux_top_track_12.tap_buf4_0_.scs8hd_inv_1 mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _207_/A vgnd vpwr scs8hd_inv_1
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XANTENNA__142__C _139_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_199 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_166 vgnd vpwr scs8hd_decap_12
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_25_34 vgnd vpwr scs8hd_decap_3
XFILLER_32_114 vgnd vpwr scs8hd_decap_12
XFILLER_17_144 vpwr vgnd scs8hd_fill_2
XANTENNA__153__B _154_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _106_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _090_/A mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _099_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_14_125 vpwr vgnd scs8hd_fill_2
X_173_ address[3] address[2] address[4] _148_/B _175_/B vgnd vpwr scs8hd_or4_4
XANTENNA__148__B _148_/B vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_180 vgnd vpwr scs8hd_fill_1
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
X_087_ _087_/A _087_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_161 vgnd vpwr scs8hd_decap_12
X_156_ _131_/A _157_/B _156_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__159__A _131_/A vgnd vpwr scs8hd_diode_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_9_ mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _094_/Y mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_3
XFILLER_3_113 vgnd vpwr scs8hd_decap_8
XANTENNA__145__C _139_/C vgnd vpwr scs8hd_diode_2
XANTENNA__161__B address[2] vgnd vpwr scs8hd_diode_2
X_139_ _139_/A address[2] _139_/C _139_/D _140_/B vgnd vpwr scs8hd_or4_4
X_208_ _208_/A chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_31_3 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _202_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_0_138 vgnd vpwr scs8hd_decap_4
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_212 vpwr vgnd scs8hd_fill_2
XANTENNA__156__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA__172__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _086_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_47 vpwr vgnd scs8hd_fill_2
XFILLER_14_58 vpwr vgnd scs8hd_fill_2
XFILLER_5_219 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_29_131 vpwr vgnd scs8hd_fill_2
XANTENNA__142__D _155_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_156 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_178 vgnd vpwr scs8hd_decap_12
XFILLER_26_134 vpwr vgnd scs8hd_fill_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XFILLER_17_112 vpwr vgnd scs8hd_fill_2
XFILLER_32_126 vgnd vpwr scs8hd_decap_12
XFILLER_17_123 vpwr vgnd scs8hd_fill_2
Xmux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _098_/Y mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_148 vpwr vgnd scs8hd_fill_2
XFILLER_23_159 vpwr vgnd scs8hd_fill_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_6
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _111_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_172_ address[0] _172_/B _172_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__164__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_13_170 vgnd vpwr scs8hd_decap_4
XFILLER_20_107 vgnd vpwr scs8hd_decap_3
XFILLER_28_218 vgnd vpwr scs8hd_decap_12
XANTENNA__090__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_218 vpwr vgnd scs8hd_fill_2
XFILLER_8_16 vpwr vgnd scs8hd_fill_2
X_086_ _086_/A _086_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_173 vgnd vpwr scs8hd_decap_12
XFILLER_12_80 vpwr vgnd scs8hd_fill_2
X_155_ address[3] _155_/B _155_/C _155_/D _157_/B vgnd vpwr scs8hd_or4_4
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XFILLER_26_6 vgnd vpwr scs8hd_decap_8
XANTENNA__159__B _160_/B vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _155_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_14 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_1_.latch data_in _101_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
XANTENNA__145__D _139_/D vgnd vpwr scs8hd_diode_2
X_207_ _207_/A chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_138_ address[0] _137_/B _138_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__C _155_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_191 vgnd vpwr scs8hd_decap_12
XFILLER_0_72 vgnd vpwr scs8hd_decap_8
XFILLER_9_92 vpwr vgnd scs8hd_fill_2
XFILLER_28_57 vgnd vpwr scs8hd_decap_12
XFILLER_28_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_39 vpwr vgnd scs8hd_fill_2
Xmem_right_track_12.LATCH_0_.latch data_in _116_/A _172_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__172__B _172_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_80 vgnd vpwr scs8hd_decap_6
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _119_/A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_168 vgnd vpwr scs8hd_decap_12
XANTENNA__167__B _155_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _086_/A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_6_82 vgnd vpwr scs8hd_decap_4
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _213_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_124 vgnd vpwr scs8hd_fill_1
XFILLER_26_102 vpwr vgnd scs8hd_fill_2
XFILLER_25_58 vgnd vpwr scs8hd_fill_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_18 vgnd vpwr scs8hd_decap_12
XFILLER_32_138 vgnd vpwr scs8hd_decap_12
XFILLER_32_105 vgnd vpwr scs8hd_decap_6
XFILLER_23_105 vgnd vpwr scs8hd_decap_6
XFILLER_31_182 vgnd vpwr scs8hd_fill_1
XANTENNA__088__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_149 vgnd vpwr scs8hd_decap_4
X_171_ _131_/A _172_/B _171_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__164__C _155_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_153 vgnd vpwr scs8hd_fill_1
XFILLER_3_94 vpwr vgnd scs8hd_fill_2
XFILLER_11_119 vgnd vpwr scs8hd_decap_3
Xmux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _193_/HI _089_/Y mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_152 vgnd vpwr scs8hd_fill_1
X_085_ _085_/A _085_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_134 vpwr vgnd scs8hd_fill_2
XFILLER_6_189 vgnd vpwr scs8hd_decap_12
XFILLER_10_185 vgnd vpwr scs8hd_decap_12
X_154_ address[0] _154_/B _154_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__175__B _175_/B vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.LATCH_0_.latch data_in _112_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_137_ _131_/A _137_/B _137_/Y vgnd vpwr scs8hd_nor2_4
X_206_ _206_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA__161__D _155_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_107 vpwr vgnd scs8hd_fill_2
XFILLER_28_69 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _114_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__096__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_5_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_155 vpwr vgnd scs8hd_fill_2
XFILLER_29_144 vpwr vgnd scs8hd_fill_2
XFILLER_4_232 vgnd vpwr scs8hd_fill_1
XFILLER_35_125 vgnd vpwr scs8hd_decap_12
XANTENNA__167__C _155_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _100_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vpwr vgnd scs8hd_fill_2
XFILLER_17_169 vgnd vpwr scs8hd_decap_12
XFILLER_31_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _103_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_150 vgnd vpwr scs8hd_decap_12
X_170_ _139_/A _155_/B _155_/C _139_/D _172_/B vgnd vpwr scs8hd_or4_4
XFILLER_26_80 vgnd vpwr scs8hd_decap_12
XANTENNA__164__D _139_/D vgnd vpwr scs8hd_diode_2
XFILLER_9_132 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_16 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _193_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _088_/A mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_142 vpwr vgnd scs8hd_fill_2
X_153_ _131_/A _154_/B _153_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_197 vgnd vpwr scs8hd_decap_12
X_084_ address[0] _131_/A vgnd vpwr scs8hd_inv_8
XFILLER_12_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__175__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _102_/A vgnd vpwr
+ scs8hd_diode_2
X_136_ _139_/A address[2] _139_/C _155_/D _137_/B vgnd vpwr scs8hd_or4_4
X_205_ _205_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _085_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_30 vgnd vpwr scs8hd_fill_1
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _092_/Y mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _105_/A vgnd vpwr
+ scs8hd_diode_2
X_119_ _119_/A _119_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
Xmem_top_track_12.LATCH_1_.latch data_in _097_/A _143_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _184_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_123 vgnd vpwr scs8hd_fill_1
XFILLER_29_101 vpwr vgnd scs8hd_fill_2
XFILLER_35_137 vgnd vpwr scs8hd_decap_12
XANTENNA__167__D _155_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_17_148 vpwr vgnd scs8hd_fill_2
XFILLER_31_92 vgnd vpwr scs8hd_decap_8
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_162 vgnd vpwr scs8hd_decap_12
XFILLER_14_107 vgnd vpwr scs8hd_decap_3
XFILLER_14_129 vpwr vgnd scs8hd_fill_2
XFILLER_22_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _088_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_140 vpwr vgnd scs8hd_fill_2
XFILLER_13_184 vpwr vgnd scs8hd_fill_2
XFILLER_22_28 vgnd vpwr scs8hd_fill_1
Xmux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _096_/Y mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_083_ enable _083_/Y vgnd vpwr scs8hd_inv_8
X_152_ address[3] address[2] _155_/C _139_/D _154_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _109_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_232 vgnd vpwr scs8hd_fill_1
XFILLER_5_180 vgnd vpwr scs8hd_fill_1
XFILLER_17_28 vgnd vpwr scs8hd_decap_4
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
XFILLER_33_49 vpwr vgnd scs8hd_fill_2
XFILLER_33_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_202 vgnd vpwr scs8hd_fill_1
X_204_ _204_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
X_135_ address[0] _134_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_172 vgnd vpwr scs8hd_decap_4
XFILLER_24_6 vpwr vgnd scs8hd_fill_2
XFILLER_0_42 vgnd vpwr scs8hd_fill_1
XFILLER_9_40 vpwr vgnd scs8hd_fill_2
XFILLER_9_73 vpwr vgnd scs8hd_fill_2
XFILLER_18_60 vpwr vgnd scs8hd_fill_2
XFILLER_18_71 vgnd vpwr scs8hd_decap_12
XFILLER_7_220 vpwr vgnd scs8hd_fill_2
X_118_ _118_/A _118_/Y vgnd vpwr scs8hd_inv_8
Xmem_right_track_4.LATCH_0_.latch data_in _108_/A _160_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_149 vgnd vpwr scs8hd_decap_6
XFILLER_6_41 vgnd vpwr scs8hd_decap_4
XFILLER_26_138 vgnd vpwr scs8hd_decap_12
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_182 vgnd vpwr scs8hd_fill_1
XFILLER_17_116 vpwr vgnd scs8hd_fill_2
XFILLER_17_127 vpwr vgnd scs8hd_fill_2
XFILLER_15_83 vpwr vgnd scs8hd_fill_2
XFILLER_31_174 vgnd vpwr scs8hd_decap_8
XFILLER_31_141 vgnd vpwr scs8hd_fill_1
XFILLER_16_171 vgnd vpwr scs8hd_decap_3
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _117_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_119 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_163 vgnd vpwr scs8hd_decap_12
XFILLER_9_101 vpwr vgnd scs8hd_fill_2
XFILLER_13_163 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_156 vgnd vpwr scs8hd_decap_12
XFILLER_3_53 vgnd vpwr scs8hd_decap_8
XFILLER_3_20 vgnd vpwr scs8hd_decap_4
X_151_ address[0] _151_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_115 vpwr vgnd scs8hd_fill_2
XFILLER_12_40 vgnd vpwr scs8hd_decap_4
XFILLER_12_84 vgnd vpwr scs8hd_decap_8
X_082_ address[2] _155_/B vgnd vpwr scs8hd_inv_8
XFILLER_33_225 vpwr vgnd scs8hd_fill_2
XFILLER_33_214 vpwr vgnd scs8hd_fill_2
XFILLER_18_211 vgnd vpwr scs8hd_decap_3
XFILLER_5_170 vpwr vgnd scs8hd_fill_2
XFILLER_15_214 vgnd vpwr scs8hd_decap_8
XFILLER_15_225 vpwr vgnd scs8hd_fill_2
X_203_ _203_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _192_/HI _087_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_134_ _131_/A _134_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_10 vgnd vpwr scs8hd_decap_12
XFILLER_17_6 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_4
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_96 vgnd vpwr scs8hd_decap_3
XFILLER_18_83 vgnd vpwr scs8hd_decap_3
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_232 vgnd vpwr scs8hd_fill_1
X_117_ _117_/A _117_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_3 vgnd vpwr scs8hd_decap_4
XFILLER_30_18 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _112_/A mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_224 vgnd vpwr scs8hd_decap_8
XFILLER_4_202 vgnd vpwr scs8hd_fill_1
XFILLER_35_106 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.LATCH_1_.latch data_in _119_/A _176_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_20 vgnd vpwr scs8hd_decap_4
XFILLER_6_64 vpwr vgnd scs8hd_fill_2
XFILLER_26_106 vgnd vpwr scs8hd_decap_12
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_17_106 vgnd vpwr scs8hd_decap_4
XFILLER_15_62 vgnd vpwr scs8hd_decap_4
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_183 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_175 vgnd vpwr scs8hd_decap_12
XFILLER_13_197 vgnd vpwr scs8hd_decap_8
XFILLER_9_168 vgnd vpwr scs8hd_decap_12
XFILLER_3_65 vpwr vgnd scs8hd_fill_2
XFILLER_3_43 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _113_/A vgnd
+ vpwr scs8hd_diode_2
X_150_ _131_/A _151_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_081_ address[3] _139_/A vgnd vpwr scs8hd_inv_8
XFILLER_6_105 vgnd vpwr scs8hd_fill_1
XFILLER_6_138 vgnd vpwr scs8hd_decap_12
XFILLER_12_74 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _106_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_218 vgnd vpwr scs8hd_decap_12
X_202_ _202_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_133_ address[3] _155_/B _139_/C _139_/D _134_/B vgnd vpwr scs8hd_or4_4
XFILLER_23_73 vgnd vpwr scs8hd_decap_12
XFILLER_2_152 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _120_/A mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _099_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_22 vgnd vpwr scs8hd_decap_8
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _085_/A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_88 vgnd vpwr scs8hd_decap_3
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_12_218 vgnd vpwr scs8hd_decap_12
X_116_ _116_/A _116_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XFILLER_29_148 vgnd vpwr scs8hd_decap_4
XFILLER_20_41 vgnd vpwr scs8hd_decap_3
XFILLER_20_63 vpwr vgnd scs8hd_fill_2
XFILLER_35_118 vgnd vpwr scs8hd_decap_6
XFILLER_28_181 vgnd vpwr scs8hd_decap_12
XFILLER_26_118 vgnd vpwr scs8hd_decap_6
Xmux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _090_/Y mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in _094_/A _138_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_0_.latch data_in _104_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_206 vgnd vpwr scs8hd_decap_12
XFILLER_25_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_110 vpwr vgnd scs8hd_fill_2
XFILLER_22_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _108_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_187 vgnd vpwr scs8hd_decap_12
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _086_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _101_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_176 vgnd vpwr scs8hd_decap_4
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
X_080_ address[5] _148_/B vgnd vpwr scs8hd_inv_8
XFILLER_10_102 vgnd vpwr scs8hd_decap_3
XFILLER_10_135 vgnd vpwr scs8hd_decap_4
XFILLER_10_146 vgnd vpwr scs8hd_decap_6
XFILLER_10_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _194_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_3 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _204_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_224 vgnd vpwr scs8hd_decap_8
XANTENNA__108__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_201_ _201_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
X_132_ address[0] _131_/B _132_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_85 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _196_/A vgnd vpwr scs8hd_inv_1
XFILLER_9_65 vpwr vgnd scs8hd_fill_2
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _107_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_208 vpwr vgnd scs8hd_fill_2
XFILLER_20_230 vgnd vpwr scs8hd_decap_3
XANTENNA__211__A _211_/A vgnd vpwr scs8hd_diode_2
X_115_ _115_/A _115_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__121__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_127 vpwr vgnd scs8hd_fill_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _087_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _185_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_73 vgnd vpwr scs8hd_decap_3
XFILLER_28_193 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_88 vgnd vpwr scs8hd_decap_4
XFILLER_20_3 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _186_/HI _111_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_196 vgnd vpwr scs8hd_decap_12
XFILLER_25_152 vgnd vpwr scs8hd_decap_12
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_74 vgnd vpwr scs8hd_decap_4
XFILLER_31_100 vpwr vgnd scs8hd_fill_2
XFILLER_16_141 vpwr vgnd scs8hd_fill_2
XFILLER_16_163 vgnd vpwr scs8hd_decap_8
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

