* NGSPICE file created from cbx_1__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt cbx_1__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_grid_pin_0_ bottom_grid_pin_4_ bottom_grid_pin_8_ chanx_left_in[0]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ data_in enable top_grid_pin_0_ top_grid_pin_10_ top_grid_pin_12_ top_grid_pin_14_
+ top_grid_pin_2_ top_grid_pin_4_ top_grid_pin_6_ top_grid_pin_8_ vpwr vgnd
XFILLER_7_7 vpwr vgnd scs8hd_fill_2
XFILLER_26_41 vpwr vgnd scs8hd_fill_2
XFILLER_13_111 vpwr vgnd scs8hd_fill_2
XFILLER_9_104 vpwr vgnd scs8hd_fill_2
XFILLER_9_115 vgnd vpwr scs8hd_decap_6
XFILLER_9_126 vpwr vgnd scs8hd_fill_2
XFILLER_13_177 vgnd vpwr scs8hd_decap_4
XFILLER_3_23 vpwr vgnd scs8hd_fill_2
XANTENNA__113__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_1_.latch data_in mem_bottom_ipin_2.LATCH_1_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_32 vgnd vpwr scs8hd_decap_3
XFILLER_12_76 vgnd vpwr scs8hd_decap_3
XANTENNA__108__B _108_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_140 vpwr vgnd scs8hd_fill_2
XANTENNA__124__A _055_/D vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_4_.latch data_in mem_bottom_ipin_4.LATCH_4_.latch/Q _070_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_062_ _062_/A _088_/A _062_/Y vgnd vpwr scs8hd_nor2_4
X_131_ _131_/HI _131_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_110 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__110__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_9_22 vgnd vpwr scs8hd_decap_4
XANTENNA__119__A _086_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_53 vgnd vpwr scs8hd_decap_3
XFILLER_7_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_045_ _045_/A _045_/Y vgnd vpwr scs8hd_inv_8
X_114_ _088_/A _111_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__121__B _123_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_2_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_106 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_21 vpwr vgnd scs8hd_fill_2
XFILLER_20_32 vpwr vgnd scs8hd_fill_2
XFILLER_29_52 vpwr vgnd scs8hd_fill_2
XFILLER_28_194 vgnd vpwr scs8hd_decap_12
XANTENNA__116__B _111_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _131_/HI mem_bottom_ipin_0.LATCH_5_.latch/Q
+ mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__042__A address[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_120 vpwr vgnd scs8hd_fill_2
XFILLER_25_197 vgnd vpwr scs8hd_decap_12
XFILLER_31_97 vpwr vgnd scs8hd_fill_2
XFILLER_31_156 vgnd vpwr scs8hd_decap_12
XFILLER_31_112 vgnd vpwr scs8hd_decap_12
XFILLER_31_101 vgnd vpwr scs8hd_decap_4
XANTENNA__127__A _127_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_112 vgnd vpwr scs8hd_decap_3
XFILLER_26_64 vgnd vpwr scs8hd_decap_3
XFILLER_26_20 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_5.LATCH_0_.latch data_in mem_bottom_ipin_5.LATCH_0_.latch/Q _082_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_123 vgnd vpwr scs8hd_decap_3
XFILLER_13_156 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_137 vpwr vgnd scs8hd_fill_2
XFILLER_10_148 vpwr vgnd scs8hd_fill_2
XFILLER_12_55 vpwr vgnd scs8hd_fill_2
XFILLER_12_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_7.LATCH_3_.latch data_in mem_bottom_ipin_7.LATCH_3_.latch/Q _094_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_SLEEPB _064_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__108__C _108_/C vgnd vpwr scs8hd_diode_2
XFILLER_5_174 vpwr vgnd scs8hd_fill_2
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XANTENNA__050__A address[6] vgnd vpwr scs8hd_diode_2
X_130_ _090_/A _127_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_21 vgnd vpwr scs8hd_decap_3
X_061_ _059_/A address[2] address[0] _088_/A vgnd vpwr scs8hd_or3_4
XFILLER_23_76 vpwr vgnd scs8hd_fill_2
XANTENNA__110__D _055_/D vgnd vpwr scs8hd_diode_2
XFILLER_0_25 vpwr vgnd scs8hd_fill_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_45 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_210 vpwr vgnd scs8hd_fill_2
XANTENNA__045__A _045_/A vgnd vpwr scs8hd_diode_2
X_113_ _127_/A _111_/B _113_/Y vgnd vpwr scs8hd_nor2_4
X_044_ _044_/A _044_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_7 vpwr vgnd scs8hd_fill_2
XFILLER_22_8 vgnd vpwr scs8hd_decap_3
XFILLER_29_129 vgnd vpwr scs8hd_fill_1
XFILLER_20_55 vgnd vpwr scs8hd_decap_3
XFILLER_29_75 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_173 vpwr vgnd scs8hd_fill_2
XFILLER_15_11 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_54 vgnd vpwr scs8hd_decap_8
XFILLER_31_21 vgnd vpwr scs8hd_decap_8
XFILLER_31_10 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_168 vgnd vpwr scs8hd_decap_12
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA__143__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XANTENNA__053__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_26_32 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_0.LATCH_4_.latch data_in mem_top_ipin_0.LATCH_4_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_76 vpwr vgnd scs8hd_fill_2
XFILLER_3_69 vpwr vgnd scs8hd_fill_2
XFILLER_3_36 vpwr vgnd scs8hd_fill_2
XFILLER_3_14 vpwr vgnd scs8hd_fill_2
XANTENNA__048__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_10_105 vgnd vpwr scs8hd_decap_4
XFILLER_10_116 vpwr vgnd scs8hd_fill_2
XFILLER_12_12 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _043_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_153 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_060_ _062_/A _127_/A _060_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_99 vgnd vpwr scs8hd_decap_3
XFILLER_2_167 vgnd vpwr scs8hd_decap_4
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__151__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__061__A _059_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_4_.latch data_in mem_bottom_ipin_0.LATCH_4_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_88 vgnd vpwr scs8hd_fill_1
X_043_ _043_/A _043_/Y vgnd vpwr scs8hd_inv_8
X_112_ _086_/A _111_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__056__A _056_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_36 vgnd vpwr scs8hd_fill_1
Xmem_top_ipin_1.LATCH_0_.latch data_in _044_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_25_166 vpwr vgnd scs8hd_fill_2
XFILLER_25_155 vpwr vgnd scs8hd_fill_2
XFILLER_25_144 vpwr vgnd scs8hd_fill_2
XFILLER_31_77 vpwr vgnd scs8hd_fill_2
XFILLER_31_66 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_31_125 vgnd vpwr scs8hd_decap_12
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_199 vgnd vpwr scs8hd_decap_12
XFILLER_22_125 vgnd vpwr scs8hd_fill_1
XFILLER_22_147 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__053__B _048_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_191 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__154__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_8_195 vpwr vgnd scs8hd_fill_2
XFILLER_12_180 vgnd vpwr scs8hd_decap_4
XFILLER_12_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__064__A _062_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_187 vpwr vgnd scs8hd_fill_2
XFILLER_5_198 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.LATCH_0_.latch data_in mem_bottom_ipin_1.LATCH_0_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XANTENNA__059__A _059_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_45 vpwr vgnd scs8hd_fill_2
XFILLER_23_56 vgnd vpwr scs8hd_decap_3
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_3.LATCH_3_.latch data_in mem_bottom_ipin_3.LATCH_3_.latch/Q _060_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _045_/A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__061__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_23 vgnd vpwr scs8hd_decap_8
XFILLER_18_45 vgnd vpwr scs8hd_decap_8
XFILLER_18_67 vpwr vgnd scs8hd_fill_2
X_042_ address[0] _108_/C vgnd vpwr scs8hd_inv_8
Xmux_top_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_111_ _056_/A _111_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__056__B _062_/A vgnd vpwr scs8hd_diode_2
XANTENNA__072__A _088_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_SLEEPB _071_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_99 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_26 vgnd vpwr scs8hd_decap_3
XANTENNA__157__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_2_.latch/Q mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_4
XFILLER_25_112 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_79 vgnd vpwr scs8hd_decap_4
XFILLER_16_145 vgnd vpwr scs8hd_decap_6
XFILLER_31_137 vgnd vpwr scs8hd_decap_12
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_137 vgnd vpwr scs8hd_decap_3
XANTENNA__053__C _108_/C vgnd vpwr scs8hd_diode_2
XFILLER_26_56 vgnd vpwr scs8hd_decap_6
XFILLER_13_115 vpwr vgnd scs8hd_fill_2
XFILLER_9_108 vgnd vpwr scs8hd_decap_4
XFILLER_21_170 vgnd vpwr scs8hd_fill_1
XFILLER_8_163 vgnd vpwr scs8hd_decap_8
XANTENNA__064__B _089_/A vgnd vpwr scs8hd_diode_2
XANTENNA__080__A _088_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_70 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_6.LATCH_2_.latch data_in mem_bottom_ipin_6.LATCH_2_.latch/Q _088_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__059__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__075__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_114 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_202 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__061__C address[0] vgnd vpwr scs8hd_diode_2
X_110_ _091_/A address[4] address[3] _055_/D _111_/B vgnd vpwr scs8hd_or4_4
XFILLER_7_206 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _131_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__072__B _071_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_25 vpwr vgnd scs8hd_fill_2
XFILLER_20_36 vpwr vgnd scs8hd_fill_2
XFILLER_20_47 vgnd vpwr scs8hd_decap_8
XFILLER_29_56 vgnd vpwr scs8hd_decap_3
XFILLER_29_12 vpwr vgnd scs8hd_fill_2
XFILLER_28_154 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_80 vpwr vgnd scs8hd_fill_2
XFILLER_19_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_187 vpwr vgnd scs8hd_fill_2
XFILLER_19_198 vpwr vgnd scs8hd_fill_2
XFILLER_31_35 vgnd vpwr scs8hd_decap_8
XANTENNA__067__B _098_/B vgnd vpwr scs8hd_diode_2
XANTENNA__083__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_25 vpwr vgnd scs8hd_fill_2
XFILLER_15_36 vpwr vgnd scs8hd_fill_2
XFILLER_31_149 vgnd vpwr scs8hd_decap_6
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_92 vpwr vgnd scs8hd_fill_2
XFILLER_26_24 vgnd vpwr scs8hd_decap_4
XANTENNA__078__A _086_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _043_/A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_208 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_59 vpwr vgnd scs8hd_fill_2
XANTENNA__080__B _081_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_123 vpwr vgnd scs8hd_fill_2
XFILLER_5_112 vpwr vgnd scs8hd_fill_2
XFILLER_5_178 vgnd vpwr scs8hd_decap_4
XANTENNA__059__C _108_/C vgnd vpwr scs8hd_diode_2
XANTENNA__075__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_23_211 vgnd vpwr scs8hd_fill_1
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_126 vgnd vpwr scs8hd_decap_3
XFILLER_0_29 vpwr vgnd scs8hd_fill_2
XFILLER_9_16 vgnd vpwr scs8hd_decap_4
XFILLER_1_170 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_0_.latch/Q mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_100 vpwr vgnd scs8hd_fill_2
XFILLER_19_166 vgnd vpwr scs8hd_decap_4
XFILLER_19_177 vgnd vpwr scs8hd_decap_6
XFILLER_15_15 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__083__B _091_/B vgnd vpwr scs8hd_diode_2
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_80 vgnd vpwr scs8hd_decap_4
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_15_180 vgnd vpwr scs8hd_fill_1
XFILLER_22_117 vpwr vgnd scs8hd_fill_2
XANTENNA__078__B _081_/B vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_139 vpwr vgnd scs8hd_fill_2
XFILLER_3_18 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_SLEEPB _077_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_109 vgnd vpwr scs8hd_fill_1
XFILLER_12_16 vpwr vgnd scs8hd_fill_2
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XFILLER_12_38 vpwr vgnd scs8hd_fill_2
XANTENNA__089__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_209 vgnd vpwr scs8hd_decap_3
XFILLER_5_157 vpwr vgnd scs8hd_fill_2
XFILLER_27_90 vgnd vpwr scs8hd_decap_3
XFILLER_4_83 vpwr vgnd scs8hd_fill_2
XANTENNA__075__C _091_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_26 vpwr vgnd scs8hd_fill_2
XANTENNA__091__B _091_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XFILLER_9_28 vpwr vgnd scs8hd_fill_2
XFILLER_13_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_193 vpwr vgnd scs8hd_fill_2
XFILLER_18_15 vpwr vgnd scs8hd_fill_2
XANTENNA__086__B _088_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_204 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_2.LATCH_2_.latch data_in mem_bottom_ipin_2.LATCH_2_.latch/Q _128_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_27_3 vpwr vgnd scs8hd_fill_2
X_099_ _091_/A address[4] address[3] _108_/B _102_/B vgnd vpwr scs8hd_or4_4
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XFILLER_1_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _132_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_5_.latch data_in mem_bottom_ipin_4.LATCH_5_.latch/Q _069_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__097__A _090_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_3_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_10_93 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_159 vpwr vgnd scs8hd_fill_2
XFILLER_25_148 vgnd vpwr scs8hd_decap_4
XFILLER_25_104 vpwr vgnd scs8hd_fill_2
XANTENNA__083__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_16_126 vpwr vgnd scs8hd_fill_2
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_30_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_37 vpwr vgnd scs8hd_fill_2
XANTENNA__094__B _093_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_107 vpwr vgnd scs8hd_fill_2
XFILLER_21_173 vgnd vpwr scs8hd_decap_8
XFILLER_8_144 vpwr vgnd scs8hd_fill_2
XFILLER_12_195 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__089__B _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_136 vpwr vgnd scs8hd_fill_2
XFILLER_4_180 vgnd vpwr scs8hd_decap_8
XFILLER_4_62 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_0_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__091__C _091_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_106 vpwr vgnd scs8hd_fill_2
XFILLER_13_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_5.LATCH_1_.latch data_in mem_bottom_ipin_5.LATCH_1_.latch/Q _081_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_SLEEPB _074_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_24_81 vgnd vpwr scs8hd_decap_8
XFILLER_24_70 vpwr vgnd scs8hd_fill_2
X_098_ address[5] _098_/B _108_/B vgnd vpwr scs8hd_or2_4
Xmem_bottom_ipin_7.LATCH_4_.latch data_in mem_bottom_ipin_7.LATCH_4_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_20_17 vpwr vgnd scs8hd_fill_2
XFILLER_29_48 vpwr vgnd scs8hd_fill_2
XFILLER_28_135 vgnd vpwr scs8hd_decap_12
XFILLER_28_124 vgnd vpwr scs8hd_decap_8
XFILLER_28_113 vgnd vpwr scs8hd_decap_8
XFILLER_28_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XANTENNA__097__B _093_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_116 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_108 vpwr vgnd scs8hd_fill_2
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_193 vpwr vgnd scs8hd_fill_2
XFILLER_7_51 vpwr vgnd scs8hd_fill_2
XFILLER_7_73 vpwr vgnd scs8hd_fill_2
XFILLER_26_16 vpwr vgnd scs8hd_fill_2
XFILLER_13_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_71 vpwr vgnd scs8hd_fill_2
XFILLER_16_93 vgnd vpwr scs8hd_decap_4
XFILLER_8_134 vgnd vpwr scs8hd_fill_1
XFILLER_12_130 vgnd vpwr scs8hd_decap_4
XFILLER_12_163 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ _046_/A mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_211 vgnd vpwr scs8hd_fill_1
XFILLER_5_104 vpwr vgnd scs8hd_fill_2
XFILLER_17_211 vgnd vpwr scs8hd_fill_1
XFILLER_4_192 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_203 vgnd vpwr scs8hd_decap_8
XFILLER_23_17 vpwr vgnd scs8hd_fill_2
XANTENNA__091__D _091_/D vgnd vpwr scs8hd_diode_2
XFILLER_1_140 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_0.LATCH_5_.latch data_in mem_top_ipin_0.LATCH_5_.latch/Q _100_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
XFILLER_6_210 vpwr vgnd scs8hd_fill_2
X_097_ _090_/A _093_/B _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_1_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _133_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_29 vpwr vgnd scs8hd_fill_2
XFILLER_29_16 vpwr vgnd scs8hd_fill_2
XFILLER_28_158 vgnd vpwr scs8hd_decap_12
XFILLER_28_147 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_40 vpwr vgnd scs8hd_fill_2
XFILLER_10_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_136 vpwr vgnd scs8hd_fill_2
X_149_ chanx_right_in[1] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_17 vpwr vgnd scs8hd_fill_2
XFILLER_15_29 vpwr vgnd scs8hd_fill_2
XFILLER_18_180 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_0.LATCH_5_.latch data_in mem_bottom_ipin_0.LATCH_5_.latch/Q _111_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_0_.latch/Q mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_161 vpwr vgnd scs8hd_fill_2
XFILLER_15_172 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_30 vpwr vgnd scs8hd_fill_2
XFILLER_26_28 vgnd vpwr scs8hd_fill_1
XFILLER_21_153 vpwr vgnd scs8hd_fill_2
XFILLER_8_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_50 vpwr vgnd scs8hd_fill_2
XFILLER_12_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_1.LATCH_1_.latch data_in _043_/A _106_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_116 vgnd vpwr scs8hd_decap_4
XFILLER_27_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_20 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_95 vgnd vpwr scs8hd_fill_1
XFILLER_1_174 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _056_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_7 vgnd vpwr scs8hd_fill_1
X_096_ _089_/A _093_/B _096_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_98 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.LATCH_1_.latch data_in mem_bottom_ipin_1.LATCH_1_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _044_/A mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_19_104 vpwr vgnd scs8hd_fill_2
X_148_ chanx_right_in[2] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
X_079_ _127_/A _081_/B _079_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_129 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_3.LATCH_4_.latch data_in mem_bottom_ipin_3.LATCH_4_.latch/Q _058_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_29 vpwr vgnd scs8hd_fill_2
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_decap_3
XFILLER_21_84 vgnd vpwr scs8hd_fill_1
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_21_110 vgnd vpwr scs8hd_fill_1
XFILLER_21_132 vpwr vgnd scs8hd_fill_2
XFILLER_21_187 vpwr vgnd scs8hd_fill_2
XFILLER_21_198 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_125 vgnd vpwr scs8hd_fill_1
XFILLER_16_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_191 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_150 vgnd vpwr scs8hd_fill_1
XFILLER_4_87 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _141_/HI _045_/Y mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_197 vgnd vpwr scs8hd_decap_4
XFILLER_1_153 vpwr vgnd scs8hd_fill_2
XANTENNA__100__B _102_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_19 vpwr vgnd scs8hd_fill_2
XFILLER_11_208 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_0_.latch/Q mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_0_.latch data_in mem_bottom_ipin_4.LATCH_0_.latch/Q _074_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_095_ _088_/A _093_/B _095_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_SLEEPB _060_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_7 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _056_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _134_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_29_29 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_6.LATCH_3_.latch data_in mem_bottom_ipin_6.LATCH_3_.latch/Q _087_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_204 vpwr vgnd scs8hd_fill_2
XFILLER_10_64 vgnd vpwr scs8hd_decap_3
XFILLER_19_73 vpwr vgnd scs8hd_fill_2
XFILLER_19_149 vpwr vgnd scs8hd_fill_2
XFILLER_27_182 vgnd vpwr scs8hd_fill_1
XANTENNA__106__A _117_/B vgnd vpwr scs8hd_diode_2
X_078_ _086_/A _081_/B _078_/Y vgnd vpwr scs8hd_nor2_4
X_147_ chanx_right_in[3] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_18_3 vgnd vpwr scs8hd_fill_1
XFILLER_25_108 vpwr vgnd scs8hd_fill_2
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_174 vgnd vpwr scs8hd_decap_12
XFILLER_24_163 vgnd vpwr scs8hd_decap_8
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_21_166 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_148 vgnd vpwr scs8hd_decap_3
XANTENNA__103__B _102_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_203 vgnd vpwr scs8hd_decap_8
XFILLER_27_95 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_66 vpwr vgnd scs8hd_fill_2
XANTENNA__114__A _088_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_13_75 vpwr vgnd scs8hd_fill_2
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_74 vgnd vpwr scs8hd_decap_4
XFILLER_24_41 vgnd vpwr scs8hd_decap_4
X_094_ _127_/A _093_/B _094_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_202 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_23 vpwr vgnd scs8hd_fill_2
XANTENNA__111__B _111_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_8_ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_106 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_7.LATCH_3_.latch/Q mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_32 vgnd vpwr scs8hd_fill_1
XFILLER_10_76 vpwr vgnd scs8hd_fill_2
XFILLER_19_41 vpwr vgnd scs8hd_fill_2
XFILLER_19_52 vpwr vgnd scs8hd_fill_2
XFILLER_19_85 vpwr vgnd scs8hd_fill_2
XANTENNA__106__B _108_/B vgnd vpwr scs8hd_diode_2
X_077_ _056_/A _081_/B _077_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__A _089_/A vgnd vpwr scs8hd_diode_2
X_146_ chanx_right_in[4] chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_0_208 vgnd vpwr scs8hd_decap_4
XFILLER_16_109 vgnd vpwr scs8hd_decap_8
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_186 vgnd vpwr scs8hd_decap_12
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_42 vpwr vgnd scs8hd_fill_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _140_/HI _043_/Y mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XFILLER_7_22 vpwr vgnd scs8hd_fill_2
XFILLER_7_55 vgnd vpwr scs8hd_decap_4
XANTENNA__117__A _055_/D vgnd vpwr scs8hd_diode_2
XFILLER_7_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_197 vgnd vpwr scs8hd_decap_4
XFILLER_30_3 vpwr vgnd scs8hd_fill_2
X_129_ _089_/A _127_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_145 vpwr vgnd scs8hd_fill_2
XFILLER_12_167 vpwr vgnd scs8hd_fill_2
XFILLER_16_97 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_0_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_108 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_163 vgnd vpwr scs8hd_decap_8
XFILLER_4_45 vpwr vgnd scs8hd_fill_2
XANTENNA__130__A _090_/A vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_0_.latch data_in mem_top_ipin_0.LATCH_0_.latch/Q _105_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_21 vpwr vgnd scs8hd_fill_2
XFILLER_1_111 vgnd vpwr scs8hd_decap_4
XFILLER_8_3 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _108_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _056_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_1_.latch/Q mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_093_ _086_/A _093_/B _093_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _135_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_44 vpwr vgnd scs8hd_fill_2
XFILLER_10_88 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
X_145_ chanx_right_in[5] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__106__C _108_/C vgnd vpwr scs8hd_diode_2
X_076_ _091_/D _117_/B _081_/B vgnd vpwr scs8hd_or2_4
XANTENNA__122__B _123_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_0_.latch data_in mem_bottom_ipin_0.LATCH_0_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_198 vgnd vpwr scs8hd_decap_12
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_10 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_76 vpwr vgnd scs8hd_fill_2
XFILLER_21_87 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_165 vpwr vgnd scs8hd_fill_2
XFILLER_15_176 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_2.LATCH_3_.latch data_in mem_bottom_ipin_2.LATCH_3_.latch/Q _127_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_34 vpwr vgnd scs8hd_fill_2
XANTENNA__117__B _117_/B vgnd vpwr scs8hd_diode_2
X_128_ _088_/A _127_/B _128_/Y vgnd vpwr scs8hd_nor2_4
X_059_ _059_/A address[2] _108_/C _127_/A vgnd vpwr scs8hd_or3_4
XFILLER_23_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_102 vpwr vgnd scs8hd_fill_2
XANTENNA__043__A _043_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_SLEEPB _069_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_21 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XFILLER_16_54 vpwr vgnd scs8hd_fill_2
XFILLER_8_106 vpwr vgnd scs8hd_fill_2
XFILLER_8_128 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _088_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XFILLER_27_42 vpwr vgnd scs8hd_fill_2
XFILLER_4_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__130__B _127_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_6.LATCH_3_.latch/Q mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_33 vgnd vpwr scs8hd_decap_3
XFILLER_13_88 vgnd vpwr scs8hd_decap_4
XFILLER_1_178 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA__109__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__051__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_4_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
X_092_ _056_/A _093_/B _092_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _046_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__046__A _046_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_12 vpwr vgnd scs8hd_fill_2
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_19_108 vgnd vpwr scs8hd_decap_3
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
X_075_ _091_/A address[4] _091_/C _117_/B vgnd vpwr scs8hd_or3_4
X_144_ chanx_right_in[6] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XFILLER_24_133 vgnd vpwr scs8hd_fill_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_5.LATCH_2_.latch data_in mem_bottom_ipin_5.LATCH_2_.latch/Q _080_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_144 vpwr vgnd scs8hd_fill_2
X_127_ _127_/A _127_/B _127_/Y vgnd vpwr scs8hd_nor2_4
X_058_ _062_/A _086_/A _058_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_3 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_7.LATCH_5_.latch data_in mem_bottom_ipin_7.LATCH_5_.latch/Q _092_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_21_136 vpwr vgnd scs8hd_fill_2
XFILLER_20_180 vgnd vpwr scs8hd_decap_8
XFILLER_20_191 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_180 vgnd vpwr scs8hd_fill_1
XANTENNA__144__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_173 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_1_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__054__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_21 vpwr vgnd scs8hd_fill_2
XFILLER_4_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__049__A enable vgnd vpwr scs8hd_diode_2
XFILLER_14_209 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_SLEEPB _066_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_091_ _091_/A _091_/B _091_/C _091_/D _093_/B vgnd vpwr scs8hd_or4_4
XFILLER_24_55 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__152__A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _136_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__062__A _062_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_208 vpwr vgnd scs8hd_fill_2
XFILLER_27_153 vpwr vgnd scs8hd_fill_2
XFILLER_19_77 vgnd vpwr scs8hd_decap_8
XFILLER_27_164 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_074_ _090_/A _071_/B _074_/Y vgnd vpwr scs8hd_nor2_4
X_143_ chanx_right_in[7] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_120 vpwr vgnd scs8hd_fill_2
XFILLER_18_197 vgnd vpwr scs8hd_decap_12
XANTENNA__147__A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_145 vgnd vpwr scs8hd_decap_8
XFILLER_24_112 vgnd vpwr scs8hd_decap_4
XANTENNA__057__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_23 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_123 vgnd vpwr scs8hd_decap_4
XFILLER_30_115 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_5.LATCH_3_.latch/Q mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_057_ address[1] _048_/Y address[0] _086_/A vgnd vpwr scs8hd_or3_4
XFILLER_7_69 vpwr vgnd scs8hd_fill_2
X_126_ _086_/A _127_/B _126_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ _046_/Y mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_119 vgnd vpwr scs8hd_decap_6
XFILLER_16_67 vpwr vgnd scs8hd_fill_2
X_109_ _124_/B _108_/B address[0] _109_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__054__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_27_11 vgnd vpwr scs8hd_fill_1
XANTENNA__070__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_77 vpwr vgnd scs8hd_fill_2
XFILLER_4_26 vgnd vpwr scs8hd_decap_3
XANTENNA__155__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__065__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_136 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_0_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XFILLER_5_91 vpwr vgnd scs8hd_fill_2
XFILLER_24_23 vgnd vpwr scs8hd_decap_8
X_090_ _090_/A _088_/B _090_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_89 vgnd vpwr scs8hd_decap_3
XFILLER_6_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__062__B _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_176 vgnd vpwr scs8hd_decap_6
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_23 vgnd vpwr scs8hd_decap_4
XFILLER_19_45 vpwr vgnd scs8hd_fill_2
XFILLER_19_56 vgnd vpwr scs8hd_decap_3
X_142_ chanx_right_in[8] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
X_073_ _089_/A _071_/B _073_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_1_.latch/Q mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_143 vgnd vpwr scs8hd_decap_4
XANTENNA__057__B _048_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_46 vpwr vgnd scs8hd_fill_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XFILLER_15_102 vpwr vgnd scs8hd_fill_2
XFILLER_15_113 vgnd vpwr scs8hd_decap_4
XFILLER_30_127 vgnd vpwr scs8hd_decap_12
X_125_ _056_/A _127_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_7 vpwr vgnd scs8hd_fill_2
X_056_ _056_/A _062_/A _056_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__158__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_21_149 vpwr vgnd scs8hd_fill_2
XANTENNA__068__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_127 vgnd vpwr scs8hd_fill_1
XFILLER_12_149 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.LATCH_2_.latch data_in mem_bottom_ipin_1.LATCH_2_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_108_ _124_/B _108_/B _108_/C _108_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_11_193 vpwr vgnd scs8hd_fill_2
XANTENNA__070__B _071_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_3.LATCH_5_.latch data_in mem_bottom_ipin_3.LATCH_5_.latch/Q _056_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_49 vpwr vgnd scs8hd_fill_2
XFILLER_4_16 vpwr vgnd scs8hd_fill_2
XFILLER_31_211 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__065__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_0_.latch/Q mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__081__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_115 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_204 vgnd vpwr scs8hd_decap_8
XFILLER_0_181 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__076__A _091_/D vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_4.LATCH_3_.latch/Q mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _044_/Y mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _137_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_59 vgnd vpwr scs8hd_decap_3
X_141_ _141_/HI _141_/LO vgnd vpwr scs8hd_conb_1
X_072_ _088_/A _071_/B _072_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _140_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_125 vgnd vpwr scs8hd_decap_6
XFILLER_2_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__057__C address[0] vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__B _071_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_139 vgnd vpwr scs8hd_decap_12
X_124_ _055_/D _124_/B _127_/B vgnd vpwr scs8hd_or2_4
X_055_ _091_/A _091_/B _091_/C _055_/D _062_/A vgnd vpwr scs8hd_or4_4
XFILLER_23_191 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_SLEEPB _072_/Y vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_1_.latch data_in mem_bottom_ipin_4.LATCH_1_.latch/Q _073_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_180 vgnd vpwr scs8hd_decap_4
XFILLER_21_106 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__068__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_12_106 vpwr vgnd scs8hd_fill_2
XFILLER_16_25 vpwr vgnd scs8hd_fill_2
XFILLER_16_36 vgnd vpwr scs8hd_decap_3
XANTENNA__084__A _091_/D vgnd vpwr scs8hd_diode_2
X_107_ _117_/B _108_/B address[0] _107_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_7_187 vpwr vgnd scs8hd_fill_2
XFILLER_7_198 vpwr vgnd scs8hd_fill_2
XFILLER_11_172 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_6.LATCH_4_.latch data_in mem_bottom_ipin_6.LATCH_4_.latch/Q _086_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_46 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_146 vgnd vpwr scs8hd_decap_4
XFILLER_4_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _045_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__081__B _081_/B vgnd vpwr scs8hd_diode_2
XANTENNA__065__C address[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_1_.latch/Q mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_60 vgnd vpwr scs8hd_fill_1
XFILLER_24_47 vgnd vpwr scs8hd_decap_8
XANTENNA__076__B _117_/B vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _056_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_80 vgnd vpwr scs8hd_decap_4
XFILLER_10_16 vpwr vgnd scs8hd_fill_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_27_112 vgnd vpwr scs8hd_decap_4
XANTENNA__087__A _127_/A vgnd vpwr scs8hd_diode_2
X_140_ _140_/HI _140_/LO vgnd vpwr scs8hd_conb_1
X_071_ _127_/A _071_/B _071_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_167 vgnd vpwr scs8hd_decap_4
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_7.LATCH_0_.latch data_in mem_bottom_ipin_7.LATCH_0_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_148 vpwr vgnd scs8hd_fill_2
XFILLER_23_170 vpwr vgnd scs8hd_fill_2
X_054_ address[5] address[6] _055_/D vgnd vpwr scs8hd_or2_4
X_123_ _090_/A _123_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_7 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_0_.latch/Q mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA__068__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__084__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
X_106_ _117_/B _108_/B _108_/C _106_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_7_155 vpwr vgnd scs8hd_fill_2
XFILLER_7_177 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_80 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_60 vpwr vgnd scs8hd_fill_2
XFILLER_8_82 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_3.LATCH_3_.latch/Q mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_25 vpwr vgnd scs8hd_fill_2
XANTENNA__079__B _081_/B vgnd vpwr scs8hd_diode_2
XANTENNA__095__A _088_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_13_49 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_0_ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_72 vpwr vgnd scs8hd_fill_2
XANTENNA__092__B _093_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_7.LATCH_4_.latch/Q mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _138_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_157 vgnd vpwr scs8hd_decap_4
XANTENNA__087__B _088_/B vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_1_.latch data_in mem_top_ipin_0.LATCH_1_.latch/Q _104_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_070_ _086_/A _071_/B _070_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XFILLER_18_113 vgnd vpwr scs8hd_decap_4
XFILLER_18_124 vpwr vgnd scs8hd_fill_2
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _141_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XFILLER_21_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__098__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_30_108 vgnd vpwr scs8hd_decap_4
XFILLER_7_18 vpwr vgnd scs8hd_fill_2
XFILLER_23_182 vgnd vpwr scs8hd_fill_1
X_053_ address[1] _048_/Y _108_/C _056_/A vgnd vpwr scs8hd_or3_4
X_122_ _089_/A _123_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_71 vgnd vpwr scs8hd_decap_4
XFILLER_11_93 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_1_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_208 vgnd vpwr scs8hd_decap_4
XANTENNA__068__D _091_/D vgnd vpwr scs8hd_diode_2
XFILLER_12_119 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_163 vgnd vpwr scs8hd_decap_8
X_105_ _090_/A _102_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_112 vgnd vpwr scs8hd_decap_4
XFILLER_7_134 vpwr vgnd scs8hd_fill_2
XFILLER_21_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_1_.latch data_in mem_bottom_ipin_0.LATCH_1_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__095__B _093_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_211 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_2.LATCH_4_.latch data_in mem_bottom_ipin_2.LATCH_4_.latch/Q _126_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_17 vpwr vgnd scs8hd_fill_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_2_.latch/Q mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_3
XFILLER_6_7 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_0_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_136 vgnd vpwr scs8hd_decap_6
XFILLER_19_27 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_70 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_2.LATCH_3_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_52 vpwr vgnd scs8hd_fill_2
XFILLER_17_191 vpwr vgnd scs8hd_fill_2
XANTENNA__098__B _098_/B vgnd vpwr scs8hd_diode_2
X_121_ _088_/A _123_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_50 vgnd vpwr scs8hd_decap_4
X_052_ address[3] _091_/C vgnd vpwr scs8hd_inv_8
XANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_SLEEPB _056_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _046_/Y vgnd vpwr
+ scs8hd_diode_2
X_104_ _089_/A _102_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_168 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_142 vpwr vgnd scs8hd_fill_2
XFILLER_11_197 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_3.LATCH_0_.latch data_in mem_bottom_ipin_3.LATCH_0_.latch/Q _066_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_93 vgnd vpwr scs8hd_decap_4
XFILLER_14_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_6.LATCH_4_.latch/Q mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_38 vpwr vgnd scs8hd_fill_2
XFILLER_4_138 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_5.LATCH_3_.latch data_in mem_bottom_ipin_5.LATCH_3_.latch/Q _079_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_93 vgnd vpwr scs8hd_fill_1
XFILLER_3_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_29 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _139_/HI mem_top_ipin_0.LATCH_5_.latch/Q
+ mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_204 vpwr vgnd scs8hd_fill_2
XFILLER_0_196 vgnd vpwr scs8hd_decap_12
XFILLER_5_52 vpwr vgnd scs8hd_fill_2
XFILLER_5_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_26_181 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_71 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_129 vpwr vgnd scs8hd_fill_2
XFILLER_23_140 vgnd vpwr scs8hd_decap_3
X_051_ address[4] _091_/B vgnd vpwr scs8hd_inv_8
X_120_ _127_/A _123_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_2_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_29 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_121 vgnd vpwr scs8hd_fill_1
XFILLER_20_143 vgnd vpwr scs8hd_decap_8
X_103_ _088_/A _102_/B _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_176 vgnd vpwr scs8hd_decap_4
XFILLER_8_41 vpwr vgnd scs8hd_fill_2
XFILLER_6_180 vgnd vpwr scs8hd_decap_8
XFILLER_6_191 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_0_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_1.LATCH_3_.latch/Q mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_14_84 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__101__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_105 vpwr vgnd scs8hd_fill_2
XFILLER_18_149 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_193 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_5.LATCH_4_.latch/Q mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_119 vgnd vpwr scs8hd_decap_3
XFILLER_23_174 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_050_ address[6] _098_/B vgnd vpwr scs8hd_inv_8
XFILLER_2_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_163 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_155 vpwr vgnd scs8hd_fill_2
X_102_ _127_/A _102_/B _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_73 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_64 vgnd vpwr scs8hd_decap_3
XFILLER_8_86 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_1_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_62 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XANTENNA__104__A _089_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
XFILLER_5_21 vgnd vpwr scs8hd_fill_1
XFILLER_8_210 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.LATCH_3_.latch data_in mem_bottom_ipin_1.LATCH_3_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_209 vgnd vpwr scs8hd_decap_3
XFILLER_5_202 vpwr vgnd scs8hd_fill_2
XFILLER_14_41 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_2_.latch/Q mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__101__B _102_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_73 vpwr vgnd scs8hd_fill_2
XFILLER_25_51 vgnd vpwr scs8hd_decap_4
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_2_22 vgnd vpwr scs8hd_decap_4
XANTENNA__112__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_0_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_75 vgnd vpwr scs8hd_fill_1
XFILLER_11_97 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__107__A _117_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_186 vpwr vgnd scs8hd_fill_2
XFILLER_14_197 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_0.LATCH_3_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_101_ _086_/A _102_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_105 vgnd vpwr scs8hd_decap_4
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
XFILLER_11_101 vgnd vpwr scs8hd_fill_1
XFILLER_11_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_1_.latch/Q mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_74 vpwr vgnd scs8hd_fill_2
XFILLER_17_85 vpwr vgnd scs8hd_fill_2
XFILLER_17_96 vpwr vgnd scs8hd_fill_2
XFILLER_3_174 vpwr vgnd scs8hd_fill_2
XFILLER_3_163 vpwr vgnd scs8hd_fill_2
XFILLER_3_130 vgnd vpwr scs8hd_decap_3
XANTENNA__104__B _102_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_SLEEPB _081_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _127_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_2_.latch data_in mem_bottom_ipin_4.LATCH_2_.latch/Q _072_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_4.LATCH_4_.latch/Q mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_144 vgnd vpwr scs8hd_decap_4
XFILLER_0_111 vgnd vpwr scs8hd_fill_1
XFILLER_28_84 vpwr vgnd scs8hd_fill_2
XFILLER_28_73 vpwr vgnd scs8hd_fill_2
XFILLER_0_177 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A _089_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_6.LATCH_5_.latch data_in mem_bottom_ipin_6.LATCH_5_.latch/Q _085_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
XFILLER_14_64 vpwr vgnd scs8hd_fill_2
XFILLER_30_96 vgnd vpwr scs8hd_decap_12
XFILLER_29_170 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_27_107 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _045_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_85 vpwr vgnd scs8hd_fill_2
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_67 vpwr vgnd scs8hd_fill_2
XFILLER_2_56 vpwr vgnd scs8hd_fill_2
XFILLER_2_12 vgnd vpwr scs8hd_fill_1
XANTENNA__112__B _111_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_162 vpwr vgnd scs8hd_fill_2
XFILLER_17_173 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_SLEEPB _062_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
XFILLER_23_154 vpwr vgnd scs8hd_fill_2
XFILLER_23_187 vpwr vgnd scs8hd_fill_2
XFILLER_11_54 vgnd vpwr scs8hd_fill_1
XFILLER_14_121 vpwr vgnd scs8hd_fill_2
XANTENNA__107__B _108_/B vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_113 vgnd vpwr scs8hd_decap_8
XFILLER_20_124 vpwr vgnd scs8hd_fill_2
X_100_ _056_/A _102_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_113 vpwr vgnd scs8hd_fill_2
XFILLER_22_86 vgnd vpwr scs8hd_decap_6
XFILLER_19_202 vpwr vgnd scs8hd_fill_2
XFILLER_8_22 vpwr vgnd scs8hd_fill_2
XANTENNA__118__A _056_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_150 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_2_.latch/Q mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_3_197 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_7.LATCH_1_.latch data_in mem_bottom_ipin_7.LATCH_1_.latch/Q _096_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__120__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_13_208 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_41 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_56 vpwr vgnd scs8hd_fill_2
XANTENNA__115__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_10 vpwr vgnd scs8hd_fill_2
XFILLER_14_87 vgnd vpwr scs8hd_decap_3
XFILLER_30_42 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_160 vpwr vgnd scs8hd_fill_2
XANTENNA__126__A _086_/A vgnd vpwr scs8hd_diode_2
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_152 vgnd vpwr scs8hd_fill_1
XPHY_64 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_35 vpwr vgnd scs8hd_fill_2
XFILLER_17_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_1_.latch/Q mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_166 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_33 vpwr vgnd scs8hd_fill_2
XFILLER_14_133 vgnd vpwr scs8hd_fill_1
XANTENNA__107__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__123__B _123_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_3.LATCH_4_.latch/Q mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
XFILLER_22_43 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vgnd vpwr scs8hd_decap_3
Xmem_top_ipin_0.LATCH_2_.latch data_in mem_top_ipin_0.LATCH_2_.latch/Q _103_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_45 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
X_159_ chanx_left_in[0] chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_8_78 vpwr vgnd scs8hd_fill_2
XFILLER_10_180 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__044__A _044_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_54 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_209 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _138_/HI mem_bottom_ipin_7.LATCH_5_.latch/Q
+ mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_28_64 vgnd vpwr scs8hd_decap_3
XFILLER_8_202 vgnd vpwr scs8hd_decap_8
XFILLER_5_68 vpwr vgnd scs8hd_fill_2
XFILLER_5_13 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_76 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_2_.latch data_in mem_bottom_ipin_0.LATCH_2_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_150 vgnd vpwr scs8hd_decap_6
XANTENNA__126__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA__142__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__052__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_18_109 vpwr vgnd scs8hd_fill_2
XFILLER_26_142 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_2.LATCH_5_.latch data_in mem_bottom_ipin_2.LATCH_5_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_32 vpwr vgnd scs8hd_fill_2
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_65 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_2_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__047__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_12 vpwr vgnd scs8hd_fill_2
XFILLER_2_7 vgnd vpwr scs8hd_decap_3
XFILLER_11_78 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vpwr vgnd scs8hd_fill_2
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_0_.latch/Q mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_159 vpwr vgnd scs8hd_fill_2
XFILLER_22_22 vpwr vgnd scs8hd_fill_2
XFILLER_22_55 vgnd vpwr scs8hd_decap_3
XFILLER_22_99 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_089_ _089_/A _088_/B _089_/Y vgnd vpwr scs8hd_nor2_4
X_158_ chanx_left_in[1] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_6_163 vpwr vgnd scs8hd_fill_2
XFILLER_26_3 vpwr vgnd scs8hd_fill_2
XANTENNA__150__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_12_ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__060__A _062_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_11 vpwr vgnd scs8hd_fill_2
XFILLER_30_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_SLEEPB _070_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _127_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__145__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_80 vgnd vpwr scs8hd_fill_1
XANTENNA__055__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_210 vpwr vgnd scs8hd_fill_2
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_0_169 vgnd vpwr scs8hd_decap_4
XFILLER_0_125 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_1_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_210 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_3.LATCH_1_.latch data_in mem_bottom_ipin_3.LATCH_1_.latch/Q _064_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_30_22 vgnd vpwr scs8hd_decap_8
XFILLER_5_206 vgnd vpwr scs8hd_decap_6
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_45 vpwr vgnd scs8hd_fill_2
XFILLER_30_88 vgnd vpwr scs8hd_decap_4
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_2.LATCH_4_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_ipin_5.LATCH_4_.latch data_in mem_bottom_ipin_5.LATCH_4_.latch/Q _078_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_209 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_25_77 vpwr vgnd scs8hd_fill_2
XFILLER_25_11 vpwr vgnd scs8hd_fill_2
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_66 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_2_26 vgnd vpwr scs8hd_fill_1
XFILLER_17_187 vpwr vgnd scs8hd_fill_2
XANTENNA__153__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_113 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__063__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_46 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__148__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _137_/HI mem_bottom_ipin_6.LATCH_5_.latch/Q
+ mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_9_150 vpwr vgnd scs8hd_fill_2
XANTENNA__058__A _062_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_109 vgnd vpwr scs8hd_fill_1
XFILLER_11_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_157_ chanx_left_in[2] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_8_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_088_ _088_/A _088_/B _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__060__B _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_34 vpwr vgnd scs8hd_fill_2
XFILLER_17_45 vpwr vgnd scs8hd_fill_2
XFILLER_17_78 vpwr vgnd scs8hd_fill_2
XFILLER_17_89 vgnd vpwr scs8hd_decap_4
XFILLER_3_178 vgnd vpwr scs8hd_decap_3
XFILLER_3_167 vpwr vgnd scs8hd_fill_2
XFILLER_3_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__055__B _091_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_90 vgnd vpwr scs8hd_decap_3
XANTENNA__071__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_88 vgnd vpwr scs8hd_decap_4
XFILLER_0_148 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_6.LATCH_0_.latch data_in mem_bottom_ipin_6.LATCH_0_.latch/Q _090_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_37 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__156__A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__066__A _062_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_68 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_199 vgnd vpwr scs8hd_decap_12
XFILLER_25_89 vpwr vgnd scs8hd_fill_2
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_67 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_111 vgnd vpwr scs8hd_decap_6
XFILLER_17_166 vpwr vgnd scs8hd_fill_2
XFILLER_17_177 vpwr vgnd scs8hd_fill_2
XFILLER_17_199 vpwr vgnd scs8hd_fill_2
XFILLER_23_136 vpwr vgnd scs8hd_fill_2
XFILLER_23_158 vpwr vgnd scs8hd_fill_2
XFILLER_31_180 vgnd vpwr scs8hd_decap_6
XANTENNA__063__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_14_125 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_206 vgnd vpwr scs8hd_decap_6
XANTENNA__058__B _086_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_1_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _044_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_117 vgnd vpwr scs8hd_decap_3
XANTENNA__074__A _090_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_206 vgnd vpwr scs8hd_decap_6
X_156_ chanx_left_in[3] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
X_087_ _127_/A _088_/B _087_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_26 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_25_209 vgnd vpwr scs8hd_decap_3
XANTENNA__159__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _056_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_1.LATCH_4_.latch/Q mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_146 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
X_139_ _139_/HI _139_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__055__C _091_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XANTENNA__071__B _071_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_45 vgnd vpwr scs8hd_decap_4
XFILLER_28_23 vpwr vgnd scs8hd_fill_2
XFILLER_28_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _139_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_58 vgnd vpwr scs8hd_decap_4
XANTENNA__066__B _090_/A vgnd vpwr scs8hd_diode_2
XANTENNA__082__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_175 vpwr vgnd scs8hd_fill_2
XFILLER_29_164 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _136_/HI mem_bottom_ipin_5.LATCH_5_.latch/Q
+ mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_123 vpwr vgnd scs8hd_fill_2
XANTENNA__077__A _056_/A vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_68 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_39 vpwr vgnd scs8hd_fill_2
XFILLER_17_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_1.LATCH_4_.latch data_in mem_bottom_ipin_1.LATCH_4_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__063__C _108_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_130 vpwr vgnd scs8hd_fill_2
XFILLER_9_163 vpwr vgnd scs8hd_fill_2
XFILLER_9_174 vpwr vgnd scs8hd_fill_2
XFILLER_3_93 vpwr vgnd scs8hd_fill_2
XANTENNA__074__B _071_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_2_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_69 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A _090_/A vgnd vpwr scs8hd_diode_2
X_086_ _086_/A _088_/B _086_/Y vgnd vpwr scs8hd_nor2_4
X_155_ chanx_left_in[4] chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_6_144 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_0_.latch data_in _046_/A _109_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__069__B _071_/B vgnd vpwr scs8hd_diode_2
XANTENNA__085__A _056_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_210 vpwr vgnd scs8hd_fill_2
XFILLER_17_58 vgnd vpwr scs8hd_decap_3
XFILLER_30_202 vgnd vpwr scs8hd_decap_8
X_138_ _138_/HI _138_/LO vgnd vpwr scs8hd_conb_1
X_069_ _056_/A _071_/B _069_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_180 vgnd vpwr scs8hd_decap_8
XFILLER_24_3 vgnd vpwr scs8hd_decap_3
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_202 vgnd vpwr scs8hd_decap_8
XANTENNA__055__D _055_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_202 vgnd vpwr scs8hd_decap_8
XFILLER_5_17 vgnd vpwr scs8hd_decap_4
XFILLER_30_47 vgnd vpwr scs8hd_decap_3
XANTENNA__082__B _081_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_0_.latch data_in mem_bottom_ipin_2.LATCH_0_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_1_.latch/Q mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_71 vpwr vgnd scs8hd_fill_2
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_157 vgnd vpwr scs8hd_decap_12
XFILLER_26_146 vgnd vpwr scs8hd_decap_6
XFILLER_25_47 vpwr vgnd scs8hd_fill_2
XFILLER_25_36 vpwr vgnd scs8hd_fill_2
XPHY_69 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__077__B _081_/B vgnd vpwr scs8hd_diode_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XANTENNA__093__A _086_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_2_29 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_4.LATCH_3_.latch data_in mem_bottom_ipin_4.LATCH_3_.latch/Q _071_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_0.LATCH_4_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_16 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A _088_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_149 vpwr vgnd scs8hd_fill_2
XFILLER_13_160 vpwr vgnd scs8hd_fill_2
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_9_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_2_.latch/Q mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_26 vgnd vpwr scs8hd_decap_3
XANTENNA__090__B _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_8 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_141 vgnd vpwr scs8hd_decap_4
XFILLER_10_152 vgnd vpwr scs8hd_fill_1
X_085_ _056_/A _088_/B _085_/Y vgnd vpwr scs8hd_nor2_4
X_154_ chanx_left_in[5] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_6_123 vgnd vpwr scs8hd_fill_1
XFILLER_6_167 vgnd vpwr scs8hd_decap_4
XFILLER_10_163 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_SLEEPB _073_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_15 vpwr vgnd scs8hd_fill_2
XANTENNA__085__B _088_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _135_/HI mem_bottom_ipin_4.LATCH_5_.latch/Q
+ mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_137_ _137_/HI _137_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
X_068_ _091_/A address[4] address[3] _091_/D _071_/B vgnd vpwr scs8hd_or4_4
XFILLER_9_71 vpwr vgnd scs8hd_fill_2
XFILLER_0_107 vpwr vgnd scs8hd_fill_2
XFILLER_0_129 vpwr vgnd scs8hd_fill_2
XFILLER_28_69 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XFILLER_30_59 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_50 vpwr vgnd scs8hd_fill_2
XFILLER_6_61 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_7.LATCH_2_.latch data_in mem_bottom_ipin_7.LATCH_2_.latch/Q _095_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_169 vgnd vpwr scs8hd_decap_12
XFILLER_25_15 vpwr vgnd scs8hd_fill_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _093_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_180 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_80 vpwr vgnd scs8hd_fill_2
XFILLER_9_121 vgnd vpwr scs8hd_fill_1
XFILLER_3_40 vpwr vgnd scs8hd_fill_2
XFILLER_3_73 vgnd vpwr scs8hd_decap_3
XANTENNA__099__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
X_153_ chanx_left_in[6] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_102 vpwr vgnd scs8hd_fill_2
XFILLER_6_113 vpwr vgnd scs8hd_fill_2
XFILLER_6_135 vpwr vgnd scs8hd_fill_2
XFILLER_8_18 vpwr vgnd scs8hd_fill_2
XFILLER_10_120 vgnd vpwr scs8hd_decap_6
X_084_ _091_/D _124_/B _088_/B vgnd vpwr scs8hd_or2_4
XFILLER_10_197 vgnd vpwr scs8hd_decap_12
XFILLER_17_49 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_116 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_136_ _136_/HI _136_/LO vgnd vpwr scs8hd_conb_1
XFILLER_31_6 vpwr vgnd scs8hd_fill_2
X_067_ address[5] _098_/B _091_/D vgnd vpwr scs8hd_nand2_4
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_59 vgnd vpwr scs8hd_decap_3
XANTENNA__096__B _093_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_119_ _086_/A _123_/B _119_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_ipin_0.LATCH_3_.latch data_in mem_top_ipin_0.LATCH_3_.latch/Q _102_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_38 vgnd vpwr scs8hd_fill_1
XFILLER_29_134 vpwr vgnd scs8hd_fill_2
XFILLER_29_123 vgnd vpwr scs8hd_decap_6
XFILLER_4_211 vgnd vpwr scs8hd_fill_1
XFILLER_20_60 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_2_.latch/Q mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XFILLER_26_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _043_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_17_126 vpwr vgnd scs8hd_fill_2
XFILLER_25_192 vgnd vpwr scs8hd_decap_3
XFILLER_25_170 vgnd vpwr scs8hd_decap_12
XFILLER_31_81 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _134_/HI mem_bottom_ipin_3.LATCH_5_.latch/Q
+ mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_16_192 vgnd vpwr scs8hd_decap_3
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_11_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_13_173 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_0.LATCH_3_.latch data_in mem_bottom_ipin_0.LATCH_3_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__099__B address[4] vgnd vpwr scs8hd_diode_2
X_152_ chanx_left_in[7] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
X_083_ _091_/A _091_/B address[3] _124_/B vgnd vpwr scs8hd_or3_4
XFILLER_12_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_8 vpwr vgnd scs8hd_fill_2
XFILLER_5_191 vpwr vgnd scs8hd_fill_2
XFILLER_17_28 vgnd vpwr scs8hd_decap_4
XFILLER_3_106 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_135_ _135_/HI _135_/LO vgnd vpwr scs8hd_conb_1
X_066_ _062_/A _090_/A _066_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_93 vgnd vpwr scs8hd_decap_4
XFILLER_28_49 vgnd vpwr scs8hd_fill_1
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_16 vpwr vgnd scs8hd_fill_2
XFILLER_18_71 vpwr vgnd scs8hd_fill_2
XFILLER_18_93 vgnd vpwr scs8hd_fill_1
X_049_ enable _091_/A vgnd vpwr scs8hd_inv_8
X_118_ _056_/A _123_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_127 vgnd vpwr scs8hd_decap_4
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_25_28 vpwr vgnd scs8hd_fill_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_1_204 vgnd vpwr scs8hd_decap_8
XFILLER_25_182 vgnd vpwr scs8hd_fill_1
XFILLER_17_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_14_108 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_1_.latch/Q mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_ipin_3.LATCH_2_.latch data_in mem_bottom_ipin_3.LATCH_2_.latch/Q _062_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_163 vgnd vpwr scs8hd_decap_8
XFILLER_22_174 vgnd vpwr scs8hd_decap_8
XFILLER_22_185 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_9_112 vgnd vpwr scs8hd_fill_1
XFILLER_9_134 vgnd vpwr scs8hd_decap_3
XFILLER_9_167 vpwr vgnd scs8hd_fill_2
XFILLER_9_178 vgnd vpwr scs8hd_decap_3
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_5.LATCH_5_.latch data_in mem_bottom_ipin_5.LATCH_5_.latch/Q _077_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__099__C address[3] vgnd vpwr scs8hd_diode_2
X_082_ _090_/A _081_/B _082_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
X_151_ chanx_left_in[8] chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_5_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_SLEEPB _058_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_2_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_134_ _134_/HI _134_/LO vgnd vpwr scs8hd_conb_1
X_065_ address[1] address[2] address[0] _090_/A vgnd vpwr scs8hd_or3_4
XFILLER_0_21 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_fill_1
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_76 vpwr vgnd scs8hd_fill_2
XFILLER_9_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _133_/HI mem_bottom_ipin_2.LATCH_5_.latch/Q
+ mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_117_ _055_/D _117_/B _123_/B vgnd vpwr scs8hd_or2_4
X_048_ address[2] _048_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_18 vpwr vgnd scs8hd_fill_2
XFILLER_29_114 vgnd vpwr scs8hd_decap_8
XFILLER_29_71 vpwr vgnd scs8hd_fill_2
XFILLER_6_20 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_19_191 vpwr vgnd scs8hd_fill_2
XFILLER_15_40 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _127_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_6.LATCH_1_.latch data_in mem_bottom_ipin_6.LATCH_1_.latch/Q _089_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_142 vgnd vpwr scs8hd_decap_3
XFILLER_22_197 vgnd vpwr scs8hd_decap_12
XFILLER_9_146 vpwr vgnd scs8hd_fill_2
XFILLER_13_197 vgnd vpwr scs8hd_decap_4
XANTENNA__099__D _108_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_112 vgnd vpwr scs8hd_fill_1
X_150_ chanx_right_in[0] chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_081_ _089_/A _081_/B _081_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_145 vgnd vpwr scs8hd_fill_1
XFILLER_10_167 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_204 vgnd vpwr scs8hd_decap_8
X_133_ _133_/HI _133_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_62 vgnd vpwr scs8hd_decap_3
XFILLER_2_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_064_ _062_/A _089_/A _064_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__110__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XFILLER_24_8 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
XFILLER_9_86 vpwr vgnd scs8hd_fill_2
XFILLER_18_84 vgnd vpwr scs8hd_decap_4
XANTENNA__105__A _090_/A vgnd vpwr scs8hd_diode_2
X_116_ _090_/A _111_/B _116_/Y vgnd vpwr scs8hd_nor2_4
X_047_ address[1] _059_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _044_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_203 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_74 vgnd vpwr scs8hd_decap_12
XFILLER_20_96 vgnd vpwr scs8hd_decap_8
XFILLER_29_83 vgnd vpwr scs8hd_fill_1
XFILLER_28_170 vgnd vpwr scs8hd_decap_12
XFILLER_6_32 vpwr vgnd scs8hd_fill_2
XFILLER_6_54 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_19_170 vgnd vpwr scs8hd_fill_1
XFILLER_17_107 vpwr vgnd scs8hd_fill_2
XFILLER_25_184 vgnd vpwr scs8hd_decap_8
XFILLER_15_96 vgnd vpwr scs8hd_decap_4
XANTENNA__102__B _102_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_187 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_2_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_6
XFILLER_13_143 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _127_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_180 vgnd vpwr scs8hd_decap_8
XFILLER_8_191 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _132_/HI mem_bottom_ipin_1.LATCH_5_.latch/Q
+ mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_080_ _088_/A _081_/B _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_106 vpwr vgnd scs8hd_fill_2
XFILLER_6_117 vgnd vpwr scs8hd_decap_6
XFILLER_5_3 vgnd vpwr scs8hd_fill_1
XFILLER_6_139 vgnd vpwr scs8hd_decap_3
XFILLER_12_42 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
X_132_ _132_/HI _132_/LO vgnd vpwr scs8hd_conb_1
X_063_ address[1] address[2] _108_/C _089_/A vgnd vpwr scs8hd_or3_4
Xmem_bottom_ipin_1.LATCH_5_.latch data_in mem_bottom_ipin_1.LATCH_5_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_41 vpwr vgnd scs8hd_fill_2
XFILLER_23_52 vpwr vgnd scs8hd_fill_2
XFILLER_2_197 vgnd vpwr scs8hd_decap_12
XFILLER_2_131 vgnd vpwr scs8hd_decap_3
XANTENNA__110__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_41 vpwr vgnd scs8hd_fill_2
XANTENNA__105__B _102_/B vgnd vpwr scs8hd_diode_2
X_115_ _089_/A _111_/B _115_/Y vgnd vpwr scs8hd_nor2_4
X_046_ _046_/A _046_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__121__A _088_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_138 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_2.LATCH_1_.latch data_in _045_/A _108_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_64 vgnd vpwr scs8hd_fill_1
XFILLER_20_86 vgnd vpwr scs8hd_decap_6
XFILLER_29_95 vpwr vgnd scs8hd_fill_2
XFILLER_28_182 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_66 vgnd vpwr scs8hd_decap_3
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_26_108 vgnd vpwr scs8hd_decap_6
XFILLER_20_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_17_119 vgnd vpwr scs8hd_decap_3
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_130 vpwr vgnd scs8hd_fill_2
XFILLER_16_163 vgnd vpwr scs8hd_decap_8
XFILLER_31_199 vgnd vpwr scs8hd_decap_12
.ends

