magic
tech sky130A
magscale 1 2
timestamp 1606224408
<< locali >>
rect 5733 4063 5767 4233
rect 9689 3519 9723 3689
<< viali >>
rect 3893 14025 3927 14059
rect 5365 14025 5399 14059
rect 9229 14025 9263 14059
rect 4629 13957 4663 13991
rect 7205 13957 7239 13991
rect 3709 13821 3743 13855
rect 4445 13821 4479 13855
rect 5181 13821 5215 13855
rect 7021 13821 7055 13855
rect 9045 13821 9079 13855
rect 5610 11237 5644 11271
rect 5365 11101 5399 11135
rect 6745 10965 6779 10999
rect 8309 10625 8343 10659
rect 8401 10625 8435 10659
rect 9321 10625 9355 10659
rect 8217 10557 8251 10591
rect 9045 10489 9079 10523
rect 7849 10421 7883 10455
rect 8677 10421 8711 10455
rect 9137 10421 9171 10455
rect 11253 10217 11287 10251
rect 6745 10149 6779 10183
rect 5181 10081 5215 10115
rect 6653 10081 6687 10115
rect 7665 10081 7699 10115
rect 10129 10081 10163 10115
rect 6837 10013 6871 10047
rect 9873 10013 9907 10047
rect 8953 9945 8987 9979
rect 4997 9877 5031 9911
rect 6285 9877 6319 9911
rect 5917 9605 5951 9639
rect 11345 9605 11379 9639
rect 6561 9537 6595 9571
rect 7757 9537 7791 9571
rect 7941 9537 7975 9571
rect 10885 9537 10919 9571
rect 8677 9469 8711 9503
rect 11529 9469 11563 9503
rect 8922 9401 8956 9435
rect 6285 9333 6319 9367
rect 6377 9333 6411 9367
rect 7297 9333 7331 9367
rect 7665 9333 7699 9367
rect 10057 9333 10091 9367
rect 10333 9333 10367 9367
rect 10701 9333 10735 9367
rect 10793 9333 10827 9367
rect 6745 9129 6779 9163
rect 9137 9129 9171 9163
rect 9689 9129 9723 9163
rect 10149 9129 10183 9163
rect 10701 9129 10735 9163
rect 7205 9061 7239 9095
rect 10057 9061 10091 9095
rect 7113 8993 7147 9027
rect 8013 8993 8047 9027
rect 11069 8993 11103 9027
rect 7297 8925 7331 8959
rect 7757 8925 7791 8959
rect 10241 8925 10275 8959
rect 11161 8925 11195 8959
rect 11253 8925 11287 8959
rect 8401 8585 8435 8619
rect 8861 8449 8895 8483
rect 9045 8449 9079 8483
rect 10425 8449 10459 8483
rect 8769 8313 8803 8347
rect 4077 6817 4111 6851
rect 4261 6749 4295 6783
rect 6837 4777 6871 4811
rect 7389 4777 7423 4811
rect 5181 4641 5215 4675
rect 6653 4641 6687 4675
rect 7205 4641 7239 4675
rect 7757 4641 7791 4675
rect 8309 4641 8343 4675
rect 8953 4641 8987 4675
rect 9689 4641 9723 4675
rect 10241 4641 10275 4675
rect 11897 4641 11931 4675
rect 7941 4505 7975 4539
rect 8493 4505 8527 4539
rect 5365 4437 5399 4471
rect 9137 4437 9171 4471
rect 9873 4437 9907 4471
rect 10425 4437 10459 4471
rect 12081 4437 12115 4471
rect 5733 4233 5767 4267
rect 7021 4165 7055 4199
rect 3709 4029 3743 4063
rect 4721 4029 4755 4063
rect 5273 4029 5307 4063
rect 5733 4029 5767 4063
rect 5825 4029 5859 4063
rect 6837 4029 6871 4063
rect 7665 4029 7699 4063
rect 8217 4029 8251 4063
rect 8953 4029 8987 4063
rect 9505 4029 9539 4063
rect 10057 4029 10091 4063
rect 10609 4029 10643 4063
rect 11529 4029 11563 4063
rect 12449 4029 12483 4063
rect 13001 4029 13035 4063
rect 3893 3893 3927 3927
rect 4905 3893 4939 3927
rect 5457 3893 5491 3927
rect 6009 3893 6043 3927
rect 7849 3893 7883 3927
rect 8401 3893 8435 3927
rect 9137 3893 9171 3927
rect 9689 3893 9723 3927
rect 10241 3893 10275 3927
rect 10793 3893 10827 3927
rect 11713 3893 11747 3927
rect 12633 3893 12667 3927
rect 13185 3893 13219 3927
rect 5733 3689 5767 3723
rect 7573 3689 7607 3723
rect 8125 3689 8159 3723
rect 9137 3689 9171 3723
rect 9689 3689 9723 3723
rect 9965 3689 9999 3723
rect 4721 3553 4755 3587
rect 5549 3553 5583 3587
rect 6285 3553 6319 3587
rect 6837 3553 6871 3587
rect 7389 3553 7423 3587
rect 7941 3553 7975 3587
rect 8953 3553 8987 3587
rect 9781 3553 9815 3587
rect 10609 3553 10643 3587
rect 11529 3553 11563 3587
rect 12357 3553 12391 3587
rect 9689 3485 9723 3519
rect 4905 3417 4939 3451
rect 10793 3417 10827 3451
rect 12541 3417 12575 3451
rect 6469 3349 6503 3383
rect 7021 3349 7055 3383
rect 11713 3349 11747 3383
rect 9413 2941 9447 2975
rect 9597 2805 9631 2839
<< metal1 >>
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 3786 15104 3792 15156
rect 3844 15144 3850 15156
rect 3844 15116 4016 15144
rect 3844 15104 3850 15116
rect 566 14968 572 15020
rect 624 15008 630 15020
rect 1302 15008 1308 15020
rect 624 14980 1308 15008
rect 624 14968 630 14980
rect 1302 14968 1308 14980
rect 1360 14968 1366 15020
rect 3988 14952 4016 15116
rect 7098 15104 7104 15156
rect 7156 15144 7162 15156
rect 9490 15144 9496 15156
rect 7156 15116 9496 15144
rect 7156 15104 7162 15116
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 6546 15036 6552 15088
rect 6604 15076 6610 15088
rect 8662 15076 8668 15088
rect 6604 15048 8668 15076
rect 6604 15036 6610 15048
rect 8662 15036 8668 15048
rect 8720 15036 8726 15088
rect 8754 15036 8760 15088
rect 8812 15076 8818 15088
rect 11606 15076 11612 15088
rect 8812 15048 11612 15076
rect 8812 15036 8818 15048
rect 11606 15036 11612 15048
rect 11664 15036 11670 15088
rect 7190 14968 7196 15020
rect 7248 15008 7254 15020
rect 9122 15008 9128 15020
rect 7248 14980 9128 15008
rect 7248 14968 7254 14980
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 3142 14900 3148 14952
rect 3200 14940 3206 14952
rect 3878 14940 3884 14952
rect 3200 14912 3884 14940
rect 3200 14900 3206 14912
rect 3878 14900 3884 14912
rect 3936 14900 3942 14952
rect 3970 14900 3976 14952
rect 4028 14900 4034 14952
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 7742 14940 7748 14952
rect 6972 14912 7748 14940
rect 6972 14900 6978 14912
rect 7742 14900 7748 14912
rect 7800 14900 7806 14952
rect 7926 14900 7932 14952
rect 7984 14940 7990 14952
rect 9950 14940 9956 14952
rect 7984 14912 9956 14940
rect 7984 14900 7990 14912
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 8846 14832 8852 14884
rect 8904 14872 8910 14884
rect 10686 14872 10692 14884
rect 8904 14844 10692 14872
rect 8904 14832 8910 14844
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 5258 14764 5264 14816
rect 5316 14804 5322 14816
rect 9030 14804 9036 14816
rect 5316 14776 9036 14804
rect 5316 14764 5322 14776
rect 9030 14764 9036 14776
rect 9088 14764 9094 14816
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 11698 14600 11704 14612
rect 7432 14572 11704 14600
rect 7432 14560 7438 14572
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 13630 14560 13636 14612
rect 13688 14600 13694 14612
rect 16758 14600 16764 14612
rect 13688 14572 16764 14600
rect 13688 14560 13694 14572
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 6270 14492 6276 14544
rect 6328 14532 6334 14544
rect 10318 14532 10324 14544
rect 6328 14504 10324 14532
rect 6328 14492 6334 14504
rect 10318 14492 10324 14504
rect 10376 14492 10382 14544
rect 4798 14424 4804 14476
rect 4856 14464 4862 14476
rect 8938 14464 8944 14476
rect 4856 14436 8944 14464
rect 4856 14424 4862 14436
rect 8938 14424 8944 14436
rect 8996 14424 9002 14476
rect 9122 14424 9128 14476
rect 9180 14464 9186 14476
rect 11238 14464 11244 14476
rect 9180 14436 11244 14464
rect 9180 14424 9186 14436
rect 11238 14424 11244 14436
rect 11296 14424 11302 14476
rect 13078 14424 13084 14476
rect 13136 14464 13142 14476
rect 15930 14464 15936 14476
rect 13136 14436 15936 14464
rect 13136 14424 13142 14436
rect 15930 14424 15936 14436
rect 15988 14424 15994 14476
rect 5718 14356 5724 14408
rect 5776 14396 5782 14408
rect 9858 14396 9864 14408
rect 5776 14368 9864 14396
rect 5776 14356 5782 14368
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 12066 14396 12072 14408
rect 10336 14368 12072 14396
rect 1854 14288 1860 14340
rect 1912 14328 1918 14340
rect 5350 14328 5356 14340
rect 1912 14300 5356 14328
rect 1912 14288 1918 14300
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 7374 14288 7380 14340
rect 7432 14328 7438 14340
rect 10336 14328 10364 14368
rect 12066 14356 12072 14368
rect 12124 14356 12130 14408
rect 7432 14300 10364 14328
rect 7432 14288 7438 14300
rect 10686 14288 10692 14340
rect 10744 14328 10750 14340
rect 15470 14328 15476 14340
rect 10744 14300 15476 14328
rect 10744 14288 10750 14300
rect 15470 14288 15476 14300
rect 15528 14288 15534 14340
rect 2682 14220 2688 14272
rect 2740 14260 2746 14272
rect 6454 14260 6460 14272
rect 2740 14232 6460 14260
rect 2740 14220 2746 14232
rect 6454 14220 6460 14232
rect 6512 14220 6518 14272
rect 6822 14220 6828 14272
rect 6880 14260 6886 14272
rect 9122 14260 9128 14272
rect 6880 14232 9128 14260
rect 6880 14220 6886 14232
rect 9122 14220 9128 14232
rect 9180 14220 9186 14272
rect 9306 14220 9312 14272
rect 9364 14260 9370 14272
rect 13814 14260 13820 14272
rect 9364 14232 13820 14260
rect 9364 14220 9370 14232
rect 13814 14220 13820 14232
rect 13872 14220 13878 14272
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 198 14016 204 14068
rect 256 14056 262 14068
rect 3881 14059 3939 14065
rect 3881 14056 3893 14059
rect 256 14028 3893 14056
rect 256 14016 262 14028
rect 3881 14025 3893 14028
rect 3927 14025 3939 14059
rect 3881 14019 3939 14025
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 5350 14056 5356 14068
rect 4488 14028 5212 14056
rect 5311 14028 5356 14056
rect 4488 14016 4494 14028
rect 1026 13948 1032 14000
rect 1084 13988 1090 14000
rect 4617 13991 4675 13997
rect 4617 13988 4629 13991
rect 1084 13960 4629 13988
rect 1084 13948 1090 13960
rect 4617 13957 4629 13960
rect 4663 13957 4675 13991
rect 5184 13988 5212 14028
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 7006 14016 7012 14068
rect 7064 14056 7070 14068
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 7064 14028 9229 14056
rect 7064 14016 7070 14028
rect 9217 14025 9229 14028
rect 9263 14025 9275 14059
rect 9217 14019 9275 14025
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 13170 14056 13176 14068
rect 10652 14028 13176 14056
rect 10652 14016 10658 14028
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 7193 13991 7251 13997
rect 7193 13988 7205 13991
rect 5184 13960 7205 13988
rect 4617 13951 4675 13957
rect 7193 13957 7205 13960
rect 7239 13957 7251 13991
rect 7193 13951 7251 13957
rect 8018 13948 8024 14000
rect 8076 13988 8082 14000
rect 10410 13988 10416 14000
rect 8076 13960 10416 13988
rect 8076 13948 8082 13960
rect 10410 13948 10416 13960
rect 10468 13948 10474 14000
rect 11882 13948 11888 14000
rect 11940 13988 11946 14000
rect 16298 13988 16304 14000
rect 11940 13960 16304 13988
rect 11940 13948 11946 13960
rect 16298 13948 16304 13960
rect 16356 13948 16362 14000
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 2682 13920 2688 13932
rect 1452 13892 2688 13920
rect 1452 13880 1458 13892
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 5626 13920 5632 13932
rect 4448 13892 5632 13920
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13852 3755 13855
rect 4338 13852 4344 13864
rect 3743 13824 4344 13852
rect 3743 13821 3755 13824
rect 3697 13815 3755 13821
rect 4338 13812 4344 13824
rect 4396 13812 4402 13864
rect 4448 13861 4476 13892
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 6638 13880 6644 13932
rect 6696 13920 6702 13932
rect 6696 13892 10456 13920
rect 6696 13880 6702 13892
rect 10428 13864 10456 13892
rect 10502 13880 10508 13932
rect 10560 13920 10566 13932
rect 12526 13920 12532 13932
rect 10560 13892 12532 13920
rect 10560 13880 10566 13892
rect 12526 13880 12532 13892
rect 12584 13880 12590 13932
rect 4433 13855 4491 13861
rect 4433 13821 4445 13855
rect 4479 13821 4491 13855
rect 5166 13852 5172 13864
rect 5127 13824 5172 13852
rect 4433 13815 4491 13821
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 6822 13852 6828 13864
rect 6656 13824 6828 13852
rect 6656 13796 6684 13824
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7009 13855 7067 13861
rect 7009 13821 7021 13855
rect 7055 13852 7067 13855
rect 8754 13852 8760 13864
rect 7055 13824 8760 13852
rect 7055 13821 7067 13824
rect 7009 13815 7067 13821
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13852 9091 13855
rect 9766 13852 9772 13864
rect 9079 13824 9772 13852
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 10410 13812 10416 13864
rect 10468 13812 10474 13864
rect 11146 13812 11152 13864
rect 11204 13852 11210 13864
rect 12894 13852 12900 13864
rect 11204 13824 12900 13852
rect 11204 13812 11210 13824
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 6638 13744 6644 13796
rect 6696 13744 6702 13796
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 3510 13200 3516 13252
rect 3568 13240 3574 13252
rect 5534 13240 5540 13252
rect 3568 13212 5540 13240
rect 3568 13200 3574 13212
rect 5534 13200 5540 13212
rect 5592 13200 5598 13252
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 13998 11704 14004 11756
rect 14056 11744 14062 11756
rect 14642 11744 14648 11756
rect 14056 11716 14648 11744
rect 14056 11704 14062 11716
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 13906 11636 13912 11688
rect 13964 11676 13970 11688
rect 15010 11676 15016 11688
rect 13964 11648 15016 11676
rect 13964 11636 13970 11648
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 5534 11228 5540 11280
rect 5592 11277 5598 11280
rect 5592 11271 5656 11277
rect 5592 11237 5610 11271
rect 5644 11237 5656 11271
rect 5592 11231 5656 11237
rect 5592 11228 5598 11231
rect 4982 11092 4988 11144
rect 5040 11132 5046 11144
rect 5353 11135 5411 11141
rect 5353 11132 5365 11135
rect 5040 11104 5365 11132
rect 5040 11092 5046 11104
rect 5353 11101 5365 11104
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 6730 10996 6736 11008
rect 6691 10968 6736 10996
rect 6730 10956 6736 10968
rect 6788 10956 6794 11008
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 5166 10752 5172 10804
rect 5224 10792 5230 10804
rect 7742 10792 7748 10804
rect 5224 10764 7748 10792
rect 5224 10752 5230 10764
rect 7742 10752 7748 10764
rect 7800 10792 7806 10804
rect 7800 10764 8340 10792
rect 7800 10752 7806 10764
rect 7190 10684 7196 10736
rect 7248 10724 7254 10736
rect 7466 10724 7472 10736
rect 7248 10696 7472 10724
rect 7248 10684 7254 10696
rect 7466 10684 7472 10696
rect 7524 10684 7530 10736
rect 8312 10665 8340 10764
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10625 8355 10659
rect 8297 10619 8355 10625
rect 8386 10616 8392 10668
rect 8444 10656 8450 10668
rect 9309 10659 9367 10665
rect 8444 10628 8489 10656
rect 8444 10616 8450 10628
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 12434 10656 12440 10668
rect 9355 10628 12440 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 8128 10560 8217 10588
rect 5166 10480 5172 10532
rect 5224 10520 5230 10532
rect 8018 10520 8024 10532
rect 5224 10492 8024 10520
rect 5224 10480 5230 10492
rect 8018 10480 8024 10492
rect 8076 10520 8082 10532
rect 8128 10520 8156 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 8076 10492 8156 10520
rect 8076 10480 8082 10492
rect 8386 10480 8392 10532
rect 8444 10520 8450 10532
rect 9033 10523 9091 10529
rect 8444 10492 8708 10520
rect 8444 10480 8450 10492
rect 7834 10452 7840 10464
rect 7795 10424 7840 10452
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 8680 10461 8708 10492
rect 9033 10489 9045 10523
rect 9079 10520 9091 10523
rect 9674 10520 9680 10532
rect 9079 10492 9680 10520
rect 9079 10489 9091 10492
rect 9033 10483 9091 10489
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 8665 10455 8723 10461
rect 8665 10421 8677 10455
rect 8711 10421 8723 10455
rect 9122 10452 9128 10464
rect 9083 10424 9128 10452
rect 8665 10415 8723 10421
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 7800 10220 7972 10248
rect 7800 10208 7806 10220
rect 4338 10140 4344 10192
rect 4396 10180 4402 10192
rect 6733 10183 6791 10189
rect 6733 10180 6745 10183
rect 4396 10152 6745 10180
rect 4396 10140 4402 10152
rect 6733 10149 6745 10152
rect 6779 10180 6791 10183
rect 7834 10180 7840 10192
rect 6779 10152 7840 10180
rect 6779 10149 6791 10152
rect 6733 10143 6791 10149
rect 7834 10140 7840 10152
rect 7892 10140 7898 10192
rect 7944 10180 7972 10220
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 8202 10248 8208 10260
rect 8076 10220 8208 10248
rect 8076 10208 8082 10220
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 11241 10251 11299 10257
rect 11241 10217 11253 10251
rect 11287 10248 11299 10251
rect 12434 10248 12440 10260
rect 11287 10220 12440 10248
rect 11287 10217 11299 10220
rect 11241 10211 11299 10217
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 9582 10180 9588 10192
rect 7944 10152 9588 10180
rect 9582 10140 9588 10152
rect 9640 10140 9646 10192
rect 5169 10115 5227 10121
rect 5169 10081 5181 10115
rect 5215 10081 5227 10115
rect 5169 10075 5227 10081
rect 5184 9976 5212 10075
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 6546 10112 6552 10124
rect 5592 10084 6552 10112
rect 5592 10072 5598 10084
rect 6546 10072 6552 10084
rect 6604 10112 6610 10124
rect 6641 10115 6699 10121
rect 6641 10112 6653 10115
rect 6604 10084 6653 10112
rect 6604 10072 6610 10084
rect 6641 10081 6653 10084
rect 6687 10081 6699 10115
rect 6641 10075 6699 10081
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7653 10115 7711 10121
rect 7248 10084 7420 10112
rect 7248 10072 7254 10084
rect 6730 10004 6736 10056
rect 6788 10044 6794 10056
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6788 10016 6837 10044
rect 6788 10004 6794 10016
rect 6825 10013 6837 10016
rect 6871 10044 6883 10047
rect 7282 10044 7288 10056
rect 6871 10016 7288 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 7392 10044 7420 10084
rect 7653 10081 7665 10115
rect 7699 10112 7711 10115
rect 8202 10112 8208 10124
rect 7699 10084 8208 10112
rect 7699 10081 7711 10084
rect 7653 10075 7711 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10117 10115 10175 10121
rect 10117 10112 10129 10115
rect 10008 10084 10129 10112
rect 10008 10072 10014 10084
rect 10117 10081 10129 10084
rect 10163 10081 10175 10115
rect 10117 10075 10175 10081
rect 8386 10044 8392 10056
rect 7392 10016 8392 10044
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 9858 10044 9864 10056
rect 9819 10016 9864 10044
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 8941 9979 8999 9985
rect 8941 9976 8953 9979
rect 5184 9948 8953 9976
rect 8941 9945 8953 9948
rect 8987 9945 8999 9979
rect 8941 9939 8999 9945
rect 4982 9908 4988 9920
rect 4943 9880 4988 9908
rect 4982 9868 4988 9880
rect 5040 9868 5046 9920
rect 6273 9911 6331 9917
rect 6273 9877 6285 9911
rect 6319 9908 6331 9911
rect 7742 9908 7748 9920
rect 6319 9880 7748 9908
rect 6319 9877 6331 9880
rect 6273 9871 6331 9877
rect 7742 9868 7748 9880
rect 7800 9868 7806 9920
rect 8956 9908 8984 9939
rect 11514 9908 11520 9920
rect 8956 9880 11520 9908
rect 11514 9868 11520 9880
rect 11572 9868 11578 9920
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 8846 9704 8852 9716
rect 7616 9676 8852 9704
rect 7616 9664 7622 9676
rect 8846 9664 8852 9676
rect 8904 9664 8910 9716
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 10778 9704 10784 9716
rect 10560 9676 10784 9704
rect 10560 9664 10566 9676
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 5905 9639 5963 9645
rect 5905 9605 5917 9639
rect 5951 9636 5963 9639
rect 7006 9636 7012 9648
rect 5951 9608 7012 9636
rect 5951 9605 5963 9608
rect 5905 9599 5963 9605
rect 7006 9596 7012 9608
rect 7064 9596 7070 9648
rect 9858 9596 9864 9648
rect 9916 9636 9922 9648
rect 11333 9639 11391 9645
rect 11333 9636 11345 9639
rect 9916 9608 11345 9636
rect 9916 9596 9922 9608
rect 11333 9605 11345 9608
rect 11379 9605 11391 9639
rect 11333 9599 11391 9605
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6564 9500 6592 9531
rect 6822 9528 6828 9580
rect 6880 9568 6886 9580
rect 7558 9568 7564 9580
rect 6880 9540 7564 9568
rect 6880 9528 6886 9540
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 7742 9568 7748 9580
rect 7703 9540 7748 9568
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 7929 9571 7987 9577
rect 7929 9537 7941 9571
rect 7975 9537 7987 9571
rect 7929 9531 7987 9537
rect 6564 9472 7880 9500
rect 6270 9364 6276 9376
rect 6231 9336 6276 9364
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 6411 9336 7297 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 7650 9364 7656 9376
rect 7611 9336 7656 9364
rect 7285 9327 7343 9333
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 7852 9364 7880 9472
rect 7944 9432 7972 9531
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 9876 9500 9904 9596
rect 10873 9571 10931 9577
rect 10873 9568 10885 9571
rect 8711 9472 9904 9500
rect 9968 9540 10885 9568
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 8910 9435 8968 9441
rect 8910 9432 8922 9435
rect 7944 9404 8922 9432
rect 8910 9401 8922 9404
rect 8956 9432 8968 9435
rect 9122 9432 9128 9444
rect 8956 9404 9128 9432
rect 8956 9401 8968 9404
rect 8910 9395 8968 9401
rect 9122 9392 9128 9404
rect 9180 9432 9186 9444
rect 9968 9432 9996 9540
rect 10873 9537 10885 9540
rect 10919 9537 10931 9571
rect 10873 9531 10931 9537
rect 11514 9500 11520 9512
rect 11475 9472 11520 9500
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 9180 9404 9996 9432
rect 9180 9392 9186 9404
rect 9858 9364 9864 9376
rect 7852 9336 9864 9364
rect 9858 9324 9864 9336
rect 9916 9364 9922 9376
rect 10045 9367 10103 9373
rect 10045 9364 10057 9367
rect 9916 9336 10057 9364
rect 9916 9324 9922 9336
rect 10045 9333 10057 9336
rect 10091 9333 10103 9367
rect 10318 9364 10324 9376
rect 10279 9336 10324 9364
rect 10045 9327 10103 9333
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 10689 9367 10747 9373
rect 10689 9364 10701 9367
rect 10468 9336 10701 9364
rect 10468 9324 10474 9336
rect 10689 9333 10701 9336
rect 10735 9333 10747 9367
rect 10689 9327 10747 9333
rect 10781 9367 10839 9373
rect 10781 9333 10793 9367
rect 10827 9364 10839 9367
rect 11238 9364 11244 9376
rect 10827 9336 11244 9364
rect 10827 9333 10839 9336
rect 10781 9327 10839 9333
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 6733 9163 6791 9169
rect 6733 9129 6745 9163
rect 6779 9160 6791 9163
rect 7650 9160 7656 9172
rect 6779 9132 7656 9160
rect 6779 9129 6791 9132
rect 6733 9123 6791 9129
rect 7650 9120 7656 9132
rect 7708 9120 7714 9172
rect 9122 9160 9128 9172
rect 9083 9132 9128 9160
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 9674 9160 9680 9172
rect 9635 9132 9680 9160
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10137 9163 10195 9169
rect 10137 9129 10149 9163
rect 10183 9160 10195 9163
rect 10689 9163 10747 9169
rect 10689 9160 10701 9163
rect 10183 9132 10701 9160
rect 10183 9129 10195 9132
rect 10137 9123 10195 9129
rect 10689 9129 10701 9132
rect 10735 9129 10747 9163
rect 10689 9123 10747 9129
rect 5626 9052 5632 9104
rect 5684 9092 5690 9104
rect 7193 9095 7251 9101
rect 7193 9092 7205 9095
rect 5684 9064 7205 9092
rect 5684 9052 5690 9064
rect 7193 9061 7205 9064
rect 7239 9092 7251 9095
rect 7742 9092 7748 9104
rect 7239 9064 7748 9092
rect 7239 9061 7251 9064
rect 7193 9055 7251 9061
rect 7742 9052 7748 9064
rect 7800 9052 7806 9104
rect 9766 9052 9772 9104
rect 9824 9052 9830 9104
rect 10045 9095 10103 9101
rect 10045 9061 10057 9095
rect 10091 9092 10103 9095
rect 10318 9092 10324 9104
rect 10091 9064 10324 9092
rect 10091 9061 10103 9064
rect 10045 9055 10103 9061
rect 10318 9052 10324 9064
rect 10376 9052 10382 9104
rect 5258 8984 5264 9036
rect 5316 9024 5322 9036
rect 7098 9024 7104 9036
rect 5316 8996 7104 9024
rect 5316 8984 5322 8996
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 8001 9027 8059 9033
rect 8001 9024 8013 9027
rect 7300 8996 8013 9024
rect 7300 8968 7328 8996
rect 8001 8993 8013 8996
rect 8047 8993 8059 9027
rect 9784 9024 9812 9052
rect 11057 9027 11115 9033
rect 11057 9024 11069 9027
rect 9784 8996 11069 9024
rect 8001 8987 8059 8993
rect 11057 8993 11069 8996
rect 11103 9024 11115 9027
rect 15470 9024 15476 9036
rect 11103 8996 15476 9024
rect 11103 8993 11115 8996
rect 11057 8987 11115 8993
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 7282 8916 7288 8968
rect 7340 8956 7346 8968
rect 7745 8959 7803 8965
rect 7340 8928 7385 8956
rect 7340 8916 7346 8928
rect 7745 8925 7757 8959
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 4982 8848 4988 8900
rect 5040 8888 5046 8900
rect 7760 8888 7788 8919
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 9916 8928 10241 8956
rect 9916 8916 9922 8928
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 11146 8956 11152 8968
rect 11107 8928 11152 8956
rect 10229 8919 10287 8925
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 5040 8860 7788 8888
rect 5040 8848 5046 8860
rect 9122 8848 9128 8900
rect 9180 8888 9186 8900
rect 11256 8888 11284 8919
rect 9180 8860 11284 8888
rect 9180 8848 9186 8860
rect 10042 8780 10048 8832
rect 10100 8820 10106 8832
rect 11238 8820 11244 8832
rect 10100 8792 11244 8820
rect 10100 8780 10106 8792
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 6270 8576 6276 8628
rect 6328 8616 6334 8628
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 6328 8588 8401 8616
rect 6328 8576 6334 8588
rect 8389 8585 8401 8588
rect 8435 8585 8447 8619
rect 8389 8579 8447 8585
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 8720 8452 8861 8480
rect 8720 8440 8726 8452
rect 8849 8449 8861 8452
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8480 9091 8483
rect 9122 8480 9128 8492
rect 9079 8452 9128 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 10410 8480 10416 8492
rect 10371 8452 10416 8480
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 8754 8344 8760 8356
rect 8667 8316 8760 8344
rect 8754 8304 8760 8316
rect 8812 8344 8818 8356
rect 11974 8344 11980 8356
rect 8812 8316 11980 8344
rect 8812 8304 8818 8316
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 7190 6848 7196 6860
rect 4111 6820 7196 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 7190 6808 7196 6820
rect 7248 6808 7254 6860
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4249 6783 4307 6789
rect 4249 6780 4261 6783
rect 4212 6752 4261 6780
rect 4212 6740 4218 6752
rect 4249 6749 4261 6752
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 8202 5312 8208 5364
rect 8260 5352 8266 5364
rect 12434 5352 12440 5364
rect 8260 5324 12440 5352
rect 8260 5312 8266 5324
rect 12434 5312 12440 5324
rect 12492 5312 12498 5364
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10318 5148 10324 5160
rect 9732 5120 10324 5148
rect 9732 5108 9738 5120
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 7742 5040 7748 5092
rect 7800 5080 7806 5092
rect 11146 5080 11152 5092
rect 7800 5052 11152 5080
rect 7800 5040 7806 5052
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 7098 4972 7104 5024
rect 7156 5012 7162 5024
rect 11238 5012 11244 5024
rect 7156 4984 11244 5012
rect 7156 4972 7162 4984
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 6825 4811 6883 4817
rect 6825 4808 6837 4811
rect 6512 4780 6837 4808
rect 6512 4768 6518 4780
rect 6825 4777 6837 4780
rect 6871 4777 6883 4811
rect 6825 4771 6883 4777
rect 7377 4811 7435 4817
rect 7377 4777 7389 4811
rect 7423 4777 7435 4811
rect 10594 4808 10600 4820
rect 7377 4771 7435 4777
rect 8956 4780 10600 4808
rect 3878 4700 3884 4752
rect 3936 4740 3942 4752
rect 7392 4740 7420 4771
rect 8846 4740 8852 4752
rect 3936 4712 7420 4740
rect 7668 4712 8852 4740
rect 3936 4700 3942 4712
rect 5166 4672 5172 4684
rect 5127 4644 5172 4672
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 6641 4675 6699 4681
rect 6641 4641 6653 4675
rect 6687 4672 6699 4675
rect 7098 4672 7104 4684
rect 6687 4644 7104 4672
rect 6687 4641 6699 4644
rect 6641 4635 6699 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7193 4675 7251 4681
rect 7193 4641 7205 4675
rect 7239 4672 7251 4675
rect 7668 4672 7696 4712
rect 8846 4700 8852 4712
rect 8904 4700 8910 4752
rect 7239 4644 7696 4672
rect 7239 4641 7251 4644
rect 7193 4635 7251 4641
rect 7742 4632 7748 4684
rect 7800 4672 7806 4684
rect 8956 4681 8984 4780
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 13998 4740 14004 4752
rect 10244 4712 14004 4740
rect 8297 4675 8355 4681
rect 7800 4644 7845 4672
rect 7800 4632 7806 4644
rect 8297 4641 8309 4675
rect 8343 4641 8355 4675
rect 8297 4635 8355 4641
rect 8941 4675 8999 4681
rect 8941 4641 8953 4675
rect 8987 4641 8999 4675
rect 8941 4635 8999 4641
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4672 9735 4675
rect 10042 4672 10048 4684
rect 9723 4644 10048 4672
rect 9723 4641 9735 4644
rect 9677 4635 9735 4641
rect 6362 4564 6368 4616
rect 6420 4604 6426 4616
rect 8312 4604 8340 4635
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10244 4681 10272 4712
rect 13998 4700 14004 4712
rect 14056 4700 14062 4752
rect 10229 4675 10287 4681
rect 10229 4641 10241 4675
rect 10275 4641 10287 4675
rect 11882 4672 11888 4684
rect 11843 4644 11888 4672
rect 10229 4635 10287 4641
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 10686 4604 10692 4616
rect 6420 4576 8044 4604
rect 8312 4576 10692 4604
rect 6420 4564 6426 4576
rect 4798 4496 4804 4548
rect 4856 4536 4862 4548
rect 4856 4508 5580 4536
rect 4856 4496 4862 4508
rect 5350 4468 5356 4480
rect 5311 4440 5356 4468
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 5552 4468 5580 4508
rect 5810 4496 5816 4548
rect 5868 4536 5874 4548
rect 7929 4539 7987 4545
rect 7929 4536 7941 4539
rect 5868 4508 7941 4536
rect 5868 4496 5874 4508
rect 7929 4505 7941 4508
rect 7975 4505 7987 4539
rect 8016 4536 8044 4576
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 8481 4539 8539 4545
rect 8481 4536 8493 4539
rect 8016 4508 8493 4536
rect 7929 4499 7987 4505
rect 8481 4505 8493 4508
rect 8527 4505 8539 4539
rect 8481 4499 8539 4505
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 11606 4536 11612 4548
rect 8904 4508 11612 4536
rect 8904 4496 8910 4508
rect 11606 4496 11612 4508
rect 11664 4496 11670 4548
rect 9125 4471 9183 4477
rect 9125 4468 9137 4471
rect 5552 4440 9137 4468
rect 9125 4437 9137 4440
rect 9171 4437 9183 4471
rect 9125 4431 9183 4437
rect 9398 4428 9404 4480
rect 9456 4468 9462 4480
rect 9861 4471 9919 4477
rect 9861 4468 9873 4471
rect 9456 4440 9873 4468
rect 9456 4428 9462 4440
rect 9861 4437 9873 4440
rect 9907 4437 9919 4471
rect 10410 4468 10416 4480
rect 10371 4440 10416 4468
rect 9861 4431 9919 4437
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 11514 4428 11520 4480
rect 11572 4468 11578 4480
rect 12069 4471 12127 4477
rect 12069 4468 12081 4471
rect 11572 4440 12081 4468
rect 11572 4428 11578 4440
rect 12069 4437 12081 4440
rect 12115 4437 12127 4471
rect 12069 4431 12127 4437
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 5721 4267 5779 4273
rect 5721 4233 5733 4267
rect 5767 4264 5779 4267
rect 7926 4264 7932 4276
rect 5767 4236 7932 4264
rect 5767 4233 5779 4236
rect 5721 4227 5779 4233
rect 7926 4224 7932 4236
rect 7984 4224 7990 4276
rect 10410 4264 10416 4276
rect 8772 4236 10416 4264
rect 7009 4199 7067 4205
rect 7009 4196 7021 4199
rect 6748 4168 7021 4196
rect 3786 4088 3792 4140
rect 3844 4128 3850 4140
rect 3844 4100 5948 4128
rect 3844 4088 3850 4100
rect 3697 4063 3755 4069
rect 3697 4029 3709 4063
rect 3743 4060 3755 4063
rect 4614 4060 4620 4072
rect 3743 4032 4620 4060
rect 3743 4029 3755 4032
rect 3697 4023 3755 4029
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 4709 4063 4767 4069
rect 4709 4029 4721 4063
rect 4755 4060 4767 4063
rect 4755 4032 5212 4060
rect 4755 4029 4767 4032
rect 4709 4023 4767 4029
rect 566 3952 572 4004
rect 624 3992 630 4004
rect 5184 3992 5212 4032
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 5721 4063 5779 4069
rect 5316 4032 5361 4060
rect 5316 4020 5322 4032
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 5813 4063 5871 4069
rect 5813 4060 5825 4063
rect 5767 4032 5825 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 5813 4029 5825 4032
rect 5859 4029 5871 4063
rect 5920 4060 5948 4100
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 6748 4128 6776 4168
rect 7009 4165 7021 4168
rect 7055 4165 7067 4199
rect 7009 4159 7067 4165
rect 6328 4100 6776 4128
rect 6328 4088 6334 4100
rect 7742 4088 7748 4140
rect 7800 4128 7806 4140
rect 8772 4128 8800 4236
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 12526 4196 12532 4208
rect 7800 4100 8800 4128
rect 8864 4168 12532 4196
rect 7800 4088 7806 4100
rect 6822 4060 6828 4072
rect 5920 4032 6224 4060
rect 6783 4032 6828 4060
rect 5813 4023 5871 4029
rect 6086 3992 6092 4004
rect 624 3964 4936 3992
rect 5184 3964 6092 3992
rect 624 3952 630 3964
rect 198 3884 204 3936
rect 256 3924 262 3936
rect 4908 3933 4936 3964
rect 6086 3952 6092 3964
rect 6144 3952 6150 4004
rect 3881 3927 3939 3933
rect 3881 3924 3893 3927
rect 256 3896 3893 3924
rect 256 3884 262 3896
rect 3881 3893 3893 3896
rect 3927 3893 3939 3927
rect 3881 3887 3939 3893
rect 4893 3927 4951 3933
rect 4893 3893 4905 3927
rect 4939 3893 4951 3927
rect 5442 3924 5448 3936
rect 5403 3896 5448 3924
rect 4893 3887 4951 3893
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 5997 3927 6055 3933
rect 5997 3924 6009 3927
rect 5592 3896 6009 3924
rect 5592 3884 5598 3896
rect 5997 3893 6009 3896
rect 6043 3893 6055 3927
rect 6196 3924 6224 4032
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 7374 4020 7380 4072
rect 7432 4060 7438 4072
rect 7653 4063 7711 4069
rect 7653 4060 7665 4063
rect 7432 4032 7665 4060
rect 7432 4020 7438 4032
rect 7653 4029 7665 4032
rect 7699 4029 7711 4063
rect 7653 4023 7711 4029
rect 8205 4063 8263 4069
rect 8205 4029 8217 4063
rect 8251 4060 8263 4063
rect 8864 4060 8892 4168
rect 12526 4156 12532 4168
rect 12584 4156 12590 4208
rect 9674 4128 9680 4140
rect 8956 4100 9680 4128
rect 8956 4069 8984 4100
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 15930 4128 15936 4140
rect 11532 4100 15936 4128
rect 8251 4032 8892 4060
rect 8941 4063 8999 4069
rect 8251 4029 8263 4032
rect 8205 4023 8263 4029
rect 8941 4029 8953 4063
rect 8987 4029 8999 4063
rect 9490 4060 9496 4072
rect 9451 4032 9496 4060
rect 8941 4023 8999 4029
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 10042 4060 10048 4072
rect 10003 4032 10048 4060
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 10594 4060 10600 4072
rect 10555 4032 10600 4060
rect 10594 4020 10600 4032
rect 10652 4020 10658 4072
rect 11532 4069 11560 4100
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 11517 4063 11575 4069
rect 11517 4029 11529 4063
rect 11563 4029 11575 4063
rect 11517 4023 11575 4029
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 12989 4063 13047 4069
rect 12989 4029 13001 4063
rect 13035 4060 13047 4063
rect 16758 4060 16764 4072
rect 13035 4032 16764 4060
rect 13035 4029 13047 4032
rect 12989 4023 13047 4029
rect 12452 3992 12480 4023
rect 16758 4020 16764 4032
rect 16816 4020 16822 4072
rect 16298 3992 16304 4004
rect 12452 3964 16304 3992
rect 16298 3952 16304 3964
rect 16356 3952 16362 4004
rect 7837 3927 7895 3933
rect 7837 3924 7849 3927
rect 6196 3896 7849 3924
rect 5997 3887 6055 3893
rect 7837 3893 7849 3896
rect 7883 3893 7895 3927
rect 8386 3924 8392 3936
rect 8347 3896 8392 3924
rect 7837 3887 7895 3893
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 9030 3884 9036 3936
rect 9088 3924 9094 3936
rect 9125 3927 9183 3933
rect 9125 3924 9137 3927
rect 9088 3896 9137 3924
rect 9088 3884 9094 3896
rect 9125 3893 9137 3896
rect 9171 3893 9183 3927
rect 9125 3887 9183 3893
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3924 9735 3927
rect 9766 3924 9772 3936
rect 9723 3896 9772 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 10226 3924 10232 3936
rect 10187 3896 10232 3924
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10502 3884 10508 3936
rect 10560 3924 10566 3936
rect 10781 3927 10839 3933
rect 10781 3924 10793 3927
rect 10560 3896 10793 3924
rect 10560 3884 10566 3896
rect 10781 3893 10793 3896
rect 10827 3893 10839 3927
rect 11698 3924 11704 3936
rect 11659 3896 11704 3924
rect 10781 3887 10839 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 12618 3924 12624 3936
rect 12579 3896 12624 3924
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 13170 3924 13176 3936
rect 13131 3896 13176 3924
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 2682 3680 2688 3732
rect 2740 3720 2746 3732
rect 5721 3723 5779 3729
rect 5721 3720 5733 3723
rect 2740 3692 5733 3720
rect 2740 3680 2746 3692
rect 5721 3689 5733 3692
rect 5767 3689 5779 3723
rect 7561 3723 7619 3729
rect 7561 3720 7573 3723
rect 5721 3683 5779 3689
rect 5828 3692 7573 3720
rect 3142 3612 3148 3664
rect 3200 3652 3206 3664
rect 5828 3652 5856 3692
rect 7561 3689 7573 3692
rect 7607 3689 7619 3723
rect 7561 3683 7619 3689
rect 8113 3723 8171 3729
rect 8113 3689 8125 3723
rect 8159 3689 8171 3723
rect 8113 3683 8171 3689
rect 3200 3624 5856 3652
rect 3200 3612 3206 3624
rect 8018 3612 8024 3664
rect 8076 3652 8082 3664
rect 8128 3652 8156 3683
rect 8938 3680 8944 3732
rect 8996 3720 9002 3732
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 8996 3692 9137 3720
rect 8996 3680 9002 3692
rect 9125 3689 9137 3692
rect 9171 3689 9183 3723
rect 9125 3683 9183 3689
rect 9677 3723 9735 3729
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 9953 3723 10011 3729
rect 9953 3720 9965 3723
rect 9723 3692 9965 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 9953 3689 9965 3692
rect 9999 3689 10011 3723
rect 9953 3683 10011 3689
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 15010 3720 15016 3732
rect 10652 3692 15016 3720
rect 10652 3680 10658 3692
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 8076 3624 8156 3652
rect 8076 3612 8082 3624
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 10686 3652 10692 3664
rect 8260 3624 10692 3652
rect 8260 3612 8266 3624
rect 10686 3612 10692 3624
rect 10744 3612 10750 3664
rect 13078 3652 13084 3664
rect 11532 3624 13084 3652
rect 4706 3584 4712 3596
rect 4667 3556 4712 3584
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3584 5595 3587
rect 6178 3584 6184 3596
rect 5583 3556 6184 3584
rect 5583 3553 5595 3556
rect 5537 3547 5595 3553
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3584 6331 3587
rect 6546 3584 6552 3596
rect 6319 3556 6552 3584
rect 6319 3553 6331 3556
rect 6273 3547 6331 3553
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 6638 3544 6644 3596
rect 6696 3584 6702 3596
rect 6825 3587 6883 3593
rect 6825 3584 6837 3587
rect 6696 3556 6837 3584
rect 6696 3544 6702 3556
rect 6825 3553 6837 3556
rect 6871 3553 6883 3587
rect 6825 3547 6883 3553
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 7377 3587 7435 3593
rect 7377 3584 7389 3587
rect 6972 3556 7389 3584
rect 6972 3544 6978 3556
rect 7377 3553 7389 3556
rect 7423 3553 7435 3587
rect 7377 3547 7435 3553
rect 7926 3544 7932 3596
rect 7984 3584 7990 3596
rect 8938 3584 8944 3596
rect 7984 3556 8029 3584
rect 8899 3556 8944 3584
rect 7984 3544 7990 3556
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 9766 3584 9772 3596
rect 9727 3556 9772 3584
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 11532 3593 11560 3624
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 10597 3587 10655 3593
rect 10597 3553 10609 3587
rect 10643 3553 10655 3587
rect 10597 3547 10655 3553
rect 11517 3587 11575 3593
rect 11517 3553 11529 3587
rect 11563 3553 11575 3587
rect 11517 3547 11575 3553
rect 12345 3587 12403 3593
rect 12345 3553 12357 3587
rect 12391 3584 12403 3587
rect 13630 3584 13636 3596
rect 12391 3556 13636 3584
rect 12391 3553 12403 3556
rect 12345 3547 12403 3553
rect 1026 3476 1032 3528
rect 1084 3516 1090 3528
rect 5442 3516 5448 3528
rect 1084 3488 5448 3516
rect 1084 3476 1090 3488
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 5776 3488 9689 3516
rect 5776 3476 5782 3488
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 10612 3516 10640 3547
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 13906 3516 13912 3528
rect 10612 3488 13912 3516
rect 9677 3479 9735 3485
rect 13906 3476 13912 3488
rect 13964 3476 13970 3528
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 4893 3451 4951 3457
rect 4893 3448 4905 3451
rect 1360 3420 4905 3448
rect 1360 3408 1366 3420
rect 4893 3417 4905 3420
rect 4939 3417 4951 3451
rect 4893 3411 4951 3417
rect 4982 3408 4988 3460
rect 5040 3448 5046 3460
rect 6270 3448 6276 3460
rect 5040 3420 6276 3448
rect 5040 3408 5046 3420
rect 6270 3408 6276 3420
rect 6328 3408 6334 3460
rect 6546 3408 6552 3460
rect 6604 3448 6610 3460
rect 10781 3451 10839 3457
rect 10781 3448 10793 3451
rect 6604 3420 10793 3448
rect 6604 3408 6610 3420
rect 10781 3417 10793 3420
rect 10827 3417 10839 3451
rect 10781 3411 10839 3417
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 12529 3451 12587 3457
rect 12529 3448 12541 3451
rect 11204 3420 12541 3448
rect 11204 3408 11210 3420
rect 12529 3417 12541 3420
rect 12575 3417 12587 3451
rect 12529 3411 12587 3417
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 5534 3380 5540 3392
rect 1452 3352 5540 3380
rect 1452 3340 1458 3352
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 6454 3380 6460 3392
rect 6415 3352 6460 3380
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 7006 3380 7012 3392
rect 6967 3352 7012 3380
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 11701 3383 11759 3389
rect 11701 3380 11713 3383
rect 7524 3352 11713 3380
rect 7524 3340 7530 3352
rect 11701 3349 11713 3352
rect 11747 3349 11759 3383
rect 11701 3343 11759 3349
rect 11790 3340 11796 3392
rect 11848 3380 11854 3392
rect 14182 3380 14188 3392
rect 11848 3352 14188 3380
rect 11848 3340 11854 3352
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 5810 3176 5816 3188
rect 4488 3148 5816 3176
rect 4488 3136 4494 3148
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 6178 3136 6184 3188
rect 6236 3176 6242 3188
rect 9214 3176 9220 3188
rect 6236 3148 9220 3176
rect 6236 3136 6242 3148
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 11790 3176 11796 3188
rect 9548 3148 11796 3176
rect 9548 3136 9554 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 12894 3176 12900 3188
rect 12032 3148 12900 3176
rect 12032 3136 12038 3148
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 4706 3068 4712 3120
rect 4764 3108 4770 3120
rect 4764 3080 7880 3108
rect 4764 3068 4770 3080
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 6454 3040 6460 3052
rect 2556 3012 6460 3040
rect 2556 3000 2562 3012
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 2682 2932 2688 2984
rect 2740 2972 2746 2984
rect 7006 2972 7012 2984
rect 2740 2944 7012 2972
rect 2740 2932 2746 2944
rect 7006 2932 7012 2944
rect 7064 2932 7070 2984
rect 7852 2972 7880 3080
rect 8018 3068 8024 3120
rect 8076 3108 8082 3120
rect 8662 3108 8668 3120
rect 8076 3080 8668 3108
rect 8076 3068 8082 3080
rect 8662 3068 8668 3080
rect 8720 3068 8726 3120
rect 8938 3068 8944 3120
rect 8996 3108 9002 3120
rect 13170 3108 13176 3120
rect 8996 3080 13176 3108
rect 8996 3068 9002 3080
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 7926 3000 7932 3052
rect 7984 3040 7990 3052
rect 7984 3012 9996 3040
rect 7984 3000 7990 3012
rect 9122 2972 9128 2984
rect 7852 2944 9128 2972
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 9401 2975 9459 2981
rect 9401 2972 9413 2975
rect 9364 2944 9413 2972
rect 9364 2932 9370 2944
rect 9401 2941 9413 2944
rect 9447 2941 9459 2975
rect 9968 2972 9996 3012
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 14642 3040 14648 3052
rect 10100 3012 14648 3040
rect 10100 3000 10106 3012
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 12066 2972 12072 2984
rect 9968 2944 12072 2972
rect 9401 2935 9459 2941
rect 12066 2932 12072 2944
rect 12124 2932 12130 2984
rect 1854 2864 1860 2916
rect 1912 2904 1918 2916
rect 5350 2904 5356 2916
rect 1912 2876 5356 2904
rect 1912 2864 1918 2876
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 6270 2864 6276 2916
rect 6328 2904 6334 2916
rect 7742 2904 7748 2916
rect 6328 2876 7748 2904
rect 6328 2864 6334 2876
rect 7742 2864 7748 2876
rect 7800 2864 7806 2916
rect 8202 2864 8208 2916
rect 8260 2904 8266 2916
rect 8260 2876 9720 2904
rect 8260 2864 8266 2876
rect 2314 2796 2320 2848
rect 2372 2836 2378 2848
rect 4982 2836 4988 2848
rect 2372 2808 4988 2836
rect 2372 2796 2378 2808
rect 4982 2796 4988 2808
rect 5040 2796 5046 2848
rect 5258 2796 5264 2848
rect 5316 2836 5322 2848
rect 9585 2839 9643 2845
rect 9585 2836 9597 2839
rect 5316 2808 9597 2836
rect 5316 2796 5322 2808
rect 9585 2805 9597 2808
rect 9631 2805 9643 2839
rect 9692 2836 9720 2876
rect 9766 2864 9772 2916
rect 9824 2904 9830 2916
rect 14090 2904 14096 2916
rect 9824 2876 14096 2904
rect 9824 2864 9830 2876
rect 14090 2864 14096 2876
rect 14148 2864 14154 2916
rect 11146 2836 11152 2848
rect 9692 2808 11152 2836
rect 9585 2799 9643 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 11514 2632 11520 2644
rect 7892 2604 11520 2632
rect 7892 2592 7898 2604
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 9214 2524 9220 2576
rect 9272 2564 9278 2576
rect 9950 2564 9956 2576
rect 9272 2536 9956 2564
rect 9272 2524 9278 2536
rect 9950 2524 9956 2536
rect 10008 2524 10014 2576
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 9674 2048 9680 2100
rect 9732 2088 9738 2100
rect 13814 2088 13820 2100
rect 9732 2060 13820 2088
rect 9732 2048 9738 2060
rect 13814 2048 13820 2060
rect 13872 2048 13878 2100
rect 3970 552 3976 604
rect 4028 592 4034 604
rect 6362 592 6368 604
rect 4028 564 6368 592
rect 4028 552 4034 564
rect 6362 552 6368 564
rect 6420 552 6426 604
rect 7006 552 7012 604
rect 7064 592 7070 604
rect 9398 592 9404 604
rect 7064 564 9404 592
rect 7064 552 7070 564
rect 9398 552 9404 564
rect 9456 552 9462 604
<< via1 >>
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 3792 15104 3844 15156
rect 572 14968 624 15020
rect 1308 14968 1360 15020
rect 7104 15104 7156 15156
rect 9496 15104 9548 15156
rect 6552 15036 6604 15088
rect 8668 15036 8720 15088
rect 8760 15036 8812 15088
rect 11612 15036 11664 15088
rect 7196 14968 7248 15020
rect 9128 14968 9180 15020
rect 3148 14900 3200 14952
rect 3884 14900 3936 14952
rect 3976 14900 4028 14952
rect 6920 14900 6972 14952
rect 7748 14900 7800 14952
rect 7932 14900 7984 14952
rect 9956 14900 10008 14952
rect 8852 14832 8904 14884
rect 10692 14832 10744 14884
rect 5264 14764 5316 14816
rect 9036 14764 9088 14816
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 7380 14560 7432 14612
rect 11704 14560 11756 14612
rect 13636 14560 13688 14612
rect 16764 14560 16816 14612
rect 6276 14492 6328 14544
rect 10324 14492 10376 14544
rect 4804 14424 4856 14476
rect 8944 14424 8996 14476
rect 9128 14424 9180 14476
rect 11244 14424 11296 14476
rect 13084 14424 13136 14476
rect 15936 14424 15988 14476
rect 5724 14356 5776 14408
rect 9864 14356 9916 14408
rect 1860 14288 1912 14340
rect 5356 14288 5408 14340
rect 7380 14288 7432 14340
rect 12072 14356 12124 14408
rect 10692 14288 10744 14340
rect 15476 14288 15528 14340
rect 2688 14220 2740 14272
rect 6460 14220 6512 14272
rect 6828 14220 6880 14272
rect 9128 14220 9180 14272
rect 9312 14220 9364 14272
rect 13820 14220 13872 14272
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 204 14016 256 14068
rect 4436 14016 4488 14068
rect 5356 14059 5408 14068
rect 1032 13948 1084 14000
rect 5356 14025 5365 14059
rect 5365 14025 5399 14059
rect 5399 14025 5408 14059
rect 5356 14016 5408 14025
rect 7012 14016 7064 14068
rect 10600 14016 10652 14068
rect 13176 14016 13228 14068
rect 8024 13948 8076 14000
rect 10416 13948 10468 14000
rect 11888 13948 11940 14000
rect 16304 13948 16356 14000
rect 1400 13880 1452 13932
rect 2688 13880 2740 13932
rect 4344 13812 4396 13864
rect 5632 13880 5684 13932
rect 6644 13880 6696 13932
rect 10508 13880 10560 13932
rect 12532 13880 12584 13932
rect 5172 13855 5224 13864
rect 5172 13821 5181 13855
rect 5181 13821 5215 13855
rect 5215 13821 5224 13855
rect 5172 13812 5224 13821
rect 6828 13812 6880 13864
rect 8760 13812 8812 13864
rect 9772 13812 9824 13864
rect 10416 13812 10468 13864
rect 11152 13812 11204 13864
rect 12900 13812 12952 13864
rect 6644 13744 6696 13796
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 3516 13200 3568 13252
rect 5540 13200 5592 13252
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 14004 11704 14056 11756
rect 14648 11704 14700 11756
rect 13912 11636 13964 11688
rect 15016 11636 15068 11688
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 5540 11228 5592 11280
rect 4988 11092 5040 11144
rect 6736 10999 6788 11008
rect 6736 10965 6745 10999
rect 6745 10965 6779 10999
rect 6779 10965 6788 10999
rect 6736 10956 6788 10965
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 5172 10752 5224 10804
rect 7748 10752 7800 10804
rect 7196 10684 7248 10736
rect 7472 10684 7524 10736
rect 8392 10659 8444 10668
rect 8392 10625 8401 10659
rect 8401 10625 8435 10659
rect 8435 10625 8444 10659
rect 8392 10616 8444 10625
rect 12440 10616 12492 10668
rect 5172 10480 5224 10532
rect 8024 10480 8076 10532
rect 8392 10480 8444 10532
rect 7840 10455 7892 10464
rect 7840 10421 7849 10455
rect 7849 10421 7883 10455
rect 7883 10421 7892 10455
rect 7840 10412 7892 10421
rect 9680 10480 9732 10532
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9128 10412 9180 10421
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 7748 10208 7800 10260
rect 4344 10140 4396 10192
rect 7840 10140 7892 10192
rect 8024 10208 8076 10260
rect 8208 10208 8260 10260
rect 12440 10208 12492 10260
rect 9588 10140 9640 10192
rect 5540 10072 5592 10124
rect 6552 10072 6604 10124
rect 7196 10072 7248 10124
rect 6736 10004 6788 10056
rect 7288 10004 7340 10056
rect 8208 10072 8260 10124
rect 9956 10072 10008 10124
rect 8392 10004 8444 10056
rect 9864 10047 9916 10056
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 4988 9911 5040 9920
rect 4988 9877 4997 9911
rect 4997 9877 5031 9911
rect 5031 9877 5040 9911
rect 4988 9868 5040 9877
rect 7748 9868 7800 9920
rect 11520 9868 11572 9920
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 7564 9664 7616 9716
rect 8852 9664 8904 9716
rect 10508 9664 10560 9716
rect 10784 9664 10836 9716
rect 7012 9596 7064 9648
rect 9864 9596 9916 9648
rect 6828 9528 6880 9580
rect 7564 9528 7616 9580
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 6276 9367 6328 9376
rect 6276 9333 6285 9367
rect 6285 9333 6319 9367
rect 6319 9333 6328 9367
rect 6276 9324 6328 9333
rect 7656 9367 7708 9376
rect 7656 9333 7665 9367
rect 7665 9333 7699 9367
rect 7699 9333 7708 9367
rect 7656 9324 7708 9333
rect 9128 9392 9180 9444
rect 11520 9503 11572 9512
rect 11520 9469 11529 9503
rect 11529 9469 11563 9503
rect 11563 9469 11572 9503
rect 11520 9460 11572 9469
rect 9864 9324 9916 9376
rect 10324 9367 10376 9376
rect 10324 9333 10333 9367
rect 10333 9333 10367 9367
rect 10367 9333 10376 9367
rect 10324 9324 10376 9333
rect 10416 9324 10468 9376
rect 11244 9324 11296 9376
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 7656 9120 7708 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9128 9120 9180 9129
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 5632 9052 5684 9104
rect 7748 9052 7800 9104
rect 9772 9052 9824 9104
rect 10324 9052 10376 9104
rect 5264 8984 5316 9036
rect 7104 9027 7156 9036
rect 7104 8993 7113 9027
rect 7113 8993 7147 9027
rect 7147 8993 7156 9027
rect 7104 8984 7156 8993
rect 15476 8984 15528 9036
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 4988 8848 5040 8900
rect 9864 8916 9916 8968
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 9128 8848 9180 8900
rect 10048 8780 10100 8832
rect 11244 8780 11296 8832
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 6276 8576 6328 8628
rect 8668 8440 8720 8492
rect 9128 8440 9180 8492
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 8760 8347 8812 8356
rect 8760 8313 8769 8347
rect 8769 8313 8803 8347
rect 8803 8313 8812 8347
rect 8760 8304 8812 8313
rect 11980 8304 12032 8356
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 7196 6808 7248 6860
rect 4160 6740 4212 6792
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 8208 5312 8260 5364
rect 12440 5312 12492 5364
rect 9680 5108 9732 5160
rect 10324 5108 10376 5160
rect 7748 5040 7800 5092
rect 11152 5040 11204 5092
rect 7104 4972 7156 5024
rect 11244 4972 11296 5024
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 6460 4768 6512 4820
rect 3884 4700 3936 4752
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 7104 4632 7156 4684
rect 8852 4700 8904 4752
rect 7748 4675 7800 4684
rect 7748 4641 7757 4675
rect 7757 4641 7791 4675
rect 7791 4641 7800 4675
rect 10600 4768 10652 4820
rect 7748 4632 7800 4641
rect 6368 4564 6420 4616
rect 10048 4632 10100 4684
rect 14004 4700 14056 4752
rect 11888 4675 11940 4684
rect 11888 4641 11897 4675
rect 11897 4641 11931 4675
rect 11931 4641 11940 4675
rect 11888 4632 11940 4641
rect 4804 4496 4856 4548
rect 5356 4471 5408 4480
rect 5356 4437 5365 4471
rect 5365 4437 5399 4471
rect 5399 4437 5408 4471
rect 5356 4428 5408 4437
rect 5816 4496 5868 4548
rect 10692 4564 10744 4616
rect 8852 4496 8904 4548
rect 11612 4496 11664 4548
rect 9404 4428 9456 4480
rect 10416 4471 10468 4480
rect 10416 4437 10425 4471
rect 10425 4437 10459 4471
rect 10459 4437 10468 4471
rect 10416 4428 10468 4437
rect 11520 4428 11572 4480
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 7932 4224 7984 4276
rect 3792 4088 3844 4140
rect 4620 4020 4672 4072
rect 572 3952 624 4004
rect 5264 4063 5316 4072
rect 5264 4029 5273 4063
rect 5273 4029 5307 4063
rect 5307 4029 5316 4063
rect 5264 4020 5316 4029
rect 6276 4088 6328 4140
rect 7748 4088 7800 4140
rect 10416 4224 10468 4276
rect 6828 4063 6880 4072
rect 204 3884 256 3936
rect 6092 3952 6144 4004
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 5540 3884 5592 3936
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 7380 4020 7432 4072
rect 12532 4156 12584 4208
rect 9680 4088 9732 4140
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 9496 4020 9548 4029
rect 10048 4063 10100 4072
rect 10048 4029 10057 4063
rect 10057 4029 10091 4063
rect 10091 4029 10100 4063
rect 10048 4020 10100 4029
rect 10600 4063 10652 4072
rect 10600 4029 10609 4063
rect 10609 4029 10643 4063
rect 10643 4029 10652 4063
rect 10600 4020 10652 4029
rect 15936 4088 15988 4140
rect 16764 4020 16816 4072
rect 16304 3952 16356 4004
rect 8392 3927 8444 3936
rect 8392 3893 8401 3927
rect 8401 3893 8435 3927
rect 8435 3893 8444 3927
rect 8392 3884 8444 3893
rect 9036 3884 9088 3936
rect 9772 3884 9824 3936
rect 10232 3927 10284 3936
rect 10232 3893 10241 3927
rect 10241 3893 10275 3927
rect 10275 3893 10284 3927
rect 10232 3884 10284 3893
rect 10508 3884 10560 3936
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 12624 3927 12676 3936
rect 12624 3893 12633 3927
rect 12633 3893 12667 3927
rect 12667 3893 12676 3927
rect 12624 3884 12676 3893
rect 13176 3927 13228 3936
rect 13176 3893 13185 3927
rect 13185 3893 13219 3927
rect 13219 3893 13228 3927
rect 13176 3884 13228 3893
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 2688 3680 2740 3732
rect 3148 3612 3200 3664
rect 8024 3612 8076 3664
rect 8944 3680 8996 3732
rect 10600 3680 10652 3732
rect 15016 3680 15068 3732
rect 8208 3612 8260 3664
rect 10692 3612 10744 3664
rect 4712 3587 4764 3596
rect 4712 3553 4721 3587
rect 4721 3553 4755 3587
rect 4755 3553 4764 3587
rect 4712 3544 4764 3553
rect 6184 3544 6236 3596
rect 6552 3544 6604 3596
rect 6644 3544 6696 3596
rect 6920 3544 6972 3596
rect 7932 3587 7984 3596
rect 7932 3553 7941 3587
rect 7941 3553 7975 3587
rect 7975 3553 7984 3587
rect 8944 3587 8996 3596
rect 7932 3544 7984 3553
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 9772 3587 9824 3596
rect 9772 3553 9781 3587
rect 9781 3553 9815 3587
rect 9815 3553 9824 3587
rect 9772 3544 9824 3553
rect 13084 3612 13136 3664
rect 1032 3476 1084 3528
rect 5448 3476 5500 3528
rect 5724 3476 5776 3528
rect 13636 3544 13688 3596
rect 13912 3476 13964 3528
rect 1308 3408 1360 3460
rect 4988 3408 5040 3460
rect 6276 3408 6328 3460
rect 6552 3408 6604 3460
rect 11152 3408 11204 3460
rect 1400 3340 1452 3392
rect 5540 3340 5592 3392
rect 6460 3383 6512 3392
rect 6460 3349 6469 3383
rect 6469 3349 6503 3383
rect 6503 3349 6512 3383
rect 6460 3340 6512 3349
rect 7012 3383 7064 3392
rect 7012 3349 7021 3383
rect 7021 3349 7055 3383
rect 7055 3349 7064 3383
rect 7012 3340 7064 3349
rect 7472 3340 7524 3392
rect 11796 3340 11848 3392
rect 14188 3340 14240 3392
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 4436 3136 4488 3188
rect 5816 3136 5868 3188
rect 6184 3136 6236 3188
rect 9220 3136 9272 3188
rect 9496 3136 9548 3188
rect 11796 3136 11848 3188
rect 11980 3136 12032 3188
rect 12900 3136 12952 3188
rect 4712 3068 4764 3120
rect 2504 3000 2556 3052
rect 6460 3000 6512 3052
rect 2688 2932 2740 2984
rect 7012 2932 7064 2984
rect 8024 3068 8076 3120
rect 8668 3068 8720 3120
rect 8944 3068 8996 3120
rect 13176 3068 13228 3120
rect 7932 3000 7984 3052
rect 9128 2932 9180 2984
rect 9312 2932 9364 2984
rect 10048 3000 10100 3052
rect 14648 3000 14700 3052
rect 12072 2932 12124 2984
rect 1860 2864 1912 2916
rect 5356 2864 5408 2916
rect 6276 2864 6328 2916
rect 7748 2864 7800 2916
rect 8208 2864 8260 2916
rect 2320 2796 2372 2848
rect 4988 2796 5040 2848
rect 5264 2796 5316 2848
rect 9772 2864 9824 2916
rect 14096 2864 14148 2916
rect 11152 2796 11204 2848
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 7840 2592 7892 2644
rect 11520 2592 11572 2644
rect 9220 2524 9272 2576
rect 9956 2524 10008 2576
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 9680 2048 9732 2100
rect 13820 2048 13872 2100
rect 3976 552 4028 604
rect 6368 552 6420 604
rect 7012 552 7064 604
rect 9404 552 9456 604
<< metal2 >>
rect 202 17520 258 18000
rect 570 17520 626 18000
rect 1030 17520 1086 18000
rect 1398 17520 1454 18000
rect 1858 17520 1914 18000
rect 2318 17520 2374 18000
rect 2686 17520 2742 18000
rect 3146 17520 3202 18000
rect 3606 17520 3662 18000
rect 3974 17520 4030 18000
rect 4434 17520 4490 18000
rect 4802 17520 4858 18000
rect 5262 17520 5318 18000
rect 5722 17520 5778 18000
rect 6090 17520 6146 18000
rect 6550 17520 6606 18000
rect 7010 17520 7066 18000
rect 7378 17520 7434 18000
rect 7838 17520 7894 18000
rect 8206 17520 8262 18000
rect 8666 17520 8722 18000
rect 9126 17520 9182 18000
rect 9494 17520 9550 18000
rect 9954 17520 10010 18000
rect 10414 17520 10470 18000
rect 10782 17520 10838 18000
rect 11242 17520 11298 18000
rect 11610 17520 11666 18000
rect 12070 17520 12126 18000
rect 12530 17520 12586 18000
rect 12898 17520 12954 18000
rect 13358 17520 13414 18000
rect 13818 17520 13874 18000
rect 14186 17520 14242 18000
rect 14646 17520 14702 18000
rect 15014 17520 15070 18000
rect 15474 17520 15530 18000
rect 15934 17520 15990 18000
rect 16302 17520 16358 18000
rect 16762 17520 16818 18000
rect 216 14074 244 17520
rect 584 15026 612 17520
rect 572 15020 624 15026
rect 572 14962 624 14968
rect 204 14068 256 14074
rect 204 14010 256 14016
rect 1044 14006 1072 17520
rect 1308 15020 1360 15026
rect 1308 14962 1360 14968
rect 1032 14000 1084 14006
rect 1032 13942 1084 13948
rect 572 4004 624 4010
rect 572 3946 624 3952
rect 204 3936 256 3942
rect 204 3878 256 3884
rect 216 480 244 3878
rect 584 480 612 3946
rect 1032 3528 1084 3534
rect 1032 3470 1084 3476
rect 1044 480 1072 3470
rect 1320 3466 1348 14962
rect 1412 13938 1440 17520
rect 1872 14346 1900 17520
rect 2332 15178 2360 17520
rect 2332 15150 2544 15178
rect 1860 14340 1912 14346
rect 1860 14282 1912 14288
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1412 480 1440 3334
rect 2516 3058 2544 15150
rect 2700 14278 2728 17520
rect 3160 14958 3188 17520
rect 3620 15450 3648 17520
rect 3620 15422 3832 15450
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 3804 15162 3832 15422
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3988 15042 4016 17520
rect 3804 15014 4016 15042
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2700 3738 2728 13874
rect 3514 13560 3570 13569
rect 3514 13495 3570 13504
rect 3528 13258 3556 13495
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3804 4298 3832 15014
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3896 4758 3924 14894
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3804 4270 3924 4298
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1872 480 1900 2858
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 2332 480 2360 2790
rect 2700 480 2728 2926
rect 3160 480 3188 3606
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 3804 1578 3832 4082
rect 3896 4049 3924 4270
rect 3882 4040 3938 4049
rect 3882 3975 3938 3984
rect 3988 3641 4016 14894
rect 4448 14074 4476 17520
rect 4816 14482 4844 17520
rect 5276 14822 5304 17520
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 5736 14414 5764 17520
rect 6104 15994 6132 17520
rect 6104 15966 6316 15994
rect 5886 15804 6182 15824
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 5886 14716 6182 14736
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 6288 14550 6316 15966
rect 6564 15178 6592 17520
rect 6564 15150 6684 15178
rect 6552 15088 6604 15094
rect 6552 15030 6604 15036
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5368 14074 5396 14282
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 4356 10198 4384 13806
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 5000 9926 5028 11086
rect 5184 10810 5212 13806
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5552 11286 5580 13194
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 5000 8906 5028 9862
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4066 4584 4122 4593
rect 4172 4570 4200 6734
rect 5184 4690 5212 10474
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 4122 4542 4200 4570
rect 4804 4548 4856 4554
rect 4066 4519 4122 4528
rect 4804 4490 4856 4496
rect 4618 4176 4674 4185
rect 4618 4111 4674 4120
rect 4632 4078 4660 4111
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 3974 3632 4030 3641
rect 3974 3567 4030 3576
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 3620 1550 3832 1578
rect 3620 480 3648 1550
rect 3976 604 4028 610
rect 3976 546 4028 552
rect 3988 480 4016 546
rect 4448 480 4476 3130
rect 4724 3126 4752 3538
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4816 480 4844 4490
rect 5276 4078 5304 8978
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 5000 2854 5028 3402
rect 5368 2922 5396 4422
rect 5552 4185 5580 10066
rect 5644 9110 5672 13874
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 5886 12540 6182 12560
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 5886 11452 6182 11472
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 5886 9276 6182 9296
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 6288 8634 6316 9318
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 5886 8188 6182 8208
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 5886 7100 6182 7120
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 6472 4826 6500 14214
rect 6564 10130 6592 15030
rect 6656 13938 6684 15150
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6840 13870 6868 14214
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5538 4176 5594 4185
rect 5538 4111 5594 4120
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5460 3534 5488 3878
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5552 3398 5580 3878
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5276 480 5304 2790
rect 5736 480 5764 3470
rect 5828 3194 5856 4490
rect 6090 4176 6146 4185
rect 6090 4111 6146 4120
rect 6276 4140 6328 4146
rect 6104 4010 6132 4111
rect 6276 4082 6328 4088
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 5886 3836 6182 3856
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6196 3194 6224 3538
rect 6288 3466 6316 4082
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 6288 1442 6316 2858
rect 6104 1414 6316 1442
rect 6104 480 6132 1414
rect 6380 610 6408 4558
rect 6550 3768 6606 3777
rect 6550 3703 6606 3712
rect 6564 3602 6592 3703
rect 6656 3602 6684 13738
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6748 10713 6776 10950
rect 6734 10704 6790 10713
rect 6734 10639 6790 10648
rect 6748 10062 6776 10639
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6840 4078 6868 9522
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6932 3602 6960 14894
rect 7024 14074 7052 17520
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7010 10024 7066 10033
rect 7010 9959 7066 9968
rect 7024 9654 7052 9959
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 7116 9042 7144 15098
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7208 10742 7236 14962
rect 7392 14618 7420 17520
rect 7746 15056 7802 15065
rect 7852 15042 7880 17520
rect 7852 15014 8156 15042
rect 7746 14991 7802 15000
rect 7760 14958 7788 14991
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7208 6866 7236 10066
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7300 8974 7328 9998
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 7116 4690 7144 4966
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7392 4078 7420 14282
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 7484 4185 7512 10678
rect 7760 10266 7788 10746
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7852 10305 7880 10406
rect 7838 10296 7894 10305
rect 7748 10260 7800 10266
rect 7838 10231 7894 10240
rect 7748 10202 7800 10208
rect 7840 10192 7892 10198
rect 7840 10134 7892 10140
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7576 9586 7604 9658
rect 7760 9586 7788 9862
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 9178 7696 9318
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7748 9104 7800 9110
rect 7668 9052 7748 9058
rect 7668 9046 7800 9052
rect 7668 9030 7788 9046
rect 7470 4176 7526 4185
rect 7470 4111 7526 4120
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 3058 6500 3334
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6368 604 6420 610
rect 6368 546 6420 552
rect 6564 480 6592 3402
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7024 2990 7052 3334
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7484 1714 7512 3334
rect 7668 3097 7696 9030
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7760 4690 7788 5034
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7654 3088 7710 3097
rect 7654 3023 7710 3032
rect 7760 2922 7788 4082
rect 7852 2938 7880 10134
rect 7944 4282 7972 14894
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 8036 10538 8064 13942
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 8036 3754 8064 10202
rect 8128 3913 8156 15014
rect 8220 10266 8248 17520
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8352 15184 8648 15204
rect 8680 15094 8708 17520
rect 8668 15088 8720 15094
rect 8760 15088 8812 15094
rect 8668 15030 8720 15036
rect 8758 15056 8760 15065
rect 8812 15056 8814 15065
rect 9140 15026 9168 17520
rect 9508 15162 9536 17520
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 8758 14991 8814 15000
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9968 14958 9996 17520
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8352 14096 8648 14116
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8352 13084 8648 13104
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8352 11920 8648 11940
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 8390 10704 8446 10713
rect 8390 10639 8392 10648
rect 8444 10639 8446 10648
rect 8392 10610 8444 10616
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8220 5370 8248 10066
rect 8404 10062 8432 10474
rect 8666 10296 8722 10305
rect 8666 10231 8722 10240
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8680 8498 8708 10231
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8772 8362 8800 13806
rect 8864 9722 8892 14826
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8352 7644 8648 7664
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8352 7568 8648 7588
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8352 6480 8648 6500
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8864 4554 8892 4694
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8390 4040 8446 4049
rect 8390 3975 8446 3984
rect 8404 3942 8432 3975
rect 8392 3936 8444 3942
rect 8114 3904 8170 3913
rect 8392 3878 8444 3884
rect 8114 3839 8170 3848
rect 8206 3768 8262 3777
rect 8036 3726 8156 3754
rect 8024 3664 8076 3670
rect 8022 3632 8024 3641
rect 8076 3632 8078 3641
rect 7932 3596 7984 3602
rect 8022 3567 8078 3576
rect 7932 3538 7984 3544
rect 7944 3058 7972 3538
rect 8128 3505 8156 3726
rect 8956 3738 8984 14418
rect 9048 3942 9076 14758
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 9140 14278 9168 14418
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 10033 9168 10406
rect 9126 10024 9182 10033
rect 9126 9959 9182 9968
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9140 9178 9168 9386
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9140 8906 9168 9114
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9140 8498 9168 8842
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 8206 3703 8262 3712
rect 8944 3732 8996 3738
rect 8220 3670 8248 3703
rect 8944 3674 8996 3680
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8114 3496 8170 3505
rect 8114 3431 8170 3440
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8352 3216 8648 3236
rect 8956 3126 8984 3538
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8036 2938 8064 3062
rect 7748 2916 7800 2922
rect 7852 2910 8064 2938
rect 8208 2916 8260 2922
rect 7748 2858 7800 2864
rect 8208 2858 8260 2864
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7392 1686 7512 1714
rect 7012 604 7064 610
rect 7012 546 7064 552
rect 7024 480 7052 546
rect 7392 480 7420 1686
rect 7852 480 7880 2586
rect 8220 480 8248 2858
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 8680 480 8708 3062
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9140 480 9168 2926
rect 9232 2582 9260 3130
rect 9324 2990 9352 14214
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9600 9058 9628 10134
rect 9692 9178 9720 10474
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9784 9110 9812 13806
rect 9876 10169 9904 14350
rect 9862 10160 9918 10169
rect 9862 10095 9918 10104
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9876 9654 9904 9998
rect 9864 9648 9916 9654
rect 9968 9625 9996 10066
rect 10138 9752 10194 9761
rect 10138 9687 10194 9696
rect 10152 9636 10180 9687
rect 10152 9625 10272 9636
rect 9864 9590 9916 9596
rect 9954 9616 10010 9625
rect 10152 9616 10286 9625
rect 10152 9608 10230 9616
rect 9954 9551 10010 9560
rect 10230 9551 10286 9560
rect 9862 9480 9918 9489
rect 10336 9466 10364 14486
rect 10428 14006 10456 17520
rect 10796 15994 10824 17520
rect 10704 15966 10824 15994
rect 10704 14890 10732 15966
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 11256 14482 11284 17520
rect 11624 15094 11652 17520
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10416 14000 10468 14006
rect 10416 13942 10468 13948
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 9862 9415 9918 9424
rect 10244 9438 10364 9466
rect 10428 9466 10456 13806
rect 10520 9722 10548 13874
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10428 9438 10548 9466
rect 9876 9382 9904 9415
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9772 9104 9824 9110
rect 9600 9030 9720 9058
rect 9772 9046 9824 9052
rect 9692 5166 9720 9030
rect 9876 8974 9904 9318
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 10060 4690 10088 8774
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 9416 610 9444 4422
rect 9770 4176 9826 4185
rect 9680 4140 9732 4146
rect 9770 4111 9826 4120
rect 9680 4082 9732 4088
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9508 3194 9536 4014
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9494 3088 9550 3097
rect 9494 3023 9550 3032
rect 9404 604 9456 610
rect 9404 546 9456 552
rect 9508 480 9536 3023
rect 9692 2106 9720 4082
rect 9784 3942 9812 4111
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9784 2922 9812 3538
rect 10060 3058 10088 4014
rect 10244 3942 10272 9438
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10336 9110 10364 9318
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10428 8498 10456 9318
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 9968 480 9996 2518
rect 10336 592 10364 5102
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10428 4282 10456 4422
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10520 3942 10548 9438
rect 10612 4826 10640 14010
rect 10704 9625 10732 14282
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 10817 13628 11113 13648
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10817 10288 11113 10308
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10690 9616 10746 9625
rect 10690 9551 10746 9560
rect 10796 9466 10824 9658
rect 10704 9438 10824 9466
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10704 4622 10732 9438
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 11164 8974 11192 13806
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11242 9616 11298 9625
rect 11242 9551 11298 9560
rect 11256 9382 11284 9551
rect 11532 9518 11560 9862
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 10817 8188 11113 8208
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 11164 5098 11192 8910
rect 11256 8838 11284 9318
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10612 3738 10640 4014
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10704 2530 10732 3606
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 2854 11192 3402
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 10704 2502 10824 2530
rect 10336 564 10456 592
rect 10428 480 10456 564
rect 10796 480 10824 2502
rect 11256 480 11284 4966
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 11532 2650 11560 4422
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11624 480 11652 4490
rect 11716 3942 11744 14554
rect 12084 14414 12112 17520
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11900 4690 11928 13942
rect 12544 13938 12572 17520
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12912 13870 12940 17520
rect 13372 15450 13400 17520
rect 13188 15422 13400 15450
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12438 13560 12494 13569
rect 12438 13495 12494 13504
rect 12452 10674 12480 13495
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12452 10266 12480 10610
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11808 3194 11836 3334
rect 11992 3194 12020 8298
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12452 4593 12480 5306
rect 12438 4584 12494 4593
rect 12438 4519 12494 4528
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12084 480 12112 2926
rect 12544 480 12572 4150
rect 12622 4040 12678 4049
rect 12622 3975 12678 3984
rect 12636 3942 12664 3975
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 13096 3670 13124 14418
rect 13188 14074 13216 15422
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 13188 3505 13216 3878
rect 13648 3602 13676 14554
rect 13832 14278 13860 17520
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13924 3534 13952 11630
rect 14016 4758 14044 11698
rect 14200 5250 14228 17520
rect 14660 11762 14688 17520
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 15028 11694 15056 17520
rect 15488 14346 15516 17520
rect 15948 14482 15976 17520
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 16316 14006 16344 17520
rect 16776 14618 16804 17520
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 14108 5222 14228 5250
rect 14004 4752 14056 4758
rect 14004 4694 14056 4700
rect 13912 3528 13964 3534
rect 13174 3496 13230 3505
rect 13912 3470 13964 3476
rect 13174 3431 13230 3440
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 12912 480 12940 3130
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13188 1850 13216 3062
rect 14108 2922 14136 5222
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14096 2916 14148 2922
rect 14096 2858 14148 2864
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 13820 2100 13872 2106
rect 13820 2042 13872 2048
rect 13188 1822 13400 1850
rect 13372 480 13400 1822
rect 13832 480 13860 2042
rect 14200 480 14228 3334
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14660 480 14688 2994
rect 15028 480 15056 3674
rect 15488 480 15516 8978
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15948 480 15976 4082
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16316 480 16344 3946
rect 16776 480 16804 4014
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1398 0 1454 480
rect 1858 0 1914 480
rect 2318 0 2374 480
rect 2686 0 2742 480
rect 3146 0 3202 480
rect 3606 0 3662 480
rect 3974 0 4030 480
rect 4434 0 4490 480
rect 4802 0 4858 480
rect 5262 0 5318 480
rect 5722 0 5778 480
rect 6090 0 6146 480
rect 6550 0 6606 480
rect 7010 0 7066 480
rect 7378 0 7434 480
rect 7838 0 7894 480
rect 8206 0 8262 480
rect 8666 0 8722 480
rect 9126 0 9182 480
rect 9494 0 9550 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10782 0 10838 480
rect 11242 0 11298 480
rect 11610 0 11666 480
rect 12070 0 12126 480
rect 12530 0 12586 480
rect 12898 0 12954 480
rect 13358 0 13414 480
rect 13818 0 13874 480
rect 14186 0 14242 480
rect 14646 0 14702 480
rect 15014 0 15070 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16302 0 16358 480
rect 16762 0 16818 480
<< via2 >>
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3514 13504 3570 13560
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 3882 3984 3938 4040
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 4066 4528 4122 4584
rect 4618 4120 4674 4176
rect 3974 3576 4030 3632
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 5538 4120 5594 4176
rect 6090 4120 6146 4176
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 6550 3712 6606 3768
rect 6734 10648 6790 10704
rect 7010 9968 7066 10024
rect 7746 15000 7802 15056
rect 7838 10240 7894 10296
rect 7470 4120 7526 4176
rect 7654 3032 7710 3088
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 8758 15036 8760 15056
rect 8760 15036 8812 15056
rect 8812 15036 8814 15056
rect 8758 15000 8814 15036
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 8390 10668 8446 10704
rect 8390 10648 8392 10668
rect 8392 10648 8444 10668
rect 8444 10648 8446 10668
rect 8666 10240 8722 10296
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 8390 3984 8446 4040
rect 8114 3848 8170 3904
rect 8022 3612 8024 3632
rect 8024 3612 8076 3632
rect 8076 3612 8078 3632
rect 8022 3576 8078 3612
rect 8206 3712 8262 3768
rect 9126 9968 9182 10024
rect 8114 3440 8170 3496
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 9862 10104 9918 10160
rect 10138 9696 10194 9752
rect 9954 9560 10010 9616
rect 10230 9560 10286 9616
rect 9862 9424 9918 9480
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 9770 4120 9826 4176
rect 9494 3032 9550 3088
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 10690 9560 10746 9616
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 11242 9560 11298 9616
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 12438 13504 12494 13560
rect 12438 4528 12494 4584
rect 12622 3984 12678 4040
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13174 3440 13230 3496
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
<< metal3 >>
rect 5874 15808 6194 15809
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 3409 15264 3729 15265
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 7741 15058 7807 15061
rect 8753 15058 8819 15061
rect 7741 15056 8819 15058
rect 7741 15000 7746 15056
rect 7802 15000 8758 15056
rect 8814 15000 8819 15056
rect 7741 14998 8819 15000
rect 7741 14995 7807 14998
rect 8753 14995 8819 14998
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 3409 14176 3729 14177
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 5874 13632 6194 13633
rect 0 13562 480 13592
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 3509 13562 3575 13565
rect 0 13560 3575 13562
rect 0 13504 3514 13560
rect 3570 13504 3575 13560
rect 0 13502 3575 13504
rect 0 13472 480 13502
rect 3509 13499 3575 13502
rect 12433 13562 12499 13565
rect 16520 13562 17000 13592
rect 12433 13560 17000 13562
rect 12433 13504 12438 13560
rect 12494 13504 17000 13560
rect 12433 13502 17000 13504
rect 12433 13499 12499 13502
rect 16520 13472 17000 13502
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 5874 12544 6194 12545
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 3409 12000 3729 12001
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 5874 11456 6194 11457
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 6729 10706 6795 10709
rect 8385 10706 8451 10709
rect 6729 10704 8451 10706
rect 6729 10648 6734 10704
rect 6790 10648 8390 10704
rect 8446 10648 8451 10704
rect 6729 10646 8451 10648
rect 6729 10643 6795 10646
rect 8385 10643 8451 10646
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 7833 10298 7899 10301
rect 8661 10298 8727 10301
rect 7833 10296 8727 10298
rect 7833 10240 7838 10296
rect 7894 10240 8666 10296
rect 8722 10240 8727 10296
rect 7833 10238 8727 10240
rect 7833 10235 7899 10238
rect 8661 10235 8727 10238
rect 9857 10160 9923 10165
rect 9857 10104 9862 10160
rect 9918 10104 9923 10160
rect 9857 10099 9923 10104
rect 7005 10026 7071 10029
rect 9121 10026 9187 10029
rect 7005 10024 9187 10026
rect 7005 9968 7010 10024
rect 7066 9968 9126 10024
rect 9182 9968 9187 10024
rect 7005 9966 9187 9968
rect 7005 9963 7071 9966
rect 9121 9963 9187 9966
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 9860 9754 9920 10099
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 9759 13590 9760
rect 10133 9754 10199 9757
rect 9860 9752 10199 9754
rect 9860 9696 10138 9752
rect 10194 9696 10199 9752
rect 9860 9694 10199 9696
rect 10133 9691 10199 9694
rect 9949 9618 10015 9621
rect 9814 9616 10015 9618
rect 9814 9560 9954 9616
rect 10010 9560 10015 9616
rect 9814 9558 10015 9560
rect 9814 9485 9874 9558
rect 9949 9555 10015 9558
rect 10225 9618 10291 9621
rect 10358 9618 10364 9620
rect 10225 9616 10364 9618
rect 10225 9560 10230 9616
rect 10286 9560 10364 9616
rect 10225 9558 10364 9560
rect 10225 9555 10291 9558
rect 10358 9556 10364 9558
rect 10428 9556 10434 9620
rect 10685 9618 10751 9621
rect 11237 9618 11303 9621
rect 10685 9616 11303 9618
rect 10685 9560 10690 9616
rect 10746 9560 11242 9616
rect 11298 9560 11303 9616
rect 10685 9558 11303 9560
rect 10685 9555 10751 9558
rect 11237 9555 11303 9558
rect 9814 9480 9923 9485
rect 9814 9424 9862 9480
rect 9918 9424 9923 9480
rect 9814 9422 9923 9424
rect 9857 9419 9923 9422
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 5874 8192 6194 8193
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 3409 6560 3729 6561
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 3409 5472 3729 5473
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 0 4586 480 4616
rect 4061 4586 4127 4589
rect 0 4584 4127 4586
rect 0 4528 4066 4584
rect 4122 4528 4127 4584
rect 0 4526 4127 4528
rect 0 4496 480 4526
rect 4061 4523 4127 4526
rect 12433 4586 12499 4589
rect 16520 4586 17000 4616
rect 12433 4584 17000 4586
rect 12433 4528 12438 4584
rect 12494 4528 17000 4584
rect 12433 4526 17000 4528
rect 12433 4523 12499 4526
rect 16520 4496 17000 4526
rect 3409 4384 3729 4385
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 4613 4178 4679 4181
rect 5533 4178 5599 4181
rect 4613 4176 5599 4178
rect 4613 4120 4618 4176
rect 4674 4120 5538 4176
rect 5594 4120 5599 4176
rect 4613 4118 5599 4120
rect 4613 4115 4679 4118
rect 5533 4115 5599 4118
rect 6085 4178 6151 4181
rect 7465 4178 7531 4181
rect 6085 4176 7531 4178
rect 6085 4120 6090 4176
rect 6146 4120 7470 4176
rect 7526 4120 7531 4176
rect 6085 4118 7531 4120
rect 6085 4115 6151 4118
rect 7465 4115 7531 4118
rect 9765 4178 9831 4181
rect 10358 4178 10364 4180
rect 9765 4176 10364 4178
rect 9765 4120 9770 4176
rect 9826 4120 10364 4176
rect 9765 4118 10364 4120
rect 9765 4115 9831 4118
rect 10358 4116 10364 4118
rect 10428 4116 10434 4180
rect 3877 4042 3943 4045
rect 8385 4042 8451 4045
rect 12617 4042 12683 4045
rect 3877 4040 8451 4042
rect 3877 3984 3882 4040
rect 3938 3984 8390 4040
rect 8446 3984 8451 4040
rect 3877 3982 8451 3984
rect 3877 3979 3943 3982
rect 8385 3979 8451 3982
rect 8526 4040 12683 4042
rect 8526 3984 12622 4040
rect 12678 3984 12683 4040
rect 8526 3982 12683 3984
rect 8109 3906 8175 3909
rect 8526 3906 8586 3982
rect 12617 3979 12683 3982
rect 8109 3904 8586 3906
rect 8109 3848 8114 3904
rect 8170 3848 8586 3904
rect 8109 3846 8586 3848
rect 8109 3843 8175 3846
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 6545 3770 6611 3773
rect 8201 3770 8267 3773
rect 6545 3768 8267 3770
rect 6545 3712 6550 3768
rect 6606 3712 8206 3768
rect 8262 3712 8267 3768
rect 6545 3710 8267 3712
rect 6545 3707 6611 3710
rect 8201 3707 8267 3710
rect 3969 3634 4035 3637
rect 8017 3634 8083 3637
rect 3969 3632 8083 3634
rect 3969 3576 3974 3632
rect 4030 3576 8022 3632
rect 8078 3576 8083 3632
rect 3969 3574 8083 3576
rect 3969 3571 4035 3574
rect 8017 3571 8083 3574
rect 8109 3498 8175 3501
rect 13169 3498 13235 3501
rect 8109 3496 13235 3498
rect 8109 3440 8114 3496
rect 8170 3440 13174 3496
rect 13230 3440 13235 3496
rect 8109 3438 13235 3440
rect 8109 3435 8175 3438
rect 13169 3435 13235 3438
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 3231 13590 3232
rect 7649 3090 7715 3093
rect 9489 3090 9555 3093
rect 7649 3088 9555 3090
rect 7649 3032 7654 3088
rect 7710 3032 9494 3088
rect 9550 3032 9555 3088
rect 7649 3030 9555 3032
rect 7649 3027 7715 3030
rect 9489 3027 9555 3030
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
<< via3 >>
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 10364 9556 10428 9620
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 10364 4116 10428 4180
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
<< metal4 >>
rect 3409 15264 3729 15824
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 14176 3729 15200
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 13088 3729 14112
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 12000 3729 13024
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 10912 3729 11936
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 9824 3729 10848
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 3296 3729 4320
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 5874 15808 6195 15824
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 5874 14720 6195 15744
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5874 13632 6195 14656
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5874 12544 6195 13568
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5874 11456 6195 12480
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5874 10368 6195 11392
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 5874 8192 6195 9216
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 5874 7104 6195 8128
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5874 6016 6195 7040
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5874 2752 6195 3776
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 5874 2128 6195 2688
rect 8340 15264 8660 15824
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 14176 8660 15200
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 13088 8660 14112
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 12000 8660 13024
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 10912 8660 11936
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 9824 8660 10848
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 8736 8660 9760
rect 10805 15808 11125 15824
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 14720 11125 15744
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 13632 11125 14656
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 12544 11125 13568
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 11456 11125 12480
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 10368 11125 11392
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10363 9620 10429 9621
rect 10363 9556 10364 9620
rect 10428 9556 10429 9620
rect 10363 9555 10429 9556
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 7648 8660 8672
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 5472 8660 6496
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 10366 4181 10426 9555
rect 10805 9280 11125 10304
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 8192 11125 9216
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 7104 11125 8128
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 6016 11125 7040
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10363 4180 10429 4181
rect 10363 4116 10364 4180
rect 10428 4116 10429 4180
rect 10363 4115 10429 4116
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 2208 8660 3232
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 10805 3840 11125 4864
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 2752 11125 3776
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2128 11125 2688
rect 13270 15264 13590 15824
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 14176 13590 15200
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 13088 13590 14112
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 12000 13590 13024
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 10912 13590 11936
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 9824 13590 10848
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 8736 13590 9760
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 6560 13590 7584
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 5472 13590 6496
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 2208 13590 3232
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1605641404
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1605641404
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1605641404
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1605641404
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1605641404
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1605641404
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _25_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 9384 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1605641404
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1605641404
transform 1 0 9016 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1605641404
transform 1 0 9752 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1605641404
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1605641404
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_106
timestamp 1605641404
transform 1 0 10856 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1605641404
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1605641404
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1605641404
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1605641404
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_147
timestamp 1605641404
transform 1 0 14628 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1605641404
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1605641404
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1605641404
transform 1 0 4692 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1605641404
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_32
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_38
timestamp 1605641404
transform 1 0 4600 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1605641404
transform 1 0 6256 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1605641404
transform 1 0 5520 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1605641404
transform 1 0 6808 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_43
timestamp 1605641404
transform 1 0 5060 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_47
timestamp 1605641404
transform 1 0 5428 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_52
timestamp 1605641404
transform 1 0 5888 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_60
timestamp 1605641404
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _09_
timestamp 1605641404
transform 1 0 7912 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1605641404
transform 1 0 7360 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1605641404
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_72
timestamp 1605641404
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1605641404
transform 1 0 8280 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _06_
timestamp 1605641404
transform 1 0 8924 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1605641404
transform 1 0 10580 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1605641404
transform 1 0 9752 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_84
timestamp 1605641404
transform 1 0 8832 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1605641404
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_98
timestamp 1605641404
transform 1 0 10120 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_102
timestamp 1605641404
transform 1 0 10488 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1605641404
transform 1 0 12328 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1605641404
transform 1 0 11500 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_107
timestamp 1605641404
transform 1 0 10948 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1605641404
transform 1 0 11868 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1605641404
transform 1 0 12236 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_126
timestamp 1605641404
transform 1 0 12696 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_138
timestamp 1605641404
transform 1 0 13800 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1605641404
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1605641404
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1605641404
transform 1 0 4692 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1605641404
transform 1 0 3680 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_27
timestamp 1605641404
transform 1 0 3588 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_32
timestamp 1605641404
transform 1 0 4048 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_38
timestamp 1605641404
transform 1 0 4600 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1605641404
transform 1 0 5796 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1605641404
transform 1 0 5244 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 1605641404
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_49
timestamp 1605641404
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_55
timestamp 1605641404
transform 1 0 6164 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1605641404
transform 1 0 8188 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1605641404
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_66
timestamp 1605641404
transform 1 0 7176 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_70
timestamp 1605641404
transform 1 0 7544 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1605641404
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_81
timestamp 1605641404
transform 1 0 8556 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _02_
timestamp 1605641404
transform 1 0 10580 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _03_
timestamp 1605641404
transform 1 0 10028 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _04_
timestamp 1605641404
transform 1 0 9476 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1605641404
transform 1 0 8924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1605641404
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_95
timestamp 1605641404
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1605641404
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1605641404
transform 1 0 11500 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_107
timestamp 1605641404
transform 1 0 10948 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1605641404
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1605641404
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1605641404
transform 1 0 12972 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1605641404
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_133
timestamp 1605641404
transform 1 0 13340 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_145
timestamp 1605641404
transform 1 0 14444 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1605641404
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1605641404
transform 1 0 6624 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1605641404
transform 1 0 5152 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_48
timestamp 1605641404
transform 1 0 5520 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1605641404
transform 1 0 7176 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1605641404
transform 1 0 7728 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1605641404
transform 1 0 8280 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_64
timestamp 1605641404
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_70
timestamp 1605641404
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_76
timestamp 1605641404
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_82
timestamp 1605641404
transform 1 0 8648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1605641404
transform 1 0 10212 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1605641404
transform 1 0 8924 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1605641404
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1605641404
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_103
timestamp 1605641404
transform 1 0 10580 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1605641404
transform 1 0 11868 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_115
timestamp 1605641404
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1605641404
transform 1 0 12236 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_133
timestamp 1605641404
transform 1 0 13340 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_145
timestamp 1605641404
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1605641404
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1605641404
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1605641404
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1605641404
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1605641404
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1605641404
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1605641404
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1605641404
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1605641404
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_147
timestamp 1605641404
transform 1 0 14628 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_155
timestamp 1605641404
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1605641404
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1605641404
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1605641404
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1605641404
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1605641404
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1605641404
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1605641404
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1605641404
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1605641404
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1605641404
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1605641404
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1605641404
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1605641404
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1605641404
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1605641404
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1605641404
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1605641404
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1605641404
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1605641404
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1605641404
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_147
timestamp 1605641404
transform 1 0 14628 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1605641404
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1605641404
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1605641404
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_38
timestamp 1605641404
transform 1 0 4600 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_50
timestamp 1605641404
transform 1 0 5704 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1605641404
transform 1 0 6808 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_74
timestamp 1605641404
transform 1 0 7912 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_86
timestamp 1605641404
transform 1 0 9016 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1605641404
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1605641404
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1605641404
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1605641404
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1605641404
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1605641404
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1605641404
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1605641404
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1605641404
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1605641404
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1605641404
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1605641404
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1605641404
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1605641404
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_147
timestamp 1605641404
transform 1 0 14628 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_155
timestamp 1605641404
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1605641404
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1605641404
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1605641404
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1605641404
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1605641404
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1605641404
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1605641404
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1605641404
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1605641404
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1605641404
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1605641404
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1605641404
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1605641404
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1605641404
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1605641404
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_74
timestamp 1605641404
transform 1 0 7912 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_78
timestamp 1605641404
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _01_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_88
timestamp 1605641404
transform 1 0 9200 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_100
timestamp 1605641404
transform 1 0 10304 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_104
timestamp 1605641404
transform 1 0 10672 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_116
timestamp 1605641404
transform 1 0 11776 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1605641404
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_147
timestamp 1605641404
transform 1 0 14628 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1605641404
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1605641404
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1605641404
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6716 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1605641404
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_56
timestamp 1605641404
transform 1 0 6256 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_60
timestamp 1605641404
transform 1 0 6624 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7728 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_70
timestamp 1605641404
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10672 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1605641404
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1605641404
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_113
timestamp 1605641404
transform 1 0 11500 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_125
timestamp 1605641404
transform 1 0 12604 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_137
timestamp 1605641404
transform 1 0 13708 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1605641404
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1605641404
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1605641404
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1605641404
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1605641404
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1605641404
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_40
timestamp 1605641404
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6256 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5888 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4968 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_51
timestamp 1605641404
transform 1 0 5796 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_45
timestamp 1605641404
transform 1 0 5244 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_53
timestamp 1605641404
transform 1 0 5980 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8648 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7268 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7636 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_13_66
timestamp 1605641404
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_76
timestamp 1605641404
transform 1 0 8096 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1605641404
transform 1 0 7084 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 9844 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10304 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_98
timestamp 1605641404
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1605641404
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_109
timestamp 1605641404
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1605641404
transform 1 0 11592 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_111
timestamp 1605641404
transform 1 0 11316 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1605641404
transform 1 0 12420 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1605641404
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_135
timestamp 1605641404
transform 1 0 13524 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_147
timestamp 1605641404
transform 1 0 14628 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1605641404
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_147
timestamp 1605641404
transform 1 0 14628 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1605641404
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1605641404
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1605641404
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1605641404
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1605641404
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 7820 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 8648 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_70
timestamp 1605641404
transform 1 0 7544 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_91
timestamp 1605641404
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_103
timestamp 1605641404
transform 1 0 10580 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_115
timestamp 1605641404
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1605641404
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1605641404
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_147
timestamp 1605641404
transform 1 0 14628 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1605641404
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1605641404
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1605641404
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5336 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_44
timestamp 1605641404
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_62
timestamp 1605641404
transform 1 0 6808 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_74
timestamp 1605641404
transform 1 0 7912 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_86
timestamp 1605641404
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1605641404
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1605641404
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1605641404
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1605641404
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1605641404
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1605641404
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1605641404
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1605641404
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1605641404
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1605641404
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1605641404
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1605641404
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1605641404
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1605641404
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_147
timestamp 1605641404
transform 1 0 14628 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1605641404
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1605641404
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1605641404
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1605641404
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1605641404
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1605641404
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1605641404
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1605641404
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1605641404
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1605641404
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1605641404
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1605641404
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1605641404
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1605641404
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1605641404
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1605641404
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1605641404
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1605641404
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1605641404
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1605641404
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1605641404
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1605641404
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1605641404
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1605641404
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1605641404
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1605641404
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1605641404
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1605641404
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1605641404
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1605641404
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_147
timestamp 1605641404
transform 1 0 14628 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1605641404
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1605641404
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1605641404
transform 1 0 4416 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1605641404
transform 1 0 3680 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_27
timestamp 1605641404
transform 1 0 3588 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_32
timestamp 1605641404
transform 1 0 4048 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_40
timestamp 1605641404
transform 1 0 4784 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1605641404
transform 1 0 5152 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_48
timestamp 1605641404
transform 1 0 5520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1605641404
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _07_
timestamp 1605641404
transform 1 0 6992 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_68
timestamp 1605641404
transform 1 0 7360 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_80
timestamp 1605641404
transform 1 0 8464 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1605641404
transform 1 0 9016 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_90
timestamp 1605641404
transform 1 0 9384 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_102
timestamp 1605641404
transform 1 0 10488 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1605641404
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1605641404
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_147
timestamp 1605641404
transform 1 0 14628 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_155
timestamp 1605641404
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1605641404
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1605641404
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1605641404
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1605641404
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1605641404
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1605641404
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1605641404
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1605641404
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1605641404
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1605641404
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1605641404
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1605641404
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1605641404
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1605641404
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1605641404
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1605641404
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1605641404
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1605641404
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1605641404
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1605641404
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1605641404
transform 1 0 14628 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1605641404
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1605641404
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1605641404
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 6808 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1605641404
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_56
timestamp 1605641404
transform 1 0 6256 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_63
timestamp 1605641404
transform 1 0 6900 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_75
timestamp 1605641404
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_87
timestamp 1605641404
transform 1 0 9108 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_94
timestamp 1605641404
transform 1 0 9752 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 12512 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_106
timestamp 1605641404
transform 1 0 10856 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_118
timestamp 1605641404
transform 1 0 11960 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_125
timestamp 1605641404
transform 1 0 12604 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_137
timestamp 1605641404
transform 1 0 13708 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 15364 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_149
timestamp 1605641404
transform 1 0 14812 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_156
timestamp 1605641404
transform 1 0 15456 0 -1 15776
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 13472 480 13592 6 ccff_head
port 0 nsew default input
rlabel metal3 s 16520 13472 17000 13592 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 13818 0 13874 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 11242 0 11298 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 12070 0 12126 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4434 0 4490 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 7010 0 7066 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 1030 0 1086 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1858 0 1914 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2686 0 2742 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 3146 0 3202 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3974 0 4030 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8666 17520 8722 18000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12898 17520 12954 18000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 13358 17520 13414 18000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 13818 17520 13874 18000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 14186 17520 14242 18000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 14646 17520 14702 18000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 15014 17520 15070 18000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 15474 17520 15530 18000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 15934 17520 15990 18000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 16302 17520 16358 18000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 16762 17520 16818 18000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 9126 17520 9182 18000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 9494 17520 9550 18000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9954 17520 10010 18000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 10414 17520 10470 18000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10782 17520 10838 18000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 11242 17520 11298 18000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 11610 17520 11666 18000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 12070 17520 12126 18000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 12530 17520 12586 18000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 17520 258 18000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4434 17520 4490 18000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4802 17520 4858 18000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 5262 17520 5318 18000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5722 17520 5778 18000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 6090 17520 6146 18000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6550 17520 6606 18000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 7010 17520 7066 18000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 7378 17520 7434 18000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7838 17520 7894 18000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 8206 17520 8262 18000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 17520 626 18000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 1030 17520 1086 18000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 17520 1454 18000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1858 17520 1914 18000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2318 17520 2374 18000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2686 17520 2742 18000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 3146 17520 3202 18000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3606 17520 3662 18000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3974 17520 4030 18000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 4496 480 4616 6 left_grid_pin_0_
port 82 nsew default tristate
rlabel metal3 s 16520 4496 17000 4616 6 prog_clk
port 83 nsew default input
rlabel metal4 s 3409 2128 3729 15824 6 VPWR
port 84 nsew default input
rlabel metal4 s 5875 2128 6195 15824 6 VGND
port 85 nsew default input
<< properties >>
string FIXED_BBOX 0 0 17000 18000
<< end >>
