magic
tech EFS8A
magscale 1 2
timestamp 1602873129
<< locali >>
rect 5779 8041 5825 8075
rect 9781 7905 9942 7939
rect 14231 7905 14266 7939
rect 9781 7871 9815 7905
rect 16635 7497 16773 7531
rect 20223 7157 20361 7191
rect 12575 6817 12702 6851
rect 18279 6817 18314 6851
rect 18567 6409 18705 6443
rect 14007 6103 14041 6171
rect 14007 6069 14013 6103
rect 4439 5865 4445 5899
rect 6279 5865 6285 5899
rect 21275 5865 21281 5899
rect 4439 5797 4473 5865
rect 6279 5797 6313 5865
rect 21275 5797 21309 5865
rect 11621 5015 11655 5185
rect 11563 4981 11655 5015
rect 8211 4777 8217 4811
rect 24955 4777 24961 4811
rect 8211 4709 8245 4777
rect 11713 4675 11747 4777
rect 14105 4607 14139 4777
rect 24955 4709 24989 4777
rect 17693 3927 17727 4029
rect 2547 3553 2582 3587
rect 19441 3383 19475 3689
rect 27255 2601 27261 2635
rect 25973 2431 26007 2601
rect 27255 2533 27289 2601
rect 17417 2397 17543 2431
rect 17509 2295 17543 2397
rect 32229 2295 32263 2465
<< viali >>
rect 1593 11305 1627 11339
rect 35633 11305 35667 11339
rect 1409 11169 1443 11203
rect 35449 11169 35483 11203
rect 1685 10421 1719 10455
rect 35449 10421 35483 10455
rect 1593 10217 1627 10251
rect 35633 10217 35667 10251
rect 1409 10081 1443 10115
rect 35449 10081 35483 10115
rect 1685 9333 1719 9367
rect 35449 9333 35483 9367
rect 1593 9129 1627 9163
rect 35633 9129 35667 9163
rect 1409 8993 1443 9027
rect 2580 8993 2614 9027
rect 35449 8993 35483 9027
rect 2651 8789 2685 8823
rect 1593 8585 1627 8619
rect 35633 8585 35667 8619
rect 2421 8449 2455 8483
rect 1409 8381 1443 8415
rect 2564 8381 2598 8415
rect 3576 8381 3610 8415
rect 4077 8381 4111 8415
rect 4604 8381 4638 8415
rect 35449 8381 35483 8415
rect 36001 8381 36035 8415
rect 2651 8313 2685 8347
rect 3663 8313 3697 8347
rect 2053 8245 2087 8279
rect 2973 8245 3007 8279
rect 3341 8245 3375 8279
rect 4675 8245 4709 8279
rect 5089 8245 5123 8279
rect 35265 8245 35299 8279
rect 1593 8041 1627 8075
rect 5089 8041 5123 8075
rect 5825 8041 5859 8075
rect 35633 8041 35667 8075
rect 4261 7973 4295 8007
rect 1409 7905 1443 7939
rect 2513 7905 2547 7939
rect 5676 7905 5710 7939
rect 14197 7905 14231 7939
rect 19165 7905 19199 7939
rect 35449 7905 35483 7939
rect 4169 7837 4203 7871
rect 4813 7837 4847 7871
rect 9781 7837 9815 7871
rect 2697 7769 2731 7803
rect 3157 7701 3191 7735
rect 10011 7701 10045 7735
rect 14335 7701 14369 7735
rect 14657 7701 14691 7735
rect 19349 7701 19383 7735
rect 1593 7497 1627 7531
rect 5641 7497 5675 7531
rect 16773 7497 16807 7531
rect 35357 7497 35391 7531
rect 35633 7497 35667 7531
rect 36737 7497 36771 7531
rect 2605 7429 2639 7463
rect 4169 7429 4203 7463
rect 13507 7429 13541 7463
rect 2973 7361 3007 7395
rect 4721 7361 4755 7395
rect 4997 7361 5031 7395
rect 14473 7361 14507 7395
rect 36001 7361 36035 7395
rect 1409 7293 1443 7327
rect 10276 7293 10310 7327
rect 10701 7293 10735 7327
rect 13436 7293 13470 7327
rect 13829 7293 13863 7327
rect 16532 7293 16566 7327
rect 16957 7293 16991 7327
rect 19108 7293 19142 7327
rect 19901 7293 19935 7327
rect 20152 7293 20186 7327
rect 20545 7293 20579 7327
rect 21465 7293 21499 7327
rect 22201 7293 22235 7327
rect 35449 7293 35483 7327
rect 36553 7293 36587 7327
rect 2053 7225 2087 7259
rect 3157 7225 3191 7259
rect 3249 7225 3283 7259
rect 3801 7225 3835 7259
rect 4813 7225 4847 7259
rect 14565 7225 14599 7259
rect 15117 7225 15151 7259
rect 19211 7225 19245 7259
rect 22293 7225 22327 7259
rect 37105 7225 37139 7259
rect 4445 7157 4479 7191
rect 6009 7157 6043 7191
rect 9965 7157 9999 7191
rect 10379 7157 10413 7191
rect 14197 7157 14231 7191
rect 15485 7157 15519 7191
rect 18981 7157 19015 7191
rect 19625 7157 19659 7191
rect 20361 7157 20395 7191
rect 20913 7157 20947 7191
rect 23443 6953 23477 6987
rect 35633 6953 35667 6987
rect 2558 6885 2592 6919
rect 4261 6885 4295 6919
rect 5733 6885 5767 6919
rect 5825 6885 5859 6919
rect 10333 6885 10367 6919
rect 10425 6885 10459 6919
rect 13829 6885 13863 6919
rect 15485 6885 15519 6919
rect 19441 6885 19475 6919
rect 21097 6885 21131 6919
rect 12541 6817 12575 6851
rect 16865 6817 16899 6851
rect 18245 6817 18279 6851
rect 23372 6817 23406 6851
rect 24501 6817 24535 6851
rect 35449 6817 35483 6851
rect 2237 6749 2271 6783
rect 4169 6749 4203 6783
rect 4629 6749 4663 6783
rect 6009 6749 6043 6783
rect 6837 6749 6871 6783
rect 8585 6749 8619 6783
rect 12771 6749 12805 6783
rect 13185 6749 13219 6783
rect 13737 6749 13771 6783
rect 14381 6749 14415 6783
rect 15393 6749 15427 6783
rect 15669 6749 15703 6783
rect 19349 6749 19383 6783
rect 20637 6749 20671 6783
rect 21005 6749 21039 6783
rect 3433 6681 3467 6715
rect 10885 6681 10919 6715
rect 11345 6681 11379 6715
rect 18383 6681 18417 6715
rect 19901 6681 19935 6715
rect 21557 6681 21591 6715
rect 21925 6681 21959 6715
rect 1685 6613 1719 6647
rect 2145 6613 2179 6647
rect 3157 6613 3191 6647
rect 5089 6613 5123 6647
rect 13553 6613 13587 6647
rect 14749 6613 14783 6647
rect 15117 6613 15151 6647
rect 17049 6613 17083 6647
rect 18705 6613 18739 6647
rect 19073 6613 19107 6647
rect 20269 6613 20303 6647
rect 24593 6613 24627 6647
rect 25329 6613 25363 6647
rect 1593 6409 1627 6443
rect 2053 6409 2087 6443
rect 3433 6409 3467 6443
rect 4077 6409 4111 6443
rect 6009 6409 6043 6443
rect 8769 6409 8803 6443
rect 10333 6409 10367 6443
rect 15301 6409 15335 6443
rect 18337 6409 18371 6443
rect 18705 6409 18739 6443
rect 22385 6409 22419 6443
rect 23489 6409 23523 6443
rect 24501 6409 24535 6443
rect 2421 6341 2455 6375
rect 3801 6341 3835 6375
rect 5273 6341 5307 6375
rect 5641 6341 5675 6375
rect 9597 6341 9631 6375
rect 11161 6341 11195 6375
rect 12909 6341 12943 6375
rect 16037 6341 16071 6375
rect 20085 6341 20119 6375
rect 21649 6341 21683 6375
rect 4353 6273 4387 6307
rect 4629 6273 4663 6307
rect 6929 6273 6963 6307
rect 7205 6273 7239 6307
rect 9045 6273 9079 6307
rect 10609 6273 10643 6307
rect 15485 6273 15519 6307
rect 17095 6273 17129 6307
rect 19533 6273 19567 6307
rect 22017 6273 22051 6307
rect 23029 6273 23063 6307
rect 25421 6273 25455 6307
rect 35449 6273 35483 6307
rect 1409 6205 1443 6239
rect 2513 6205 2547 6239
rect 12265 6205 12299 6239
rect 12449 6205 12483 6239
rect 13645 6205 13679 6239
rect 17008 6205 17042 6239
rect 18496 6205 18530 6239
rect 18889 6205 18923 6239
rect 22636 6205 22670 6239
rect 2875 6137 2909 6171
rect 4445 6137 4479 6171
rect 7021 6137 7055 6171
rect 9137 6137 9171 6171
rect 10701 6137 10735 6171
rect 11529 6137 11563 6171
rect 13553 6137 13587 6171
rect 14933 6137 14967 6171
rect 15577 6137 15611 6171
rect 19625 6137 19659 6171
rect 20545 6137 20579 6171
rect 21097 6137 21131 6171
rect 21189 6137 21223 6171
rect 25145 6137 25179 6171
rect 25237 6137 25271 6171
rect 6561 6069 6595 6103
rect 12633 6069 12667 6103
rect 14013 6069 14047 6103
rect 14565 6069 14599 6103
rect 16405 6069 16439 6103
rect 16773 6069 16807 6103
rect 17509 6069 17543 6103
rect 17785 6069 17819 6103
rect 19257 6069 19291 6103
rect 20821 6069 20855 6103
rect 22707 6069 22741 6103
rect 24041 6069 24075 6103
rect 24961 6069 24995 6103
rect 3157 5865 3191 5899
rect 4445 5865 4479 5899
rect 6285 5865 6319 5899
rect 6837 5865 6871 5899
rect 9045 5865 9079 5899
rect 10333 5865 10367 5899
rect 14013 5865 14047 5899
rect 14289 5865 14323 5899
rect 18429 5865 18463 5899
rect 19165 5865 19199 5899
rect 21281 5865 21315 5899
rect 25421 5865 25455 5899
rect 2558 5797 2592 5831
rect 7849 5797 7883 5831
rect 10793 5797 10827 5831
rect 13455 5797 13489 5831
rect 15485 5797 15519 5831
rect 16313 5797 16347 5831
rect 17871 5797 17905 5831
rect 19349 5797 19383 5831
rect 19441 5797 19475 5831
rect 22569 5797 22603 5831
rect 22753 5797 22787 5831
rect 22845 5797 22879 5831
rect 24593 5797 24627 5831
rect 12541 5729 12575 5763
rect 19993 5729 20027 5763
rect 26617 5729 26651 5763
rect 2237 5661 2271 5695
rect 4077 5661 4111 5695
rect 5917 5661 5951 5695
rect 7757 5661 7791 5695
rect 8033 5661 8067 5695
rect 10701 5661 10735 5695
rect 13093 5661 13127 5695
rect 14657 5661 14691 5695
rect 15393 5661 15427 5695
rect 15669 5661 15703 5695
rect 17509 5661 17543 5695
rect 20913 5661 20947 5695
rect 23029 5661 23063 5695
rect 24501 5661 24535 5695
rect 24777 5661 24811 5695
rect 26525 5661 26559 5695
rect 11253 5593 11287 5627
rect 1777 5525 1811 5559
rect 2145 5525 2179 5559
rect 3433 5525 3467 5559
rect 3801 5525 3835 5559
rect 4997 5525 5031 5559
rect 7573 5525 7607 5559
rect 12817 5525 12851 5559
rect 15025 5525 15059 5559
rect 16773 5525 16807 5559
rect 17417 5525 17451 5559
rect 18797 5525 18831 5559
rect 20361 5525 20395 5559
rect 21833 5525 21867 5559
rect 22109 5525 22143 5559
rect 23673 5525 23707 5559
rect 27537 5525 27571 5559
rect 27905 5525 27939 5559
rect 1593 5321 1627 5355
rect 2421 5321 2455 5355
rect 5917 5321 5951 5355
rect 7389 5321 7423 5355
rect 8769 5321 8803 5355
rect 10517 5321 10551 5355
rect 10793 5321 10827 5355
rect 12265 5321 12299 5355
rect 15669 5321 15703 5355
rect 18981 5321 19015 5355
rect 20729 5321 20763 5355
rect 22937 5321 22971 5355
rect 23811 5321 23845 5355
rect 24593 5321 24627 5355
rect 27261 5321 27295 5355
rect 35633 5321 35667 5355
rect 9505 5253 9539 5287
rect 13829 5253 13863 5287
rect 14657 5253 14691 5287
rect 24225 5253 24259 5287
rect 25329 5253 25363 5287
rect 6837 5185 6871 5219
rect 7849 5185 7883 5219
rect 11161 5185 11195 5219
rect 11621 5185 11655 5219
rect 18061 5185 18095 5219
rect 21649 5185 21683 5219
rect 22293 5185 22327 5219
rect 24777 5185 24811 5219
rect 27537 5185 27571 5219
rect 1409 5117 1443 5151
rect 2053 5117 2087 5151
rect 2789 5117 2823 5151
rect 3065 5117 3099 5151
rect 3433 5117 3467 5151
rect 3893 5117 3927 5151
rect 4997 5117 5031 5151
rect 9137 5117 9171 5151
rect 9597 5117 9631 5151
rect 11345 5117 11379 5151
rect 5359 5049 5393 5083
rect 6285 5049 6319 5083
rect 7757 5049 7791 5083
rect 8211 5049 8245 5083
rect 9918 5049 9952 5083
rect 12449 5117 12483 5151
rect 12909 5117 12943 5151
rect 13277 5117 13311 5151
rect 13645 5117 13679 5151
rect 14749 5117 14783 5151
rect 16681 5117 16715 5151
rect 17325 5117 17359 5151
rect 19809 5117 19843 5151
rect 23740 5117 23774 5151
rect 26484 5117 26518 5151
rect 35449 5117 35483 5151
rect 36001 5117 36035 5151
rect 14197 5049 14231 5083
rect 15111 5049 15145 5083
rect 16313 5049 16347 5083
rect 16497 5049 16531 5083
rect 17049 5049 17083 5083
rect 18423 5049 18457 5083
rect 20171 5049 20205 5083
rect 21373 5049 21407 5083
rect 21741 5049 21775 5083
rect 24869 5049 24903 5083
rect 26571 5049 26605 5083
rect 27629 5049 27663 5083
rect 28181 5049 28215 5083
rect 2605 4981 2639 5015
rect 4353 4981 4387 5015
rect 4905 4981 4939 5015
rect 6653 4981 6687 5015
rect 11529 4981 11563 5015
rect 11805 4981 11839 5015
rect 15945 4981 15979 5015
rect 17877 4981 17911 5015
rect 19349 4981 19383 5015
rect 19717 4981 19751 5015
rect 21097 4981 21131 5015
rect 22661 4981 22695 5015
rect 23489 4981 23523 5015
rect 25697 4981 25731 5015
rect 26985 4981 27019 5015
rect 1961 4777 1995 4811
rect 3801 4777 3835 4811
rect 4537 4777 4571 4811
rect 5089 4777 5123 4811
rect 5273 4777 5307 4811
rect 7665 4777 7699 4811
rect 8217 4777 8251 4811
rect 8769 4777 8803 4811
rect 9781 4777 9815 4811
rect 11713 4777 11747 4811
rect 12265 4777 12299 4811
rect 13829 4777 13863 4811
rect 14105 4777 14139 4811
rect 14289 4777 14323 4811
rect 17601 4777 17635 4811
rect 20729 4777 20763 4811
rect 22109 4777 22143 4811
rect 23489 4777 23523 4811
rect 24041 4777 24075 4811
rect 24501 4777 24535 4811
rect 24961 4777 24995 4811
rect 25513 4777 25547 4811
rect 4215 4709 4249 4743
rect 1869 4641 1903 4675
rect 2421 4641 2455 4675
rect 2697 4641 2731 4675
rect 3065 4641 3099 4675
rect 4123 4641 4157 4675
rect 5181 4641 5215 4675
rect 5733 4641 5767 4675
rect 6193 4641 6227 4675
rect 6469 4641 6503 4675
rect 9781 4641 9815 4675
rect 10425 4641 10459 4675
rect 10609 4641 10643 4675
rect 11069 4641 11103 4675
rect 11713 4641 11747 4675
rect 12449 4641 12483 4675
rect 12909 4641 12943 4675
rect 13277 4641 13311 4675
rect 13737 4641 13771 4675
rect 15117 4709 15151 4743
rect 15761 4709 15795 4743
rect 19993 4709 20027 4743
rect 20269 4709 20303 4743
rect 21051 4709 21085 4743
rect 21373 4709 21407 4743
rect 27721 4709 27755 4743
rect 28273 4709 28307 4743
rect 16221 4641 16255 4675
rect 16957 4641 16991 4675
rect 17233 4641 17267 4675
rect 17417 4641 17451 4675
rect 18521 4641 18555 4675
rect 18981 4641 19015 4675
rect 19349 4641 19383 4675
rect 19717 4641 19751 4675
rect 20948 4641 20982 4675
rect 22293 4641 22327 4675
rect 22753 4641 22787 4675
rect 23121 4641 23155 4675
rect 23489 4641 23523 4675
rect 26560 4641 26594 4675
rect 29193 4641 29227 4675
rect 30732 4641 30766 4675
rect 7849 4573 7883 4607
rect 14105 4573 14139 4607
rect 16129 4573 16163 4607
rect 21833 4573 21867 4607
rect 24593 4573 24627 4607
rect 27629 4573 27663 4607
rect 3525 4505 3559 4539
rect 18061 4505 18095 4539
rect 18429 4505 18463 4539
rect 27353 4505 27387 4539
rect 9137 4437 9171 4471
rect 11529 4437 11563 4471
rect 11897 4437 11931 4471
rect 14657 4437 14691 4471
rect 26663 4437 26697 4471
rect 27077 4437 27111 4471
rect 29561 4437 29595 4471
rect 30803 4437 30837 4471
rect 2237 4233 2271 4267
rect 5733 4233 5767 4267
rect 6561 4233 6595 4267
rect 10517 4233 10551 4267
rect 10977 4233 11011 4267
rect 11529 4233 11563 4267
rect 21281 4233 21315 4267
rect 22017 4233 22051 4267
rect 24593 4233 24627 4267
rect 26433 4233 26467 4267
rect 28089 4233 28123 4267
rect 29101 4233 29135 4267
rect 29837 4233 29871 4267
rect 7205 4165 7239 4199
rect 12173 4165 12207 4199
rect 13829 4165 13863 4199
rect 14749 4165 14783 4199
rect 4813 4097 4847 4131
rect 5457 4097 5491 4131
rect 15485 4097 15519 4131
rect 17141 4097 17175 4131
rect 19901 4097 19935 4131
rect 23673 4097 23707 4131
rect 2421 4029 2455 4063
rect 3065 4029 3099 4063
rect 3249 4029 3283 4063
rect 3801 4029 3835 4063
rect 7941 4029 7975 4063
rect 8401 4029 8435 4063
rect 8861 4029 8895 4063
rect 9413 4029 9447 4063
rect 9597 4029 9631 4063
rect 11345 4029 11379 4063
rect 12449 4029 12483 4063
rect 12909 4029 12943 4063
rect 13277 4029 13311 4063
rect 13737 4029 13771 4063
rect 15669 4029 15703 4063
rect 16405 4029 16439 4063
rect 16681 4029 16715 4063
rect 16957 4029 16991 4063
rect 17693 4029 17727 4063
rect 18061 4029 18095 4063
rect 18797 4029 18831 4063
rect 19073 4029 19107 4063
rect 19441 4029 19475 4063
rect 20361 4029 20395 4063
rect 22109 4029 22143 4063
rect 25456 4029 25490 4063
rect 25559 4029 25593 4063
rect 26525 4029 26559 4063
rect 27445 4029 27479 4063
rect 29336 4029 29370 4063
rect 31401 4029 31435 4063
rect 4905 3961 4939 3995
rect 7481 3961 7515 3995
rect 20269 3961 20303 3995
rect 20723 3961 20757 3995
rect 22661 3961 22695 3995
rect 23489 3961 23523 3995
rect 24035 3961 24069 3995
rect 25237 3961 25271 3995
rect 26887 3961 26921 3995
rect 29423 3961 29457 3995
rect 30389 3961 30423 3995
rect 30481 3961 30515 3995
rect 31033 3961 31067 3995
rect 1961 3893 1995 3927
rect 2513 3893 2547 3927
rect 4261 3893 4295 3927
rect 4629 3893 4663 3927
rect 6101 3893 6135 3927
rect 8217 3893 8251 3927
rect 8493 3893 8527 3927
rect 10241 3893 10275 3927
rect 11805 3893 11839 3927
rect 14473 3893 14507 3927
rect 15209 3893 15243 3927
rect 17417 3893 17451 3927
rect 17693 3893 17727 3927
rect 17785 3893 17819 3927
rect 18153 3893 18187 3927
rect 21649 3893 21683 3927
rect 22293 3893 22327 3927
rect 23029 3893 23063 3927
rect 24961 3893 24995 3927
rect 25973 3893 26007 3927
rect 27813 3893 27847 3927
rect 30113 3893 30147 3927
rect 2651 3689 2685 3723
rect 4813 3689 4847 3723
rect 5089 3689 5123 3723
rect 6653 3689 6687 3723
rect 9137 3689 9171 3723
rect 9873 3689 9907 3723
rect 12541 3689 12575 3723
rect 13277 3689 13311 3723
rect 16313 3689 16347 3723
rect 16681 3689 16715 3723
rect 17417 3689 17451 3723
rect 19257 3689 19291 3723
rect 19441 3689 19475 3723
rect 25881 3689 25915 3723
rect 27445 3689 27479 3723
rect 28181 3689 28215 3723
rect 30389 3689 30423 3723
rect 2145 3621 2179 3655
rect 2973 3621 3007 3655
rect 12909 3621 12943 3655
rect 16037 3621 16071 3655
rect 18981 3621 19015 3655
rect 2513 3553 2547 3587
rect 3433 3553 3467 3587
rect 5273 3553 5307 3587
rect 5733 3553 5767 3587
rect 6101 3553 6135 3587
rect 6469 3553 6503 3587
rect 8677 3553 8711 3587
rect 9689 3553 9723 3587
rect 10149 3553 10183 3587
rect 11805 3553 11839 3587
rect 14289 3553 14323 3587
rect 15117 3553 15151 3587
rect 15301 3553 15335 3587
rect 17509 3553 17543 3587
rect 17969 3553 18003 3587
rect 18521 3553 18555 3587
rect 18889 3553 18923 3587
rect 7849 3485 7883 3519
rect 8769 3485 8803 3519
rect 11897 3485 11931 3519
rect 14381 3485 14415 3519
rect 15669 3485 15703 3519
rect 1777 3417 1811 3451
rect 11069 3417 11103 3451
rect 15466 3417 15500 3451
rect 21097 3621 21131 3655
rect 21649 3621 21683 3655
rect 23949 3621 23983 3655
rect 24961 3621 24995 3655
rect 25053 3621 25087 3655
rect 26887 3621 26921 3655
rect 28365 3621 28399 3655
rect 28457 3621 28491 3655
rect 30021 3621 30055 3655
rect 30573 3621 30607 3655
rect 30665 3621 30699 3655
rect 32137 3621 32171 3655
rect 22017 3553 22051 3587
rect 22477 3553 22511 3587
rect 23213 3553 23247 3587
rect 23305 3553 23339 3587
rect 23673 3553 23707 3587
rect 32229 3553 32263 3587
rect 19809 3485 19843 3519
rect 21005 3485 21039 3519
rect 24593 3485 24627 3519
rect 25237 3485 25271 3519
rect 26525 3485 26559 3519
rect 31033 3485 31067 3519
rect 20361 3417 20395 3451
rect 28917 3417 28951 3451
rect 14749 3349 14783 3383
rect 15577 3349 15611 3383
rect 19441 3349 19475 3383
rect 19717 3349 19751 3383
rect 20637 3349 20671 3383
rect 22293 3349 22327 3383
rect 24225 3349 24259 3383
rect 26249 3349 26283 3383
rect 29285 3349 29319 3383
rect 33149 3349 33183 3383
rect 4813 3145 4847 3179
rect 5181 3145 5215 3179
rect 7205 3145 7239 3179
rect 17141 3145 17175 3179
rect 17509 3145 17543 3179
rect 20269 3145 20303 3179
rect 20545 3145 20579 3179
rect 25421 3145 25455 3179
rect 27169 3145 27203 3179
rect 28549 3145 28583 3179
rect 30573 3145 30607 3179
rect 32229 3145 32263 3179
rect 13737 3077 13771 3111
rect 14657 3077 14691 3111
rect 15485 3077 15519 3111
rect 21097 3077 21131 3111
rect 22661 3077 22695 3111
rect 29009 3077 29043 3111
rect 4169 3009 4203 3043
rect 5825 3009 5859 3043
rect 7481 3009 7515 3043
rect 11529 3009 11563 3043
rect 12449 3009 12483 3043
rect 14289 3009 14323 3043
rect 14749 3009 14783 3043
rect 15945 3009 15979 3043
rect 25145 3009 25179 3043
rect 27813 3009 27847 3043
rect 29285 3009 29319 3043
rect 31585 3009 31619 3043
rect 32781 3009 32815 3043
rect 1777 2941 1811 2975
rect 2973 2941 3007 2975
rect 3341 2941 3375 2975
rect 3525 2941 3559 2975
rect 4077 2941 4111 2975
rect 4445 2941 4479 2975
rect 4997 2941 5031 2975
rect 6653 2941 6687 2975
rect 7021 2941 7055 2975
rect 8033 2941 8067 2975
rect 8493 2941 8527 2975
rect 8861 2941 8895 2975
rect 9229 2941 9263 2975
rect 11161 2941 11195 2975
rect 11897 2941 11931 2975
rect 12725 2941 12759 2975
rect 14528 2941 14562 2975
rect 15853 2941 15887 2975
rect 16589 2941 16623 2975
rect 18061 2941 18095 2975
rect 18521 2941 18555 2975
rect 19073 2941 19107 2975
rect 19441 2941 19475 2975
rect 21557 2941 21591 2975
rect 21741 2941 21775 2975
rect 22109 2941 22143 2975
rect 22477 2941 22511 2975
rect 23397 2941 23431 2975
rect 23673 2941 23707 2975
rect 24133 2941 24167 2975
rect 24501 2941 24535 2975
rect 24869 2941 24903 2975
rect 26249 2941 26283 2975
rect 29377 2941 29411 2975
rect 2237 2873 2271 2907
rect 10885 2873 10919 2907
rect 10977 2873 11011 2907
rect 14381 2873 14415 2907
rect 15117 2873 15151 2907
rect 19809 2873 19843 2907
rect 26570 2873 26604 2907
rect 30941 2873 30975 2907
rect 31033 2873 31067 2907
rect 32505 2873 32539 2907
rect 32597 2873 32631 2907
rect 33425 2873 33459 2907
rect 2605 2805 2639 2839
rect 5457 2805 5491 2839
rect 7941 2805 7975 2839
rect 8125 2805 8159 2839
rect 9781 2805 9815 2839
rect 12173 2805 12207 2839
rect 18337 2805 18371 2839
rect 23121 2805 23155 2839
rect 26157 2805 26191 2839
rect 27445 2805 27479 2839
rect 28089 2805 28123 2839
rect 3065 2601 3099 2635
rect 3525 2601 3559 2635
rect 7573 2601 7607 2635
rect 7849 2601 7883 2635
rect 8493 2601 8527 2635
rect 8861 2601 8895 2635
rect 12449 2601 12483 2635
rect 12817 2601 12851 2635
rect 13737 2601 13771 2635
rect 14933 2601 14967 2635
rect 15301 2601 15335 2635
rect 15669 2601 15703 2635
rect 17693 2601 17727 2635
rect 18153 2601 18187 2635
rect 19901 2601 19935 2635
rect 20637 2601 20671 2635
rect 21005 2601 21039 2635
rect 21557 2601 21591 2635
rect 25789 2601 25823 2635
rect 25973 2601 26007 2635
rect 26157 2601 26191 2635
rect 26617 2601 26651 2635
rect 27261 2601 27295 2635
rect 29101 2601 29135 2635
rect 29561 2601 29595 2635
rect 32045 2601 32079 2635
rect 2789 2533 2823 2567
rect 5273 2533 5307 2567
rect 15945 2533 15979 2567
rect 16313 2533 16347 2567
rect 16865 2533 16899 2567
rect 18658 2533 18692 2567
rect 19625 2533 19659 2567
rect 23121 2533 23155 2567
rect 1777 2465 1811 2499
rect 7665 2465 7699 2499
rect 8677 2465 8711 2499
rect 9137 2465 9171 2499
rect 10793 2465 10827 2499
rect 12633 2465 12667 2499
rect 13369 2465 13403 2499
rect 13829 2465 13863 2499
rect 13976 2465 14010 2499
rect 15485 2465 15519 2499
rect 18337 2465 18371 2499
rect 20152 2465 20186 2499
rect 21925 2465 21959 2499
rect 22109 2465 22143 2499
rect 22477 2465 22511 2499
rect 23029 2465 23063 2499
rect 24041 2465 24075 2499
rect 24501 2465 24535 2499
rect 24961 2465 24995 2499
rect 25237 2465 25271 2499
rect 25513 2465 25547 2499
rect 29837 2533 29871 2567
rect 29929 2533 29963 2567
rect 31309 2533 31343 2567
rect 34161 2533 34195 2567
rect 26893 2465 26927 2499
rect 27813 2465 27847 2499
rect 28708 2465 28742 2499
rect 31560 2465 31594 2499
rect 32229 2465 32263 2499
rect 32689 2465 32723 2499
rect 11437 2397 11471 2431
rect 12081 2397 12115 2431
rect 14194 2397 14228 2431
rect 14289 2397 14323 2431
rect 16773 2397 16807 2431
rect 23857 2397 23891 2431
rect 25973 2397 26007 2431
rect 28089 2397 28123 2431
rect 30113 2397 30147 2431
rect 30941 2397 30975 2431
rect 8217 2329 8251 2363
rect 19257 2329 19291 2363
rect 20223 2329 20257 2363
rect 28457 2329 28491 2363
rect 31631 2329 31665 2363
rect 32597 2397 32631 2431
rect 10517 2261 10551 2295
rect 14105 2261 14139 2295
rect 17509 2261 17543 2295
rect 23397 2261 23431 2295
rect 28779 2261 28813 2295
rect 32229 2261 32263 2295
rect 32321 2261 32355 2295
<< metal1 >>
rect 5810 15512 5816 15564
rect 5868 15552 5874 15564
rect 6638 15552 6644 15564
rect 5868 15524 6644 15552
rect 5868 15512 5874 15524
rect 6638 15512 6644 15524
rect 6696 15512 6702 15564
rect 19978 15512 19984 15564
rect 20036 15552 20042 15564
rect 20622 15552 20628 15564
rect 20036 15524 20628 15552
rect 20036 15512 20042 15524
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 35618 11336 35624 11348
rect 35579 11308 35624 11336
rect 35618 11296 35624 11308
rect 35676 11296 35682 11348
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 35434 11200 35440 11212
rect 35395 11172 35440 11200
rect 35434 11160 35440 11172
rect 35492 11160 35498 11212
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 1394 10412 1400 10464
rect 1452 10452 1458 10464
rect 1673 10455 1731 10461
rect 1673 10452 1685 10455
rect 1452 10424 1685 10452
rect 1452 10412 1458 10424
rect 1673 10421 1685 10424
rect 1719 10452 1731 10455
rect 2222 10452 2228 10464
rect 1719 10424 2228 10452
rect 1719 10421 1731 10424
rect 1673 10415 1731 10421
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 29822 10412 29828 10464
rect 29880 10452 29886 10464
rect 35434 10452 35440 10464
rect 29880 10424 35440 10452
rect 29880 10412 29886 10424
rect 35434 10412 35440 10424
rect 35492 10412 35498 10464
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 35618 10248 35624 10260
rect 35579 10220 35624 10248
rect 35618 10208 35624 10220
rect 35676 10208 35682 10260
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1670 10112 1676 10124
rect 1443 10084 1676 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 35434 10112 35440 10124
rect 35395 10084 35440 10112
rect 35434 10072 35440 10084
rect 35492 10072 35498 10124
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 1670 9364 1676 9376
rect 1631 9336 1676 9364
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 35434 9364 35440 9376
rect 35395 9336 35440 9364
rect 35434 9324 35440 9336
rect 35492 9324 35498 9376
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 35618 9160 35624 9172
rect 35579 9132 35624 9160
rect 35618 9120 35624 9132
rect 35676 9120 35682 9172
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2130 9024 2136 9036
rect 1443 8996 2136 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2130 8984 2136 8996
rect 2188 8984 2194 9036
rect 2222 8984 2228 9036
rect 2280 9024 2286 9036
rect 2568 9027 2626 9033
rect 2568 9024 2580 9027
rect 2280 8996 2580 9024
rect 2280 8984 2286 8996
rect 2568 8993 2580 8996
rect 2614 9024 2626 9027
rect 3326 9024 3332 9036
rect 2614 8996 3332 9024
rect 2614 8993 2626 8996
rect 2568 8987 2626 8993
rect 3326 8984 3332 8996
rect 3384 8984 3390 9036
rect 35250 8984 35256 9036
rect 35308 9024 35314 9036
rect 35437 9027 35495 9033
rect 35437 9024 35449 9027
rect 35308 8996 35449 9024
rect 35308 8984 35314 8996
rect 35437 8993 35449 8996
rect 35483 8993 35495 9027
rect 35437 8987 35495 8993
rect 2639 8823 2697 8829
rect 2639 8789 2651 8823
rect 2685 8820 2697 8823
rect 4982 8820 4988 8832
rect 2685 8792 4988 8820
rect 2685 8789 2697 8792
rect 2639 8783 2697 8789
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 1210 8576 1216 8628
rect 1268 8616 1274 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1268 8588 1593 8616
rect 1268 8576 1274 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 35618 8616 35624 8628
rect 35579 8588 35624 8616
rect 1581 8579 1639 8585
rect 35618 8576 35624 8588
rect 35676 8576 35682 8628
rect 2409 8483 2467 8489
rect 2409 8480 2421 8483
rect 1412 8452 2421 8480
rect 1412 8421 1440 8452
rect 2409 8449 2421 8452
rect 2455 8480 2467 8483
rect 2455 8452 4635 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 2552 8415 2610 8421
rect 2552 8381 2564 8415
rect 2598 8412 2610 8415
rect 3564 8415 3622 8421
rect 2598 8381 2611 8412
rect 2552 8375 2611 8381
rect 3564 8381 3576 8415
rect 3610 8412 3622 8415
rect 4062 8412 4068 8424
rect 3610 8384 4068 8412
rect 3610 8381 3622 8384
rect 3564 8375 3622 8381
rect 2041 8279 2099 8285
rect 2041 8245 2053 8279
rect 2087 8276 2099 8279
rect 2130 8276 2136 8288
rect 2087 8248 2136 8276
rect 2087 8245 2099 8248
rect 2041 8239 2099 8245
rect 2130 8236 2136 8248
rect 2188 8236 2194 8288
rect 2583 8276 2611 8375
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4607 8421 4635 8452
rect 4592 8415 4650 8421
rect 4592 8381 4604 8415
rect 4638 8412 4650 8415
rect 4638 8384 5120 8412
rect 4638 8381 4650 8384
rect 4592 8375 4650 8381
rect 2639 8347 2697 8353
rect 2639 8313 2651 8347
rect 2685 8344 2697 8347
rect 3418 8344 3424 8356
rect 2685 8316 3424 8344
rect 2685 8313 2697 8316
rect 2639 8307 2697 8313
rect 3418 8304 3424 8316
rect 3476 8304 3482 8356
rect 3651 8347 3709 8353
rect 3651 8313 3663 8347
rect 3697 8344 3709 8347
rect 4338 8344 4344 8356
rect 3697 8316 4344 8344
rect 3697 8313 3709 8316
rect 3651 8307 3709 8313
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 5092 8288 5120 8384
rect 34054 8372 34060 8424
rect 34112 8412 34118 8424
rect 35437 8415 35495 8421
rect 35437 8412 35449 8415
rect 34112 8384 35449 8412
rect 34112 8372 34118 8384
rect 35437 8381 35449 8384
rect 35483 8412 35495 8415
rect 35989 8415 36047 8421
rect 35989 8412 36001 8415
rect 35483 8384 36001 8412
rect 35483 8381 35495 8384
rect 35437 8375 35495 8381
rect 35989 8381 36001 8384
rect 36035 8381 36047 8415
rect 35989 8375 36047 8381
rect 2958 8276 2964 8288
rect 2583 8248 2964 8276
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 3326 8276 3332 8288
rect 3287 8248 3332 8276
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 4663 8279 4721 8285
rect 4663 8245 4675 8279
rect 4709 8276 4721 8279
rect 4798 8276 4804 8288
rect 4709 8248 4804 8276
rect 4709 8245 4721 8248
rect 4663 8239 4721 8245
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 5074 8276 5080 8288
rect 5035 8248 5080 8276
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 34146 8236 34152 8288
rect 34204 8276 34210 8288
rect 35250 8276 35256 8288
rect 34204 8248 35256 8276
rect 34204 8236 34210 8248
rect 35250 8236 35256 8248
rect 35308 8236 35314 8288
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 5040 8044 5089 8072
rect 5040 8032 5046 8044
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 5810 8072 5816 8084
rect 5771 8044 5816 8072
rect 5077 8035 5135 8041
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 35621 8075 35679 8081
rect 35621 8041 35633 8075
rect 35667 8072 35679 8075
rect 35710 8072 35716 8084
rect 35667 8044 35716 8072
rect 35667 8041 35679 8044
rect 35621 8035 35679 8041
rect 35710 8032 35716 8044
rect 35768 8032 35774 8084
rect 4154 7964 4160 8016
rect 4212 8004 4218 8016
rect 4249 8007 4307 8013
rect 4249 8004 4261 8007
rect 4212 7976 4261 8004
rect 4212 7964 4218 7976
rect 4249 7973 4261 7976
rect 4295 7973 4307 8007
rect 4249 7967 4307 7973
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 2038 7936 2044 7948
rect 1443 7908 2044 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 2498 7936 2504 7948
rect 2459 7908 2504 7936
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 5664 7939 5722 7945
rect 5664 7936 5676 7939
rect 5500 7908 5676 7936
rect 5500 7896 5506 7908
rect 5664 7905 5676 7908
rect 5710 7905 5722 7939
rect 14182 7936 14188 7948
rect 14143 7908 14188 7936
rect 5664 7899 5722 7905
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 19153 7939 19211 7945
rect 19153 7905 19165 7939
rect 19199 7936 19211 7939
rect 19610 7936 19616 7948
rect 19199 7908 19616 7936
rect 19199 7905 19211 7908
rect 19153 7899 19211 7905
rect 19610 7896 19616 7908
rect 19668 7896 19674 7948
rect 35434 7936 35440 7948
rect 35395 7908 35440 7936
rect 35434 7896 35440 7908
rect 35492 7896 35498 7948
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 4338 7868 4344 7880
rect 4203 7840 4344 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 4982 7868 4988 7880
rect 4847 7840 4988 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7868 9827 7871
rect 9950 7868 9956 7880
rect 9815 7840 9956 7868
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 2682 7800 2688 7812
rect 2643 7772 2688 7800
rect 2682 7760 2688 7772
rect 2740 7760 2746 7812
rect 3142 7732 3148 7744
rect 3103 7704 3148 7732
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 9999 7735 10057 7741
rect 9999 7701 10011 7735
rect 10045 7732 10057 7735
rect 10318 7732 10324 7744
rect 10045 7704 10324 7732
rect 10045 7701 10057 7704
rect 9999 7695 10057 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 14323 7735 14381 7741
rect 14323 7701 14335 7735
rect 14369 7732 14381 7735
rect 14458 7732 14464 7744
rect 14369 7704 14464 7732
rect 14369 7701 14381 7704
rect 14323 7695 14381 7701
rect 14458 7692 14464 7704
rect 14516 7732 14522 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 14516 7704 14657 7732
rect 14516 7692 14522 7704
rect 14645 7701 14657 7704
rect 14691 7701 14703 7735
rect 14645 7695 14703 7701
rect 19337 7735 19395 7741
rect 19337 7701 19349 7735
rect 19383 7732 19395 7735
rect 22002 7732 22008 7744
rect 19383 7704 22008 7732
rect 19383 7701 19395 7704
rect 19337 7695 19395 7701
rect 22002 7692 22008 7704
rect 22060 7692 22066 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 1486 7488 1492 7540
rect 1544 7528 1550 7540
rect 1581 7531 1639 7537
rect 1581 7528 1593 7531
rect 1544 7500 1593 7528
rect 1544 7488 1550 7500
rect 1581 7497 1593 7500
rect 1627 7497 1639 7531
rect 1581 7491 1639 7497
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 5629 7531 5687 7537
rect 5629 7528 5641 7531
rect 4396 7500 5641 7528
rect 4396 7488 4402 7500
rect 5629 7497 5641 7500
rect 5675 7497 5687 7531
rect 16758 7528 16764 7540
rect 16719 7500 16764 7528
rect 5629 7491 5687 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 35345 7531 35403 7537
rect 35345 7497 35357 7531
rect 35391 7528 35403 7531
rect 35434 7528 35440 7540
rect 35391 7500 35440 7528
rect 35391 7497 35403 7500
rect 35345 7491 35403 7497
rect 35434 7488 35440 7500
rect 35492 7488 35498 7540
rect 35526 7488 35532 7540
rect 35584 7528 35590 7540
rect 35621 7531 35679 7537
rect 35621 7528 35633 7531
rect 35584 7500 35633 7528
rect 35584 7488 35590 7500
rect 35621 7497 35633 7500
rect 35667 7497 35679 7531
rect 36722 7528 36728 7540
rect 36683 7500 36728 7528
rect 35621 7491 35679 7497
rect 36722 7488 36728 7500
rect 36780 7488 36786 7540
rect 2498 7420 2504 7472
rect 2556 7460 2562 7472
rect 2593 7463 2651 7469
rect 2593 7460 2605 7463
rect 2556 7432 2605 7460
rect 2556 7420 2562 7432
rect 2593 7429 2605 7432
rect 2639 7460 2651 7463
rect 3602 7460 3608 7472
rect 2639 7432 3608 7460
rect 2639 7429 2651 7432
rect 2593 7423 2651 7429
rect 3602 7420 3608 7432
rect 3660 7420 3666 7472
rect 4154 7420 4160 7472
rect 4212 7460 4218 7472
rect 4890 7460 4896 7472
rect 4212 7432 4257 7460
rect 4724 7432 4896 7460
rect 4212 7420 4218 7432
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3234 7392 3240 7404
rect 3007 7364 3240 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3234 7352 3240 7364
rect 3292 7392 3298 7404
rect 4172 7392 4200 7420
rect 4724 7401 4752 7432
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 13495 7463 13553 7469
rect 13495 7429 13507 7463
rect 13541 7460 13553 7463
rect 15378 7460 15384 7472
rect 13541 7432 15384 7460
rect 13541 7429 13553 7432
rect 13495 7423 13553 7429
rect 15378 7420 15384 7432
rect 15436 7420 15442 7472
rect 3292 7364 4200 7392
rect 4709 7395 4767 7401
rect 3292 7352 3298 7364
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4982 7392 4988 7404
rect 4943 7364 4988 7392
rect 4709 7355 4767 7361
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 14458 7392 14464 7404
rect 14419 7364 14464 7392
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 14918 7352 14924 7404
rect 14976 7392 14982 7404
rect 35986 7392 35992 7404
rect 14976 7364 20208 7392
rect 14976 7352 14982 7364
rect 20180 7336 20208 7364
rect 35452 7364 35992 7392
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 1670 7324 1676 7336
rect 1443 7296 1676 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 5350 7284 5356 7336
rect 5408 7324 5414 7336
rect 10264 7327 10322 7333
rect 10264 7324 10276 7327
rect 5408 7296 10276 7324
rect 5408 7284 5414 7296
rect 10264 7293 10276 7296
rect 10310 7324 10322 7327
rect 10686 7324 10692 7336
rect 10310 7296 10692 7324
rect 10310 7293 10322 7296
rect 10264 7287 10322 7293
rect 10686 7284 10692 7296
rect 10744 7284 10750 7336
rect 13424 7327 13482 7333
rect 13424 7293 13436 7327
rect 13470 7324 13482 7327
rect 13630 7324 13636 7336
rect 13470 7296 13636 7324
rect 13470 7293 13482 7296
rect 13424 7287 13482 7293
rect 13630 7284 13636 7296
rect 13688 7324 13694 7336
rect 13817 7327 13875 7333
rect 13817 7324 13829 7327
rect 13688 7296 13829 7324
rect 13688 7284 13694 7296
rect 13817 7293 13829 7296
rect 13863 7293 13875 7327
rect 13817 7287 13875 7293
rect 15194 7284 15200 7336
rect 15252 7324 15258 7336
rect 16520 7327 16578 7333
rect 16520 7324 16532 7327
rect 15252 7296 16532 7324
rect 15252 7284 15258 7296
rect 16520 7293 16532 7296
rect 16566 7324 16578 7327
rect 16945 7327 17003 7333
rect 16945 7324 16957 7327
rect 16566 7296 16957 7324
rect 16566 7293 16578 7296
rect 16520 7287 16578 7293
rect 16945 7293 16957 7296
rect 16991 7293 17003 7327
rect 16945 7287 17003 7293
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 19096 7327 19154 7333
rect 19096 7324 19108 7327
rect 18932 7296 19108 7324
rect 18932 7284 18938 7296
rect 19096 7293 19108 7296
rect 19142 7324 19154 7327
rect 19889 7327 19947 7333
rect 19889 7324 19901 7327
rect 19142 7296 19901 7324
rect 19142 7293 19154 7296
rect 19096 7287 19154 7293
rect 19889 7293 19901 7296
rect 19935 7324 19947 7327
rect 19978 7324 19984 7336
rect 19935 7296 19984 7324
rect 19935 7293 19947 7296
rect 19889 7287 19947 7293
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 20162 7333 20168 7336
rect 20140 7327 20168 7333
rect 20140 7324 20152 7327
rect 20075 7296 20152 7324
rect 20140 7293 20152 7296
rect 20220 7324 20226 7336
rect 20533 7327 20591 7333
rect 20533 7324 20545 7327
rect 20220 7296 20545 7324
rect 20140 7287 20168 7293
rect 20162 7284 20168 7287
rect 20220 7284 20226 7296
rect 20533 7293 20545 7296
rect 20579 7293 20591 7327
rect 20533 7287 20591 7293
rect 21453 7327 21511 7333
rect 21453 7293 21465 7327
rect 21499 7324 21511 7327
rect 22189 7327 22247 7333
rect 22189 7324 22201 7327
rect 21499 7296 22201 7324
rect 21499 7293 21511 7296
rect 21453 7287 21511 7293
rect 22189 7293 22201 7296
rect 22235 7324 22247 7327
rect 22738 7324 22744 7336
rect 22235 7296 22744 7324
rect 22235 7293 22247 7296
rect 22189 7287 22247 7293
rect 22738 7284 22744 7296
rect 22796 7284 22802 7336
rect 35452 7333 35480 7364
rect 35986 7352 35992 7364
rect 36044 7352 36050 7404
rect 35437 7327 35495 7333
rect 35437 7293 35449 7327
rect 35483 7293 35495 7327
rect 35437 7287 35495 7293
rect 36541 7327 36599 7333
rect 36541 7293 36553 7327
rect 36587 7293 36599 7327
rect 36541 7287 36599 7293
rect 2038 7256 2044 7268
rect 1999 7228 2044 7256
rect 2038 7216 2044 7228
rect 2096 7216 2102 7268
rect 3142 7256 3148 7268
rect 3055 7228 3148 7256
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 3234 7216 3240 7268
rect 3292 7256 3298 7268
rect 3789 7259 3847 7265
rect 3292 7228 3337 7256
rect 3292 7216 3298 7228
rect 3789 7225 3801 7259
rect 3835 7256 3847 7259
rect 4522 7256 4528 7268
rect 3835 7228 4528 7256
rect 3835 7225 3847 7228
rect 3789 7219 3847 7225
rect 4522 7216 4528 7228
rect 4580 7216 4586 7268
rect 4801 7259 4859 7265
rect 4801 7225 4813 7259
rect 4847 7225 4859 7259
rect 4801 7219 4859 7225
rect 14553 7259 14611 7265
rect 14553 7225 14565 7259
rect 14599 7256 14611 7259
rect 14826 7256 14832 7268
rect 14599 7228 14832 7256
rect 14599 7225 14611 7228
rect 14553 7219 14611 7225
rect 3160 7188 3188 7216
rect 3510 7188 3516 7200
rect 3160 7160 3516 7188
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 4062 7148 4068 7200
rect 4120 7188 4126 7200
rect 4433 7191 4491 7197
rect 4433 7188 4445 7191
rect 4120 7160 4445 7188
rect 4120 7148 4126 7160
rect 4433 7157 4445 7160
rect 4479 7188 4491 7191
rect 4816 7188 4844 7219
rect 14826 7216 14832 7228
rect 14884 7216 14890 7268
rect 15105 7259 15163 7265
rect 15105 7225 15117 7259
rect 15151 7225 15163 7259
rect 15105 7219 15163 7225
rect 19199 7259 19257 7265
rect 19199 7225 19211 7259
rect 19245 7256 19257 7259
rect 21266 7256 21272 7268
rect 19245 7228 21272 7256
rect 19245 7225 19257 7228
rect 19199 7219 19257 7225
rect 4479 7160 4844 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 5442 7148 5448 7200
rect 5500 7188 5506 7200
rect 5997 7191 6055 7197
rect 5997 7188 6009 7191
rect 5500 7160 6009 7188
rect 5500 7148 5506 7160
rect 5997 7157 6009 7160
rect 6043 7188 6055 7191
rect 7190 7188 7196 7200
rect 6043 7160 7196 7188
rect 6043 7157 6055 7160
rect 5997 7151 6055 7157
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 9950 7188 9956 7200
rect 9911 7160 9956 7188
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 10367 7191 10425 7197
rect 10367 7157 10379 7191
rect 10413 7188 10425 7191
rect 10502 7188 10508 7200
rect 10413 7160 10508 7188
rect 10413 7157 10425 7160
rect 10367 7151 10425 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 14182 7188 14188 7200
rect 14143 7160 14188 7188
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 15120 7188 15148 7219
rect 21266 7216 21272 7228
rect 21324 7216 21330 7268
rect 22281 7259 22339 7265
rect 22281 7225 22293 7259
rect 22327 7256 22339 7259
rect 23934 7256 23940 7268
rect 22327 7228 23940 7256
rect 22327 7225 22339 7228
rect 22281 7219 22339 7225
rect 23934 7216 23940 7228
rect 23992 7216 23998 7268
rect 26142 7216 26148 7268
rect 26200 7256 26206 7268
rect 36556 7256 36584 7287
rect 37093 7259 37151 7265
rect 37093 7256 37105 7259
rect 26200 7228 37105 7256
rect 26200 7216 26206 7228
rect 37093 7225 37105 7228
rect 37139 7225 37151 7259
rect 37093 7219 37151 7225
rect 15473 7191 15531 7197
rect 15473 7188 15485 7191
rect 15120 7160 15485 7188
rect 15473 7157 15485 7160
rect 15519 7188 15531 7191
rect 15562 7188 15568 7200
rect 15519 7160 15568 7188
rect 15519 7157 15531 7160
rect 15473 7151 15531 7157
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 18966 7188 18972 7200
rect 18927 7160 18972 7188
rect 18966 7148 18972 7160
rect 19024 7148 19030 7200
rect 19610 7188 19616 7200
rect 19571 7160 19616 7188
rect 19610 7148 19616 7160
rect 19668 7148 19674 7200
rect 20346 7188 20352 7200
rect 20307 7160 20352 7188
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 20898 7188 20904 7200
rect 20859 7160 20904 7188
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 20622 6944 20628 6996
rect 20680 6984 20686 6996
rect 23431 6987 23489 6993
rect 23431 6984 23443 6987
rect 20680 6956 23443 6984
rect 20680 6944 20686 6956
rect 23431 6953 23443 6956
rect 23477 6953 23489 6987
rect 23431 6947 23489 6953
rect 35621 6987 35679 6993
rect 35621 6953 35633 6987
rect 35667 6984 35679 6987
rect 39574 6984 39580 6996
rect 35667 6956 39580 6984
rect 35667 6953 35679 6956
rect 35621 6947 35679 6953
rect 39574 6944 39580 6956
rect 39632 6944 39638 6996
rect 2406 6876 2412 6928
rect 2464 6916 2470 6928
rect 2546 6919 2604 6925
rect 2546 6916 2558 6919
rect 2464 6888 2558 6916
rect 2464 6876 2470 6888
rect 2546 6885 2558 6888
rect 2592 6885 2604 6919
rect 4246 6916 4252 6928
rect 4207 6888 4252 6916
rect 2546 6879 2604 6885
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 4798 6876 4804 6928
rect 4856 6916 4862 6928
rect 5718 6916 5724 6928
rect 4856 6888 5724 6916
rect 4856 6876 4862 6888
rect 5718 6876 5724 6888
rect 5776 6876 5782 6928
rect 5810 6876 5816 6928
rect 5868 6916 5874 6928
rect 10318 6916 10324 6928
rect 5868 6888 5913 6916
rect 10279 6888 10324 6916
rect 5868 6876 5874 6888
rect 10318 6876 10324 6888
rect 10376 6876 10382 6928
rect 10410 6876 10416 6928
rect 10468 6916 10474 6928
rect 13817 6919 13875 6925
rect 10468 6888 10513 6916
rect 10468 6876 10474 6888
rect 13817 6885 13829 6919
rect 13863 6916 13875 6919
rect 13998 6916 14004 6928
rect 13863 6888 14004 6916
rect 13863 6885 13875 6888
rect 13817 6879 13875 6885
rect 13998 6876 14004 6888
rect 14056 6916 14062 6928
rect 15470 6916 15476 6928
rect 14056 6888 15476 6916
rect 14056 6876 14062 6888
rect 15470 6876 15476 6888
rect 15528 6876 15534 6928
rect 19058 6876 19064 6928
rect 19116 6916 19122 6928
rect 19429 6919 19487 6925
rect 19429 6916 19441 6919
rect 19116 6888 19441 6916
rect 19116 6876 19122 6888
rect 19429 6885 19441 6888
rect 19475 6885 19487 6919
rect 19429 6879 19487 6885
rect 20714 6876 20720 6928
rect 20772 6916 20778 6928
rect 21085 6919 21143 6925
rect 21085 6916 21097 6919
rect 20772 6888 21097 6916
rect 20772 6876 20778 6888
rect 21085 6885 21097 6888
rect 21131 6885 21143 6919
rect 21085 6879 21143 6885
rect 12526 6848 12532 6860
rect 12487 6820 12532 6848
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 16758 6808 16764 6860
rect 16816 6848 16822 6860
rect 16853 6851 16911 6857
rect 16853 6848 16865 6851
rect 16816 6820 16865 6848
rect 16816 6808 16822 6820
rect 16853 6817 16865 6820
rect 16899 6817 16911 6851
rect 16853 6811 16911 6817
rect 18233 6851 18291 6857
rect 18233 6817 18245 6851
rect 18279 6848 18291 6851
rect 18322 6848 18328 6860
rect 18279 6820 18328 6848
rect 18279 6817 18291 6820
rect 18233 6811 18291 6817
rect 18322 6808 18328 6820
rect 18380 6808 18386 6860
rect 23360 6851 23418 6857
rect 23360 6817 23372 6851
rect 23406 6848 23418 6851
rect 23474 6848 23480 6860
rect 23406 6820 23480 6848
rect 23406 6817 23418 6820
rect 23360 6811 23418 6817
rect 23474 6808 23480 6820
rect 23532 6808 23538 6860
rect 24486 6848 24492 6860
rect 24447 6820 24492 6848
rect 24486 6808 24492 6820
rect 24544 6808 24550 6860
rect 35434 6848 35440 6860
rect 35395 6820 35440 6848
rect 35434 6808 35440 6820
rect 35492 6808 35498 6860
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 1670 6644 1676 6656
rect 1631 6616 1676 6644
rect 1670 6604 1676 6616
rect 1728 6604 1734 6656
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 2240 6644 2268 6743
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 3844 6752 4169 6780
rect 3844 6740 3850 6752
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4614 6780 4620 6792
rect 4575 6752 4620 6780
rect 4157 6743 4215 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6780 6055 6783
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 6043 6752 6837 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6825 6749 6837 6752
rect 6871 6780 6883 6783
rect 6914 6780 6920 6792
rect 6871 6752 6920 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 2590 6672 2596 6724
rect 2648 6712 2654 6724
rect 3421 6715 3479 6721
rect 3421 6712 3433 6715
rect 2648 6684 3433 6712
rect 2648 6672 2654 6684
rect 3421 6681 3433 6684
rect 3467 6681 3479 6715
rect 3421 6675 3479 6681
rect 4982 6672 4988 6724
rect 5040 6712 5046 6724
rect 6012 6712 6040 6743
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 8570 6780 8576 6792
rect 8531 6752 8576 6780
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 12759 6783 12817 6789
rect 12759 6749 12771 6783
rect 12805 6780 12817 6783
rect 13173 6783 13231 6789
rect 13173 6780 13185 6783
rect 12805 6752 13185 6780
rect 12805 6749 12817 6752
rect 12759 6743 12817 6749
rect 13173 6749 13185 6752
rect 13219 6780 13231 6783
rect 13725 6783 13783 6789
rect 13725 6780 13737 6783
rect 13219 6752 13737 6780
rect 13219 6749 13231 6752
rect 13173 6743 13231 6749
rect 13725 6749 13737 6752
rect 13771 6749 13783 6783
rect 14366 6780 14372 6792
rect 14327 6752 14372 6780
rect 13725 6743 13783 6749
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 15378 6780 15384 6792
rect 15339 6752 15384 6780
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 15562 6740 15568 6792
rect 15620 6780 15626 6792
rect 15657 6783 15715 6789
rect 15657 6780 15669 6783
rect 15620 6752 15669 6780
rect 15620 6740 15626 6752
rect 15657 6749 15669 6752
rect 15703 6749 15715 6783
rect 15657 6743 15715 6749
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 19337 6783 19395 6789
rect 19337 6780 19349 6783
rect 18840 6752 19349 6780
rect 18840 6740 18846 6752
rect 19337 6749 19349 6752
rect 19383 6780 19395 6783
rect 20625 6783 20683 6789
rect 20625 6780 20637 6783
rect 19383 6752 20637 6780
rect 19383 6749 19395 6752
rect 19337 6743 19395 6749
rect 20625 6749 20637 6752
rect 20671 6749 20683 6783
rect 20625 6743 20683 6749
rect 20806 6740 20812 6792
rect 20864 6780 20870 6792
rect 20993 6783 21051 6789
rect 20993 6780 21005 6783
rect 20864 6752 21005 6780
rect 20864 6740 20870 6752
rect 20993 6749 21005 6752
rect 21039 6749 21051 6783
rect 20993 6743 21051 6749
rect 5040 6684 6040 6712
rect 5040 6672 5046 6684
rect 10594 6672 10600 6724
rect 10652 6712 10658 6724
rect 10873 6715 10931 6721
rect 10873 6712 10885 6715
rect 10652 6684 10885 6712
rect 10652 6672 10658 6684
rect 10873 6681 10885 6684
rect 10919 6712 10931 6715
rect 11333 6715 11391 6721
rect 11333 6712 11345 6715
rect 10919 6684 11345 6712
rect 10919 6681 10931 6684
rect 10873 6675 10931 6681
rect 11333 6681 11345 6684
rect 11379 6712 11391 6715
rect 14384 6712 14412 6740
rect 11379 6684 14412 6712
rect 18371 6715 18429 6721
rect 11379 6681 11391 6684
rect 11333 6675 11391 6681
rect 18371 6681 18383 6715
rect 18417 6712 18429 6715
rect 18966 6712 18972 6724
rect 18417 6684 18972 6712
rect 18417 6681 18429 6684
rect 18371 6675 18429 6681
rect 18966 6672 18972 6684
rect 19024 6672 19030 6724
rect 19889 6715 19947 6721
rect 19889 6681 19901 6715
rect 19935 6712 19947 6715
rect 19978 6712 19984 6724
rect 19935 6684 19984 6712
rect 19935 6681 19947 6684
rect 19889 6675 19947 6681
rect 19978 6672 19984 6684
rect 20036 6712 20042 6724
rect 20898 6712 20904 6724
rect 20036 6684 20904 6712
rect 20036 6672 20042 6684
rect 20898 6672 20904 6684
rect 20956 6672 20962 6724
rect 21542 6712 21548 6724
rect 21503 6684 21548 6712
rect 21542 6672 21548 6684
rect 21600 6712 21606 6724
rect 21913 6715 21971 6721
rect 21913 6712 21925 6715
rect 21600 6684 21925 6712
rect 21600 6672 21606 6684
rect 21913 6681 21925 6684
rect 21959 6681 21971 6715
rect 21913 6675 21971 6681
rect 2498 6644 2504 6656
rect 2179 6616 2504 6644
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 3145 6647 3203 6653
rect 3145 6613 3157 6647
rect 3191 6644 3203 6647
rect 4062 6644 4068 6656
rect 3191 6616 4068 6644
rect 3191 6613 3203 6616
rect 3145 6607 3203 6613
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 5077 6647 5135 6653
rect 5077 6644 5089 6647
rect 4396 6616 5089 6644
rect 4396 6604 4402 6616
rect 5077 6613 5089 6616
rect 5123 6613 5135 6647
rect 5077 6607 5135 6613
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 13814 6644 13820 6656
rect 13587 6616 13820 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 14737 6647 14795 6653
rect 14737 6613 14749 6647
rect 14783 6644 14795 6647
rect 14826 6644 14832 6656
rect 14783 6616 14832 6644
rect 14783 6613 14795 6616
rect 14737 6607 14795 6613
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 15102 6644 15108 6656
rect 15063 6616 15108 6644
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 17000 6616 17049 6644
rect 17000 6604 17006 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 18690 6644 18696 6656
rect 18651 6616 18696 6644
rect 17037 6607 17095 6613
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 19058 6644 19064 6656
rect 19019 6616 19064 6644
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 20257 6647 20315 6653
rect 20257 6644 20269 6647
rect 19392 6616 20269 6644
rect 19392 6604 19398 6616
rect 20257 6613 20269 6616
rect 20303 6644 20315 6647
rect 20346 6644 20352 6656
rect 20303 6616 20352 6644
rect 20303 6613 20315 6616
rect 20257 6607 20315 6613
rect 20346 6604 20352 6616
rect 20404 6604 20410 6656
rect 24578 6644 24584 6656
rect 24539 6616 24584 6644
rect 24578 6604 24584 6616
rect 24636 6604 24642 6656
rect 25130 6604 25136 6656
rect 25188 6644 25194 6656
rect 25317 6647 25375 6653
rect 25317 6644 25329 6647
rect 25188 6616 25329 6644
rect 25188 6604 25194 6616
rect 25317 6613 25329 6616
rect 25363 6613 25375 6647
rect 25317 6607 25375 6613
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 14 6400 20 6452
rect 72 6440 78 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 72 6412 1593 6440
rect 72 6400 78 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 1581 6403 1639 6409
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 3234 6400 3240 6452
rect 3292 6440 3298 6452
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 3292 6412 3433 6440
rect 3292 6400 3298 6412
rect 3421 6409 3433 6412
rect 3467 6409 3479 6443
rect 4062 6440 4068 6452
rect 4023 6412 4068 6440
rect 3421 6403 3479 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4430 6440 4436 6452
rect 4172 6412 4436 6440
rect 2406 6372 2412 6384
rect 2319 6344 2412 6372
rect 2406 6332 2412 6344
rect 2464 6372 2470 6384
rect 3789 6375 3847 6381
rect 3789 6372 3801 6375
rect 2464 6344 3801 6372
rect 2464 6332 2470 6344
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2038 6236 2044 6248
rect 1443 6208 2044 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 2590 6236 2596 6248
rect 2547 6208 2596 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 2878 6177 2906 6344
rect 3789 6341 3801 6344
rect 3835 6372 3847 6375
rect 4172 6372 4200 6412
rect 4430 6400 4436 6412
rect 4488 6400 4494 6452
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5776 6412 6009 6440
rect 5776 6400 5782 6412
rect 5997 6409 6009 6412
rect 6043 6409 6055 6443
rect 5997 6403 6055 6409
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 8628 6412 8769 6440
rect 8628 6400 8634 6412
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 8757 6403 8815 6409
rect 10321 6443 10379 6449
rect 10321 6409 10333 6443
rect 10367 6440 10379 6443
rect 10410 6440 10416 6452
rect 10367 6412 10416 6440
rect 10367 6409 10379 6412
rect 10321 6403 10379 6409
rect 3835 6344 4200 6372
rect 3835 6341 3847 6344
rect 3789 6335 3847 6341
rect 4246 6332 4252 6384
rect 4304 6372 4310 6384
rect 5261 6375 5319 6381
rect 5261 6372 5273 6375
rect 4304 6344 5273 6372
rect 4304 6332 4310 6344
rect 5261 6341 5273 6344
rect 5307 6372 5319 6375
rect 5629 6375 5687 6381
rect 5629 6372 5641 6375
rect 5307 6344 5641 6372
rect 5307 6341 5319 6344
rect 5261 6335 5319 6341
rect 5629 6341 5641 6344
rect 5675 6372 5687 6375
rect 5810 6372 5816 6384
rect 5675 6344 5816 6372
rect 5675 6341 5687 6344
rect 5629 6335 5687 6341
rect 5810 6332 5816 6344
rect 5868 6332 5874 6384
rect 4338 6304 4344 6316
rect 4126 6276 4344 6304
rect 2863 6171 2921 6177
rect 2863 6137 2875 6171
rect 2909 6137 2921 6171
rect 2863 6131 2921 6137
rect 3418 6128 3424 6180
rect 3476 6168 3482 6180
rect 4126 6168 4154 6276
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 4614 6304 4620 6316
rect 4575 6276 4620 6304
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 6914 6304 6920 6316
rect 6875 6276 6920 6304
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 7190 6304 7196 6316
rect 7151 6276 7196 6304
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 8772 6304 8800 6403
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 15194 6440 15200 6452
rect 11164 6412 15200 6440
rect 11164 6381 11192 6412
rect 15194 6400 15200 6412
rect 15252 6400 15258 6452
rect 15289 6443 15347 6449
rect 15289 6409 15301 6443
rect 15335 6440 15347 6443
rect 15470 6440 15476 6452
rect 15335 6412 15476 6440
rect 15335 6409 15347 6412
rect 15289 6403 15347 6409
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 18322 6440 18328 6452
rect 18283 6412 18328 6440
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 18693 6443 18751 6449
rect 18693 6409 18705 6443
rect 18739 6440 18751 6443
rect 18782 6440 18788 6452
rect 18739 6412 18788 6440
rect 18739 6409 18751 6412
rect 18693 6403 18751 6409
rect 18782 6400 18788 6412
rect 18840 6400 18846 6452
rect 21266 6400 21272 6452
rect 21324 6440 21330 6452
rect 22373 6443 22431 6449
rect 22373 6440 22385 6443
rect 21324 6412 22385 6440
rect 21324 6400 21330 6412
rect 22373 6409 22385 6412
rect 22419 6409 22431 6443
rect 22373 6403 22431 6409
rect 23474 6400 23480 6452
rect 23532 6440 23538 6452
rect 24486 6440 24492 6452
rect 23532 6412 23577 6440
rect 24447 6412 24492 6440
rect 23532 6400 23538 6412
rect 24486 6400 24492 6412
rect 24544 6440 24550 6452
rect 24854 6440 24860 6452
rect 24544 6412 24860 6440
rect 24544 6400 24550 6412
rect 24854 6400 24860 6412
rect 24912 6400 24918 6452
rect 9585 6375 9643 6381
rect 9585 6341 9597 6375
rect 9631 6372 9643 6375
rect 11149 6375 11207 6381
rect 11149 6372 11161 6375
rect 9631 6344 11161 6372
rect 9631 6341 9643 6344
rect 9585 6335 9643 6341
rect 11149 6341 11161 6344
rect 11195 6341 11207 6375
rect 11149 6335 11207 6341
rect 12526 6332 12532 6384
rect 12584 6372 12590 6384
rect 12897 6375 12955 6381
rect 12897 6372 12909 6375
rect 12584 6344 12909 6372
rect 12584 6332 12590 6344
rect 12897 6341 12909 6344
rect 12943 6372 12955 6375
rect 12943 6344 13814 6372
rect 12943 6341 12955 6344
rect 12897 6335 12955 6341
rect 9033 6307 9091 6313
rect 9033 6304 9045 6307
rect 8772 6276 9045 6304
rect 9033 6273 9045 6276
rect 9079 6273 9091 6307
rect 10594 6304 10600 6316
rect 10555 6276 10600 6304
rect 9033 6267 9091 6273
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 13786 6304 13814 6344
rect 14366 6332 14372 6384
rect 14424 6372 14430 6384
rect 16025 6375 16083 6381
rect 16025 6372 16037 6375
rect 14424 6344 16037 6372
rect 14424 6332 14430 6344
rect 16025 6341 16037 6344
rect 16071 6341 16083 6375
rect 16025 6335 16083 6341
rect 20073 6375 20131 6381
rect 20073 6341 20085 6375
rect 20119 6372 20131 6375
rect 21542 6372 21548 6384
rect 20119 6344 21548 6372
rect 20119 6341 20131 6344
rect 20073 6335 20131 6341
rect 21542 6332 21548 6344
rect 21600 6372 21606 6384
rect 21637 6375 21695 6381
rect 21637 6372 21649 6375
rect 21600 6344 21649 6372
rect 21600 6332 21606 6344
rect 21637 6341 21649 6344
rect 21683 6341 21695 6375
rect 21637 6335 21695 6341
rect 14918 6304 14924 6316
rect 13786 6276 14924 6304
rect 14918 6264 14924 6276
rect 14976 6264 14982 6316
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 15473 6307 15531 6313
rect 15473 6304 15485 6307
rect 15160 6276 15485 6304
rect 15160 6264 15166 6276
rect 15473 6273 15485 6276
rect 15519 6304 15531 6307
rect 17083 6307 17141 6313
rect 17083 6304 17095 6307
rect 15519 6276 17095 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 17083 6273 17095 6276
rect 17129 6273 17141 6307
rect 17083 6267 17141 6273
rect 18966 6264 18972 6316
rect 19024 6304 19030 6316
rect 19521 6307 19579 6313
rect 19521 6304 19533 6307
rect 19024 6276 19533 6304
rect 19024 6264 19030 6276
rect 19521 6273 19533 6276
rect 19567 6273 19579 6307
rect 19521 6267 19579 6273
rect 20806 6264 20812 6316
rect 20864 6304 20870 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 20864 6276 22017 6304
rect 20864 6264 20870 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22370 6264 22376 6316
rect 22428 6304 22434 6316
rect 23017 6307 23075 6313
rect 23017 6304 23029 6307
rect 22428 6276 23029 6304
rect 22428 6264 22434 6276
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6236 12311 6239
rect 12434 6236 12440 6248
rect 12299 6208 12440 6236
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 13633 6239 13691 6245
rect 13633 6205 13645 6239
rect 13679 6236 13691 6239
rect 13814 6236 13820 6248
rect 13679 6208 13820 6236
rect 13679 6205 13691 6208
rect 13633 6199 13691 6205
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 16996 6239 17054 6245
rect 16996 6205 17008 6239
rect 17042 6236 17054 6239
rect 17494 6236 17500 6248
rect 17042 6208 17500 6236
rect 17042 6205 17054 6208
rect 16996 6199 17054 6205
rect 17494 6196 17500 6208
rect 17552 6196 17558 6248
rect 18484 6239 18542 6245
rect 18484 6205 18496 6239
rect 18530 6236 18542 6239
rect 18598 6236 18604 6248
rect 18530 6208 18604 6236
rect 18530 6205 18542 6208
rect 18484 6199 18542 6205
rect 18598 6196 18604 6208
rect 18656 6236 18662 6248
rect 22639 6245 22667 6276
rect 23017 6273 23029 6276
rect 23063 6273 23075 6307
rect 25406 6304 25412 6316
rect 25367 6276 25412 6304
rect 23017 6267 23075 6273
rect 25406 6264 25412 6276
rect 25464 6264 25470 6316
rect 35434 6304 35440 6316
rect 35395 6276 35440 6304
rect 35434 6264 35440 6276
rect 35492 6264 35498 6316
rect 18877 6239 18935 6245
rect 18877 6236 18889 6239
rect 18656 6208 18889 6236
rect 18656 6196 18662 6208
rect 18877 6205 18889 6208
rect 18923 6205 18935 6239
rect 18877 6199 18935 6205
rect 22624 6239 22682 6245
rect 22624 6205 22636 6239
rect 22670 6205 22682 6239
rect 22624 6199 22682 6205
rect 3476 6140 4154 6168
rect 4433 6171 4491 6177
rect 3476 6128 3482 6140
rect 4433 6137 4445 6171
rect 4479 6137 4491 6171
rect 4433 6131 4491 6137
rect 7009 6171 7067 6177
rect 7009 6137 7021 6171
rect 7055 6137 7067 6171
rect 9122 6168 9128 6180
rect 9083 6140 9128 6168
rect 7009 6131 7067 6137
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 4448 6100 4476 6131
rect 6546 6100 6552 6112
rect 4120 6072 4476 6100
rect 6507 6072 6552 6100
rect 4120 6060 4126 6072
rect 6546 6060 6552 6072
rect 6604 6100 6610 6112
rect 7024 6100 7052 6131
rect 9122 6128 9128 6140
rect 9180 6128 9186 6180
rect 9490 6128 9496 6180
rect 9548 6168 9554 6180
rect 10689 6171 10747 6177
rect 10689 6168 10701 6171
rect 9548 6140 10701 6168
rect 9548 6128 9554 6140
rect 10689 6137 10701 6140
rect 10735 6168 10747 6171
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 10735 6140 11529 6168
rect 10735 6137 10747 6140
rect 10689 6131 10747 6137
rect 11517 6137 11529 6140
rect 11563 6137 11575 6171
rect 13538 6168 13544 6180
rect 13451 6140 13544 6168
rect 11517 6131 11575 6137
rect 13538 6128 13544 6140
rect 13596 6168 13602 6180
rect 13596 6140 13814 6168
rect 13596 6128 13602 6140
rect 12618 6100 12624 6112
rect 6604 6072 7052 6100
rect 12579 6072 12624 6100
rect 6604 6060 6610 6072
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 13786 6100 13814 6140
rect 14826 6128 14832 6180
rect 14884 6168 14890 6180
rect 14921 6171 14979 6177
rect 14921 6168 14933 6171
rect 14884 6140 14933 6168
rect 14884 6128 14890 6140
rect 14921 6137 14933 6140
rect 14967 6168 14979 6171
rect 15565 6171 15623 6177
rect 15565 6168 15577 6171
rect 14967 6140 15577 6168
rect 14967 6137 14979 6140
rect 14921 6131 14979 6137
rect 15565 6137 15577 6140
rect 15611 6168 15623 6171
rect 15654 6168 15660 6180
rect 15611 6140 15660 6168
rect 15611 6137 15623 6140
rect 15565 6131 15623 6137
rect 15654 6128 15660 6140
rect 15712 6128 15718 6180
rect 19613 6171 19671 6177
rect 19613 6137 19625 6171
rect 19659 6137 19671 6171
rect 20530 6168 20536 6180
rect 20443 6140 20536 6168
rect 19613 6131 19671 6137
rect 14001 6103 14059 6109
rect 14001 6100 14013 6103
rect 13786 6072 14013 6100
rect 14001 6069 14013 6072
rect 14047 6069 14059 6103
rect 14001 6063 14059 6069
rect 14553 6103 14611 6109
rect 14553 6069 14565 6103
rect 14599 6100 14611 6103
rect 14734 6100 14740 6112
rect 14599 6072 14740 6100
rect 14599 6069 14611 6072
rect 14553 6063 14611 6069
rect 14734 6060 14740 6072
rect 14792 6060 14798 6112
rect 15378 6060 15384 6112
rect 15436 6100 15442 6112
rect 16393 6103 16451 6109
rect 16393 6100 16405 6103
rect 15436 6072 16405 6100
rect 15436 6060 15442 6072
rect 16393 6069 16405 6072
rect 16439 6069 16451 6103
rect 16758 6100 16764 6112
rect 16719 6072 16764 6100
rect 16393 6063 16451 6069
rect 16758 6060 16764 6072
rect 16816 6060 16822 6112
rect 17494 6100 17500 6112
rect 17455 6072 17500 6100
rect 17494 6060 17500 6072
rect 17552 6060 17558 6112
rect 17770 6100 17776 6112
rect 17731 6072 17776 6100
rect 17770 6060 17776 6072
rect 17828 6060 17834 6112
rect 18966 6060 18972 6112
rect 19024 6100 19030 6112
rect 19245 6103 19303 6109
rect 19245 6100 19257 6103
rect 19024 6072 19257 6100
rect 19024 6060 19030 6072
rect 19245 6069 19257 6072
rect 19291 6100 19303 6103
rect 19628 6100 19656 6131
rect 20530 6128 20536 6140
rect 20588 6168 20594 6180
rect 21082 6168 21088 6180
rect 20588 6140 20944 6168
rect 21043 6140 21088 6168
rect 20588 6128 20594 6140
rect 19291 6072 19656 6100
rect 19291 6069 19303 6072
rect 19245 6063 19303 6069
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 20809 6103 20867 6109
rect 20809 6100 20821 6103
rect 20772 6072 20821 6100
rect 20772 6060 20778 6072
rect 20809 6069 20821 6072
rect 20855 6069 20867 6103
rect 20916 6100 20944 6140
rect 21082 6128 21088 6140
rect 21140 6128 21146 6180
rect 21177 6171 21235 6177
rect 21177 6137 21189 6171
rect 21223 6137 21235 6171
rect 21177 6131 21235 6137
rect 21192 6100 21220 6131
rect 24394 6128 24400 6180
rect 24452 6168 24458 6180
rect 25130 6168 25136 6180
rect 24452 6140 25136 6168
rect 24452 6128 24458 6140
rect 25130 6128 25136 6140
rect 25188 6128 25194 6180
rect 25225 6171 25283 6177
rect 25225 6137 25237 6171
rect 25271 6137 25283 6171
rect 25225 6131 25283 6137
rect 20916 6072 21220 6100
rect 20809 6063 20867 6069
rect 22554 6060 22560 6112
rect 22612 6100 22618 6112
rect 22695 6103 22753 6109
rect 22695 6100 22707 6103
rect 22612 6072 22707 6100
rect 22612 6060 22618 6072
rect 22695 6069 22707 6072
rect 22741 6069 22753 6103
rect 24026 6100 24032 6112
rect 23987 6072 24032 6100
rect 22695 6063 22753 6069
rect 24026 6060 24032 6072
rect 24084 6060 24090 6112
rect 24949 6103 25007 6109
rect 24949 6069 24961 6103
rect 24995 6100 25007 6103
rect 25240 6100 25268 6131
rect 25498 6100 25504 6112
rect 24995 6072 25504 6100
rect 24995 6069 25007 6072
rect 24949 6063 25007 6069
rect 25498 6060 25504 6072
rect 25556 6060 25562 6112
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 3145 5899 3203 5905
rect 3145 5865 3157 5899
rect 3191 5896 3203 5899
rect 4246 5896 4252 5908
rect 3191 5868 4252 5896
rect 3191 5865 3203 5868
rect 3145 5859 3203 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 4430 5896 4436 5908
rect 4391 5868 4436 5896
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 6270 5896 6276 5908
rect 6231 5868 6276 5896
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 6825 5899 6883 5905
rect 6825 5865 6837 5899
rect 6871 5896 6883 5899
rect 7466 5896 7472 5908
rect 6871 5868 7472 5896
rect 6871 5865 6883 5868
rect 6825 5859 6883 5865
rect 7466 5856 7472 5868
rect 7524 5896 7530 5908
rect 9033 5899 9091 5905
rect 7524 5868 7880 5896
rect 7524 5856 7530 5868
rect 2406 5788 2412 5840
rect 2464 5828 2470 5840
rect 7852 5837 7880 5868
rect 9033 5865 9045 5899
rect 9079 5896 9091 5899
rect 9122 5896 9128 5908
rect 9079 5868 9128 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 10318 5896 10324 5908
rect 10279 5868 10324 5896
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 13998 5896 14004 5908
rect 13959 5868 14004 5896
rect 13998 5856 14004 5868
rect 14056 5896 14062 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 14056 5868 14289 5896
rect 14056 5856 14062 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14277 5859 14335 5865
rect 18417 5899 18475 5905
rect 18417 5865 18429 5899
rect 18463 5896 18475 5899
rect 19153 5899 19211 5905
rect 19153 5896 19165 5899
rect 18463 5868 19165 5896
rect 18463 5865 18475 5868
rect 18417 5859 18475 5865
rect 19153 5865 19165 5868
rect 19199 5896 19211 5899
rect 21266 5896 21272 5908
rect 19199 5868 19472 5896
rect 21227 5868 21272 5896
rect 19199 5865 19211 5868
rect 19153 5859 19211 5865
rect 2546 5831 2604 5837
rect 2546 5828 2558 5831
rect 2464 5800 2558 5828
rect 2464 5788 2470 5800
rect 2546 5797 2558 5800
rect 2592 5797 2604 5831
rect 2546 5791 2604 5797
rect 7837 5831 7895 5837
rect 7837 5797 7849 5831
rect 7883 5797 7895 5831
rect 7837 5791 7895 5797
rect 10410 5788 10416 5840
rect 10468 5828 10474 5840
rect 10781 5831 10839 5837
rect 10781 5828 10793 5831
rect 10468 5800 10793 5828
rect 10468 5788 10474 5800
rect 10781 5797 10793 5800
rect 10827 5797 10839 5831
rect 10781 5791 10839 5797
rect 13443 5831 13501 5837
rect 13443 5797 13455 5831
rect 13489 5828 13501 5831
rect 13538 5828 13544 5840
rect 13489 5800 13544 5828
rect 13489 5797 13501 5800
rect 13443 5791 13501 5797
rect 13538 5788 13544 5800
rect 13596 5788 13602 5840
rect 14734 5788 14740 5840
rect 14792 5828 14798 5840
rect 15473 5831 15531 5837
rect 15473 5828 15485 5831
rect 14792 5800 15485 5828
rect 14792 5788 14798 5800
rect 15473 5797 15485 5800
rect 15519 5828 15531 5831
rect 16301 5831 16359 5837
rect 16301 5828 16313 5831
rect 15519 5800 16313 5828
rect 15519 5797 15531 5800
rect 15473 5791 15531 5797
rect 16301 5797 16313 5800
rect 16347 5797 16359 5831
rect 16301 5791 16359 5797
rect 17859 5831 17917 5837
rect 17859 5797 17871 5831
rect 17905 5828 17917 5831
rect 18138 5828 18144 5840
rect 17905 5800 18144 5828
rect 17905 5797 17917 5800
rect 17859 5791 17917 5797
rect 18138 5788 18144 5800
rect 18196 5788 18202 5840
rect 19334 5828 19340 5840
rect 19295 5800 19340 5828
rect 19334 5788 19340 5800
rect 19392 5788 19398 5840
rect 19444 5837 19472 5868
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 25406 5896 25412 5908
rect 25367 5868 25412 5896
rect 25406 5856 25412 5868
rect 25464 5856 25470 5908
rect 19429 5831 19487 5837
rect 19429 5797 19441 5831
rect 19475 5828 19487 5831
rect 20530 5828 20536 5840
rect 19475 5800 20536 5828
rect 19475 5797 19487 5800
rect 19429 5791 19487 5797
rect 20530 5788 20536 5800
rect 20588 5788 20594 5840
rect 22554 5828 22560 5840
rect 22515 5800 22560 5828
rect 22554 5788 22560 5800
rect 22612 5828 22618 5840
rect 22741 5831 22799 5837
rect 22741 5828 22753 5831
rect 22612 5800 22753 5828
rect 22612 5788 22618 5800
rect 22741 5797 22753 5800
rect 22787 5797 22799 5831
rect 22741 5791 22799 5797
rect 22833 5831 22891 5837
rect 22833 5797 22845 5831
rect 22879 5828 22891 5831
rect 22922 5828 22928 5840
rect 22879 5800 22928 5828
rect 22879 5797 22891 5800
rect 22833 5791 22891 5797
rect 22922 5788 22928 5800
rect 22980 5788 22986 5840
rect 24578 5828 24584 5840
rect 24539 5800 24584 5828
rect 24578 5788 24584 5800
rect 24636 5788 24642 5840
rect 12529 5763 12587 5769
rect 12529 5729 12541 5763
rect 12575 5760 12587 5763
rect 12618 5760 12624 5772
rect 12575 5732 12624 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 12618 5720 12624 5732
rect 12676 5760 12682 5772
rect 13262 5760 13268 5772
rect 12676 5732 13268 5760
rect 12676 5720 12682 5732
rect 13262 5720 13268 5732
rect 13320 5720 13326 5772
rect 19978 5720 19984 5772
rect 20036 5760 20042 5772
rect 20036 5732 21312 5760
rect 20036 5720 20042 5732
rect 2222 5692 2228 5704
rect 2183 5664 2228 5692
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5692 4123 5695
rect 4522 5692 4528 5704
rect 4111 5664 4528 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5692 5963 5695
rect 6638 5692 6644 5704
rect 5951 5664 6644 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 7745 5695 7803 5701
rect 7745 5692 7757 5695
rect 7432 5664 7757 5692
rect 7432 5652 7438 5664
rect 7745 5661 7757 5664
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 7190 5584 7196 5636
rect 7248 5624 7254 5636
rect 8036 5624 8064 5655
rect 10502 5652 10508 5704
rect 10560 5692 10566 5704
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 10560 5664 10701 5692
rect 10560 5652 10566 5664
rect 10689 5661 10701 5664
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 13722 5692 13728 5704
rect 13127 5664 13728 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 13722 5652 13728 5664
rect 13780 5692 13786 5704
rect 14645 5695 14703 5701
rect 14645 5692 14657 5695
rect 13780 5664 14657 5692
rect 13780 5652 13786 5664
rect 14645 5661 14657 5664
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5692 15439 5695
rect 15562 5692 15568 5704
rect 15427 5664 15568 5692
rect 15427 5661 15439 5664
rect 15381 5655 15439 5661
rect 7248 5596 8064 5624
rect 11241 5627 11299 5633
rect 7248 5584 7254 5596
rect 11241 5593 11253 5627
rect 11287 5624 11299 5627
rect 15396 5624 15424 5655
rect 15562 5652 15568 5664
rect 15620 5652 15626 5704
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5661 15715 5695
rect 15657 5655 15715 5661
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 11287 5596 15424 5624
rect 11287 5593 11299 5596
rect 11241 5587 11299 5593
rect 1762 5556 1768 5568
rect 1723 5528 1768 5556
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 2130 5556 2136 5568
rect 2091 5528 2136 5556
rect 2130 5516 2136 5528
rect 2188 5516 2194 5568
rect 3050 5516 3056 5568
rect 3108 5556 3114 5568
rect 3421 5559 3479 5565
rect 3421 5556 3433 5559
rect 3108 5528 3433 5556
rect 3108 5516 3114 5528
rect 3421 5525 3433 5528
rect 3467 5525 3479 5559
rect 3786 5556 3792 5568
rect 3747 5528 3792 5556
rect 3421 5519 3479 5525
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 4982 5556 4988 5568
rect 4943 5528 4988 5556
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 7561 5559 7619 5565
rect 7561 5525 7573 5559
rect 7607 5556 7619 5559
rect 8110 5556 8116 5568
rect 7607 5528 8116 5556
rect 7607 5525 7619 5528
rect 7561 5519 7619 5525
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 12342 5516 12348 5568
rect 12400 5556 12406 5568
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 12400 5528 12817 5556
rect 12400 5516 12406 5528
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 15010 5556 15016 5568
rect 14971 5528 15016 5556
rect 12805 5519 12863 5525
rect 15010 5516 15016 5528
rect 15068 5516 15074 5568
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 15672 5556 15700 5655
rect 15252 5528 15700 5556
rect 16761 5559 16819 5565
rect 15252 5516 15258 5528
rect 16761 5525 16773 5559
rect 16807 5556 16819 5559
rect 16850 5556 16856 5568
rect 16807 5528 16856 5556
rect 16807 5525 16819 5528
rect 16761 5519 16819 5525
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 17405 5559 17463 5565
rect 17405 5525 17417 5559
rect 17451 5556 17463 5559
rect 17512 5556 17540 5655
rect 20622 5652 20628 5704
rect 20680 5692 20686 5704
rect 20901 5695 20959 5701
rect 20901 5692 20913 5695
rect 20680 5664 20913 5692
rect 20680 5652 20686 5664
rect 20901 5661 20913 5664
rect 20947 5661 20959 5695
rect 21284 5692 21312 5732
rect 25498 5720 25504 5772
rect 25556 5760 25562 5772
rect 26605 5763 26663 5769
rect 26605 5760 26617 5763
rect 25556 5732 26617 5760
rect 25556 5720 25562 5732
rect 26605 5729 26617 5732
rect 26651 5760 26663 5763
rect 27246 5760 27252 5772
rect 26651 5732 27252 5760
rect 26651 5729 26663 5732
rect 26605 5723 26663 5729
rect 27246 5720 27252 5732
rect 27304 5720 27310 5772
rect 21450 5692 21456 5704
rect 21284 5664 21456 5692
rect 20901 5655 20959 5661
rect 21450 5652 21456 5664
rect 21508 5692 21514 5704
rect 23017 5695 23075 5701
rect 23017 5692 23029 5695
rect 21508 5664 23029 5692
rect 21508 5652 21514 5664
rect 23017 5661 23029 5664
rect 23063 5661 23075 5695
rect 23017 5655 23075 5661
rect 24026 5652 24032 5704
rect 24084 5692 24090 5704
rect 24486 5692 24492 5704
rect 24084 5664 24492 5692
rect 24084 5652 24090 5664
rect 24486 5652 24492 5664
rect 24544 5652 24550 5704
rect 24765 5695 24823 5701
rect 24765 5661 24777 5695
rect 24811 5661 24823 5695
rect 26510 5692 26516 5704
rect 26471 5664 26516 5692
rect 24765 5655 24823 5661
rect 23474 5584 23480 5636
rect 23532 5624 23538 5636
rect 24780 5624 24808 5655
rect 26510 5652 26516 5664
rect 26568 5652 26574 5704
rect 25314 5624 25320 5636
rect 23532 5596 25320 5624
rect 23532 5584 23538 5596
rect 25314 5584 25320 5596
rect 25372 5584 25378 5636
rect 17862 5556 17868 5568
rect 17451 5528 17868 5556
rect 17451 5525 17463 5528
rect 17405 5519 17463 5525
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 18785 5559 18843 5565
rect 18785 5525 18797 5559
rect 18831 5556 18843 5559
rect 18874 5556 18880 5568
rect 18831 5528 18880 5556
rect 18831 5525 18843 5528
rect 18785 5519 18843 5525
rect 18874 5516 18880 5528
rect 18932 5516 18938 5568
rect 20346 5556 20352 5568
rect 20307 5528 20352 5556
rect 20346 5516 20352 5528
rect 20404 5516 20410 5568
rect 21818 5556 21824 5568
rect 21779 5528 21824 5556
rect 21818 5516 21824 5528
rect 21876 5516 21882 5568
rect 22094 5556 22100 5568
rect 22055 5528 22100 5556
rect 22094 5516 22100 5528
rect 22152 5516 22158 5568
rect 22278 5516 22284 5568
rect 22336 5556 22342 5568
rect 23661 5559 23719 5565
rect 23661 5556 23673 5559
rect 22336 5528 23673 5556
rect 22336 5516 22342 5528
rect 23661 5525 23673 5528
rect 23707 5525 23719 5559
rect 23661 5519 23719 5525
rect 27430 5516 27436 5568
rect 27488 5556 27494 5568
rect 27525 5559 27583 5565
rect 27525 5556 27537 5559
rect 27488 5528 27537 5556
rect 27488 5516 27494 5528
rect 27525 5525 27537 5528
rect 27571 5525 27583 5559
rect 27890 5556 27896 5568
rect 27851 5528 27896 5556
rect 27525 5519 27583 5525
rect 27890 5516 27896 5528
rect 27948 5516 27954 5568
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 1026 5312 1032 5364
rect 1084 5352 1090 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1084 5324 1593 5352
rect 1084 5312 1090 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 2406 5352 2412 5364
rect 2367 5324 2412 5352
rect 1581 5315 1639 5321
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 6546 5352 6552 5364
rect 5951 5324 6552 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 7374 5352 7380 5364
rect 6840 5324 7380 5352
rect 1762 5176 1768 5228
rect 1820 5216 1826 5228
rect 6840 5225 6868 5324
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 9122 5352 9128 5364
rect 8803 5324 9128 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 10505 5355 10563 5361
rect 10505 5352 10517 5355
rect 10468 5324 10517 5352
rect 10468 5312 10474 5324
rect 10505 5321 10517 5324
rect 10551 5352 10563 5355
rect 10781 5355 10839 5361
rect 10781 5352 10793 5355
rect 10551 5324 10793 5352
rect 10551 5321 10563 5324
rect 10505 5315 10563 5321
rect 10781 5321 10793 5324
rect 10827 5321 10839 5355
rect 10781 5315 10839 5321
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 13538 5352 13544 5364
rect 12299 5324 13544 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 9493 5287 9551 5293
rect 9493 5253 9505 5287
rect 9539 5284 9551 5287
rect 12268 5284 12296 5315
rect 13538 5312 13544 5324
rect 13596 5352 13602 5364
rect 15654 5352 15660 5364
rect 13596 5324 14688 5352
rect 15615 5324 15660 5352
rect 13596 5312 13602 5324
rect 9539 5256 12296 5284
rect 9539 5253 9551 5256
rect 9493 5247 9551 5253
rect 6825 5219 6883 5225
rect 1820 5188 3464 5216
rect 1820 5176 1826 5188
rect 3436 5160 3464 5188
rect 6825 5185 6837 5219
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 7837 5219 7895 5225
rect 7837 5185 7849 5219
rect 7883 5216 7895 5219
rect 8110 5216 8116 5228
rect 7883 5188 8116 5216
rect 7883 5185 7895 5188
rect 7837 5179 7895 5185
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 2038 5148 2044 5160
rect 1443 5120 2044 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 2130 5108 2136 5160
rect 2188 5148 2194 5160
rect 2777 5151 2835 5157
rect 2777 5148 2789 5151
rect 2188 5120 2789 5148
rect 2188 5108 2194 5120
rect 2777 5117 2789 5120
rect 2823 5117 2835 5151
rect 3050 5148 3056 5160
rect 3011 5120 3056 5148
rect 2777 5111 2835 5117
rect 2792 5080 2820 5111
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 3418 5108 3424 5160
rect 3476 5148 3482 5160
rect 3881 5151 3939 5157
rect 3476 5120 3569 5148
rect 3476 5108 3482 5120
rect 3881 5117 3893 5151
rect 3927 5148 3939 5151
rect 4062 5148 4068 5160
rect 3927 5120 4068 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5148 5043 5151
rect 5074 5148 5080 5160
rect 5031 5120 5080 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 9125 5151 9183 5157
rect 9125 5117 9137 5151
rect 9171 5148 9183 5151
rect 9582 5148 9588 5160
rect 9171 5120 9588 5148
rect 9171 5117 9183 5120
rect 9125 5111 9183 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 5166 5080 5172 5092
rect 2792 5052 5172 5080
rect 5166 5040 5172 5052
rect 5224 5040 5230 5092
rect 5347 5083 5405 5089
rect 5347 5049 5359 5083
rect 5393 5080 5405 5083
rect 6270 5080 6276 5092
rect 5393 5052 6276 5080
rect 5393 5049 5405 5052
rect 5347 5043 5405 5049
rect 2590 5012 2596 5024
rect 2551 4984 2596 5012
rect 2590 4972 2596 4984
rect 2648 4972 2654 5024
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 4430 5012 4436 5024
rect 4387 4984 4436 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 4430 4972 4436 4984
rect 4488 5012 4494 5024
rect 4893 5015 4951 5021
rect 4893 5012 4905 5015
rect 4488 4984 4905 5012
rect 4488 4972 4494 4984
rect 4893 4981 4905 4984
rect 4939 5012 4951 5015
rect 5362 5012 5390 5043
rect 6270 5040 6276 5052
rect 6328 5080 6334 5092
rect 8202 5089 8208 5092
rect 7745 5083 7803 5089
rect 7745 5080 7757 5083
rect 6328 5052 7757 5080
rect 6328 5040 6334 5052
rect 7745 5049 7757 5052
rect 7791 5080 7803 5083
rect 8199 5080 8208 5089
rect 7791 5052 8208 5080
rect 7791 5049 7803 5052
rect 7745 5043 7803 5049
rect 8199 5043 8208 5052
rect 8260 5080 8266 5092
rect 9921 5089 9949 5256
rect 13814 5244 13820 5296
rect 13872 5284 13878 5296
rect 14660 5293 14688 5324
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 18966 5352 18972 5364
rect 18927 5324 18972 5352
rect 18966 5312 18972 5324
rect 19024 5312 19030 5364
rect 20714 5352 20720 5364
rect 20627 5324 20720 5352
rect 20714 5312 20720 5324
rect 20772 5352 20778 5364
rect 22922 5352 22928 5364
rect 20772 5324 22928 5352
rect 20772 5312 20778 5324
rect 22922 5312 22928 5324
rect 22980 5312 22986 5364
rect 23799 5355 23857 5361
rect 23799 5321 23811 5355
rect 23845 5352 23857 5355
rect 24394 5352 24400 5364
rect 23845 5324 24400 5352
rect 23845 5321 23857 5324
rect 23799 5315 23857 5321
rect 24394 5312 24400 5324
rect 24452 5312 24458 5364
rect 24578 5352 24584 5364
rect 24539 5324 24584 5352
rect 24578 5312 24584 5324
rect 24636 5312 24642 5364
rect 27246 5352 27252 5364
rect 27207 5324 27252 5352
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 35621 5355 35679 5361
rect 35621 5321 35633 5355
rect 35667 5352 35679 5355
rect 35802 5352 35808 5364
rect 35667 5324 35808 5352
rect 35667 5321 35679 5324
rect 35621 5315 35679 5321
rect 35802 5312 35808 5324
rect 35860 5312 35866 5364
rect 14645 5287 14703 5293
rect 13872 5256 13917 5284
rect 13872 5244 13878 5256
rect 14645 5253 14657 5287
rect 14691 5284 14703 5287
rect 18138 5284 18144 5296
rect 14691 5256 18144 5284
rect 14691 5253 14703 5256
rect 14645 5247 14703 5253
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 11149 5219 11207 5225
rect 11149 5216 11161 5219
rect 10560 5188 11161 5216
rect 10560 5176 10566 5188
rect 11149 5185 11161 5188
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 11609 5219 11667 5225
rect 11609 5185 11621 5219
rect 11655 5216 11667 5219
rect 11655 5188 12940 5216
rect 11655 5185 11667 5188
rect 11609 5179 11667 5185
rect 11333 5151 11391 5157
rect 11333 5117 11345 5151
rect 11379 5148 11391 5151
rect 11379 5120 11836 5148
rect 11379 5117 11391 5120
rect 11333 5111 11391 5117
rect 9906 5083 9964 5089
rect 9906 5080 9918 5083
rect 8260 5052 9918 5080
rect 8202 5040 8208 5043
rect 8260 5040 8266 5052
rect 9906 5049 9918 5052
rect 9952 5049 9964 5083
rect 9906 5043 9964 5049
rect 11808 5024 11836 5120
rect 12342 5108 12348 5160
rect 12400 5148 12406 5160
rect 12912 5157 12940 5188
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 12400 5120 12449 5148
rect 12400 5108 12406 5120
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5117 12955 5151
rect 13262 5148 13268 5160
rect 13223 5120 13268 5148
rect 12897 5111 12955 5117
rect 12912 5080 12940 5111
rect 13262 5108 13268 5120
rect 13320 5108 13326 5160
rect 13538 5108 13544 5160
rect 13596 5148 13602 5160
rect 13633 5151 13691 5157
rect 13633 5148 13645 5151
rect 13596 5120 13645 5148
rect 13596 5108 13602 5120
rect 13633 5117 13645 5120
rect 13679 5117 13691 5151
rect 13633 5111 13691 5117
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 13872 5120 14749 5148
rect 13872 5108 13878 5120
rect 14737 5117 14749 5120
rect 14783 5148 14795 5151
rect 15010 5148 15016 5160
rect 14783 5120 15016 5148
rect 14783 5117 14795 5120
rect 14737 5111 14795 5117
rect 15010 5108 15016 5120
rect 15068 5108 15074 5160
rect 15120 5089 15148 5256
rect 18138 5244 18144 5256
rect 18196 5244 18202 5296
rect 21542 5244 21548 5296
rect 21600 5284 21606 5296
rect 24210 5284 24216 5296
rect 21600 5256 21680 5284
rect 24171 5256 24216 5284
rect 21600 5244 21606 5256
rect 17126 5176 17132 5228
rect 17184 5216 17190 5228
rect 17770 5216 17776 5228
rect 17184 5188 17776 5216
rect 17184 5176 17190 5188
rect 17770 5176 17776 5188
rect 17828 5216 17834 5228
rect 18049 5219 18107 5225
rect 18049 5216 18061 5219
rect 17828 5188 18061 5216
rect 17828 5176 17834 5188
rect 18049 5185 18061 5188
rect 18095 5185 18107 5219
rect 21358 5216 21364 5228
rect 18049 5179 18107 5185
rect 18248 5188 21364 5216
rect 16574 5108 16580 5160
rect 16632 5148 16638 5160
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 16632 5120 16681 5148
rect 16632 5108 16638 5120
rect 16669 5117 16681 5120
rect 16715 5148 16727 5151
rect 17313 5151 17371 5157
rect 17313 5148 17325 5151
rect 16715 5120 17325 5148
rect 16715 5117 16727 5120
rect 16669 5111 16727 5117
rect 17313 5117 17325 5120
rect 17359 5117 17371 5151
rect 17313 5111 17371 5117
rect 14185 5083 14243 5089
rect 14185 5080 14197 5083
rect 12912 5052 14197 5080
rect 14185 5049 14197 5052
rect 14231 5049 14243 5083
rect 14185 5043 14243 5049
rect 15099 5083 15157 5089
rect 15099 5049 15111 5083
rect 15145 5049 15157 5083
rect 15099 5043 15157 5049
rect 15286 5040 15292 5092
rect 15344 5080 15350 5092
rect 16301 5083 16359 5089
rect 16301 5080 16313 5083
rect 15344 5052 16313 5080
rect 15344 5040 15350 5052
rect 16301 5049 16313 5052
rect 16347 5080 16359 5083
rect 16485 5083 16543 5089
rect 16485 5080 16497 5083
rect 16347 5052 16497 5080
rect 16347 5049 16359 5052
rect 16301 5043 16359 5049
rect 16485 5049 16497 5052
rect 16531 5049 16543 5083
rect 16485 5043 16543 5049
rect 17037 5083 17095 5089
rect 17037 5049 17049 5083
rect 17083 5080 17095 5083
rect 18248 5080 18276 5188
rect 21358 5176 21364 5188
rect 21416 5176 21422 5228
rect 21652 5225 21680 5256
rect 24210 5244 24216 5256
rect 24268 5244 24274 5296
rect 25314 5284 25320 5296
rect 25275 5256 25320 5284
rect 25314 5244 25320 5256
rect 25372 5244 25378 5296
rect 21637 5219 21695 5225
rect 21637 5185 21649 5219
rect 21683 5185 21695 5219
rect 22278 5216 22284 5228
rect 22239 5188 22284 5216
rect 21637 5179 21695 5185
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 19794 5148 19800 5160
rect 19755 5120 19800 5148
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 23728 5151 23786 5157
rect 23728 5117 23740 5151
rect 23774 5148 23786 5151
rect 24228 5148 24256 5244
rect 24765 5219 24823 5225
rect 24765 5185 24777 5219
rect 24811 5216 24823 5219
rect 25222 5216 25228 5228
rect 24811 5188 25228 5216
rect 24811 5185 24823 5188
rect 24765 5179 24823 5185
rect 25222 5176 25228 5188
rect 25280 5216 25286 5228
rect 25406 5216 25412 5228
rect 25280 5188 25412 5216
rect 25280 5176 25286 5188
rect 25406 5176 25412 5188
rect 25464 5176 25470 5228
rect 26786 5176 26792 5228
rect 26844 5216 26850 5228
rect 27525 5219 27583 5225
rect 27525 5216 27537 5219
rect 26844 5188 27537 5216
rect 26844 5176 26850 5188
rect 27525 5185 27537 5188
rect 27571 5216 27583 5219
rect 27890 5216 27896 5228
rect 27571 5188 27896 5216
rect 27571 5185 27583 5188
rect 27525 5179 27583 5185
rect 27890 5176 27896 5188
rect 27948 5176 27954 5228
rect 23774 5120 24256 5148
rect 26472 5151 26530 5157
rect 23774 5117 23786 5120
rect 23728 5111 23786 5117
rect 26472 5117 26484 5151
rect 26518 5148 26530 5151
rect 26970 5148 26976 5160
rect 26518 5120 26976 5148
rect 26518 5117 26530 5120
rect 26472 5111 26530 5117
rect 26970 5108 26976 5120
rect 27028 5108 27034 5160
rect 35434 5148 35440 5160
rect 35395 5120 35440 5148
rect 35434 5108 35440 5120
rect 35492 5148 35498 5160
rect 35989 5151 36047 5157
rect 35989 5148 36001 5151
rect 35492 5120 36001 5148
rect 35492 5108 35498 5120
rect 35989 5117 36001 5120
rect 36035 5117 36047 5151
rect 35989 5111 36047 5117
rect 18411 5083 18469 5089
rect 18411 5080 18423 5083
rect 17083 5052 18276 5080
rect 18340 5052 18423 5080
rect 17083 5049 17095 5052
rect 17037 5043 17095 5049
rect 6638 5012 6644 5024
rect 4939 4984 5390 5012
rect 6599 4984 6644 5012
rect 4939 4981 4951 4984
rect 4893 4975 4951 4981
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 10410 4972 10416 5024
rect 10468 5012 10474 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 10468 4984 11529 5012
rect 10468 4972 10474 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11790 5012 11796 5024
rect 11751 4984 11796 5012
rect 11517 4975 11575 4981
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 15654 4972 15660 5024
rect 15712 5012 15718 5024
rect 15933 5015 15991 5021
rect 15933 5012 15945 5015
rect 15712 4984 15945 5012
rect 15712 4972 15718 4984
rect 15933 4981 15945 4984
rect 15979 5012 15991 5015
rect 16942 5012 16948 5024
rect 15979 4984 16948 5012
rect 15979 4981 15991 4984
rect 15933 4975 15991 4981
rect 16942 4972 16948 4984
rect 17000 4972 17006 5024
rect 17865 5015 17923 5021
rect 17865 4981 17877 5015
rect 17911 5012 17923 5015
rect 18138 5012 18144 5024
rect 17911 4984 18144 5012
rect 17911 4981 17923 4984
rect 17865 4975 17923 4981
rect 18138 4972 18144 4984
rect 18196 5012 18202 5024
rect 18340 5012 18368 5052
rect 18411 5049 18423 5052
rect 18457 5080 18469 5083
rect 20159 5083 20217 5089
rect 18457 5052 19748 5080
rect 18457 5049 18469 5052
rect 18411 5043 18469 5049
rect 18196 4984 18368 5012
rect 18196 4972 18202 4984
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19720 5021 19748 5052
rect 20159 5049 20171 5083
rect 20205 5049 20217 5083
rect 20159 5043 20217 5049
rect 19705 5015 19763 5021
rect 19392 4984 19437 5012
rect 19392 4972 19398 4984
rect 19705 4981 19717 5015
rect 19751 5012 19763 5015
rect 20174 5012 20202 5043
rect 20622 5040 20628 5092
rect 20680 5080 20686 5092
rect 21361 5083 21419 5089
rect 21361 5080 21373 5083
rect 20680 5052 21373 5080
rect 20680 5040 20686 5052
rect 21361 5049 21373 5052
rect 21407 5049 21419 5083
rect 21361 5043 21419 5049
rect 21726 5040 21732 5092
rect 21784 5080 21790 5092
rect 22094 5080 22100 5092
rect 21784 5052 22100 5080
rect 21784 5040 21790 5052
rect 22094 5040 22100 5052
rect 22152 5040 22158 5092
rect 24854 5080 24860 5092
rect 24815 5052 24860 5080
rect 24854 5040 24860 5052
rect 24912 5040 24918 5092
rect 26559 5083 26617 5089
rect 26559 5049 26571 5083
rect 26605 5080 26617 5083
rect 27154 5080 27160 5092
rect 26605 5052 27160 5080
rect 26605 5049 26617 5052
rect 26559 5043 26617 5049
rect 27154 5040 27160 5052
rect 27212 5040 27218 5092
rect 27617 5083 27675 5089
rect 27617 5049 27629 5083
rect 27663 5049 27675 5083
rect 27617 5043 27675 5049
rect 28169 5083 28227 5089
rect 28169 5049 28181 5083
rect 28215 5080 28227 5083
rect 28258 5080 28264 5092
rect 28215 5052 28264 5080
rect 28215 5049 28227 5052
rect 28169 5043 28227 5049
rect 21085 5015 21143 5021
rect 21085 5012 21097 5015
rect 19751 4984 21097 5012
rect 19751 4981 19763 4984
rect 19705 4975 19763 4981
rect 21085 4981 21097 4984
rect 21131 5012 21143 5015
rect 21266 5012 21272 5024
rect 21131 4984 21272 5012
rect 21131 4981 21143 4984
rect 21085 4975 21143 4981
rect 21266 4972 21272 4984
rect 21324 5012 21330 5024
rect 22278 5012 22284 5024
rect 21324 4984 22284 5012
rect 21324 4972 21330 4984
rect 22278 4972 22284 4984
rect 22336 4972 22342 5024
rect 22649 5015 22707 5021
rect 22649 4981 22661 5015
rect 22695 5012 22707 5015
rect 22830 5012 22836 5024
rect 22695 4984 22836 5012
rect 22695 4981 22707 4984
rect 22649 4975 22707 4981
rect 22830 4972 22836 4984
rect 22888 4972 22894 5024
rect 23474 4972 23480 5024
rect 23532 5012 23538 5024
rect 24872 5012 24900 5040
rect 25685 5015 25743 5021
rect 25685 5012 25697 5015
rect 23532 4984 23577 5012
rect 24872 4984 25697 5012
rect 23532 4972 23538 4984
rect 25685 4981 25697 4984
rect 25731 4981 25743 5015
rect 26970 5012 26976 5024
rect 26931 4984 26976 5012
rect 25685 4975 25743 4981
rect 26970 4972 26976 4984
rect 27028 4972 27034 5024
rect 27430 4972 27436 5024
rect 27488 5012 27494 5024
rect 27632 5012 27660 5043
rect 28258 5040 28264 5052
rect 28316 5040 28322 5092
rect 27488 4984 27660 5012
rect 27488 4972 27494 4984
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2222 4808 2228 4820
rect 1995 4780 2228 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2222 4768 2228 4780
rect 2280 4808 2286 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 2280 4780 3801 4808
rect 2280 4768 2286 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 4522 4808 4528 4820
rect 4483 4780 4528 4808
rect 3789 4771 3847 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 5074 4808 5080 4820
rect 4987 4780 5080 4808
rect 5074 4768 5080 4780
rect 5132 4808 5138 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5132 4780 5273 4808
rect 5132 4768 5138 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 5261 4771 5319 4777
rect 7466 4768 7472 4820
rect 7524 4808 7530 4820
rect 7653 4811 7711 4817
rect 7653 4808 7665 4811
rect 7524 4780 7665 4808
rect 7524 4768 7530 4780
rect 7653 4777 7665 4780
rect 7699 4777 7711 4811
rect 8202 4808 8208 4820
rect 8163 4780 8208 4808
rect 7653 4771 7711 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8757 4811 8815 4817
rect 8757 4777 8769 4811
rect 8803 4808 8815 4811
rect 9490 4808 9496 4820
rect 8803 4780 9496 4808
rect 8803 4777 8815 4780
rect 8757 4771 8815 4777
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 9769 4811 9827 4817
rect 9769 4808 9781 4811
rect 9640 4780 9781 4808
rect 9640 4768 9646 4780
rect 9769 4777 9781 4780
rect 9815 4777 9827 4811
rect 9769 4771 9827 4777
rect 11701 4811 11759 4817
rect 11701 4777 11713 4811
rect 11747 4808 11759 4811
rect 12253 4811 12311 4817
rect 12253 4808 12265 4811
rect 11747 4780 12265 4808
rect 11747 4777 11759 4780
rect 11701 4771 11759 4777
rect 12253 4777 12265 4780
rect 12299 4808 12311 4811
rect 13538 4808 13544 4820
rect 12299 4780 13544 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 13814 4808 13820 4820
rect 13775 4780 13820 4808
rect 13814 4768 13820 4780
rect 13872 4768 13878 4820
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 14277 4811 14335 4817
rect 14277 4808 14289 4811
rect 14139 4780 14289 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 14277 4777 14289 4780
rect 14323 4808 14335 4811
rect 14734 4808 14740 4820
rect 14323 4780 14740 4808
rect 14323 4777 14335 4780
rect 14277 4771 14335 4777
rect 14734 4768 14740 4780
rect 14792 4808 14798 4820
rect 17589 4811 17647 4817
rect 14792 4780 15792 4808
rect 14792 4768 14798 4780
rect 2958 4740 2964 4752
rect 2424 4712 2964 4740
rect 1854 4672 1860 4684
rect 1815 4644 1860 4672
rect 1854 4632 1860 4644
rect 1912 4632 1918 4684
rect 2424 4681 2452 4712
rect 2958 4700 2964 4712
rect 3016 4700 3022 4752
rect 3510 4700 3516 4752
rect 3568 4740 3574 4752
rect 4203 4743 4261 4749
rect 4203 4740 4215 4743
rect 3568 4712 4215 4740
rect 3568 4700 3574 4712
rect 4203 4709 4215 4712
rect 4249 4709 4261 4743
rect 12342 4740 12348 4752
rect 4203 4703 4261 4709
rect 9784 4712 12348 4740
rect 9784 4684 9812 4712
rect 12342 4700 12348 4712
rect 12400 4700 12406 4752
rect 15105 4743 15163 4749
rect 15105 4709 15117 4743
rect 15151 4740 15163 4743
rect 15654 4740 15660 4752
rect 15151 4712 15660 4740
rect 15151 4709 15163 4712
rect 15105 4703 15163 4709
rect 15654 4700 15660 4712
rect 15712 4700 15718 4752
rect 15764 4749 15792 4780
rect 17589 4777 17601 4811
rect 17635 4808 17647 4811
rect 20622 4808 20628 4820
rect 17635 4780 20628 4808
rect 17635 4777 17647 4780
rect 17589 4771 17647 4777
rect 20622 4768 20628 4780
rect 20680 4768 20686 4820
rect 20717 4811 20775 4817
rect 20717 4777 20729 4811
rect 20763 4808 20775 4811
rect 21266 4808 21272 4820
rect 20763 4780 21272 4808
rect 20763 4777 20775 4780
rect 20717 4771 20775 4777
rect 21266 4768 21272 4780
rect 21324 4808 21330 4820
rect 21818 4808 21824 4820
rect 21324 4780 21824 4808
rect 21324 4768 21330 4780
rect 21818 4768 21824 4780
rect 21876 4768 21882 4820
rect 22002 4768 22008 4820
rect 22060 4808 22066 4820
rect 22097 4811 22155 4817
rect 22097 4808 22109 4811
rect 22060 4780 22109 4808
rect 22060 4768 22066 4780
rect 22097 4777 22109 4780
rect 22143 4777 22155 4811
rect 22097 4771 22155 4777
rect 15749 4743 15807 4749
rect 15749 4709 15761 4743
rect 15795 4740 15807 4743
rect 16114 4740 16120 4752
rect 15795 4712 16120 4740
rect 15795 4709 15807 4712
rect 15749 4703 15807 4709
rect 16114 4700 16120 4712
rect 16172 4740 16178 4752
rect 18322 4740 18328 4752
rect 16172 4712 18328 4740
rect 16172 4700 16178 4712
rect 2409 4675 2467 4681
rect 2409 4641 2421 4675
rect 2455 4641 2467 4675
rect 2409 4635 2467 4641
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4641 2743 4675
rect 2685 4635 2743 4641
rect 3053 4675 3111 4681
rect 3053 4641 3065 4675
rect 3099 4672 3111 4675
rect 3099 4644 3556 4672
rect 3099 4641 3111 4644
rect 3053 4635 3111 4641
rect 2700 4604 2728 4635
rect 3234 4604 3240 4616
rect 2700 4576 3240 4604
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 3528 4545 3556 4644
rect 3602 4632 3608 4684
rect 3660 4672 3666 4684
rect 4111 4675 4169 4681
rect 4111 4672 4123 4675
rect 3660 4644 4123 4672
rect 3660 4632 3666 4644
rect 4111 4641 4123 4644
rect 4157 4641 4169 4675
rect 5166 4672 5172 4684
rect 5127 4644 5172 4672
rect 4111 4635 4169 4641
rect 4126 4604 4154 4635
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5718 4672 5724 4684
rect 5679 4644 5724 4672
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 6178 4672 6184 4684
rect 6139 4644 6184 4672
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6454 4672 6460 4684
rect 6415 4644 6460 4672
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 9766 4672 9772 4684
rect 9727 4644 9772 4672
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 10410 4672 10416 4684
rect 10371 4644 10416 4672
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 10594 4672 10600 4684
rect 10555 4644 10600 4672
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 10962 4632 10968 4684
rect 11020 4672 11026 4684
rect 11057 4675 11115 4681
rect 11057 4672 11069 4675
rect 11020 4644 11069 4672
rect 11020 4632 11026 4644
rect 11057 4641 11069 4644
rect 11103 4672 11115 4675
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 11103 4644 11713 4672
rect 11103 4641 11115 4644
rect 11057 4635 11115 4641
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 11701 4635 11759 4641
rect 11882 4632 11888 4684
rect 11940 4672 11946 4684
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 11940 4644 12449 4672
rect 11940 4632 11946 4644
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 12894 4672 12900 4684
rect 12855 4644 12900 4672
rect 12437 4635 12495 4641
rect 12894 4632 12900 4644
rect 12952 4632 12958 4684
rect 13262 4672 13268 4684
rect 13223 4644 13268 4672
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 13538 4632 13544 4684
rect 13596 4672 13602 4684
rect 13725 4675 13783 4681
rect 13725 4672 13737 4675
rect 13596 4644 13737 4672
rect 13596 4632 13602 4644
rect 13725 4641 13737 4644
rect 13771 4672 13783 4675
rect 13814 4672 13820 4684
rect 13771 4644 13820 4672
rect 13771 4641 13783 4644
rect 13725 4635 13783 4641
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 16206 4672 16212 4684
rect 16167 4644 16212 4672
rect 16206 4632 16212 4644
rect 16264 4632 16270 4684
rect 16960 4681 16988 4712
rect 18322 4700 18328 4712
rect 18380 4700 18386 4752
rect 19794 4700 19800 4752
rect 19852 4740 19858 4752
rect 19981 4743 20039 4749
rect 19981 4740 19993 4743
rect 19852 4712 19993 4740
rect 19852 4700 19858 4712
rect 19981 4709 19993 4712
rect 20027 4740 20039 4743
rect 20257 4743 20315 4749
rect 20257 4740 20269 4743
rect 20027 4712 20269 4740
rect 20027 4709 20039 4712
rect 19981 4703 20039 4709
rect 20257 4709 20269 4712
rect 20303 4709 20315 4743
rect 20257 4703 20315 4709
rect 20806 4700 20812 4752
rect 20864 4740 20870 4752
rect 21039 4743 21097 4749
rect 21039 4740 21051 4743
rect 20864 4712 21051 4740
rect 20864 4700 20870 4712
rect 21039 4709 21051 4712
rect 21085 4709 21097 4743
rect 21358 4740 21364 4752
rect 21319 4712 21364 4740
rect 21039 4703 21097 4709
rect 21358 4700 21364 4712
rect 21416 4740 21422 4752
rect 21910 4740 21916 4752
rect 21416 4712 21916 4740
rect 21416 4700 21422 4712
rect 21910 4700 21916 4712
rect 21968 4700 21974 4752
rect 16945 4675 17003 4681
rect 16945 4641 16957 4675
rect 16991 4641 17003 4675
rect 17218 4672 17224 4684
rect 17179 4644 17224 4672
rect 16945 4635 17003 4641
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 17405 4675 17463 4681
rect 17405 4641 17417 4675
rect 17451 4641 17463 4675
rect 17405 4635 17463 4641
rect 4246 4604 4252 4616
rect 4126 4576 4252 4604
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4604 7895 4607
rect 8018 4604 8024 4616
rect 7883 4576 8024 4604
rect 7883 4573 7895 4576
rect 7837 4567 7895 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 12912 4604 12940 4632
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 12912 4576 14105 4604
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4604 16175 4607
rect 17236 4604 17264 4632
rect 16163 4576 17264 4604
rect 17420 4604 17448 4635
rect 18046 4632 18052 4684
rect 18104 4672 18110 4684
rect 18509 4675 18567 4681
rect 18509 4672 18521 4675
rect 18104 4644 18521 4672
rect 18104 4632 18110 4644
rect 18509 4641 18521 4644
rect 18555 4641 18567 4675
rect 18509 4635 18567 4641
rect 18969 4675 19027 4681
rect 18969 4641 18981 4675
rect 19015 4641 19027 4675
rect 18969 4635 19027 4641
rect 18874 4604 18880 4616
rect 17420 4576 18880 4604
rect 16163 4573 16175 4576
rect 16117 4567 16175 4573
rect 3513 4539 3571 4545
rect 3513 4505 3525 4539
rect 3559 4536 3571 4539
rect 4062 4536 4068 4548
rect 3559 4508 4068 4536
rect 3559 4505 3571 4508
rect 3513 4499 3571 4505
rect 4062 4496 4068 4508
rect 4120 4496 4126 4548
rect 12802 4496 12808 4548
rect 12860 4536 12866 4548
rect 16132 4536 16160 4567
rect 12860 4508 16160 4536
rect 12860 4496 12866 4508
rect 16942 4496 16948 4548
rect 17000 4536 17006 4548
rect 17420 4536 17448 4576
rect 18874 4564 18880 4576
rect 18932 4564 18938 4616
rect 17000 4508 17448 4536
rect 18049 4539 18107 4545
rect 17000 4496 17006 4508
rect 18049 4505 18061 4539
rect 18095 4536 18107 4539
rect 18138 4536 18144 4548
rect 18095 4508 18144 4536
rect 18095 4505 18107 4508
rect 18049 4499 18107 4505
rect 18138 4496 18144 4508
rect 18196 4496 18202 4548
rect 18322 4496 18328 4548
rect 18380 4536 18386 4548
rect 18417 4539 18475 4545
rect 18417 4536 18429 4539
rect 18380 4508 18429 4536
rect 18380 4496 18386 4508
rect 18417 4505 18429 4508
rect 18463 4536 18475 4539
rect 18984 4536 19012 4635
rect 19334 4632 19340 4684
rect 19392 4672 19398 4684
rect 19702 4672 19708 4684
rect 19392 4644 19437 4672
rect 19663 4644 19708 4672
rect 19392 4632 19398 4644
rect 19702 4632 19708 4644
rect 19760 4632 19766 4684
rect 20438 4632 20444 4684
rect 20496 4672 20502 4684
rect 20936 4675 20994 4681
rect 20936 4672 20948 4675
rect 20496 4644 20948 4672
rect 20496 4632 20502 4644
rect 20936 4641 20948 4644
rect 20982 4672 20994 4675
rect 21634 4672 21640 4684
rect 20982 4644 21640 4672
rect 20982 4641 20994 4644
rect 20936 4635 20994 4641
rect 21634 4632 21640 4644
rect 21692 4632 21698 4684
rect 22112 4672 22140 4771
rect 23474 4768 23480 4820
rect 23532 4808 23538 4820
rect 23532 4780 23577 4808
rect 23532 4768 23538 4780
rect 23934 4768 23940 4820
rect 23992 4808 23998 4820
rect 24029 4811 24087 4817
rect 24029 4808 24041 4811
rect 23992 4780 24041 4808
rect 23992 4768 23998 4780
rect 24029 4777 24041 4780
rect 24075 4777 24087 4811
rect 24486 4808 24492 4820
rect 24447 4780 24492 4808
rect 24029 4771 24087 4777
rect 24486 4768 24492 4780
rect 24544 4768 24550 4820
rect 24946 4808 24952 4820
rect 24907 4780 24952 4808
rect 24946 4768 24952 4780
rect 25004 4768 25010 4820
rect 25498 4808 25504 4820
rect 25459 4780 25504 4808
rect 25498 4768 25504 4780
rect 25556 4768 25562 4820
rect 26878 4768 26884 4820
rect 26936 4768 26942 4820
rect 24302 4700 24308 4752
rect 24360 4740 24366 4752
rect 25314 4740 25320 4752
rect 24360 4712 25320 4740
rect 24360 4700 24366 4712
rect 25314 4700 25320 4712
rect 25372 4700 25378 4752
rect 26896 4740 26924 4768
rect 27706 4740 27712 4752
rect 26563 4712 26924 4740
rect 27667 4712 27712 4740
rect 22281 4675 22339 4681
rect 22281 4672 22293 4675
rect 22112 4644 22293 4672
rect 22281 4641 22293 4644
rect 22327 4641 22339 4675
rect 22738 4672 22744 4684
rect 22699 4644 22744 4672
rect 22281 4635 22339 4641
rect 22738 4632 22744 4644
rect 22796 4632 22802 4684
rect 22830 4632 22836 4684
rect 22888 4672 22894 4684
rect 23106 4672 23112 4684
rect 22888 4644 23112 4672
rect 22888 4632 22894 4644
rect 23106 4632 23112 4644
rect 23164 4632 23170 4684
rect 26563 4681 26591 4712
rect 27706 4700 27712 4712
rect 27764 4700 27770 4752
rect 28258 4740 28264 4752
rect 28219 4712 28264 4740
rect 28258 4700 28264 4712
rect 28316 4700 28322 4752
rect 30282 4700 30288 4752
rect 30340 4740 30346 4752
rect 30340 4712 30763 4740
rect 30340 4700 30346 4712
rect 23477 4675 23535 4681
rect 23477 4641 23489 4675
rect 23523 4641 23535 4675
rect 23477 4635 23535 4641
rect 26548 4675 26606 4681
rect 26548 4641 26560 4675
rect 26594 4641 26606 4675
rect 29178 4672 29184 4684
rect 29139 4644 29184 4672
rect 26548 4635 26606 4641
rect 21821 4607 21879 4613
rect 21821 4573 21833 4607
rect 21867 4604 21879 4607
rect 22094 4604 22100 4616
rect 21867 4576 22100 4604
rect 21867 4573 21879 4576
rect 21821 4567 21879 4573
rect 22094 4564 22100 4576
rect 22152 4564 22158 4616
rect 23014 4564 23020 4616
rect 23072 4604 23078 4616
rect 23492 4604 23520 4635
rect 29178 4632 29184 4644
rect 29236 4632 29242 4684
rect 30735 4681 30763 4712
rect 30720 4675 30778 4681
rect 30720 4641 30732 4675
rect 30766 4672 30778 4675
rect 31386 4672 31392 4684
rect 30766 4644 31392 4672
rect 30766 4641 30778 4644
rect 30720 4635 30778 4641
rect 31386 4632 31392 4644
rect 31444 4632 31450 4684
rect 23072 4576 23520 4604
rect 24581 4607 24639 4613
rect 23072 4564 23078 4576
rect 24581 4573 24593 4607
rect 24627 4604 24639 4607
rect 24762 4604 24768 4616
rect 24627 4576 24768 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 24762 4564 24768 4576
rect 24820 4564 24826 4616
rect 27154 4564 27160 4616
rect 27212 4604 27218 4616
rect 27617 4607 27675 4613
rect 27617 4604 27629 4607
rect 27212 4576 27629 4604
rect 27212 4564 27218 4576
rect 27617 4573 27629 4576
rect 27663 4604 27675 4607
rect 28074 4604 28080 4616
rect 27663 4576 28080 4604
rect 27663 4573 27675 4576
rect 27617 4567 27675 4573
rect 28074 4564 28080 4576
rect 28132 4564 28138 4616
rect 18463 4508 19012 4536
rect 18463 4505 18475 4508
rect 18417 4499 18475 4505
rect 26418 4496 26424 4548
rect 26476 4536 26482 4548
rect 27341 4539 27399 4545
rect 27341 4536 27353 4539
rect 26476 4508 27353 4536
rect 26476 4496 26482 4508
rect 27341 4505 27353 4508
rect 27387 4505 27399 4539
rect 27341 4499 27399 4505
rect 9125 4471 9183 4477
rect 9125 4437 9137 4471
rect 9171 4468 9183 4471
rect 9490 4468 9496 4480
rect 9171 4440 9496 4468
rect 9171 4437 9183 4440
rect 9125 4431 9183 4437
rect 9490 4428 9496 4440
rect 9548 4428 9554 4480
rect 9858 4428 9864 4480
rect 9916 4468 9922 4480
rect 11517 4471 11575 4477
rect 11517 4468 11529 4471
rect 9916 4440 11529 4468
rect 9916 4428 9922 4440
rect 11517 4437 11529 4440
rect 11563 4468 11575 4471
rect 11882 4468 11888 4480
rect 11563 4440 11888 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 14642 4468 14648 4480
rect 14603 4440 14648 4468
rect 14642 4428 14648 4440
rect 14700 4428 14706 4480
rect 26651 4471 26709 4477
rect 26651 4437 26663 4471
rect 26697 4468 26709 4471
rect 26786 4468 26792 4480
rect 26697 4440 26792 4468
rect 26697 4437 26709 4440
rect 26651 4431 26709 4437
rect 26786 4428 26792 4440
rect 26844 4428 26850 4480
rect 27065 4471 27123 4477
rect 27065 4437 27077 4471
rect 27111 4468 27123 4471
rect 27246 4468 27252 4480
rect 27111 4440 27252 4468
rect 27111 4437 27123 4440
rect 27065 4431 27123 4437
rect 27246 4428 27252 4440
rect 27304 4428 27310 4480
rect 29546 4468 29552 4480
rect 29507 4440 29552 4468
rect 29546 4428 29552 4440
rect 29604 4428 29610 4480
rect 30558 4428 30564 4480
rect 30616 4468 30622 4480
rect 30791 4471 30849 4477
rect 30791 4468 30803 4471
rect 30616 4440 30803 4468
rect 30616 4428 30622 4440
rect 30791 4437 30803 4440
rect 30837 4437 30849 4471
rect 30791 4431 30849 4437
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 2130 4224 2136 4276
rect 2188 4264 2194 4276
rect 2225 4267 2283 4273
rect 2225 4264 2237 4267
rect 2188 4236 2237 4264
rect 2188 4224 2194 4236
rect 2225 4233 2237 4236
rect 2271 4233 2283 4267
rect 2225 4227 2283 4233
rect 2240 4060 2268 4227
rect 5166 4224 5172 4276
rect 5224 4264 5230 4276
rect 5721 4267 5779 4273
rect 5721 4264 5733 4267
rect 5224 4236 5733 4264
rect 5224 4224 5230 4236
rect 5721 4233 5733 4236
rect 5767 4233 5779 4267
rect 5721 4227 5779 4233
rect 6178 4224 6184 4276
rect 6236 4264 6242 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6236 4236 6561 4264
rect 6236 4224 6242 4236
rect 6549 4233 6561 4236
rect 6595 4264 6607 4267
rect 6595 4236 9444 4264
rect 6595 4233 6607 4236
rect 6549 4227 6607 4233
rect 6196 4196 6224 4224
rect 3712 4168 6224 4196
rect 7193 4199 7251 4205
rect 3712 4128 3740 4168
rect 7193 4165 7205 4199
rect 7239 4196 7251 4199
rect 8018 4196 8024 4208
rect 7239 4168 8024 4196
rect 7239 4165 7251 4168
rect 7193 4159 7251 4165
rect 8018 4156 8024 4168
rect 8076 4196 8082 4208
rect 8076 4168 8524 4196
rect 8076 4156 8082 4168
rect 3252 4100 3740 4128
rect 3252 4072 3280 4100
rect 4338 4088 4344 4140
rect 4396 4128 4402 4140
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 4396 4100 4813 4128
rect 4396 4088 4402 4100
rect 4801 4097 4813 4100
rect 4847 4128 4859 4131
rect 5074 4128 5080 4140
rect 4847 4100 5080 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5442 4128 5448 4140
rect 5403 4100 5448 4128
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8260 4100 8432 4128
rect 8260 4088 8266 4100
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 2240 4032 2421 4060
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 3050 4060 3056 4072
rect 2963 4032 3056 4060
rect 2409 4023 2467 4029
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 3234 4060 3240 4072
rect 3195 4032 3240 4060
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 3789 4063 3847 4069
rect 3789 4029 3801 4063
rect 3835 4060 3847 4063
rect 4062 4060 4068 4072
rect 3835 4032 4068 4060
rect 3835 4029 3847 4032
rect 3789 4023 3847 4029
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4060 7987 4063
rect 8294 4060 8300 4072
rect 7975 4032 8300 4060
rect 7975 4029 7987 4032
rect 7929 4023 7987 4029
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 8404 4069 8432 4100
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4029 8447 4063
rect 8389 4023 8447 4029
rect 3068 3992 3096 4020
rect 3510 3992 3516 4004
rect 3068 3964 3516 3992
rect 3510 3952 3516 3964
rect 3568 3952 3574 4004
rect 4893 3995 4951 4001
rect 4893 3961 4905 3995
rect 4939 3992 4951 3995
rect 4982 3992 4988 4004
rect 4939 3964 4988 3992
rect 4939 3961 4951 3964
rect 4893 3955 4951 3961
rect 4982 3952 4988 3964
rect 5040 3952 5046 4004
rect 5718 3952 5724 4004
rect 5776 3992 5782 4004
rect 7469 3995 7527 4001
rect 7469 3992 7481 3995
rect 5776 3964 7481 3992
rect 5776 3952 5782 3964
rect 7469 3961 7481 3964
rect 7515 3992 7527 3995
rect 8018 3992 8024 4004
rect 7515 3964 8024 3992
rect 7515 3961 7527 3964
rect 7469 3955 7527 3961
rect 8018 3952 8024 3964
rect 8076 3952 8082 4004
rect 1946 3924 1952 3936
rect 1907 3896 1952 3924
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 2498 3924 2504 3936
rect 2459 3896 2504 3924
rect 2498 3884 2504 3896
rect 2556 3884 2562 3936
rect 4246 3924 4252 3936
rect 4207 3896 4252 3924
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 4614 3924 4620 3936
rect 4575 3896 4620 3924
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4798 3884 4804 3936
rect 4856 3924 4862 3936
rect 6089 3927 6147 3933
rect 6089 3924 6101 3927
rect 4856 3896 6101 3924
rect 4856 3884 4862 3896
rect 6089 3893 6101 3896
rect 6135 3924 6147 3927
rect 6454 3924 6460 3936
rect 6135 3896 6460 3924
rect 6135 3893 6147 3896
rect 6089 3887 6147 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 8202 3924 8208 3936
rect 8163 3896 8208 3924
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8496 3933 8524 4168
rect 8570 4020 8576 4072
rect 8628 4060 8634 4072
rect 9416 4069 9444 4236
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 10505 4267 10563 4273
rect 10505 4264 10517 4267
rect 9824 4236 10517 4264
rect 9824 4224 9830 4236
rect 10505 4233 10517 4236
rect 10551 4233 10563 4267
rect 10962 4264 10968 4276
rect 10923 4236 10968 4264
rect 10505 4227 10563 4233
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 11517 4267 11575 4273
rect 11517 4233 11529 4267
rect 11563 4264 11575 4267
rect 12894 4264 12900 4276
rect 11563 4236 12900 4264
rect 11563 4233 11575 4236
rect 11517 4227 11575 4233
rect 12894 4224 12900 4236
rect 12952 4224 12958 4276
rect 14182 4224 14188 4276
rect 14240 4264 14246 4276
rect 14642 4264 14648 4276
rect 14240 4236 14648 4264
rect 14240 4224 14246 4236
rect 14642 4224 14648 4236
rect 14700 4264 14706 4276
rect 16482 4264 16488 4276
rect 14700 4236 16488 4264
rect 14700 4224 14706 4236
rect 16482 4224 16488 4236
rect 16540 4224 16546 4276
rect 18506 4224 18512 4276
rect 18564 4264 18570 4276
rect 19334 4264 19340 4276
rect 18564 4236 19340 4264
rect 18564 4224 18570 4236
rect 19334 4224 19340 4236
rect 19392 4224 19398 4276
rect 21269 4267 21327 4273
rect 21269 4233 21281 4267
rect 21315 4264 21327 4267
rect 21726 4264 21732 4276
rect 21315 4236 21732 4264
rect 21315 4233 21327 4236
rect 21269 4227 21327 4233
rect 21726 4224 21732 4236
rect 21784 4224 21790 4276
rect 22002 4264 22008 4276
rect 21963 4236 22008 4264
rect 22002 4224 22008 4236
rect 22060 4224 22066 4276
rect 24581 4267 24639 4273
rect 24581 4233 24593 4267
rect 24627 4264 24639 4267
rect 24854 4264 24860 4276
rect 24627 4236 24860 4264
rect 24627 4233 24639 4236
rect 24581 4227 24639 4233
rect 24854 4224 24860 4236
rect 24912 4224 24918 4276
rect 26326 4224 26332 4276
rect 26384 4264 26390 4276
rect 26421 4267 26479 4273
rect 26421 4264 26433 4267
rect 26384 4236 26433 4264
rect 26384 4224 26390 4236
rect 26421 4233 26433 4236
rect 26467 4264 26479 4267
rect 26878 4264 26884 4276
rect 26467 4236 26884 4264
rect 26467 4233 26479 4236
rect 26421 4227 26479 4233
rect 26878 4224 26884 4236
rect 26936 4224 26942 4276
rect 28074 4264 28080 4276
rect 28035 4236 28080 4264
rect 28074 4224 28080 4236
rect 28132 4224 28138 4276
rect 28442 4224 28448 4276
rect 28500 4264 28506 4276
rect 29089 4267 29147 4273
rect 29089 4264 29101 4267
rect 28500 4236 29101 4264
rect 28500 4224 28506 4236
rect 29089 4233 29101 4236
rect 29135 4264 29147 4267
rect 29178 4264 29184 4276
rect 29135 4236 29184 4264
rect 29135 4233 29147 4236
rect 29089 4227 29147 4233
rect 29178 4224 29184 4236
rect 29236 4224 29242 4276
rect 29822 4264 29828 4276
rect 29783 4236 29828 4264
rect 29822 4224 29828 4236
rect 29880 4224 29886 4276
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 12161 4199 12219 4205
rect 12161 4196 12173 4199
rect 10928 4168 12173 4196
rect 10928 4156 10934 4168
rect 12161 4165 12173 4168
rect 12207 4196 12219 4199
rect 13262 4196 13268 4208
rect 12207 4168 13268 4196
rect 12207 4165 12219 4168
rect 12161 4159 12219 4165
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 13722 4156 13728 4208
rect 13780 4196 13786 4208
rect 13817 4199 13875 4205
rect 13817 4196 13829 4199
rect 13780 4168 13829 4196
rect 13780 4156 13786 4168
rect 13817 4165 13829 4168
rect 13863 4165 13875 4199
rect 14734 4196 14740 4208
rect 14695 4168 14740 4196
rect 13817 4159 13875 4165
rect 14734 4156 14740 4168
rect 14792 4156 14798 4208
rect 17218 4156 17224 4208
rect 17276 4196 17282 4208
rect 17276 4168 18920 4196
rect 17276 4156 17282 4168
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 15473 4131 15531 4137
rect 15473 4128 15485 4131
rect 12400 4100 15485 4128
rect 12400 4088 12406 4100
rect 15473 4097 15485 4100
rect 15519 4128 15531 4131
rect 16206 4128 16212 4140
rect 15519 4100 16212 4128
rect 15519 4097 15531 4100
rect 15473 4091 15531 4097
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 8628 4032 8861 4060
rect 8628 4020 8634 4032
rect 8849 4029 8861 4032
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 9401 4063 9459 4069
rect 9401 4029 9413 4063
rect 9447 4029 9459 4063
rect 9401 4023 9459 4029
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3893 8539 3927
rect 9416 3924 9444 4023
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 9585 4063 9643 4069
rect 9585 4060 9597 4063
rect 9548 4032 9597 4060
rect 9548 4020 9554 4032
rect 9585 4029 9597 4032
rect 9631 4060 9643 4063
rect 10962 4060 10968 4072
rect 9631 4032 10968 4060
rect 9631 4029 9643 4032
rect 9585 4023 9643 4029
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 11790 4060 11796 4072
rect 11379 4032 11796 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 11882 4020 11888 4072
rect 11940 4060 11946 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 11940 4032 12449 4060
rect 11940 4020 11946 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12894 4060 12900 4072
rect 12855 4032 12900 4060
rect 12437 4023 12495 4029
rect 12452 3992 12480 4023
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 12986 4020 12992 4072
rect 13044 4060 13050 4072
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 13044 4032 13277 4060
rect 13044 4020 13050 4032
rect 13265 4029 13277 4032
rect 13311 4029 13323 4063
rect 13722 4060 13728 4072
rect 13683 4032 13728 4060
rect 13265 4023 13323 4029
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 15672 4069 15700 4100
rect 16206 4088 16212 4100
rect 16264 4088 16270 4140
rect 17126 4128 17132 4140
rect 17087 4100 17132 4128
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 18892 4128 18920 4168
rect 19889 4131 19947 4137
rect 19889 4128 19901 4131
rect 18892 4100 19901 4128
rect 15657 4063 15715 4069
rect 15657 4029 15669 4063
rect 15703 4029 15715 4063
rect 15657 4023 15715 4029
rect 16114 4020 16120 4072
rect 16172 4060 16178 4072
rect 16390 4060 16396 4072
rect 16172 4032 16396 4060
rect 16172 4020 16178 4032
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 16482 4020 16488 4072
rect 16540 4060 16546 4072
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 16540 4032 16681 4060
rect 16540 4020 16546 4032
rect 16669 4029 16681 4032
rect 16715 4029 16727 4063
rect 16942 4060 16948 4072
rect 16903 4032 16948 4060
rect 16669 4023 16727 4029
rect 16684 3992 16712 4023
rect 16942 4020 16948 4032
rect 17000 4020 17006 4072
rect 17681 4063 17739 4069
rect 17681 4029 17693 4063
rect 17727 4060 17739 4063
rect 18046 4060 18052 4072
rect 17727 4032 18052 4060
rect 17727 4029 17739 4032
rect 17681 4023 17739 4029
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 18322 4020 18328 4072
rect 18380 4060 18386 4072
rect 18782 4060 18788 4072
rect 18380 4032 18788 4060
rect 18380 4020 18386 4032
rect 18782 4020 18788 4032
rect 18840 4020 18846 4072
rect 18892 4060 18920 4100
rect 19889 4097 19901 4100
rect 19935 4128 19947 4131
rect 23014 4128 23020 4140
rect 19935 4100 23020 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 23014 4088 23020 4100
rect 23072 4088 23078 4140
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 23661 4131 23719 4137
rect 23661 4128 23673 4131
rect 23532 4100 23673 4128
rect 23532 4088 23538 4100
rect 23661 4097 23673 4100
rect 23707 4097 23719 4131
rect 23661 4091 23719 4097
rect 25314 4088 25320 4140
rect 25372 4128 25378 4140
rect 25958 4128 25964 4140
rect 25372 4100 25964 4128
rect 25372 4088 25378 4100
rect 19058 4060 19064 4072
rect 18892 4032 19064 4060
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 19429 4063 19487 4069
rect 19429 4029 19441 4063
rect 19475 4060 19487 4063
rect 19702 4060 19708 4072
rect 19475 4032 19708 4060
rect 19475 4029 19487 4032
rect 19429 4023 19487 4029
rect 19702 4020 19708 4032
rect 19760 4020 19766 4072
rect 20346 4060 20352 4072
rect 20307 4032 20352 4060
rect 20346 4020 20352 4032
rect 20404 4020 20410 4072
rect 22094 4060 22100 4072
rect 22055 4032 22100 4060
rect 22094 4020 22100 4032
rect 22152 4020 22158 4072
rect 22278 4020 22284 4072
rect 22336 4060 22342 4072
rect 25459 4069 25487 4100
rect 25958 4088 25964 4100
rect 26016 4088 26022 4140
rect 25444 4063 25502 4069
rect 22336 4032 23520 4060
rect 22336 4020 22342 4032
rect 18506 3992 18512 4004
rect 12452 3964 16620 3992
rect 16684 3964 18512 3992
rect 9582 3924 9588 3936
rect 9416 3896 9588 3924
rect 8481 3887 8539 3893
rect 9582 3884 9588 3896
rect 9640 3924 9646 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 9640 3896 10241 3924
rect 9640 3884 9646 3896
rect 10229 3893 10241 3896
rect 10275 3924 10287 3927
rect 10594 3924 10600 3936
rect 10275 3896 10600 3924
rect 10275 3893 10287 3896
rect 10229 3887 10287 3893
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11790 3924 11796 3936
rect 11751 3896 11796 3924
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3924 14519 3927
rect 14642 3924 14648 3936
rect 14507 3896 14648 3924
rect 14507 3893 14519 3896
rect 14461 3887 14519 3893
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 15194 3924 15200 3936
rect 15155 3896 15200 3924
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 16592 3924 16620 3964
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 20257 3995 20315 4001
rect 20257 3961 20269 3995
rect 20303 3992 20315 3995
rect 20711 3995 20769 4001
rect 20711 3992 20723 3995
rect 20303 3964 20723 3992
rect 20303 3961 20315 3964
rect 20257 3955 20315 3961
rect 20711 3961 20723 3964
rect 20757 3992 20769 3995
rect 22296 3992 22324 4020
rect 20757 3964 22324 3992
rect 22649 3995 22707 4001
rect 20757 3961 20769 3964
rect 20711 3955 20769 3961
rect 22649 3961 22661 3995
rect 22695 3992 22707 3995
rect 22738 3992 22744 4004
rect 22695 3964 22744 3992
rect 22695 3961 22707 3964
rect 22649 3955 22707 3961
rect 22738 3952 22744 3964
rect 22796 3992 22802 4004
rect 23198 3992 23204 4004
rect 22796 3964 23204 3992
rect 22796 3952 22802 3964
rect 23198 3952 23204 3964
rect 23256 3952 23262 4004
rect 23492 4001 23520 4032
rect 25444 4029 25456 4063
rect 25490 4029 25502 4063
rect 25444 4023 25502 4029
rect 25547 4063 25605 4069
rect 25547 4029 25559 4063
rect 25593 4060 25605 4063
rect 25866 4060 25872 4072
rect 25593 4032 25872 4060
rect 25593 4029 25605 4032
rect 25547 4023 25605 4029
rect 25866 4020 25872 4032
rect 25924 4020 25930 4072
rect 26418 4020 26424 4072
rect 26476 4060 26482 4072
rect 26513 4063 26571 4069
rect 26513 4060 26525 4063
rect 26476 4032 26525 4060
rect 26476 4020 26482 4032
rect 26513 4029 26525 4032
rect 26559 4029 26571 4063
rect 26513 4023 26571 4029
rect 27433 4063 27491 4069
rect 27433 4029 27445 4063
rect 27479 4060 27491 4063
rect 27479 4032 28488 4060
rect 27479 4029 27491 4032
rect 27433 4023 27491 4029
rect 23477 3995 23535 4001
rect 23477 3961 23489 3995
rect 23523 3992 23535 3995
rect 24023 3995 24081 4001
rect 24023 3992 24035 3995
rect 23523 3964 24035 3992
rect 23523 3961 23535 3964
rect 23477 3955 23535 3961
rect 24023 3961 24035 3964
rect 24069 3961 24081 3995
rect 24023 3955 24081 3961
rect 17402 3924 17408 3936
rect 16592 3896 17408 3924
rect 17402 3884 17408 3896
rect 17460 3924 17466 3936
rect 17681 3927 17739 3933
rect 17681 3924 17693 3927
rect 17460 3896 17693 3924
rect 17460 3884 17466 3896
rect 17681 3893 17693 3896
rect 17727 3924 17739 3927
rect 17773 3927 17831 3933
rect 17773 3924 17785 3927
rect 17727 3896 17785 3924
rect 17727 3893 17739 3896
rect 17681 3887 17739 3893
rect 17773 3893 17785 3896
rect 17819 3893 17831 3927
rect 17773 3887 17831 3893
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 18141 3927 18199 3933
rect 18141 3924 18153 3927
rect 17920 3896 18153 3924
rect 17920 3884 17926 3896
rect 18141 3893 18153 3896
rect 18187 3893 18199 3927
rect 18141 3887 18199 3893
rect 18230 3884 18236 3936
rect 18288 3924 18294 3936
rect 19610 3924 19616 3936
rect 18288 3896 19616 3924
rect 18288 3884 18294 3896
rect 19610 3884 19616 3896
rect 19668 3884 19674 3936
rect 21634 3924 21640 3936
rect 21595 3896 21640 3924
rect 21634 3884 21640 3896
rect 21692 3884 21698 3936
rect 22278 3924 22284 3936
rect 22239 3896 22284 3924
rect 22278 3884 22284 3896
rect 22336 3884 22342 3936
rect 23014 3924 23020 3936
rect 22975 3896 23020 3924
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 24038 3924 24066 3955
rect 24762 3952 24768 4004
rect 24820 3992 24826 4004
rect 25225 3995 25283 4001
rect 25225 3992 25237 3995
rect 24820 3964 25237 3992
rect 24820 3952 24826 3964
rect 25225 3961 25237 3964
rect 25271 3961 25283 3995
rect 26875 3995 26933 4001
rect 26875 3992 26887 3995
rect 25225 3955 25283 3961
rect 25332 3964 26887 3992
rect 24946 3924 24952 3936
rect 24038 3896 24952 3924
rect 24946 3884 24952 3896
rect 25004 3924 25010 3936
rect 25332 3924 25360 3964
rect 26875 3961 26887 3964
rect 26921 3992 26933 3995
rect 27246 3992 27252 4004
rect 26921 3964 27252 3992
rect 26921 3961 26933 3964
rect 26875 3955 26933 3961
rect 27246 3952 27252 3964
rect 27304 3952 27310 4004
rect 27706 3952 27712 4004
rect 27764 3952 27770 4004
rect 25958 3924 25964 3936
rect 25004 3896 25360 3924
rect 25919 3896 25964 3924
rect 25004 3884 25010 3896
rect 25958 3884 25964 3896
rect 26016 3884 26022 3936
rect 27724 3924 27752 3952
rect 27801 3927 27859 3933
rect 27801 3924 27813 3927
rect 27724 3896 27813 3924
rect 27801 3893 27813 3896
rect 27847 3924 27859 3927
rect 27982 3924 27988 3936
rect 27847 3896 27988 3924
rect 27847 3893 27859 3896
rect 27801 3887 27859 3893
rect 27982 3884 27988 3896
rect 28040 3884 28046 3936
rect 28460 3924 28488 4032
rect 29178 4020 29184 4072
rect 29236 4060 29242 4072
rect 29324 4063 29382 4069
rect 29324 4060 29336 4063
rect 29236 4032 29336 4060
rect 29236 4020 29242 4032
rect 29324 4029 29336 4032
rect 29370 4060 29382 4063
rect 29822 4060 29828 4072
rect 29370 4032 29828 4060
rect 29370 4029 29382 4032
rect 29324 4023 29382 4029
rect 29822 4020 29828 4032
rect 29880 4020 29886 4072
rect 31386 4060 31392 4072
rect 31347 4032 31392 4060
rect 31386 4020 31392 4032
rect 31444 4020 31450 4072
rect 29411 3995 29469 4001
rect 29411 3961 29423 3995
rect 29457 3992 29469 3995
rect 30374 3992 30380 4004
rect 29457 3964 30380 3992
rect 29457 3961 29469 3964
rect 29411 3955 29469 3961
rect 30374 3952 30380 3964
rect 30432 3952 30438 4004
rect 30469 3995 30527 4001
rect 30469 3961 30481 3995
rect 30515 3961 30527 3995
rect 31018 3992 31024 4004
rect 30979 3964 31024 3992
rect 30469 3955 30527 3961
rect 30101 3927 30159 3933
rect 30101 3924 30113 3927
rect 28460 3896 30113 3924
rect 30101 3893 30113 3896
rect 30147 3924 30159 3927
rect 30484 3924 30512 3955
rect 31018 3952 31024 3964
rect 31076 3952 31082 4004
rect 32214 3924 32220 3936
rect 30147 3896 32220 3924
rect 30147 3893 30159 3896
rect 30101 3887 30159 3893
rect 32214 3884 32220 3896
rect 32272 3884 32278 3936
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 2639 3723 2697 3729
rect 2639 3689 2651 3723
rect 2685 3720 2697 3723
rect 3786 3720 3792 3732
rect 2685 3692 3792 3720
rect 2685 3689 2697 3692
rect 2639 3683 2697 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 4801 3723 4859 3729
rect 4801 3689 4813 3723
rect 4847 3720 4859 3723
rect 4982 3720 4988 3732
rect 4847 3692 4988 3720
rect 4847 3689 4859 3692
rect 4801 3683 4859 3689
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 6638 3720 6644 3732
rect 5132 3692 5177 3720
rect 6599 3692 6644 3720
rect 5132 3680 5138 3692
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 9125 3723 9183 3729
rect 9125 3689 9137 3723
rect 9171 3720 9183 3723
rect 9582 3720 9588 3732
rect 9171 3692 9588 3720
rect 9171 3689 9183 3692
rect 9125 3683 9183 3689
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 9858 3720 9864 3732
rect 9819 3692 9864 3720
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 12529 3723 12587 3729
rect 12529 3720 12541 3723
rect 10652 3692 12541 3720
rect 10652 3680 10658 3692
rect 12529 3689 12541 3692
rect 12575 3720 12587 3723
rect 12986 3720 12992 3732
rect 12575 3692 12992 3720
rect 12575 3689 12587 3692
rect 12529 3683 12587 3689
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 13265 3723 13323 3729
rect 13265 3689 13277 3723
rect 13311 3720 13323 3723
rect 13722 3720 13728 3732
rect 13311 3692 13728 3720
rect 13311 3689 13323 3692
rect 13265 3683 13323 3689
rect 2133 3655 2191 3661
rect 2133 3621 2145 3655
rect 2179 3652 2191 3655
rect 2961 3655 3019 3661
rect 2961 3652 2973 3655
rect 2179 3624 2973 3652
rect 2179 3621 2191 3624
rect 2133 3615 2191 3621
rect 2961 3621 2973 3624
rect 3007 3652 3019 3655
rect 3234 3652 3240 3664
rect 3007 3624 3240 3652
rect 3007 3621 3019 3624
rect 2961 3615 3019 3621
rect 3234 3612 3240 3624
rect 3292 3612 3298 3664
rect 8478 3612 8484 3664
rect 8536 3652 8542 3664
rect 12897 3655 12955 3661
rect 8536 3624 11928 3652
rect 8536 3612 8542 3624
rect 106 3544 112 3596
rect 164 3584 170 3596
rect 2501 3587 2559 3593
rect 2501 3584 2513 3587
rect 164 3556 2513 3584
rect 164 3544 170 3556
rect 2501 3553 2513 3556
rect 2547 3584 2559 3587
rect 2590 3584 2596 3596
rect 2547 3556 2596 3584
rect 2547 3553 2559 3556
rect 2501 3547 2559 3553
rect 2590 3544 2596 3556
rect 2648 3544 2654 3596
rect 3421 3587 3479 3593
rect 3421 3553 3433 3587
rect 3467 3584 3479 3587
rect 3510 3584 3516 3596
rect 3467 3556 3516 3584
rect 3467 3553 3479 3556
rect 3421 3547 3479 3553
rect 3510 3544 3516 3556
rect 3568 3544 3574 3596
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 5224 3556 5273 3584
rect 5224 3544 5230 3556
rect 5261 3553 5273 3556
rect 5307 3553 5319 3587
rect 5718 3584 5724 3596
rect 5631 3556 5724 3584
rect 5261 3547 5319 3553
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 6086 3584 6092 3596
rect 6047 3556 6092 3584
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 8662 3584 8668 3596
rect 8623 3556 8668 3584
rect 8662 3544 8668 3556
rect 8720 3584 8726 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 8720 3556 9689 3584
rect 8720 3544 8726 3556
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 10134 3584 10140 3596
rect 10095 3556 10140 3584
rect 9677 3547 9735 3553
rect 10134 3544 10140 3556
rect 10192 3584 10198 3596
rect 10410 3584 10416 3596
rect 10192 3556 10416 3584
rect 10192 3544 10198 3556
rect 10410 3544 10416 3556
rect 10468 3544 10474 3596
rect 11790 3584 11796 3596
rect 11751 3556 11796 3584
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 4614 3476 4620 3528
rect 4672 3516 4678 3528
rect 5736 3516 5764 3544
rect 4672 3488 5764 3516
rect 6104 3516 6132 3544
rect 11900 3528 11928 3624
rect 12897 3621 12909 3655
rect 12943 3652 12955 3655
rect 13280 3652 13308 3683
rect 13722 3680 13728 3692
rect 13780 3720 13786 3732
rect 15654 3720 15660 3732
rect 13780 3692 15660 3720
rect 13780 3680 13786 3692
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 16301 3723 16359 3729
rect 16301 3720 16313 3723
rect 16264 3692 16313 3720
rect 16264 3680 16270 3692
rect 16301 3689 16313 3692
rect 16347 3689 16359 3723
rect 16301 3683 16359 3689
rect 16390 3680 16396 3732
rect 16448 3720 16454 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 16448 3692 16681 3720
rect 16448 3680 16454 3692
rect 16669 3689 16681 3692
rect 16715 3689 16727 3723
rect 17402 3720 17408 3732
rect 17363 3692 17408 3720
rect 16669 3683 16727 3689
rect 17402 3680 17408 3692
rect 17460 3680 17466 3732
rect 18782 3680 18788 3732
rect 18840 3720 18846 3732
rect 19245 3723 19303 3729
rect 19245 3720 19257 3723
rect 18840 3692 19257 3720
rect 18840 3680 18846 3692
rect 19245 3689 19257 3692
rect 19291 3689 19303 3723
rect 19245 3683 19303 3689
rect 19429 3723 19487 3729
rect 19429 3689 19441 3723
rect 19475 3720 19487 3723
rect 22738 3720 22744 3732
rect 19475 3692 22744 3720
rect 19475 3689 19487 3692
rect 19429 3683 19487 3689
rect 22738 3680 22744 3692
rect 22796 3680 22802 3732
rect 25866 3720 25872 3732
rect 24964 3692 25872 3720
rect 16025 3655 16083 3661
rect 12943 3624 13308 3652
rect 14292 3624 15424 3652
rect 12943 3621 12955 3624
rect 12897 3615 12955 3621
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 14292 3593 14320 3624
rect 14277 3587 14335 3593
rect 14277 3584 14289 3587
rect 13780 3556 14289 3584
rect 13780 3544 13786 3556
rect 14277 3553 14289 3556
rect 14323 3553 14335 3587
rect 14277 3547 14335 3553
rect 15105 3587 15163 3593
rect 15105 3553 15117 3587
rect 15151 3584 15163 3587
rect 15286 3584 15292 3596
rect 15151 3556 15292 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 15396 3584 15424 3624
rect 16025 3621 16037 3655
rect 16071 3652 16083 3655
rect 16758 3652 16764 3664
rect 16071 3624 16764 3652
rect 16071 3621 16083 3624
rect 16025 3615 16083 3621
rect 16758 3612 16764 3624
rect 16816 3612 16822 3664
rect 17420 3584 17448 3680
rect 18969 3655 19027 3661
rect 18969 3621 18981 3655
rect 19015 3652 19027 3655
rect 20346 3652 20352 3664
rect 19015 3624 20352 3652
rect 19015 3621 19027 3624
rect 18969 3615 19027 3621
rect 20346 3612 20352 3624
rect 20404 3612 20410 3664
rect 21085 3655 21143 3661
rect 21085 3621 21097 3655
rect 21131 3652 21143 3655
rect 21266 3652 21272 3664
rect 21131 3624 21272 3652
rect 21131 3621 21143 3624
rect 21085 3615 21143 3621
rect 21266 3612 21272 3624
rect 21324 3612 21330 3664
rect 21450 3612 21456 3664
rect 21508 3652 21514 3664
rect 21637 3655 21695 3661
rect 21637 3652 21649 3655
rect 21508 3624 21649 3652
rect 21508 3612 21514 3624
rect 21637 3621 21649 3624
rect 21683 3652 21695 3655
rect 22186 3652 22192 3664
rect 21683 3624 22192 3652
rect 21683 3621 21695 3624
rect 21637 3615 21695 3621
rect 22186 3612 22192 3624
rect 22244 3612 22250 3664
rect 23937 3655 23995 3661
rect 23937 3621 23949 3655
rect 23983 3652 23995 3655
rect 24762 3652 24768 3664
rect 23983 3624 24768 3652
rect 23983 3621 23995 3624
rect 23937 3615 23995 3621
rect 24762 3612 24768 3624
rect 24820 3612 24826 3664
rect 24964 3661 24992 3692
rect 25866 3680 25872 3692
rect 25924 3680 25930 3732
rect 27430 3720 27436 3732
rect 27391 3692 27436 3720
rect 27430 3680 27436 3692
rect 27488 3680 27494 3732
rect 28169 3723 28227 3729
rect 28169 3689 28181 3723
rect 28215 3720 28227 3723
rect 28258 3720 28264 3732
rect 28215 3692 28264 3720
rect 28215 3689 28227 3692
rect 28169 3683 28227 3689
rect 28258 3680 28264 3692
rect 28316 3720 28322 3732
rect 30374 3720 30380 3732
rect 28316 3692 28396 3720
rect 30335 3692 30380 3720
rect 28316 3680 28322 3692
rect 24949 3655 25007 3661
rect 24949 3621 24961 3655
rect 24995 3621 25007 3655
rect 24949 3615 25007 3621
rect 25041 3655 25099 3661
rect 25041 3621 25053 3655
rect 25087 3652 25099 3655
rect 25406 3652 25412 3664
rect 25087 3624 25412 3652
rect 25087 3621 25099 3624
rect 25041 3615 25099 3621
rect 25406 3612 25412 3624
rect 25464 3652 25470 3664
rect 26510 3652 26516 3664
rect 25464 3624 26516 3652
rect 25464 3612 25470 3624
rect 26510 3612 26516 3624
rect 26568 3612 26574 3664
rect 26875 3655 26933 3661
rect 26875 3621 26887 3655
rect 26921 3652 26933 3655
rect 27246 3652 27252 3664
rect 26921 3624 27252 3652
rect 26921 3621 26933 3624
rect 26875 3615 26933 3621
rect 27246 3612 27252 3624
rect 27304 3612 27310 3664
rect 28368 3661 28396 3692
rect 30374 3680 30380 3692
rect 30432 3680 30438 3732
rect 28353 3655 28411 3661
rect 28353 3621 28365 3655
rect 28399 3621 28411 3655
rect 28353 3615 28411 3621
rect 28442 3612 28448 3664
rect 28500 3652 28506 3664
rect 30009 3655 30067 3661
rect 28500 3624 28545 3652
rect 28500 3612 28506 3624
rect 30009 3621 30021 3655
rect 30055 3652 30067 3655
rect 30558 3652 30564 3664
rect 30055 3624 30564 3652
rect 30055 3621 30067 3624
rect 30009 3615 30067 3621
rect 30558 3612 30564 3624
rect 30616 3612 30622 3664
rect 30650 3612 30656 3664
rect 30708 3652 30714 3664
rect 32125 3655 32183 3661
rect 32125 3652 32137 3655
rect 30708 3624 32137 3652
rect 30708 3612 30714 3624
rect 32125 3621 32137 3624
rect 32171 3621 32183 3655
rect 32125 3615 32183 3621
rect 17497 3587 17555 3593
rect 17497 3584 17509 3587
rect 15396 3556 16436 3584
rect 17420 3556 17509 3584
rect 7837 3519 7895 3525
rect 7837 3516 7849 3519
rect 6104 3488 7849 3516
rect 4672 3476 4678 3488
rect 7837 3485 7849 3488
rect 7883 3516 7895 3519
rect 8570 3516 8576 3528
rect 7883 3488 8576 3516
rect 7883 3485 7895 3488
rect 7837 3479 7895 3485
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3516 8815 3519
rect 9766 3516 9772 3528
rect 8803 3488 9772 3516
rect 8803 3485 8815 3488
rect 8757 3479 8815 3485
rect 1765 3451 1823 3457
rect 1765 3417 1777 3451
rect 1811 3448 1823 3451
rect 1946 3448 1952 3460
rect 1811 3420 1952 3448
rect 1811 3417 1823 3420
rect 1765 3411 1823 3417
rect 1946 3408 1952 3420
rect 2004 3408 2010 3460
rect 2958 3408 2964 3460
rect 3016 3448 3022 3460
rect 8772 3448 8800 3479
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 11882 3516 11888 3528
rect 11843 3488 11888 3516
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 14642 3516 14648 3528
rect 14415 3488 14648 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 14642 3476 14648 3488
rect 14700 3516 14706 3528
rect 15657 3519 15715 3525
rect 15657 3516 15669 3519
rect 14700 3488 15669 3516
rect 14700 3476 14706 3488
rect 15657 3485 15669 3488
rect 15703 3516 15715 3519
rect 16298 3516 16304 3528
rect 15703 3488 16304 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 3016 3420 8800 3448
rect 11057 3451 11115 3457
rect 3016 3408 3022 3420
rect 11057 3417 11069 3451
rect 11103 3448 11115 3451
rect 11146 3448 11152 3460
rect 11103 3420 11152 3448
rect 11103 3417 11115 3420
rect 11057 3411 11115 3417
rect 11146 3408 11152 3420
rect 11204 3448 11210 3460
rect 15194 3448 15200 3460
rect 11204 3420 15200 3448
rect 11204 3408 11210 3420
rect 15194 3408 15200 3420
rect 15252 3448 15258 3460
rect 15454 3451 15512 3457
rect 15454 3448 15466 3451
rect 15252 3420 15466 3448
rect 15252 3408 15258 3420
rect 15454 3417 15466 3420
rect 15500 3448 15512 3451
rect 15930 3448 15936 3460
rect 15500 3420 15936 3448
rect 15500 3417 15512 3420
rect 15454 3411 15512 3417
rect 15930 3408 15936 3420
rect 15988 3408 15994 3460
rect 16408 3448 16436 3556
rect 17497 3553 17509 3556
rect 17543 3553 17555 3587
rect 17954 3584 17960 3596
rect 17915 3556 17960 3584
rect 17497 3547 17555 3553
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 18506 3584 18512 3596
rect 18467 3556 18512 3584
rect 18506 3544 18512 3556
rect 18564 3544 18570 3596
rect 18874 3584 18880 3596
rect 18787 3556 18880 3584
rect 18874 3544 18880 3556
rect 18932 3584 18938 3596
rect 19702 3584 19708 3596
rect 18932 3556 19708 3584
rect 18932 3544 18938 3556
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 22002 3584 22008 3596
rect 21963 3556 22008 3584
rect 22002 3544 22008 3556
rect 22060 3584 22066 3596
rect 22465 3587 22523 3593
rect 22465 3584 22477 3587
rect 22060 3556 22477 3584
rect 22060 3544 22066 3556
rect 22465 3553 22477 3556
rect 22511 3553 22523 3587
rect 23198 3584 23204 3596
rect 23159 3556 23204 3584
rect 22465 3547 22523 3553
rect 23198 3544 23204 3556
rect 23256 3544 23262 3596
rect 23293 3587 23351 3593
rect 23293 3553 23305 3587
rect 23339 3553 23351 3587
rect 23293 3547 23351 3553
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 19797 3519 19855 3525
rect 19797 3516 19809 3519
rect 16816 3488 19809 3516
rect 16816 3476 16822 3488
rect 19797 3485 19809 3488
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 20993 3519 21051 3525
rect 20993 3485 21005 3519
rect 21039 3516 21051 3519
rect 21358 3516 21364 3528
rect 21039 3488 21364 3516
rect 21039 3485 21051 3488
rect 20993 3479 21051 3485
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 22278 3476 22284 3528
rect 22336 3516 22342 3528
rect 23106 3516 23112 3528
rect 22336 3488 23112 3516
rect 22336 3476 22342 3488
rect 23106 3476 23112 3488
rect 23164 3516 23170 3528
rect 23308 3516 23336 3547
rect 23382 3544 23388 3596
rect 23440 3584 23446 3596
rect 23661 3587 23719 3593
rect 23661 3584 23673 3587
rect 23440 3556 23673 3584
rect 23440 3544 23446 3556
rect 23661 3553 23673 3556
rect 23707 3584 23719 3587
rect 24670 3584 24676 3596
rect 23707 3556 24676 3584
rect 23707 3553 23719 3556
rect 23661 3547 23719 3553
rect 24670 3544 24676 3556
rect 24728 3544 24734 3596
rect 32214 3584 32220 3596
rect 32175 3556 32220 3584
rect 32214 3544 32220 3556
rect 32272 3544 32278 3596
rect 24486 3516 24492 3528
rect 23164 3488 24492 3516
rect 23164 3476 23170 3488
rect 24486 3476 24492 3488
rect 24544 3516 24550 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 24544 3488 24593 3516
rect 24544 3476 24550 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 25222 3516 25228 3528
rect 25183 3488 25228 3516
rect 24581 3479 24639 3485
rect 25222 3476 25228 3488
rect 25280 3476 25286 3528
rect 26510 3516 26516 3528
rect 26471 3488 26516 3516
rect 26510 3476 26516 3488
rect 26568 3476 26574 3528
rect 31018 3516 31024 3528
rect 30979 3488 31024 3516
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 18230 3448 18236 3460
rect 16408 3420 18236 3448
rect 18230 3408 18236 3420
rect 18288 3408 18294 3460
rect 20349 3451 20407 3457
rect 20349 3417 20361 3451
rect 20395 3448 20407 3451
rect 28905 3451 28963 3457
rect 20395 3420 20944 3448
rect 20395 3417 20407 3420
rect 20349 3411 20407 3417
rect 14737 3383 14795 3389
rect 14737 3349 14749 3383
rect 14783 3380 14795 3383
rect 14918 3380 14924 3392
rect 14783 3352 14924 3380
rect 14783 3349 14795 3352
rect 14737 3343 14795 3349
rect 14918 3340 14924 3352
rect 14976 3380 14982 3392
rect 15562 3380 15568 3392
rect 14976 3352 15568 3380
rect 14976 3340 14982 3352
rect 15562 3340 15568 3352
rect 15620 3380 15626 3392
rect 19429 3383 19487 3389
rect 19429 3380 19441 3383
rect 15620 3352 19441 3380
rect 15620 3340 15626 3352
rect 19429 3349 19441 3352
rect 19475 3349 19487 3383
rect 19702 3380 19708 3392
rect 19663 3352 19708 3380
rect 19429 3343 19487 3349
rect 19702 3340 19708 3352
rect 19760 3340 19766 3392
rect 20622 3380 20628 3392
rect 20583 3352 20628 3380
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 20916 3380 20944 3420
rect 28905 3417 28917 3451
rect 28951 3448 28963 3451
rect 28951 3420 29316 3448
rect 28951 3417 28963 3420
rect 28905 3411 28963 3417
rect 29288 3392 29316 3420
rect 21726 3380 21732 3392
rect 20916 3352 21732 3380
rect 21726 3340 21732 3352
rect 21784 3340 21790 3392
rect 22186 3340 22192 3392
rect 22244 3380 22250 3392
rect 22281 3383 22339 3389
rect 22281 3380 22293 3383
rect 22244 3352 22293 3380
rect 22244 3340 22250 3352
rect 22281 3349 22293 3352
rect 22327 3349 22339 3383
rect 22281 3343 22339 3349
rect 23658 3340 23664 3392
rect 23716 3380 23722 3392
rect 24213 3383 24271 3389
rect 24213 3380 24225 3383
rect 23716 3352 24225 3380
rect 23716 3340 23722 3352
rect 24213 3349 24225 3352
rect 24259 3349 24271 3383
rect 26234 3380 26240 3392
rect 26195 3352 26240 3380
rect 24213 3343 24271 3349
rect 26234 3340 26240 3352
rect 26292 3340 26298 3392
rect 29270 3380 29276 3392
rect 29231 3352 29276 3380
rect 29270 3340 29276 3352
rect 29328 3340 29334 3392
rect 32490 3340 32496 3392
rect 32548 3380 32554 3392
rect 33137 3383 33195 3389
rect 33137 3380 33149 3383
rect 32548 3352 33149 3380
rect 32548 3340 32554 3352
rect 33137 3349 33149 3352
rect 33183 3349 33195 3383
rect 33137 3343 33195 3349
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 4801 3179 4859 3185
rect 4801 3176 4813 3179
rect 4672 3148 4813 3176
rect 4672 3136 4678 3148
rect 4801 3145 4813 3148
rect 4847 3145 4859 3179
rect 4801 3139 4859 3145
rect 5169 3179 5227 3185
rect 5169 3145 5181 3179
rect 5215 3176 5227 3179
rect 6178 3176 6184 3188
rect 5215 3148 6184 3176
rect 5215 3145 5227 3148
rect 5169 3139 5227 3145
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 7193 3179 7251 3185
rect 7193 3176 7205 3179
rect 6512 3148 7205 3176
rect 6512 3136 6518 3148
rect 7193 3145 7205 3148
rect 7239 3145 7251 3179
rect 7193 3139 7251 3145
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 17129 3179 17187 3185
rect 17129 3176 17141 3179
rect 11940 3148 17141 3176
rect 11940 3136 11946 3148
rect 17129 3145 17141 3148
rect 17175 3176 17187 3179
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 17175 3148 17509 3176
rect 17175 3145 17187 3148
rect 17129 3139 17187 3145
rect 17497 3145 17509 3148
rect 17543 3176 17555 3179
rect 17954 3176 17960 3188
rect 17543 3148 17960 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 17954 3136 17960 3148
rect 18012 3136 18018 3188
rect 19702 3136 19708 3188
rect 19760 3176 19766 3188
rect 20257 3179 20315 3185
rect 20257 3176 20269 3179
rect 19760 3148 20269 3176
rect 19760 3136 19766 3148
rect 20257 3145 20269 3148
rect 20303 3176 20315 3179
rect 20533 3179 20591 3185
rect 20533 3176 20545 3179
rect 20303 3148 20545 3176
rect 20303 3145 20315 3148
rect 20257 3139 20315 3145
rect 20533 3145 20545 3148
rect 20579 3145 20591 3179
rect 20533 3139 20591 3145
rect 21726 3136 21732 3188
rect 21784 3176 21790 3188
rect 23934 3176 23940 3188
rect 21784 3148 23940 3176
rect 21784 3136 21790 3148
rect 23934 3136 23940 3148
rect 23992 3136 23998 3188
rect 25406 3176 25412 3188
rect 25367 3148 25412 3176
rect 25406 3136 25412 3148
rect 25464 3136 25470 3188
rect 27157 3179 27215 3185
rect 27157 3145 27169 3179
rect 27203 3176 27215 3179
rect 28442 3176 28448 3188
rect 27203 3148 28448 3176
rect 27203 3145 27215 3148
rect 27157 3139 27215 3145
rect 28442 3136 28448 3148
rect 28500 3176 28506 3188
rect 28537 3179 28595 3185
rect 28537 3176 28549 3179
rect 28500 3148 28549 3176
rect 28500 3136 28506 3148
rect 28537 3145 28549 3148
rect 28583 3145 28595 3179
rect 28537 3139 28595 3145
rect 30561 3179 30619 3185
rect 30561 3145 30573 3179
rect 30607 3176 30619 3179
rect 30650 3176 30656 3188
rect 30607 3148 30656 3176
rect 30607 3145 30619 3148
rect 30561 3139 30619 3145
rect 30650 3136 30656 3148
rect 30708 3136 30714 3188
rect 32214 3176 32220 3188
rect 32175 3148 32220 3176
rect 32214 3136 32220 3148
rect 32272 3136 32278 3188
rect 3510 3108 3516 3120
rect 3344 3080 3516 3108
rect 1765 2975 1823 2981
rect 1765 2941 1777 2975
rect 1811 2972 1823 2975
rect 1854 2972 1860 2984
rect 1811 2944 1860 2972
rect 1811 2941 1823 2944
rect 1765 2935 1823 2941
rect 1854 2932 1860 2944
rect 1912 2972 1918 2984
rect 2958 2972 2964 2984
rect 1912 2944 2964 2972
rect 1912 2932 1918 2944
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3344 2981 3372 3080
rect 3510 3068 3516 3080
rect 3568 3068 3574 3120
rect 8018 3068 8024 3120
rect 8076 3108 8082 3120
rect 13722 3108 13728 3120
rect 8076 3080 8524 3108
rect 8076 3068 8082 3080
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4212 3012 4257 3040
rect 4212 3000 4218 3012
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 5224 3012 5825 3040
rect 5224 3000 5230 3012
rect 5813 3009 5825 3012
rect 5859 3040 5871 3043
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 5859 3012 7481 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 7469 3009 7481 3012
rect 7515 3040 7527 3043
rect 7834 3040 7840 3052
rect 7515 3012 7840 3040
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 7834 3000 7840 3012
rect 7892 3040 7898 3052
rect 8202 3040 8208 3052
rect 7892 3012 8208 3040
rect 7892 3000 7898 3012
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 3418 2932 3424 2984
rect 3476 2972 3482 2984
rect 3513 2975 3571 2981
rect 3513 2972 3525 2975
rect 3476 2944 3525 2972
rect 3476 2932 3482 2944
rect 3513 2941 3525 2944
rect 3559 2941 3571 2975
rect 4062 2972 4068 2984
rect 4023 2944 4068 2972
rect 3513 2935 3571 2941
rect 4062 2932 4068 2944
rect 4120 2972 4126 2984
rect 4433 2975 4491 2981
rect 4433 2972 4445 2975
rect 4120 2944 4445 2972
rect 4120 2932 4126 2944
rect 4433 2941 4445 2944
rect 4479 2972 4491 2975
rect 4798 2972 4804 2984
rect 4479 2944 4804 2972
rect 4479 2941 4491 2944
rect 4433 2935 4491 2941
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 4985 2975 5043 2981
rect 4985 2941 4997 2975
rect 5031 2972 5043 2975
rect 6641 2975 6699 2981
rect 5031 2944 5488 2972
rect 5031 2941 5043 2944
rect 4985 2935 5043 2941
rect 1946 2864 1952 2916
rect 2004 2904 2010 2916
rect 2225 2907 2283 2913
rect 2225 2904 2237 2907
rect 2004 2876 2237 2904
rect 2004 2864 2010 2876
rect 2225 2873 2237 2876
rect 2271 2904 2283 2907
rect 4080 2904 4108 2932
rect 2271 2876 4108 2904
rect 2271 2873 2283 2876
rect 2225 2867 2283 2873
rect 5460 2848 5488 2944
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 7006 2972 7012 2984
rect 6687 2944 7012 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 7006 2932 7012 2944
rect 7064 2932 7070 2984
rect 8036 2981 8064 3012
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8496 2984 8524 3080
rect 8864 3080 9674 3108
rect 13683 3080 13728 3108
rect 8021 2975 8079 2981
rect 8021 2941 8033 2975
rect 8067 2941 8079 2975
rect 8478 2972 8484 2984
rect 8391 2944 8484 2972
rect 8021 2935 8079 2941
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8570 2932 8576 2984
rect 8628 2972 8634 2984
rect 8864 2981 8892 3080
rect 9646 3040 9674 3080
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 13906 3068 13912 3120
rect 13964 3108 13970 3120
rect 14645 3111 14703 3117
rect 14645 3108 14657 3111
rect 13964 3080 14657 3108
rect 13964 3068 13970 3080
rect 14645 3077 14657 3080
rect 14691 3108 14703 3111
rect 15286 3108 15292 3120
rect 14691 3080 15292 3108
rect 14691 3077 14703 3080
rect 14645 3071 14703 3077
rect 15286 3068 15292 3080
rect 15344 3068 15350 3120
rect 15473 3111 15531 3117
rect 15473 3077 15485 3111
rect 15519 3108 15531 3111
rect 15562 3108 15568 3120
rect 15519 3080 15568 3108
rect 15519 3077 15531 3080
rect 15473 3071 15531 3077
rect 15562 3068 15568 3080
rect 15620 3068 15626 3120
rect 10870 3040 10876 3052
rect 9646 3012 10876 3040
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 12434 3040 12440 3052
rect 12395 3012 12440 3040
rect 12434 3000 12440 3012
rect 12492 3000 12498 3052
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14277 3043 14335 3049
rect 14277 3040 14289 3043
rect 14056 3012 14289 3040
rect 14056 3000 14062 3012
rect 14277 3009 14289 3012
rect 14323 3040 14335 3043
rect 14737 3043 14795 3049
rect 14737 3040 14749 3043
rect 14323 3012 14749 3040
rect 14323 3009 14335 3012
rect 14277 3003 14335 3009
rect 14737 3009 14749 3012
rect 14783 3009 14795 3043
rect 15930 3040 15936 3052
rect 15891 3012 15936 3040
rect 14737 3003 14795 3009
rect 8849 2975 8907 2981
rect 8849 2972 8861 2975
rect 8628 2944 8861 2972
rect 8628 2932 8634 2944
rect 8849 2941 8861 2944
rect 8895 2941 8907 2975
rect 8849 2935 8907 2941
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9490 2972 9496 2984
rect 9263 2944 9496 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 7558 2864 7564 2916
rect 7616 2904 7622 2916
rect 9232 2904 9260 2935
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 11146 2972 11152 2984
rect 11107 2944 11152 2972
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 11790 2932 11796 2984
rect 11848 2972 11854 2984
rect 11885 2975 11943 2981
rect 11885 2972 11897 2975
rect 11848 2944 11897 2972
rect 11848 2932 11854 2944
rect 11885 2941 11897 2944
rect 11931 2972 11943 2975
rect 12342 2972 12348 2984
rect 11931 2944 12348 2972
rect 11931 2941 11943 2944
rect 11885 2935 11943 2941
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 12713 2975 12771 2981
rect 12713 2941 12725 2975
rect 12759 2941 12771 2975
rect 12713 2935 12771 2941
rect 14516 2975 14574 2981
rect 14516 2941 14528 2975
rect 14562 2972 14574 2975
rect 14642 2972 14648 2984
rect 14562 2944 14648 2972
rect 14562 2941 14574 2944
rect 14516 2935 14574 2941
rect 7616 2876 9260 2904
rect 10873 2907 10931 2913
rect 7616 2864 7622 2876
rect 10873 2873 10885 2907
rect 10919 2904 10931 2907
rect 10962 2904 10968 2916
rect 10919 2876 10968 2904
rect 10919 2873 10931 2876
rect 10873 2867 10931 2873
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 2590 2836 2596 2848
rect 2551 2808 2596 2836
rect 2590 2796 2596 2808
rect 2648 2796 2654 2848
rect 5442 2836 5448 2848
rect 5403 2808 5448 2836
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 7926 2836 7932 2848
rect 7887 2808 7932 2836
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 8110 2836 8116 2848
rect 8071 2808 8116 2836
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 8662 2796 8668 2848
rect 8720 2836 8726 2848
rect 9769 2839 9827 2845
rect 9769 2836 9781 2839
rect 8720 2808 9781 2836
rect 8720 2796 8726 2808
rect 9769 2805 9781 2808
rect 9815 2805 9827 2839
rect 9769 2799 9827 2805
rect 10410 2796 10416 2848
rect 10468 2836 10474 2848
rect 12161 2839 12219 2845
rect 12161 2836 12173 2839
rect 10468 2808 12173 2836
rect 10468 2796 10474 2808
rect 12161 2805 12173 2808
rect 12207 2836 12219 2839
rect 12728 2836 12756 2935
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 14752 2972 14780 3003
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 17972 3040 18000 3136
rect 19334 3068 19340 3120
rect 19392 3108 19398 3120
rect 21085 3111 21143 3117
rect 21085 3108 21097 3111
rect 19392 3080 21097 3108
rect 19392 3068 19398 3080
rect 21085 3077 21097 3080
rect 21131 3108 21143 3111
rect 22186 3108 22192 3120
rect 21131 3080 22192 3108
rect 21131 3077 21143 3080
rect 21085 3071 21143 3077
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 22649 3111 22707 3117
rect 22649 3077 22661 3111
rect 22695 3108 22707 3111
rect 26418 3108 26424 3120
rect 22695 3080 26424 3108
rect 22695 3077 22707 3080
rect 22649 3071 22707 3077
rect 26418 3068 26424 3080
rect 26476 3068 26482 3120
rect 27430 3068 27436 3120
rect 27488 3108 27494 3120
rect 28997 3111 29055 3117
rect 28997 3108 29009 3111
rect 27488 3080 29009 3108
rect 27488 3068 27494 3080
rect 28997 3077 29009 3080
rect 29043 3108 29055 3111
rect 29043 3080 29408 3108
rect 29043 3077 29055 3080
rect 28997 3071 29055 3077
rect 22002 3040 22008 3052
rect 17972 3012 18552 3040
rect 15841 2975 15899 2981
rect 15841 2972 15853 2975
rect 14752 2944 15853 2972
rect 15841 2941 15853 2944
rect 15887 2972 15899 2975
rect 16206 2972 16212 2984
rect 15887 2944 16212 2972
rect 15887 2941 15899 2944
rect 15841 2935 15899 2941
rect 16206 2932 16212 2944
rect 16264 2972 16270 2984
rect 16574 2972 16580 2984
rect 16264 2944 16580 2972
rect 16264 2932 16270 2944
rect 16574 2932 16580 2944
rect 16632 2932 16638 2984
rect 18046 2972 18052 2984
rect 18007 2944 18052 2972
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18524 2981 18552 3012
rect 21560 3012 22008 3040
rect 18509 2975 18567 2981
rect 18509 2941 18521 2975
rect 18555 2941 18567 2975
rect 19058 2972 19064 2984
rect 19019 2944 19064 2972
rect 18509 2935 18567 2941
rect 19058 2932 19064 2944
rect 19116 2932 19122 2984
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2972 19487 2975
rect 19702 2972 19708 2984
rect 19475 2944 19708 2972
rect 19475 2941 19487 2944
rect 19429 2935 19487 2941
rect 19702 2932 19708 2944
rect 19760 2932 19766 2984
rect 20990 2932 20996 2984
rect 21048 2972 21054 2984
rect 21560 2981 21588 3012
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 21545 2975 21603 2981
rect 21545 2972 21557 2975
rect 21048 2944 21557 2972
rect 21048 2932 21054 2944
rect 21545 2941 21557 2944
rect 21591 2941 21603 2975
rect 21726 2972 21732 2984
rect 21687 2944 21732 2972
rect 21545 2935 21603 2941
rect 21726 2932 21732 2944
rect 21784 2932 21790 2984
rect 21818 2932 21824 2984
rect 21876 2972 21882 2984
rect 22097 2975 22155 2981
rect 22097 2972 22109 2975
rect 21876 2944 22109 2972
rect 21876 2932 21882 2944
rect 22097 2941 22109 2944
rect 22143 2941 22155 2975
rect 22204 2972 22232 3068
rect 25133 3043 25191 3049
rect 25133 3009 25145 3043
rect 25179 3040 25191 3043
rect 26510 3040 26516 3052
rect 25179 3012 26516 3040
rect 25179 3009 25191 3012
rect 25133 3003 25191 3009
rect 26510 3000 26516 3012
rect 26568 3040 26574 3052
rect 27801 3043 27859 3049
rect 27801 3040 27813 3043
rect 26568 3012 27813 3040
rect 26568 3000 26574 3012
rect 27801 3009 27813 3012
rect 27847 3009 27859 3043
rect 27801 3003 27859 3009
rect 27982 3000 27988 3052
rect 28040 3040 28046 3052
rect 29273 3043 29331 3049
rect 29273 3040 29285 3043
rect 28040 3012 29285 3040
rect 28040 3000 28046 3012
rect 29273 3009 29285 3012
rect 29319 3009 29331 3043
rect 29273 3003 29331 3009
rect 22465 2975 22523 2981
rect 22465 2972 22477 2975
rect 22204 2944 22477 2972
rect 22097 2935 22155 2941
rect 22465 2941 22477 2944
rect 22511 2972 22523 2975
rect 23290 2972 23296 2984
rect 22511 2944 23296 2972
rect 22511 2941 22523 2944
rect 22465 2935 22523 2941
rect 14369 2907 14427 2913
rect 14369 2873 14381 2907
rect 14415 2904 14427 2907
rect 14918 2904 14924 2916
rect 14415 2876 14924 2904
rect 14415 2873 14427 2876
rect 14369 2867 14427 2873
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 15102 2904 15108 2916
rect 15063 2876 15108 2904
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 18064 2904 18092 2932
rect 19797 2907 19855 2913
rect 19797 2904 19809 2907
rect 18064 2876 19809 2904
rect 19797 2873 19809 2876
rect 19843 2873 19855 2907
rect 22112 2904 22140 2935
rect 23290 2932 23296 2944
rect 23348 2972 23354 2984
rect 23385 2975 23443 2981
rect 23385 2972 23397 2975
rect 23348 2944 23397 2972
rect 23348 2932 23354 2944
rect 23385 2941 23397 2944
rect 23431 2941 23443 2975
rect 23658 2972 23664 2984
rect 23619 2944 23664 2972
rect 23385 2935 23443 2941
rect 23658 2932 23664 2944
rect 23716 2932 23722 2984
rect 23934 2932 23940 2984
rect 23992 2972 23998 2984
rect 24118 2972 24124 2984
rect 23992 2944 24124 2972
rect 23992 2932 23998 2944
rect 24118 2932 24124 2944
rect 24176 2932 24182 2984
rect 24486 2972 24492 2984
rect 24447 2944 24492 2972
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 24670 2932 24676 2984
rect 24728 2972 24734 2984
rect 24857 2975 24915 2981
rect 24857 2972 24869 2975
rect 24728 2944 24869 2972
rect 24728 2932 24734 2944
rect 24857 2941 24869 2944
rect 24903 2941 24915 2975
rect 26234 2972 26240 2984
rect 26195 2944 26240 2972
rect 24857 2935 24915 2941
rect 26234 2932 26240 2944
rect 26292 2932 26298 2984
rect 29380 2981 29408 3080
rect 31573 3043 31631 3049
rect 31573 3009 31585 3043
rect 31619 3040 31631 3043
rect 32030 3040 32036 3052
rect 31619 3012 32036 3040
rect 31619 3009 31631 3012
rect 31573 3003 31631 3009
rect 32030 3000 32036 3012
rect 32088 3040 32094 3052
rect 32769 3043 32827 3049
rect 32769 3040 32781 3043
rect 32088 3012 32781 3040
rect 32088 3000 32094 3012
rect 32769 3009 32781 3012
rect 32815 3009 32827 3043
rect 32769 3003 32827 3009
rect 29365 2975 29423 2981
rect 29365 2941 29377 2975
rect 29411 2941 29423 2975
rect 29365 2935 29423 2941
rect 24946 2904 24952 2916
rect 22112 2876 24952 2904
rect 19797 2867 19855 2873
rect 24946 2864 24952 2876
rect 25004 2864 25010 2916
rect 26558 2907 26616 2913
rect 26558 2904 26570 2907
rect 26160 2876 26570 2904
rect 26160 2848 26188 2876
rect 26558 2873 26570 2876
rect 26604 2873 26616 2907
rect 30926 2904 30932 2916
rect 30887 2876 30932 2904
rect 26558 2867 26616 2873
rect 30926 2864 30932 2876
rect 30984 2864 30990 2916
rect 31021 2907 31079 2913
rect 31021 2873 31033 2907
rect 31067 2873 31079 2907
rect 31021 2867 31079 2873
rect 18322 2836 18328 2848
rect 12207 2808 12756 2836
rect 18235 2808 18328 2836
rect 12207 2805 12219 2808
rect 12161 2799 12219 2805
rect 18322 2796 18328 2808
rect 18380 2836 18386 2848
rect 18690 2836 18696 2848
rect 18380 2808 18696 2836
rect 18380 2796 18386 2808
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 23109 2839 23167 2845
rect 23109 2805 23121 2839
rect 23155 2836 23167 2839
rect 23198 2836 23204 2848
rect 23155 2808 23204 2836
rect 23155 2805 23167 2808
rect 23109 2799 23167 2805
rect 23198 2796 23204 2808
rect 23256 2836 23262 2848
rect 23382 2836 23388 2848
rect 23256 2808 23388 2836
rect 23256 2796 23262 2808
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 26142 2836 26148 2848
rect 26103 2808 26148 2836
rect 26142 2796 26148 2808
rect 26200 2796 26206 2848
rect 27430 2836 27436 2848
rect 27391 2808 27436 2836
rect 27430 2796 27436 2808
rect 27488 2796 27494 2848
rect 28074 2836 28080 2848
rect 28035 2808 28080 2836
rect 28074 2796 28080 2808
rect 28132 2796 28138 2848
rect 31036 2836 31064 2867
rect 31110 2864 31116 2916
rect 31168 2904 31174 2916
rect 32490 2904 32496 2916
rect 31168 2876 32496 2904
rect 31168 2864 31174 2876
rect 32490 2864 32496 2876
rect 32548 2864 32554 2916
rect 32585 2907 32643 2913
rect 32585 2873 32597 2907
rect 32631 2904 32643 2907
rect 32674 2904 32680 2916
rect 32631 2876 32680 2904
rect 32631 2873 32643 2876
rect 32585 2867 32643 2873
rect 32674 2864 32680 2876
rect 32732 2904 32738 2916
rect 33413 2907 33471 2913
rect 33413 2904 33425 2907
rect 32732 2876 33425 2904
rect 32732 2864 32738 2876
rect 33413 2873 33425 2876
rect 33459 2873 33471 2907
rect 33413 2867 33471 2873
rect 31202 2836 31208 2848
rect 31036 2808 31208 2836
rect 31202 2796 31208 2808
rect 31260 2796 31266 2848
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3053 2635 3111 2641
rect 3053 2632 3065 2635
rect 3016 2604 3065 2632
rect 3016 2592 3022 2604
rect 3053 2601 3065 2604
rect 3099 2601 3111 2635
rect 3510 2632 3516 2644
rect 3471 2604 3516 2632
rect 3053 2595 3111 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 6086 2632 6092 2644
rect 5276 2604 6092 2632
rect 2777 2567 2835 2573
rect 2777 2533 2789 2567
rect 2823 2564 2835 2567
rect 3418 2564 3424 2576
rect 2823 2536 3424 2564
rect 2823 2533 2835 2536
rect 2777 2527 2835 2533
rect 3418 2524 3424 2536
rect 3476 2564 3482 2576
rect 5276 2573 5304 2604
rect 6086 2592 6092 2604
rect 6144 2592 6150 2644
rect 7558 2632 7564 2644
rect 7519 2604 7564 2632
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 7834 2632 7840 2644
rect 7795 2604 7840 2632
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8478 2632 8484 2644
rect 8439 2604 8484 2632
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 8846 2632 8852 2644
rect 8807 2604 8852 2632
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 12802 2632 12808 2644
rect 12763 2604 12808 2632
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 13725 2635 13783 2641
rect 13725 2601 13737 2635
rect 13771 2632 13783 2635
rect 13998 2632 14004 2644
rect 13771 2604 14004 2632
rect 13771 2601 13783 2604
rect 13725 2595 13783 2601
rect 13979 2592 14004 2604
rect 14056 2592 14062 2644
rect 14918 2632 14924 2644
rect 14879 2604 14924 2632
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 15286 2632 15292 2644
rect 15247 2604 15292 2632
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 15654 2632 15660 2644
rect 15615 2604 15660 2632
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 17681 2635 17739 2641
rect 17681 2632 17693 2635
rect 16040 2604 17693 2632
rect 5261 2567 5319 2573
rect 5261 2564 5273 2567
rect 3476 2536 5273 2564
rect 3476 2524 3482 2536
rect 5261 2533 5273 2536
rect 5307 2533 5319 2567
rect 5261 2527 5319 2533
rect 5442 2524 5448 2576
rect 5500 2564 5506 2576
rect 5500 2536 8708 2564
rect 5500 2524 5506 2536
rect 1765 2499 1823 2505
rect 1765 2465 1777 2499
rect 1811 2496 1823 2499
rect 3510 2496 3516 2508
rect 1811 2468 3516 2496
rect 1811 2465 1823 2468
rect 1765 2459 1823 2465
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 7926 2496 7932 2508
rect 7699 2468 7932 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 7926 2456 7932 2468
rect 7984 2496 7990 2508
rect 8680 2505 8708 2536
rect 8665 2499 8723 2505
rect 7984 2468 8248 2496
rect 7984 2456 7990 2468
rect 8220 2369 8248 2468
rect 8665 2465 8677 2499
rect 8711 2496 8723 2499
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8711 2468 9137 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 9125 2465 9137 2468
rect 9171 2496 9183 2499
rect 10410 2496 10416 2508
rect 9171 2468 10416 2496
rect 9171 2465 9183 2468
rect 9125 2459 9183 2465
rect 10410 2456 10416 2468
rect 10468 2456 10474 2508
rect 10502 2456 10508 2508
rect 10560 2496 10566 2508
rect 10781 2499 10839 2505
rect 10781 2496 10793 2499
rect 10560 2468 10793 2496
rect 10560 2456 10566 2468
rect 10781 2465 10793 2468
rect 10827 2465 10839 2499
rect 12452 2496 12480 2592
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12452 2468 12633 2496
rect 10781 2459 10839 2465
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 13357 2499 13415 2505
rect 13357 2465 13369 2499
rect 13403 2496 13415 2499
rect 13722 2496 13728 2508
rect 13403 2468 13728 2496
rect 13403 2465 13415 2468
rect 13357 2459 13415 2465
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 13979 2505 14007 2592
rect 15304 2564 15332 2592
rect 15933 2567 15991 2573
rect 15933 2564 15945 2567
rect 15304 2536 15945 2564
rect 15933 2533 15945 2536
rect 15979 2533 15991 2567
rect 15933 2527 15991 2533
rect 13964 2499 14022 2505
rect 13872 2468 13917 2496
rect 13872 2456 13878 2468
rect 13964 2465 13976 2499
rect 14010 2465 14022 2499
rect 13964 2459 14022 2465
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15160 2468 15485 2496
rect 15160 2456 15166 2468
rect 15473 2465 15485 2468
rect 15519 2496 15531 2499
rect 16040 2496 16068 2604
rect 17681 2601 17693 2604
rect 17727 2601 17739 2635
rect 18138 2632 18144 2644
rect 18099 2604 18144 2632
rect 17681 2595 17739 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 19334 2592 19340 2644
rect 19392 2632 19398 2644
rect 19889 2635 19947 2641
rect 19889 2632 19901 2635
rect 19392 2604 19901 2632
rect 19392 2592 19398 2604
rect 19889 2601 19901 2604
rect 19935 2601 19947 2635
rect 20622 2632 20628 2644
rect 20583 2604 20628 2632
rect 19889 2595 19947 2601
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 20990 2632 20996 2644
rect 20951 2604 20996 2632
rect 20990 2592 20996 2604
rect 21048 2592 21054 2644
rect 21545 2635 21603 2641
rect 21545 2601 21557 2635
rect 21591 2632 21603 2635
rect 23014 2632 23020 2644
rect 21591 2604 23020 2632
rect 21591 2601 21603 2604
rect 21545 2595 21603 2601
rect 16298 2564 16304 2576
rect 16259 2536 16304 2564
rect 16298 2524 16304 2536
rect 16356 2524 16362 2576
rect 16850 2564 16856 2576
rect 16763 2536 16856 2564
rect 16850 2524 16856 2536
rect 16908 2564 16914 2576
rect 18156 2564 18184 2592
rect 18646 2567 18704 2573
rect 18646 2564 18658 2567
rect 16908 2536 17724 2564
rect 18156 2536 18658 2564
rect 16908 2524 16914 2536
rect 15519 2468 16068 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11425 2431 11483 2437
rect 11425 2428 11437 2431
rect 11020 2400 11437 2428
rect 11020 2388 11026 2400
rect 11425 2397 11437 2400
rect 11471 2397 11483 2431
rect 11425 2391 11483 2397
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12115 2400 14044 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 8205 2363 8263 2369
rect 8205 2329 8217 2363
rect 8251 2360 8263 2363
rect 8662 2360 8668 2372
rect 8251 2332 8668 2360
rect 8251 2329 8263 2332
rect 8205 2323 8263 2329
rect 8662 2320 8668 2332
rect 8720 2320 8726 2372
rect 11440 2360 11468 2391
rect 13814 2360 13820 2372
rect 11440 2332 13820 2360
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 14016 2360 14044 2400
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14182 2431 14240 2437
rect 14182 2428 14194 2431
rect 14148 2400 14194 2428
rect 14148 2388 14154 2400
rect 14182 2397 14194 2400
rect 14228 2397 14240 2431
rect 14182 2391 14240 2397
rect 14274 2388 14280 2440
rect 14332 2428 14338 2440
rect 16758 2428 16764 2440
rect 14332 2400 14377 2428
rect 16671 2400 16764 2428
rect 14332 2388 14338 2400
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 17696 2428 17724 2536
rect 18646 2533 18658 2536
rect 18692 2533 18704 2567
rect 18646 2527 18704 2533
rect 19613 2567 19671 2573
rect 19613 2533 19625 2567
rect 19659 2564 19671 2567
rect 21560 2564 21588 2595
rect 23014 2592 23020 2604
rect 23072 2592 23078 2644
rect 24118 2592 24124 2644
rect 24176 2632 24182 2644
rect 25777 2635 25835 2641
rect 25777 2632 25789 2635
rect 24176 2604 25789 2632
rect 24176 2592 24182 2604
rect 25777 2601 25789 2604
rect 25823 2632 25835 2635
rect 25961 2635 26019 2641
rect 25961 2632 25973 2635
rect 25823 2604 25973 2632
rect 25823 2601 25835 2604
rect 25777 2595 25835 2601
rect 25961 2601 25973 2604
rect 26007 2601 26019 2635
rect 26142 2632 26148 2644
rect 26055 2604 26148 2632
rect 25961 2595 26019 2601
rect 26142 2592 26148 2604
rect 26200 2632 26206 2644
rect 26605 2635 26663 2641
rect 26605 2632 26617 2635
rect 26200 2604 26617 2632
rect 26200 2592 26206 2604
rect 26605 2601 26617 2604
rect 26651 2632 26663 2635
rect 27246 2632 27252 2644
rect 26651 2604 27252 2632
rect 26651 2601 26663 2604
rect 26605 2595 26663 2601
rect 27246 2592 27252 2604
rect 27304 2592 27310 2644
rect 28074 2592 28080 2644
rect 28132 2632 28138 2644
rect 29089 2635 29147 2641
rect 29089 2632 29101 2635
rect 28132 2604 29101 2632
rect 28132 2592 28138 2604
rect 29089 2601 29101 2604
rect 29135 2601 29147 2635
rect 29546 2632 29552 2644
rect 29507 2604 29552 2632
rect 29089 2595 29147 2601
rect 19659 2536 21588 2564
rect 19659 2533 19671 2536
rect 19613 2527 19671 2533
rect 21726 2524 21732 2576
rect 21784 2564 21790 2576
rect 23109 2567 23167 2573
rect 21784 2536 22140 2564
rect 21784 2524 21790 2536
rect 18322 2496 18328 2508
rect 18283 2468 18328 2496
rect 18322 2456 18328 2468
rect 18380 2456 18386 2508
rect 20140 2499 20198 2505
rect 20140 2465 20152 2499
rect 20186 2496 20198 2499
rect 21450 2496 21456 2508
rect 20186 2468 21456 2496
rect 20186 2465 20198 2468
rect 20140 2459 20198 2465
rect 17696 2400 18368 2428
rect 16776 2360 16804 2388
rect 14016 2332 16804 2360
rect 18340 2360 18368 2400
rect 19245 2363 19303 2369
rect 19245 2360 19257 2363
rect 18340 2332 19257 2360
rect 19245 2329 19257 2332
rect 19291 2329 19303 2363
rect 20155 2360 20183 2459
rect 21450 2456 21456 2468
rect 21508 2456 21514 2508
rect 21913 2499 21971 2505
rect 21913 2465 21925 2499
rect 21959 2496 21971 2499
rect 22002 2496 22008 2508
rect 21959 2468 22008 2496
rect 21959 2465 21971 2468
rect 21913 2459 21971 2465
rect 22002 2456 22008 2468
rect 22060 2456 22066 2508
rect 22112 2505 22140 2536
rect 23109 2533 23121 2567
rect 23155 2564 23167 2567
rect 26234 2564 26240 2576
rect 23155 2536 26240 2564
rect 23155 2533 23167 2536
rect 23109 2527 23167 2533
rect 26234 2524 26240 2536
rect 26292 2524 26298 2576
rect 29104 2564 29132 2595
rect 29546 2592 29552 2604
rect 29604 2632 29610 2644
rect 32030 2632 32036 2644
rect 29604 2604 29960 2632
rect 29604 2592 29610 2604
rect 29932 2573 29960 2604
rect 31956 2604 32036 2632
rect 29825 2567 29883 2573
rect 29825 2564 29837 2567
rect 29104 2536 29837 2564
rect 29825 2533 29837 2536
rect 29871 2533 29883 2567
rect 29825 2527 29883 2533
rect 29917 2567 29975 2573
rect 29917 2533 29929 2567
rect 29963 2533 29975 2567
rect 29917 2527 29975 2533
rect 30926 2524 30932 2576
rect 30984 2564 30990 2576
rect 31297 2567 31355 2573
rect 31297 2564 31309 2567
rect 30984 2536 31309 2564
rect 30984 2524 30990 2536
rect 31297 2533 31309 2536
rect 31343 2564 31355 2567
rect 31846 2564 31852 2576
rect 31343 2536 31852 2564
rect 31343 2533 31355 2536
rect 31297 2527 31355 2533
rect 31846 2524 31852 2536
rect 31904 2524 31910 2576
rect 22097 2499 22155 2505
rect 22097 2465 22109 2499
rect 22143 2465 22155 2499
rect 22097 2459 22155 2465
rect 22465 2499 22523 2505
rect 22465 2465 22477 2499
rect 22511 2465 22523 2499
rect 23014 2496 23020 2508
rect 22927 2468 23020 2496
rect 22465 2459 22523 2465
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 22278 2428 22284 2440
rect 20680 2400 22284 2428
rect 20680 2388 20686 2400
rect 22278 2388 22284 2400
rect 22336 2428 22342 2440
rect 22480 2428 22508 2459
rect 23014 2456 23020 2468
rect 23072 2456 23078 2508
rect 23658 2456 23664 2508
rect 23716 2496 23722 2508
rect 24029 2499 24087 2505
rect 24029 2496 24041 2499
rect 23716 2468 24041 2496
rect 23716 2456 23722 2468
rect 24029 2465 24041 2468
rect 24075 2465 24087 2499
rect 24029 2459 24087 2465
rect 24118 2456 24124 2508
rect 24176 2496 24182 2508
rect 24489 2499 24547 2505
rect 24489 2496 24501 2499
rect 24176 2468 24501 2496
rect 24176 2456 24182 2468
rect 24489 2465 24501 2468
rect 24535 2465 24547 2499
rect 24946 2496 24952 2508
rect 24907 2468 24952 2496
rect 24489 2459 24547 2465
rect 24946 2456 24952 2468
rect 25004 2456 25010 2508
rect 25225 2499 25283 2505
rect 25225 2465 25237 2499
rect 25271 2465 25283 2499
rect 25225 2459 25283 2465
rect 25501 2499 25559 2505
rect 25501 2465 25513 2499
rect 25547 2496 25559 2499
rect 26881 2499 26939 2505
rect 26881 2496 26893 2499
rect 25547 2468 26893 2496
rect 25547 2465 25559 2468
rect 25501 2459 25559 2465
rect 26881 2465 26893 2468
rect 26927 2496 26939 2499
rect 27430 2496 27436 2508
rect 26927 2468 27436 2496
rect 26927 2465 26939 2468
rect 26881 2459 26939 2465
rect 22336 2400 22508 2428
rect 23032 2428 23060 2456
rect 23845 2431 23903 2437
rect 23845 2428 23857 2431
rect 23032 2400 23857 2428
rect 22336 2388 22342 2400
rect 23845 2397 23857 2400
rect 23891 2428 23903 2431
rect 25240 2428 25268 2459
rect 27430 2456 27436 2468
rect 27488 2456 27494 2508
rect 27801 2499 27859 2505
rect 27801 2465 27813 2499
rect 27847 2496 27859 2499
rect 28696 2499 28754 2505
rect 27847 2468 28488 2496
rect 27847 2465 27859 2468
rect 27801 2459 27859 2465
rect 23891 2400 25268 2428
rect 25961 2431 26019 2437
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 25961 2397 25973 2431
rect 26007 2428 26019 2431
rect 28077 2431 28135 2437
rect 28077 2428 28089 2431
rect 26007 2400 28089 2428
rect 26007 2397 26019 2400
rect 25961 2391 26019 2397
rect 28077 2397 28089 2400
rect 28123 2397 28135 2431
rect 28460 2428 28488 2468
rect 28696 2465 28708 2499
rect 28742 2465 28754 2499
rect 28696 2459 28754 2465
rect 31548 2499 31606 2505
rect 31548 2465 31560 2499
rect 31594 2496 31606 2499
rect 31956 2496 31984 2604
rect 32030 2592 32036 2604
rect 32088 2592 32094 2644
rect 32122 2524 32128 2576
rect 32180 2564 32186 2576
rect 34149 2567 34207 2573
rect 34149 2564 34161 2567
rect 32180 2536 34161 2564
rect 32180 2524 32186 2536
rect 34149 2533 34161 2536
rect 34195 2533 34207 2567
rect 34149 2527 34207 2533
rect 31594 2468 31984 2496
rect 32217 2499 32275 2505
rect 31594 2465 31606 2468
rect 31548 2459 31606 2465
rect 32217 2465 32229 2499
rect 32263 2496 32275 2499
rect 32674 2496 32680 2508
rect 32263 2468 32680 2496
rect 32263 2465 32275 2468
rect 32217 2459 32275 2465
rect 28711 2428 28739 2459
rect 32674 2456 32680 2468
rect 32732 2456 32738 2508
rect 29270 2428 29276 2440
rect 28460 2400 28672 2428
rect 28711 2400 29276 2428
rect 28077 2391 28135 2397
rect 19245 2323 19303 2329
rect 19812 2332 20183 2360
rect 20211 2363 20269 2369
rect 10502 2292 10508 2304
rect 10463 2264 10508 2292
rect 10502 2252 10508 2264
rect 10560 2252 10566 2304
rect 14093 2295 14151 2301
rect 14093 2261 14105 2295
rect 14139 2292 14151 2295
rect 14918 2292 14924 2304
rect 14139 2264 14924 2292
rect 14139 2261 14151 2264
rect 14093 2255 14151 2261
rect 14918 2252 14924 2264
rect 14976 2252 14982 2304
rect 17497 2295 17555 2301
rect 17497 2261 17509 2295
rect 17543 2292 17555 2295
rect 19812 2292 19840 2332
rect 20211 2329 20223 2363
rect 20257 2360 20269 2363
rect 22094 2360 22100 2372
rect 20257 2332 22100 2360
rect 20257 2329 20269 2332
rect 20211 2323 20269 2329
rect 22094 2320 22100 2332
rect 22152 2320 22158 2372
rect 24946 2320 24952 2372
rect 25004 2360 25010 2372
rect 28445 2363 28503 2369
rect 28445 2360 28457 2363
rect 25004 2332 28457 2360
rect 25004 2320 25010 2332
rect 28445 2329 28457 2332
rect 28491 2329 28503 2363
rect 28644 2360 28672 2400
rect 29270 2388 29276 2400
rect 29328 2428 29334 2440
rect 30101 2431 30159 2437
rect 30101 2428 30113 2431
rect 29328 2400 30113 2428
rect 29328 2388 29334 2400
rect 30101 2397 30113 2400
rect 30147 2397 30159 2431
rect 30101 2391 30159 2397
rect 30929 2431 30987 2437
rect 30929 2397 30941 2431
rect 30975 2428 30987 2431
rect 31202 2428 31208 2440
rect 30975 2400 31208 2428
rect 30975 2397 30987 2400
rect 30929 2391 30987 2397
rect 31202 2388 31208 2400
rect 31260 2428 31266 2440
rect 32585 2431 32643 2437
rect 32585 2428 32597 2431
rect 31260 2400 32597 2428
rect 31260 2388 31266 2400
rect 32585 2397 32597 2400
rect 32631 2397 32643 2431
rect 32585 2391 32643 2397
rect 31619 2363 31677 2369
rect 28644 2332 31591 2360
rect 28445 2323 28503 2329
rect 17543 2264 19840 2292
rect 17543 2261 17555 2264
rect 17497 2255 17555 2261
rect 22002 2252 22008 2304
rect 22060 2292 22066 2304
rect 23385 2295 23443 2301
rect 23385 2292 23397 2295
rect 22060 2264 23397 2292
rect 22060 2252 22066 2264
rect 23385 2261 23397 2264
rect 23431 2292 23443 2295
rect 23658 2292 23664 2304
rect 23431 2264 23664 2292
rect 23431 2261 23443 2264
rect 23385 2255 23443 2261
rect 23658 2252 23664 2264
rect 23716 2252 23722 2304
rect 28767 2295 28825 2301
rect 28767 2261 28779 2295
rect 28813 2292 28825 2295
rect 30742 2292 30748 2304
rect 28813 2264 30748 2292
rect 28813 2261 28825 2264
rect 28767 2255 28825 2261
rect 30742 2252 30748 2264
rect 30800 2252 30806 2304
rect 31563 2292 31591 2332
rect 31619 2329 31631 2363
rect 31665 2360 31677 2363
rect 34146 2360 34152 2372
rect 31665 2332 34152 2360
rect 31665 2329 31677 2332
rect 31619 2323 31677 2329
rect 34146 2320 34152 2332
rect 34204 2320 34210 2372
rect 32217 2295 32275 2301
rect 32217 2292 32229 2295
rect 31563 2264 32229 2292
rect 32217 2261 32229 2264
rect 32263 2292 32275 2295
rect 32309 2295 32367 2301
rect 32309 2292 32321 2295
rect 32263 2264 32321 2292
rect 32263 2261 32275 2264
rect 32217 2255 32275 2261
rect 32309 2261 32321 2264
rect 32355 2261 32367 2295
rect 32309 2255 32367 2261
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
rect 1670 2048 1676 2100
rect 1728 2088 1734 2100
rect 10502 2088 10508 2100
rect 1728 2060 10508 2088
rect 1728 2048 1734 2060
rect 10502 2048 10508 2060
rect 10560 2048 10566 2100
<< via1 >>
rect 5816 15512 5868 15564
rect 6644 15512 6696 15564
rect 19984 15512 20036 15564
rect 20628 15512 20680 15564
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 35624 11339 35676 11348
rect 35624 11305 35633 11339
rect 35633 11305 35667 11339
rect 35667 11305 35676 11339
rect 35624 11296 35676 11305
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 35440 11203 35492 11212
rect 35440 11169 35449 11203
rect 35449 11169 35483 11203
rect 35483 11169 35492 11203
rect 35440 11160 35492 11169
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 1400 10412 1452 10464
rect 2228 10412 2280 10464
rect 29828 10412 29880 10464
rect 35440 10455 35492 10464
rect 35440 10421 35449 10455
rect 35449 10421 35483 10455
rect 35483 10421 35492 10455
rect 35440 10412 35492 10421
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 35624 10251 35676 10260
rect 35624 10217 35633 10251
rect 35633 10217 35667 10251
rect 35667 10217 35676 10251
rect 35624 10208 35676 10217
rect 1676 10072 1728 10124
rect 35440 10115 35492 10124
rect 35440 10081 35449 10115
rect 35449 10081 35483 10115
rect 35483 10081 35492 10115
rect 35440 10072 35492 10081
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 35440 9367 35492 9376
rect 35440 9333 35449 9367
rect 35449 9333 35483 9367
rect 35483 9333 35492 9367
rect 35440 9324 35492 9333
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 35624 9163 35676 9172
rect 35624 9129 35633 9163
rect 35633 9129 35667 9163
rect 35667 9129 35676 9163
rect 35624 9120 35676 9129
rect 2136 8984 2188 9036
rect 2228 8984 2280 9036
rect 3332 8984 3384 9036
rect 35256 8984 35308 9036
rect 4988 8780 5040 8832
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 1216 8576 1268 8628
rect 35624 8619 35676 8628
rect 35624 8585 35633 8619
rect 35633 8585 35667 8619
rect 35667 8585 35676 8619
rect 35624 8576 35676 8585
rect 4068 8415 4120 8424
rect 2136 8236 2188 8288
rect 4068 8381 4077 8415
rect 4077 8381 4111 8415
rect 4111 8381 4120 8415
rect 4068 8372 4120 8381
rect 3424 8304 3476 8356
rect 4344 8304 4396 8356
rect 34060 8372 34112 8424
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 3332 8279 3384 8288
rect 3332 8245 3341 8279
rect 3341 8245 3375 8279
rect 3375 8245 3384 8279
rect 3332 8236 3384 8245
rect 4804 8236 4856 8288
rect 5080 8279 5132 8288
rect 5080 8245 5089 8279
rect 5089 8245 5123 8279
rect 5123 8245 5132 8279
rect 5080 8236 5132 8245
rect 34152 8236 34204 8288
rect 35256 8279 35308 8288
rect 35256 8245 35265 8279
rect 35265 8245 35299 8279
rect 35299 8245 35308 8279
rect 35256 8236 35308 8245
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 4988 8032 5040 8084
rect 5816 8075 5868 8084
rect 5816 8041 5825 8075
rect 5825 8041 5859 8075
rect 5859 8041 5868 8075
rect 5816 8032 5868 8041
rect 35716 8032 35768 8084
rect 4160 7964 4212 8016
rect 2044 7896 2096 7948
rect 2504 7939 2556 7948
rect 2504 7905 2513 7939
rect 2513 7905 2547 7939
rect 2547 7905 2556 7939
rect 2504 7896 2556 7905
rect 5448 7896 5500 7948
rect 14188 7939 14240 7948
rect 14188 7905 14197 7939
rect 14197 7905 14231 7939
rect 14231 7905 14240 7939
rect 14188 7896 14240 7905
rect 19616 7896 19668 7948
rect 35440 7939 35492 7948
rect 35440 7905 35449 7939
rect 35449 7905 35483 7939
rect 35483 7905 35492 7939
rect 35440 7896 35492 7905
rect 4344 7828 4396 7880
rect 4988 7828 5040 7880
rect 9956 7828 10008 7880
rect 2688 7803 2740 7812
rect 2688 7769 2697 7803
rect 2697 7769 2731 7803
rect 2731 7769 2740 7803
rect 2688 7760 2740 7769
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 10324 7692 10376 7744
rect 14464 7692 14516 7744
rect 22008 7692 22060 7744
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 1492 7488 1544 7540
rect 4344 7488 4396 7540
rect 16764 7531 16816 7540
rect 16764 7497 16773 7531
rect 16773 7497 16807 7531
rect 16807 7497 16816 7531
rect 16764 7488 16816 7497
rect 35440 7488 35492 7540
rect 35532 7488 35584 7540
rect 36728 7531 36780 7540
rect 36728 7497 36737 7531
rect 36737 7497 36771 7531
rect 36771 7497 36780 7531
rect 36728 7488 36780 7497
rect 2504 7420 2556 7472
rect 3608 7420 3660 7472
rect 4160 7463 4212 7472
rect 4160 7429 4169 7463
rect 4169 7429 4203 7463
rect 4203 7429 4212 7463
rect 4160 7420 4212 7429
rect 3240 7352 3292 7404
rect 4896 7420 4948 7472
rect 15384 7420 15436 7472
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 14924 7352 14976 7404
rect 35992 7395 36044 7404
rect 1676 7284 1728 7336
rect 5356 7284 5408 7336
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 13636 7284 13688 7336
rect 15200 7284 15252 7336
rect 18880 7284 18932 7336
rect 19984 7284 20036 7336
rect 20168 7327 20220 7336
rect 20168 7293 20186 7327
rect 20186 7293 20220 7327
rect 20168 7284 20220 7293
rect 22744 7284 22796 7336
rect 35992 7361 36001 7395
rect 36001 7361 36035 7395
rect 36035 7361 36044 7395
rect 35992 7352 36044 7361
rect 2044 7259 2096 7268
rect 2044 7225 2053 7259
rect 2053 7225 2087 7259
rect 2087 7225 2096 7259
rect 2044 7216 2096 7225
rect 3148 7259 3200 7268
rect 3148 7225 3157 7259
rect 3157 7225 3191 7259
rect 3191 7225 3200 7259
rect 3148 7216 3200 7225
rect 3240 7259 3292 7268
rect 3240 7225 3249 7259
rect 3249 7225 3283 7259
rect 3283 7225 3292 7259
rect 3240 7216 3292 7225
rect 4528 7216 4580 7268
rect 3516 7148 3568 7200
rect 4068 7148 4120 7200
rect 14832 7216 14884 7268
rect 5448 7148 5500 7200
rect 7196 7148 7248 7200
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 10508 7148 10560 7200
rect 14188 7191 14240 7200
rect 14188 7157 14197 7191
rect 14197 7157 14231 7191
rect 14231 7157 14240 7191
rect 14188 7148 14240 7157
rect 21272 7216 21324 7268
rect 23940 7216 23992 7268
rect 26148 7216 26200 7268
rect 15568 7148 15620 7200
rect 18972 7191 19024 7200
rect 18972 7157 18981 7191
rect 18981 7157 19015 7191
rect 19015 7157 19024 7191
rect 18972 7148 19024 7157
rect 19616 7191 19668 7200
rect 19616 7157 19625 7191
rect 19625 7157 19659 7191
rect 19659 7157 19668 7191
rect 19616 7148 19668 7157
rect 20352 7191 20404 7200
rect 20352 7157 20361 7191
rect 20361 7157 20395 7191
rect 20395 7157 20404 7191
rect 20352 7148 20404 7157
rect 20904 7191 20956 7200
rect 20904 7157 20913 7191
rect 20913 7157 20947 7191
rect 20947 7157 20956 7191
rect 20904 7148 20956 7157
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 20628 6944 20680 6996
rect 39580 6944 39632 6996
rect 2412 6876 2464 6928
rect 4252 6919 4304 6928
rect 4252 6885 4261 6919
rect 4261 6885 4295 6919
rect 4295 6885 4304 6919
rect 4252 6876 4304 6885
rect 4804 6876 4856 6928
rect 5724 6919 5776 6928
rect 5724 6885 5733 6919
rect 5733 6885 5767 6919
rect 5767 6885 5776 6919
rect 5724 6876 5776 6885
rect 5816 6919 5868 6928
rect 5816 6885 5825 6919
rect 5825 6885 5859 6919
rect 5859 6885 5868 6919
rect 10324 6919 10376 6928
rect 5816 6876 5868 6885
rect 10324 6885 10333 6919
rect 10333 6885 10367 6919
rect 10367 6885 10376 6919
rect 10324 6876 10376 6885
rect 10416 6919 10468 6928
rect 10416 6885 10425 6919
rect 10425 6885 10459 6919
rect 10459 6885 10468 6919
rect 10416 6876 10468 6885
rect 14004 6876 14056 6928
rect 15476 6919 15528 6928
rect 15476 6885 15485 6919
rect 15485 6885 15519 6919
rect 15519 6885 15528 6919
rect 15476 6876 15528 6885
rect 19064 6876 19116 6928
rect 20720 6876 20772 6928
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 16764 6808 16816 6860
rect 18328 6808 18380 6860
rect 23480 6808 23532 6860
rect 24492 6851 24544 6860
rect 24492 6817 24501 6851
rect 24501 6817 24535 6851
rect 24535 6817 24544 6851
rect 24492 6808 24544 6817
rect 35440 6851 35492 6860
rect 35440 6817 35449 6851
rect 35449 6817 35483 6851
rect 35483 6817 35492 6851
rect 35440 6808 35492 6817
rect 1676 6647 1728 6656
rect 1676 6613 1685 6647
rect 1685 6613 1719 6647
rect 1719 6613 1728 6647
rect 1676 6604 1728 6613
rect 3792 6740 3844 6792
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 2596 6672 2648 6724
rect 4988 6672 5040 6724
rect 6920 6740 6972 6792
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 15384 6783 15436 6792
rect 15384 6749 15393 6783
rect 15393 6749 15427 6783
rect 15427 6749 15436 6783
rect 15384 6740 15436 6749
rect 15568 6740 15620 6792
rect 18788 6740 18840 6792
rect 20812 6740 20864 6792
rect 10600 6672 10652 6724
rect 18972 6672 19024 6724
rect 19984 6672 20036 6724
rect 20904 6672 20956 6724
rect 21548 6715 21600 6724
rect 21548 6681 21557 6715
rect 21557 6681 21591 6715
rect 21591 6681 21600 6715
rect 21548 6672 21600 6681
rect 2504 6604 2556 6656
rect 4068 6604 4120 6656
rect 4344 6604 4396 6656
rect 13820 6604 13872 6656
rect 14832 6604 14884 6656
rect 15108 6647 15160 6656
rect 15108 6613 15117 6647
rect 15117 6613 15151 6647
rect 15151 6613 15160 6647
rect 15108 6604 15160 6613
rect 16948 6604 17000 6656
rect 18696 6647 18748 6656
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 19064 6647 19116 6656
rect 19064 6613 19073 6647
rect 19073 6613 19107 6647
rect 19107 6613 19116 6647
rect 19064 6604 19116 6613
rect 19340 6604 19392 6656
rect 20352 6604 20404 6656
rect 24584 6647 24636 6656
rect 24584 6613 24593 6647
rect 24593 6613 24627 6647
rect 24627 6613 24636 6647
rect 24584 6604 24636 6613
rect 25136 6604 25188 6656
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 20 6400 72 6452
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 3240 6400 3292 6452
rect 4068 6443 4120 6452
rect 4068 6409 4077 6443
rect 4077 6409 4111 6443
rect 4111 6409 4120 6443
rect 4068 6400 4120 6409
rect 2412 6375 2464 6384
rect 2412 6341 2421 6375
rect 2421 6341 2455 6375
rect 2455 6341 2464 6375
rect 2412 6332 2464 6341
rect 2044 6196 2096 6248
rect 2596 6196 2648 6248
rect 4436 6400 4488 6452
rect 5724 6400 5776 6452
rect 8576 6400 8628 6452
rect 4252 6332 4304 6384
rect 5816 6332 5868 6384
rect 4344 6307 4396 6316
rect 3424 6128 3476 6180
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 6920 6307 6972 6316
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 10416 6400 10468 6452
rect 15200 6400 15252 6452
rect 15476 6400 15528 6452
rect 18328 6443 18380 6452
rect 18328 6409 18337 6443
rect 18337 6409 18371 6443
rect 18371 6409 18380 6443
rect 18328 6400 18380 6409
rect 18788 6400 18840 6452
rect 21272 6400 21324 6452
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 24492 6443 24544 6452
rect 23480 6400 23532 6409
rect 24492 6409 24501 6443
rect 24501 6409 24535 6443
rect 24535 6409 24544 6443
rect 24492 6400 24544 6409
rect 24860 6400 24912 6452
rect 12532 6332 12584 6384
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 14372 6332 14424 6384
rect 21548 6332 21600 6384
rect 14924 6264 14976 6316
rect 15108 6264 15160 6316
rect 18972 6264 19024 6316
rect 20812 6264 20864 6316
rect 22376 6264 22428 6316
rect 12440 6239 12492 6248
rect 12440 6205 12449 6239
rect 12449 6205 12483 6239
rect 12483 6205 12492 6239
rect 12440 6196 12492 6205
rect 13820 6196 13872 6248
rect 17500 6196 17552 6248
rect 18604 6196 18656 6248
rect 25412 6307 25464 6316
rect 25412 6273 25421 6307
rect 25421 6273 25455 6307
rect 25455 6273 25464 6307
rect 25412 6264 25464 6273
rect 35440 6307 35492 6316
rect 35440 6273 35449 6307
rect 35449 6273 35483 6307
rect 35483 6273 35492 6307
rect 35440 6264 35492 6273
rect 9128 6171 9180 6180
rect 4068 6060 4120 6112
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 9128 6137 9137 6171
rect 9137 6137 9171 6171
rect 9171 6137 9180 6171
rect 9128 6128 9180 6137
rect 9496 6128 9548 6180
rect 13544 6171 13596 6180
rect 13544 6137 13553 6171
rect 13553 6137 13587 6171
rect 13587 6137 13596 6171
rect 13544 6128 13596 6137
rect 12624 6103 12676 6112
rect 6552 6060 6604 6069
rect 12624 6069 12633 6103
rect 12633 6069 12667 6103
rect 12667 6069 12676 6103
rect 12624 6060 12676 6069
rect 14832 6128 14884 6180
rect 15660 6128 15712 6180
rect 20536 6171 20588 6180
rect 14740 6060 14792 6112
rect 15384 6060 15436 6112
rect 16764 6103 16816 6112
rect 16764 6069 16773 6103
rect 16773 6069 16807 6103
rect 16807 6069 16816 6103
rect 16764 6060 16816 6069
rect 17500 6103 17552 6112
rect 17500 6069 17509 6103
rect 17509 6069 17543 6103
rect 17543 6069 17552 6103
rect 17500 6060 17552 6069
rect 17776 6103 17828 6112
rect 17776 6069 17785 6103
rect 17785 6069 17819 6103
rect 17819 6069 17828 6103
rect 17776 6060 17828 6069
rect 18972 6060 19024 6112
rect 20536 6137 20545 6171
rect 20545 6137 20579 6171
rect 20579 6137 20588 6171
rect 21088 6171 21140 6180
rect 20536 6128 20588 6137
rect 20720 6060 20772 6112
rect 21088 6137 21097 6171
rect 21097 6137 21131 6171
rect 21131 6137 21140 6171
rect 21088 6128 21140 6137
rect 24400 6128 24452 6180
rect 25136 6171 25188 6180
rect 25136 6137 25145 6171
rect 25145 6137 25179 6171
rect 25179 6137 25188 6171
rect 25136 6128 25188 6137
rect 22560 6060 22612 6112
rect 24032 6103 24084 6112
rect 24032 6069 24041 6103
rect 24041 6069 24075 6103
rect 24075 6069 24084 6103
rect 24032 6060 24084 6069
rect 25504 6060 25556 6112
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 4252 5856 4304 5908
rect 4436 5899 4488 5908
rect 4436 5865 4445 5899
rect 4445 5865 4479 5899
rect 4479 5865 4488 5899
rect 4436 5856 4488 5865
rect 6276 5899 6328 5908
rect 6276 5865 6285 5899
rect 6285 5865 6319 5899
rect 6319 5865 6328 5899
rect 6276 5856 6328 5865
rect 7472 5856 7524 5908
rect 2412 5788 2464 5840
rect 9128 5856 9180 5908
rect 10324 5899 10376 5908
rect 10324 5865 10333 5899
rect 10333 5865 10367 5899
rect 10367 5865 10376 5899
rect 10324 5856 10376 5865
rect 14004 5899 14056 5908
rect 14004 5865 14013 5899
rect 14013 5865 14047 5899
rect 14047 5865 14056 5899
rect 14004 5856 14056 5865
rect 21272 5899 21324 5908
rect 10416 5788 10468 5840
rect 13544 5788 13596 5840
rect 14740 5788 14792 5840
rect 18144 5788 18196 5840
rect 19340 5831 19392 5840
rect 19340 5797 19349 5831
rect 19349 5797 19383 5831
rect 19383 5797 19392 5831
rect 19340 5788 19392 5797
rect 21272 5865 21281 5899
rect 21281 5865 21315 5899
rect 21315 5865 21324 5899
rect 21272 5856 21324 5865
rect 25412 5899 25464 5908
rect 25412 5865 25421 5899
rect 25421 5865 25455 5899
rect 25455 5865 25464 5899
rect 25412 5856 25464 5865
rect 20536 5788 20588 5840
rect 22560 5831 22612 5840
rect 22560 5797 22569 5831
rect 22569 5797 22603 5831
rect 22603 5797 22612 5831
rect 22560 5788 22612 5797
rect 22928 5788 22980 5840
rect 24584 5831 24636 5840
rect 24584 5797 24593 5831
rect 24593 5797 24627 5831
rect 24627 5797 24636 5831
rect 24584 5788 24636 5797
rect 12624 5720 12676 5772
rect 13268 5720 13320 5772
rect 19984 5763 20036 5772
rect 19984 5729 19993 5763
rect 19993 5729 20027 5763
rect 20027 5729 20036 5763
rect 19984 5720 20036 5729
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 4528 5652 4580 5704
rect 6644 5652 6696 5704
rect 7380 5652 7432 5704
rect 7196 5584 7248 5636
rect 10508 5652 10560 5704
rect 13728 5652 13780 5704
rect 15568 5652 15620 5704
rect 1768 5559 1820 5568
rect 1768 5525 1777 5559
rect 1777 5525 1811 5559
rect 1811 5525 1820 5559
rect 1768 5516 1820 5525
rect 2136 5559 2188 5568
rect 2136 5525 2145 5559
rect 2145 5525 2179 5559
rect 2179 5525 2188 5559
rect 2136 5516 2188 5525
rect 3056 5516 3108 5568
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 4988 5559 5040 5568
rect 4988 5525 4997 5559
rect 4997 5525 5031 5559
rect 5031 5525 5040 5559
rect 4988 5516 5040 5525
rect 8116 5516 8168 5568
rect 12348 5516 12400 5568
rect 15016 5559 15068 5568
rect 15016 5525 15025 5559
rect 15025 5525 15059 5559
rect 15059 5525 15068 5559
rect 15016 5516 15068 5525
rect 15200 5516 15252 5568
rect 16856 5516 16908 5568
rect 20628 5652 20680 5704
rect 25504 5720 25556 5772
rect 27252 5720 27304 5772
rect 21456 5652 21508 5704
rect 24032 5652 24084 5704
rect 24492 5695 24544 5704
rect 24492 5661 24501 5695
rect 24501 5661 24535 5695
rect 24535 5661 24544 5695
rect 24492 5652 24544 5661
rect 26516 5695 26568 5704
rect 23480 5584 23532 5636
rect 26516 5661 26525 5695
rect 26525 5661 26559 5695
rect 26559 5661 26568 5695
rect 26516 5652 26568 5661
rect 25320 5584 25372 5636
rect 17868 5516 17920 5568
rect 18880 5516 18932 5568
rect 20352 5559 20404 5568
rect 20352 5525 20361 5559
rect 20361 5525 20395 5559
rect 20395 5525 20404 5559
rect 20352 5516 20404 5525
rect 21824 5559 21876 5568
rect 21824 5525 21833 5559
rect 21833 5525 21867 5559
rect 21867 5525 21876 5559
rect 21824 5516 21876 5525
rect 22100 5559 22152 5568
rect 22100 5525 22109 5559
rect 22109 5525 22143 5559
rect 22143 5525 22152 5559
rect 22100 5516 22152 5525
rect 22284 5516 22336 5568
rect 27436 5516 27488 5568
rect 27896 5559 27948 5568
rect 27896 5525 27905 5559
rect 27905 5525 27939 5559
rect 27939 5525 27948 5559
rect 27896 5516 27948 5525
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 1032 5312 1084 5364
rect 2412 5355 2464 5364
rect 2412 5321 2421 5355
rect 2421 5321 2455 5355
rect 2455 5321 2464 5355
rect 2412 5312 2464 5321
rect 6552 5312 6604 5364
rect 7380 5355 7432 5364
rect 1768 5176 1820 5228
rect 7380 5321 7389 5355
rect 7389 5321 7423 5355
rect 7423 5321 7432 5355
rect 7380 5312 7432 5321
rect 9128 5312 9180 5364
rect 10416 5312 10468 5364
rect 13544 5312 13596 5364
rect 15660 5355 15712 5364
rect 8116 5176 8168 5228
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 2136 5108 2188 5160
rect 3056 5151 3108 5160
rect 3056 5117 3065 5151
rect 3065 5117 3099 5151
rect 3099 5117 3108 5151
rect 3056 5108 3108 5117
rect 3424 5151 3476 5160
rect 3424 5117 3433 5151
rect 3433 5117 3467 5151
rect 3467 5117 3476 5151
rect 3424 5108 3476 5117
rect 4068 5108 4120 5160
rect 5080 5108 5132 5160
rect 9588 5151 9640 5160
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 5172 5040 5224 5092
rect 6276 5083 6328 5092
rect 2596 5015 2648 5024
rect 2596 4981 2605 5015
rect 2605 4981 2639 5015
rect 2639 4981 2648 5015
rect 2596 4972 2648 4981
rect 4436 4972 4488 5024
rect 6276 5049 6285 5083
rect 6285 5049 6319 5083
rect 6319 5049 6328 5083
rect 6276 5040 6328 5049
rect 8208 5083 8260 5092
rect 8208 5049 8211 5083
rect 8211 5049 8245 5083
rect 8245 5049 8260 5083
rect 13820 5287 13872 5296
rect 13820 5253 13829 5287
rect 13829 5253 13863 5287
rect 13863 5253 13872 5287
rect 15660 5321 15669 5355
rect 15669 5321 15703 5355
rect 15703 5321 15712 5355
rect 15660 5312 15712 5321
rect 18972 5355 19024 5364
rect 18972 5321 18981 5355
rect 18981 5321 19015 5355
rect 19015 5321 19024 5355
rect 18972 5312 19024 5321
rect 20720 5355 20772 5364
rect 20720 5321 20729 5355
rect 20729 5321 20763 5355
rect 20763 5321 20772 5355
rect 22928 5355 22980 5364
rect 20720 5312 20772 5321
rect 22928 5321 22937 5355
rect 22937 5321 22971 5355
rect 22971 5321 22980 5355
rect 22928 5312 22980 5321
rect 24400 5312 24452 5364
rect 24584 5355 24636 5364
rect 24584 5321 24593 5355
rect 24593 5321 24627 5355
rect 24627 5321 24636 5355
rect 24584 5312 24636 5321
rect 27252 5355 27304 5364
rect 27252 5321 27261 5355
rect 27261 5321 27295 5355
rect 27295 5321 27304 5355
rect 27252 5312 27304 5321
rect 35808 5312 35860 5364
rect 13820 5244 13872 5253
rect 10508 5176 10560 5228
rect 8208 5040 8260 5049
rect 12348 5108 12400 5160
rect 13268 5151 13320 5160
rect 13268 5117 13277 5151
rect 13277 5117 13311 5151
rect 13311 5117 13320 5151
rect 13268 5108 13320 5117
rect 13544 5108 13596 5160
rect 13820 5108 13872 5160
rect 15016 5108 15068 5160
rect 18144 5244 18196 5296
rect 21548 5244 21600 5296
rect 24216 5287 24268 5296
rect 17132 5176 17184 5228
rect 17776 5176 17828 5228
rect 16580 5108 16632 5160
rect 15292 5040 15344 5092
rect 21364 5176 21416 5228
rect 24216 5253 24225 5287
rect 24225 5253 24259 5287
rect 24259 5253 24268 5287
rect 24216 5244 24268 5253
rect 25320 5287 25372 5296
rect 25320 5253 25329 5287
rect 25329 5253 25363 5287
rect 25363 5253 25372 5287
rect 25320 5244 25372 5253
rect 22284 5219 22336 5228
rect 22284 5185 22293 5219
rect 22293 5185 22327 5219
rect 22327 5185 22336 5219
rect 22284 5176 22336 5185
rect 19800 5151 19852 5160
rect 19800 5117 19809 5151
rect 19809 5117 19843 5151
rect 19843 5117 19852 5151
rect 19800 5108 19852 5117
rect 25228 5176 25280 5228
rect 25412 5176 25464 5228
rect 26792 5176 26844 5228
rect 27896 5176 27948 5228
rect 26976 5108 27028 5160
rect 35440 5151 35492 5160
rect 35440 5117 35449 5151
rect 35449 5117 35483 5151
rect 35483 5117 35492 5151
rect 35440 5108 35492 5117
rect 6644 5015 6696 5024
rect 6644 4981 6653 5015
rect 6653 4981 6687 5015
rect 6687 4981 6696 5015
rect 6644 4972 6696 4981
rect 10416 4972 10468 5024
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 15660 4972 15712 5024
rect 16948 4972 17000 5024
rect 18144 4972 18196 5024
rect 19340 5015 19392 5024
rect 19340 4981 19349 5015
rect 19349 4981 19383 5015
rect 19383 4981 19392 5015
rect 19340 4972 19392 4981
rect 20628 5040 20680 5092
rect 21732 5083 21784 5092
rect 21732 5049 21741 5083
rect 21741 5049 21775 5083
rect 21775 5049 21784 5083
rect 21732 5040 21784 5049
rect 22100 5040 22152 5092
rect 24860 5083 24912 5092
rect 24860 5049 24869 5083
rect 24869 5049 24903 5083
rect 24903 5049 24912 5083
rect 24860 5040 24912 5049
rect 27160 5040 27212 5092
rect 21272 4972 21324 5024
rect 22284 4972 22336 5024
rect 22836 4972 22888 5024
rect 23480 5015 23532 5024
rect 23480 4981 23489 5015
rect 23489 4981 23523 5015
rect 23523 4981 23532 5015
rect 23480 4972 23532 4981
rect 26976 5015 27028 5024
rect 26976 4981 26985 5015
rect 26985 4981 27019 5015
rect 27019 4981 27028 5015
rect 26976 4972 27028 4981
rect 27436 4972 27488 5024
rect 28264 5040 28316 5092
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 2228 4768 2280 4820
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 5080 4811 5132 4820
rect 5080 4777 5089 4811
rect 5089 4777 5123 4811
rect 5123 4777 5132 4811
rect 5080 4768 5132 4777
rect 7472 4768 7524 4820
rect 8208 4811 8260 4820
rect 8208 4777 8217 4811
rect 8217 4777 8251 4811
rect 8251 4777 8260 4811
rect 8208 4768 8260 4777
rect 9496 4768 9548 4820
rect 9588 4768 9640 4820
rect 13544 4768 13596 4820
rect 13820 4811 13872 4820
rect 13820 4777 13829 4811
rect 13829 4777 13863 4811
rect 13863 4777 13872 4811
rect 13820 4768 13872 4777
rect 14740 4768 14792 4820
rect 1860 4675 1912 4684
rect 1860 4641 1869 4675
rect 1869 4641 1903 4675
rect 1903 4641 1912 4675
rect 1860 4632 1912 4641
rect 2964 4700 3016 4752
rect 3516 4700 3568 4752
rect 12348 4700 12400 4752
rect 15660 4700 15712 4752
rect 20628 4768 20680 4820
rect 21272 4768 21324 4820
rect 21824 4768 21876 4820
rect 22008 4768 22060 4820
rect 16120 4700 16172 4752
rect 3240 4564 3292 4616
rect 3608 4632 3660 4684
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 5724 4675 5776 4684
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 6460 4675 6512 4684
rect 6460 4641 6469 4675
rect 6469 4641 6503 4675
rect 6503 4641 6512 4675
rect 6460 4632 6512 4641
rect 9772 4675 9824 4684
rect 9772 4641 9781 4675
rect 9781 4641 9815 4675
rect 9815 4641 9824 4675
rect 9772 4632 9824 4641
rect 10416 4675 10468 4684
rect 10416 4641 10425 4675
rect 10425 4641 10459 4675
rect 10459 4641 10468 4675
rect 10416 4632 10468 4641
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 10968 4632 11020 4684
rect 11888 4632 11940 4684
rect 12900 4675 12952 4684
rect 12900 4641 12909 4675
rect 12909 4641 12943 4675
rect 12943 4641 12952 4675
rect 12900 4632 12952 4641
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 13544 4632 13596 4684
rect 13820 4632 13872 4684
rect 16212 4675 16264 4684
rect 16212 4641 16221 4675
rect 16221 4641 16255 4675
rect 16255 4641 16264 4675
rect 16212 4632 16264 4641
rect 18328 4700 18380 4752
rect 19800 4700 19852 4752
rect 20812 4700 20864 4752
rect 21364 4743 21416 4752
rect 21364 4709 21373 4743
rect 21373 4709 21407 4743
rect 21407 4709 21416 4743
rect 21364 4700 21416 4709
rect 21916 4700 21968 4752
rect 17224 4675 17276 4684
rect 17224 4641 17233 4675
rect 17233 4641 17267 4675
rect 17267 4641 17276 4675
rect 17224 4632 17276 4641
rect 4252 4564 4304 4616
rect 8024 4564 8076 4616
rect 18052 4632 18104 4684
rect 4068 4496 4120 4548
rect 12808 4496 12860 4548
rect 16948 4496 17000 4548
rect 18880 4564 18932 4616
rect 18144 4496 18196 4548
rect 18328 4496 18380 4548
rect 19340 4675 19392 4684
rect 19340 4641 19349 4675
rect 19349 4641 19383 4675
rect 19383 4641 19392 4675
rect 19708 4675 19760 4684
rect 19340 4632 19392 4641
rect 19708 4641 19717 4675
rect 19717 4641 19751 4675
rect 19751 4641 19760 4675
rect 19708 4632 19760 4641
rect 20444 4632 20496 4684
rect 21640 4632 21692 4684
rect 23480 4811 23532 4820
rect 23480 4777 23489 4811
rect 23489 4777 23523 4811
rect 23523 4777 23532 4811
rect 23480 4768 23532 4777
rect 23940 4768 23992 4820
rect 24492 4811 24544 4820
rect 24492 4777 24501 4811
rect 24501 4777 24535 4811
rect 24535 4777 24544 4811
rect 24492 4768 24544 4777
rect 24952 4811 25004 4820
rect 24952 4777 24961 4811
rect 24961 4777 24995 4811
rect 24995 4777 25004 4811
rect 24952 4768 25004 4777
rect 25504 4811 25556 4820
rect 25504 4777 25513 4811
rect 25513 4777 25547 4811
rect 25547 4777 25556 4811
rect 25504 4768 25556 4777
rect 26884 4768 26936 4820
rect 24308 4700 24360 4752
rect 25320 4700 25372 4752
rect 27712 4743 27764 4752
rect 22744 4675 22796 4684
rect 22744 4641 22753 4675
rect 22753 4641 22787 4675
rect 22787 4641 22796 4675
rect 22744 4632 22796 4641
rect 22836 4632 22888 4684
rect 23112 4675 23164 4684
rect 23112 4641 23121 4675
rect 23121 4641 23155 4675
rect 23155 4641 23164 4675
rect 23112 4632 23164 4641
rect 27712 4709 27721 4743
rect 27721 4709 27755 4743
rect 27755 4709 27764 4743
rect 27712 4700 27764 4709
rect 28264 4743 28316 4752
rect 28264 4709 28273 4743
rect 28273 4709 28307 4743
rect 28307 4709 28316 4743
rect 28264 4700 28316 4709
rect 30288 4700 30340 4752
rect 29184 4675 29236 4684
rect 22100 4564 22152 4616
rect 23020 4564 23072 4616
rect 29184 4641 29193 4675
rect 29193 4641 29227 4675
rect 29227 4641 29236 4675
rect 29184 4632 29236 4641
rect 31392 4632 31444 4684
rect 24768 4564 24820 4616
rect 27160 4564 27212 4616
rect 28080 4564 28132 4616
rect 26424 4496 26476 4548
rect 9496 4428 9548 4480
rect 9864 4428 9916 4480
rect 11888 4471 11940 4480
rect 11888 4437 11897 4471
rect 11897 4437 11931 4471
rect 11931 4437 11940 4471
rect 11888 4428 11940 4437
rect 14648 4471 14700 4480
rect 14648 4437 14657 4471
rect 14657 4437 14691 4471
rect 14691 4437 14700 4471
rect 14648 4428 14700 4437
rect 26792 4428 26844 4480
rect 27252 4428 27304 4480
rect 29552 4471 29604 4480
rect 29552 4437 29561 4471
rect 29561 4437 29595 4471
rect 29595 4437 29604 4471
rect 29552 4428 29604 4437
rect 30564 4428 30616 4480
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 2136 4224 2188 4276
rect 5172 4224 5224 4276
rect 6184 4224 6236 4276
rect 8024 4156 8076 4208
rect 4344 4088 4396 4140
rect 5080 4088 5132 4140
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 8208 4088 8260 4140
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 3240 4063 3292 4072
rect 3240 4029 3249 4063
rect 3249 4029 3283 4063
rect 3283 4029 3292 4063
rect 3240 4020 3292 4029
rect 4068 4020 4120 4072
rect 8300 4020 8352 4072
rect 3516 3952 3568 4004
rect 4988 3952 5040 4004
rect 5724 3952 5776 4004
rect 8024 3952 8076 4004
rect 1952 3927 2004 3936
rect 1952 3893 1961 3927
rect 1961 3893 1995 3927
rect 1995 3893 2004 3927
rect 1952 3884 2004 3893
rect 2504 3927 2556 3936
rect 2504 3893 2513 3927
rect 2513 3893 2547 3927
rect 2547 3893 2556 3927
rect 2504 3884 2556 3893
rect 4252 3927 4304 3936
rect 4252 3893 4261 3927
rect 4261 3893 4295 3927
rect 4295 3893 4304 3927
rect 4252 3884 4304 3893
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 4804 3884 4856 3936
rect 6460 3884 6512 3936
rect 8208 3927 8260 3936
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 8576 4020 8628 4072
rect 9772 4224 9824 4276
rect 10968 4267 11020 4276
rect 10968 4233 10977 4267
rect 10977 4233 11011 4267
rect 11011 4233 11020 4267
rect 10968 4224 11020 4233
rect 12900 4224 12952 4276
rect 14188 4224 14240 4276
rect 14648 4224 14700 4276
rect 16488 4224 16540 4276
rect 18512 4224 18564 4276
rect 19340 4224 19392 4276
rect 21732 4224 21784 4276
rect 22008 4267 22060 4276
rect 22008 4233 22017 4267
rect 22017 4233 22051 4267
rect 22051 4233 22060 4267
rect 22008 4224 22060 4233
rect 24860 4224 24912 4276
rect 26332 4224 26384 4276
rect 26884 4224 26936 4276
rect 28080 4267 28132 4276
rect 28080 4233 28089 4267
rect 28089 4233 28123 4267
rect 28123 4233 28132 4267
rect 28080 4224 28132 4233
rect 28448 4224 28500 4276
rect 29184 4224 29236 4276
rect 29828 4267 29880 4276
rect 29828 4233 29837 4267
rect 29837 4233 29871 4267
rect 29871 4233 29880 4267
rect 29828 4224 29880 4233
rect 10876 4156 10928 4208
rect 13268 4156 13320 4208
rect 13728 4156 13780 4208
rect 14740 4199 14792 4208
rect 14740 4165 14749 4199
rect 14749 4165 14783 4199
rect 14783 4165 14792 4199
rect 14740 4156 14792 4165
rect 17224 4156 17276 4208
rect 12348 4088 12400 4140
rect 9496 4020 9548 4072
rect 10968 4020 11020 4072
rect 11796 4020 11848 4072
rect 11888 4020 11940 4072
rect 12900 4063 12952 4072
rect 12900 4029 12909 4063
rect 12909 4029 12943 4063
rect 12943 4029 12952 4063
rect 12900 4020 12952 4029
rect 12992 4020 13044 4072
rect 13728 4063 13780 4072
rect 13728 4029 13737 4063
rect 13737 4029 13771 4063
rect 13771 4029 13780 4063
rect 13728 4020 13780 4029
rect 16212 4088 16264 4140
rect 17132 4131 17184 4140
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 16120 4020 16172 4072
rect 16396 4063 16448 4072
rect 16396 4029 16405 4063
rect 16405 4029 16439 4063
rect 16439 4029 16448 4063
rect 16396 4020 16448 4029
rect 16488 4020 16540 4072
rect 16948 4063 17000 4072
rect 16948 4029 16957 4063
rect 16957 4029 16991 4063
rect 16991 4029 17000 4063
rect 16948 4020 17000 4029
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 18328 4020 18380 4072
rect 18788 4063 18840 4072
rect 18788 4029 18797 4063
rect 18797 4029 18831 4063
rect 18831 4029 18840 4063
rect 18788 4020 18840 4029
rect 23020 4088 23072 4140
rect 23480 4088 23532 4140
rect 25320 4088 25372 4140
rect 19064 4063 19116 4072
rect 19064 4029 19073 4063
rect 19073 4029 19107 4063
rect 19107 4029 19116 4063
rect 19064 4020 19116 4029
rect 19708 4020 19760 4072
rect 20352 4063 20404 4072
rect 20352 4029 20361 4063
rect 20361 4029 20395 4063
rect 20395 4029 20404 4063
rect 20352 4020 20404 4029
rect 22100 4063 22152 4072
rect 22100 4029 22109 4063
rect 22109 4029 22143 4063
rect 22143 4029 22152 4063
rect 22100 4020 22152 4029
rect 22284 4020 22336 4072
rect 25964 4088 26016 4140
rect 9588 3884 9640 3936
rect 10600 3884 10652 3936
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 14648 3884 14700 3936
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 18512 3952 18564 4004
rect 22744 3952 22796 4004
rect 23204 3952 23256 4004
rect 25872 4020 25924 4072
rect 26424 4020 26476 4072
rect 17408 3927 17460 3936
rect 17408 3893 17417 3927
rect 17417 3893 17451 3927
rect 17451 3893 17460 3927
rect 17408 3884 17460 3893
rect 17868 3884 17920 3936
rect 18236 3884 18288 3936
rect 19616 3884 19668 3936
rect 21640 3927 21692 3936
rect 21640 3893 21649 3927
rect 21649 3893 21683 3927
rect 21683 3893 21692 3927
rect 21640 3884 21692 3893
rect 22284 3927 22336 3936
rect 22284 3893 22293 3927
rect 22293 3893 22327 3927
rect 22327 3893 22336 3927
rect 22284 3884 22336 3893
rect 23020 3927 23072 3936
rect 23020 3893 23029 3927
rect 23029 3893 23063 3927
rect 23063 3893 23072 3927
rect 23020 3884 23072 3893
rect 24768 3952 24820 4004
rect 24952 3927 25004 3936
rect 24952 3893 24961 3927
rect 24961 3893 24995 3927
rect 24995 3893 25004 3927
rect 27252 3952 27304 4004
rect 27712 3952 27764 4004
rect 25964 3927 26016 3936
rect 24952 3884 25004 3893
rect 25964 3893 25973 3927
rect 25973 3893 26007 3927
rect 26007 3893 26016 3927
rect 25964 3884 26016 3893
rect 27988 3884 28040 3936
rect 29184 4020 29236 4072
rect 29828 4020 29880 4072
rect 31392 4063 31444 4072
rect 31392 4029 31401 4063
rect 31401 4029 31435 4063
rect 31435 4029 31444 4063
rect 31392 4020 31444 4029
rect 30380 3995 30432 4004
rect 30380 3961 30389 3995
rect 30389 3961 30423 3995
rect 30423 3961 30432 3995
rect 30380 3952 30432 3961
rect 31024 3995 31076 4004
rect 31024 3961 31033 3995
rect 31033 3961 31067 3995
rect 31067 3961 31076 3995
rect 31024 3952 31076 3961
rect 32220 3884 32272 3936
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 3792 3680 3844 3732
rect 4988 3680 5040 3732
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 6644 3723 6696 3732
rect 5080 3680 5132 3689
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 9588 3680 9640 3732
rect 9864 3723 9916 3732
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 10600 3680 10652 3732
rect 12992 3680 13044 3732
rect 3240 3612 3292 3664
rect 8484 3612 8536 3664
rect 112 3544 164 3596
rect 2596 3544 2648 3596
rect 3516 3544 3568 3596
rect 5172 3544 5224 3596
rect 5724 3587 5776 3596
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 8668 3587 8720 3596
rect 8668 3553 8677 3587
rect 8677 3553 8711 3587
rect 8711 3553 8720 3587
rect 8668 3544 8720 3553
rect 10140 3587 10192 3596
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 10416 3544 10468 3596
rect 11796 3587 11848 3596
rect 11796 3553 11805 3587
rect 11805 3553 11839 3587
rect 11839 3553 11848 3587
rect 11796 3544 11848 3553
rect 4620 3476 4672 3528
rect 13728 3680 13780 3732
rect 15660 3680 15712 3732
rect 16212 3680 16264 3732
rect 16396 3680 16448 3732
rect 17408 3723 17460 3732
rect 17408 3689 17417 3723
rect 17417 3689 17451 3723
rect 17451 3689 17460 3723
rect 17408 3680 17460 3689
rect 18788 3680 18840 3732
rect 22744 3680 22796 3732
rect 25872 3723 25924 3732
rect 13728 3544 13780 3596
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 16764 3612 16816 3664
rect 20352 3612 20404 3664
rect 21272 3612 21324 3664
rect 21456 3612 21508 3664
rect 22192 3612 22244 3664
rect 24768 3612 24820 3664
rect 25872 3689 25881 3723
rect 25881 3689 25915 3723
rect 25915 3689 25924 3723
rect 25872 3680 25924 3689
rect 27436 3723 27488 3732
rect 27436 3689 27445 3723
rect 27445 3689 27479 3723
rect 27479 3689 27488 3723
rect 27436 3680 27488 3689
rect 28264 3680 28316 3732
rect 30380 3723 30432 3732
rect 25412 3612 25464 3664
rect 26516 3612 26568 3664
rect 27252 3612 27304 3664
rect 30380 3689 30389 3723
rect 30389 3689 30423 3723
rect 30423 3689 30432 3723
rect 30380 3680 30432 3689
rect 28448 3655 28500 3664
rect 28448 3621 28457 3655
rect 28457 3621 28491 3655
rect 28491 3621 28500 3655
rect 28448 3612 28500 3621
rect 30564 3655 30616 3664
rect 30564 3621 30573 3655
rect 30573 3621 30607 3655
rect 30607 3621 30616 3655
rect 30564 3612 30616 3621
rect 30656 3655 30708 3664
rect 30656 3621 30665 3655
rect 30665 3621 30699 3655
rect 30699 3621 30708 3655
rect 30656 3612 30708 3621
rect 8576 3476 8628 3528
rect 1952 3408 2004 3460
rect 2964 3408 3016 3460
rect 9772 3476 9824 3528
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 14648 3476 14700 3528
rect 16304 3476 16356 3528
rect 11152 3408 11204 3460
rect 15200 3408 15252 3460
rect 15936 3408 15988 3460
rect 17960 3587 18012 3596
rect 17960 3553 17969 3587
rect 17969 3553 18003 3587
rect 18003 3553 18012 3587
rect 17960 3544 18012 3553
rect 18512 3587 18564 3596
rect 18512 3553 18521 3587
rect 18521 3553 18555 3587
rect 18555 3553 18564 3587
rect 18512 3544 18564 3553
rect 18880 3587 18932 3596
rect 18880 3553 18889 3587
rect 18889 3553 18923 3587
rect 18923 3553 18932 3587
rect 18880 3544 18932 3553
rect 19708 3544 19760 3596
rect 22008 3587 22060 3596
rect 22008 3553 22017 3587
rect 22017 3553 22051 3587
rect 22051 3553 22060 3587
rect 22008 3544 22060 3553
rect 23204 3587 23256 3596
rect 23204 3553 23213 3587
rect 23213 3553 23247 3587
rect 23247 3553 23256 3587
rect 23204 3544 23256 3553
rect 16764 3476 16816 3528
rect 21364 3476 21416 3528
rect 22284 3476 22336 3528
rect 23112 3476 23164 3528
rect 23388 3544 23440 3596
rect 24676 3544 24728 3596
rect 32220 3587 32272 3596
rect 32220 3553 32229 3587
rect 32229 3553 32263 3587
rect 32263 3553 32272 3587
rect 32220 3544 32272 3553
rect 24492 3476 24544 3528
rect 25228 3519 25280 3528
rect 25228 3485 25237 3519
rect 25237 3485 25271 3519
rect 25271 3485 25280 3519
rect 25228 3476 25280 3485
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 31024 3519 31076 3528
rect 31024 3485 31033 3519
rect 31033 3485 31067 3519
rect 31067 3485 31076 3519
rect 31024 3476 31076 3485
rect 18236 3408 18288 3460
rect 14924 3340 14976 3392
rect 15568 3383 15620 3392
rect 15568 3349 15577 3383
rect 15577 3349 15611 3383
rect 15611 3349 15620 3383
rect 15568 3340 15620 3349
rect 19708 3383 19760 3392
rect 19708 3349 19717 3383
rect 19717 3349 19751 3383
rect 19751 3349 19760 3383
rect 19708 3340 19760 3349
rect 20628 3383 20680 3392
rect 20628 3349 20637 3383
rect 20637 3349 20671 3383
rect 20671 3349 20680 3383
rect 20628 3340 20680 3349
rect 21732 3340 21784 3392
rect 22192 3340 22244 3392
rect 23664 3340 23716 3392
rect 26240 3383 26292 3392
rect 26240 3349 26249 3383
rect 26249 3349 26283 3383
rect 26283 3349 26292 3383
rect 26240 3340 26292 3349
rect 29276 3383 29328 3392
rect 29276 3349 29285 3383
rect 29285 3349 29319 3383
rect 29319 3349 29328 3383
rect 29276 3340 29328 3349
rect 32496 3340 32548 3392
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 4620 3136 4672 3188
rect 6184 3136 6236 3188
rect 6460 3136 6512 3188
rect 11888 3136 11940 3188
rect 17960 3136 18012 3188
rect 19708 3136 19760 3188
rect 21732 3136 21784 3188
rect 23940 3136 23992 3188
rect 25412 3179 25464 3188
rect 25412 3145 25421 3179
rect 25421 3145 25455 3179
rect 25455 3145 25464 3179
rect 25412 3136 25464 3145
rect 28448 3136 28500 3188
rect 30656 3136 30708 3188
rect 32220 3179 32272 3188
rect 32220 3145 32229 3179
rect 32229 3145 32263 3179
rect 32263 3145 32272 3179
rect 32220 3136 32272 3145
rect 1860 2932 1912 2984
rect 2964 2975 3016 2984
rect 2964 2941 2973 2975
rect 2973 2941 3007 2975
rect 3007 2941 3016 2975
rect 2964 2932 3016 2941
rect 3516 3068 3568 3120
rect 8024 3068 8076 3120
rect 13728 3111 13780 3120
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 5172 3000 5224 3052
rect 7840 3000 7892 3052
rect 3424 2932 3476 2984
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 4804 2932 4856 2984
rect 1952 2864 2004 2916
rect 7012 2975 7064 2984
rect 7012 2941 7021 2975
rect 7021 2941 7055 2975
rect 7055 2941 7064 2975
rect 7012 2932 7064 2941
rect 8208 3000 8260 3052
rect 8484 2975 8536 2984
rect 8484 2941 8493 2975
rect 8493 2941 8527 2975
rect 8527 2941 8536 2975
rect 8484 2932 8536 2941
rect 8576 2932 8628 2984
rect 13728 3077 13737 3111
rect 13737 3077 13771 3111
rect 13771 3077 13780 3111
rect 13728 3068 13780 3077
rect 13912 3068 13964 3120
rect 15292 3068 15344 3120
rect 15568 3068 15620 3120
rect 10876 3000 10928 3052
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 12440 3000 12492 3009
rect 14004 3000 14056 3052
rect 15936 3043 15988 3052
rect 7564 2864 7616 2916
rect 9496 2932 9548 2984
rect 11152 2975 11204 2984
rect 11152 2941 11161 2975
rect 11161 2941 11195 2975
rect 11195 2941 11204 2975
rect 11152 2932 11204 2941
rect 11796 2932 11848 2984
rect 12348 2932 12400 2984
rect 10968 2907 11020 2916
rect 10968 2873 10977 2907
rect 10977 2873 11011 2907
rect 11011 2873 11020 2907
rect 10968 2864 11020 2873
rect 2596 2839 2648 2848
rect 2596 2805 2605 2839
rect 2605 2805 2639 2839
rect 2639 2805 2648 2839
rect 2596 2796 2648 2805
rect 5448 2839 5500 2848
rect 5448 2805 5457 2839
rect 5457 2805 5491 2839
rect 5491 2805 5500 2839
rect 5448 2796 5500 2805
rect 7932 2839 7984 2848
rect 7932 2805 7941 2839
rect 7941 2805 7975 2839
rect 7975 2805 7984 2839
rect 7932 2796 7984 2805
rect 8116 2839 8168 2848
rect 8116 2805 8125 2839
rect 8125 2805 8159 2839
rect 8159 2805 8168 2839
rect 8116 2796 8168 2805
rect 8668 2796 8720 2848
rect 10416 2796 10468 2848
rect 14648 2932 14700 2984
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 19340 3068 19392 3120
rect 22192 3068 22244 3120
rect 26424 3068 26476 3120
rect 27436 3068 27488 3120
rect 16212 2932 16264 2984
rect 16580 2975 16632 2984
rect 16580 2941 16589 2975
rect 16589 2941 16623 2975
rect 16623 2941 16632 2975
rect 16580 2932 16632 2941
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 19064 2975 19116 2984
rect 19064 2941 19073 2975
rect 19073 2941 19107 2975
rect 19107 2941 19116 2975
rect 19064 2932 19116 2941
rect 19708 2932 19760 2984
rect 20996 2932 21048 2984
rect 22008 3000 22060 3052
rect 21732 2975 21784 2984
rect 21732 2941 21741 2975
rect 21741 2941 21775 2975
rect 21775 2941 21784 2975
rect 21732 2932 21784 2941
rect 21824 2932 21876 2984
rect 26516 3000 26568 3052
rect 27988 3000 28040 3052
rect 14924 2864 14976 2916
rect 15108 2907 15160 2916
rect 15108 2873 15117 2907
rect 15117 2873 15151 2907
rect 15151 2873 15160 2907
rect 15108 2864 15160 2873
rect 23296 2932 23348 2984
rect 23664 2975 23716 2984
rect 23664 2941 23673 2975
rect 23673 2941 23707 2975
rect 23707 2941 23716 2975
rect 23664 2932 23716 2941
rect 23940 2932 23992 2984
rect 24124 2975 24176 2984
rect 24124 2941 24133 2975
rect 24133 2941 24167 2975
rect 24167 2941 24176 2975
rect 24124 2932 24176 2941
rect 24492 2975 24544 2984
rect 24492 2941 24501 2975
rect 24501 2941 24535 2975
rect 24535 2941 24544 2975
rect 24492 2932 24544 2941
rect 24676 2932 24728 2984
rect 26240 2975 26292 2984
rect 26240 2941 26249 2975
rect 26249 2941 26283 2975
rect 26283 2941 26292 2975
rect 26240 2932 26292 2941
rect 32036 3000 32088 3052
rect 24952 2864 25004 2916
rect 30932 2907 30984 2916
rect 30932 2873 30941 2907
rect 30941 2873 30975 2907
rect 30975 2873 30984 2907
rect 30932 2864 30984 2873
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 18696 2796 18748 2848
rect 23204 2796 23256 2848
rect 23388 2796 23440 2848
rect 26148 2839 26200 2848
rect 26148 2805 26157 2839
rect 26157 2805 26191 2839
rect 26191 2805 26200 2839
rect 26148 2796 26200 2805
rect 27436 2839 27488 2848
rect 27436 2805 27445 2839
rect 27445 2805 27479 2839
rect 27479 2805 27488 2839
rect 27436 2796 27488 2805
rect 28080 2839 28132 2848
rect 28080 2805 28089 2839
rect 28089 2805 28123 2839
rect 28123 2805 28132 2839
rect 28080 2796 28132 2805
rect 31116 2864 31168 2916
rect 32496 2907 32548 2916
rect 32496 2873 32505 2907
rect 32505 2873 32539 2907
rect 32539 2873 32548 2907
rect 32496 2864 32548 2873
rect 32680 2864 32732 2916
rect 31208 2796 31260 2848
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 2964 2592 3016 2644
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 3424 2524 3476 2576
rect 6092 2592 6144 2644
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 7840 2635 7892 2644
rect 7840 2601 7849 2635
rect 7849 2601 7883 2635
rect 7883 2601 7892 2635
rect 7840 2592 7892 2601
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 8852 2635 8904 2644
rect 8852 2601 8861 2635
rect 8861 2601 8895 2635
rect 8895 2601 8904 2635
rect 8852 2592 8904 2601
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 12808 2635 12860 2644
rect 12808 2601 12817 2635
rect 12817 2601 12851 2635
rect 12851 2601 12860 2635
rect 12808 2592 12860 2601
rect 14004 2592 14056 2644
rect 14924 2635 14976 2644
rect 14924 2601 14933 2635
rect 14933 2601 14967 2635
rect 14967 2601 14976 2635
rect 14924 2592 14976 2601
rect 15292 2635 15344 2644
rect 15292 2601 15301 2635
rect 15301 2601 15335 2635
rect 15335 2601 15344 2635
rect 15292 2592 15344 2601
rect 15660 2635 15712 2644
rect 15660 2601 15669 2635
rect 15669 2601 15703 2635
rect 15703 2601 15712 2635
rect 15660 2592 15712 2601
rect 5448 2524 5500 2576
rect 3516 2456 3568 2508
rect 7932 2456 7984 2508
rect 10416 2456 10468 2508
rect 10508 2456 10560 2508
rect 13728 2456 13780 2508
rect 13820 2499 13872 2508
rect 13820 2465 13829 2499
rect 13829 2465 13863 2499
rect 13863 2465 13872 2499
rect 13820 2456 13872 2465
rect 15108 2456 15160 2508
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 19340 2592 19392 2644
rect 20628 2635 20680 2644
rect 20628 2601 20637 2635
rect 20637 2601 20671 2635
rect 20671 2601 20680 2635
rect 20628 2592 20680 2601
rect 20996 2635 21048 2644
rect 20996 2601 21005 2635
rect 21005 2601 21039 2635
rect 21039 2601 21048 2635
rect 20996 2592 21048 2601
rect 16304 2567 16356 2576
rect 16304 2533 16313 2567
rect 16313 2533 16347 2567
rect 16347 2533 16356 2567
rect 16304 2524 16356 2533
rect 16856 2567 16908 2576
rect 16856 2533 16865 2567
rect 16865 2533 16899 2567
rect 16899 2533 16908 2567
rect 16856 2524 16908 2533
rect 10968 2388 11020 2440
rect 8668 2320 8720 2372
rect 13820 2320 13872 2372
rect 14096 2388 14148 2440
rect 14280 2431 14332 2440
rect 14280 2397 14289 2431
rect 14289 2397 14323 2431
rect 14323 2397 14332 2431
rect 16764 2431 16816 2440
rect 14280 2388 14332 2397
rect 16764 2397 16773 2431
rect 16773 2397 16807 2431
rect 16807 2397 16816 2431
rect 16764 2388 16816 2397
rect 23020 2592 23072 2644
rect 24124 2592 24176 2644
rect 26148 2635 26200 2644
rect 26148 2601 26157 2635
rect 26157 2601 26191 2635
rect 26191 2601 26200 2635
rect 26148 2592 26200 2601
rect 27252 2635 27304 2644
rect 27252 2601 27261 2635
rect 27261 2601 27295 2635
rect 27295 2601 27304 2635
rect 27252 2592 27304 2601
rect 28080 2592 28132 2644
rect 29552 2635 29604 2644
rect 21732 2524 21784 2576
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 21456 2456 21508 2508
rect 22008 2456 22060 2508
rect 26240 2524 26292 2576
rect 29552 2601 29561 2635
rect 29561 2601 29595 2635
rect 29595 2601 29604 2635
rect 32036 2635 32088 2644
rect 29552 2592 29604 2601
rect 30932 2524 30984 2576
rect 31852 2524 31904 2576
rect 23020 2499 23072 2508
rect 20628 2388 20680 2440
rect 22284 2388 22336 2440
rect 23020 2465 23029 2499
rect 23029 2465 23063 2499
rect 23063 2465 23072 2499
rect 23020 2456 23072 2465
rect 23664 2456 23716 2508
rect 24124 2456 24176 2508
rect 24952 2499 25004 2508
rect 24952 2465 24961 2499
rect 24961 2465 24995 2499
rect 24995 2465 25004 2499
rect 24952 2456 25004 2465
rect 27436 2456 27488 2508
rect 32036 2601 32045 2635
rect 32045 2601 32079 2635
rect 32079 2601 32088 2635
rect 32036 2592 32088 2601
rect 32128 2524 32180 2576
rect 32680 2499 32732 2508
rect 32680 2465 32689 2499
rect 32689 2465 32723 2499
rect 32723 2465 32732 2499
rect 32680 2456 32732 2465
rect 10508 2295 10560 2304
rect 10508 2261 10517 2295
rect 10517 2261 10551 2295
rect 10551 2261 10560 2295
rect 10508 2252 10560 2261
rect 14924 2252 14976 2304
rect 22100 2320 22152 2372
rect 24952 2320 25004 2372
rect 29276 2388 29328 2440
rect 31208 2388 31260 2440
rect 22008 2252 22060 2304
rect 23664 2252 23716 2304
rect 30748 2252 30800 2304
rect 34152 2320 34204 2372
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
rect 1676 2048 1728 2100
rect 10508 2048 10560 2100
<< metal2 >>
rect 5816 15564 5868 15570
rect 6642 15564 6698 16000
rect 6642 15520 6644 15564
rect 5816 15506 5868 15512
rect 6696 15520 6698 15564
rect 19982 15564 20038 16000
rect 33322 15586 33378 16000
rect 19982 15520 19984 15564
rect 6644 15506 6696 15512
rect 20036 15520 20038 15564
rect 20628 15564 20680 15570
rect 19984 15506 20036 15512
rect 33322 15558 33456 15586
rect 33322 15520 33378 15558
rect 20628 15506 20680 15512
rect 1214 15056 1270 15065
rect 1214 14991 1270 15000
rect 18 13832 74 13841
rect 18 13767 74 13776
rect 32 6458 60 13767
rect 1030 12336 1086 12345
rect 1030 12271 1086 12280
rect 20 6452 72 6458
rect 20 6394 72 6400
rect 1044 5370 1072 12271
rect 1228 8634 1256 14991
rect 1490 14240 1546 14249
rect 1490 14175 1546 14184
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 10470 1440 11154
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1216 8628 1268 8634
rect 1216 8570 1268 8576
rect 1504 7546 1532 14175
rect 1582 11520 1638 11529
rect 1582 11455 1638 11464
rect 1596 11354 1624 11455
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1582 10568 1638 10577
rect 1582 10503 1638 10512
rect 1596 10266 1624 10503
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1596 9178 1624 9687
rect 1688 9382 1716 10066
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1688 8945 1716 9318
rect 2240 9042 2268 10406
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 1674 8936 1730 8945
rect 1674 8871 1730 8880
rect 1582 8800 1638 8809
rect 1582 8735 1638 8744
rect 1596 8090 1624 8735
rect 2148 8294 2176 8978
rect 3344 8294 3372 8978
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 2136 8288 2188 8294
rect 2136 8230 2188 8236
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1688 6662 1716 7278
rect 2056 7274 2084 7890
rect 2148 7313 2176 8230
rect 2686 8120 2742 8129
rect 2686 8055 2742 8064
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2516 7478 2544 7890
rect 2700 7818 2728 8055
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2134 7304 2190 7313
rect 2044 7268 2096 7274
rect 2134 7239 2190 7248
rect 2044 7210 2096 7216
rect 2056 7177 2084 7210
rect 2042 7168 2098 7177
rect 2042 7103 2098 7112
rect 2412 6928 2464 6934
rect 2042 6896 2098 6905
rect 2412 6870 2464 6876
rect 2042 6831 2098 6840
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1688 6089 1716 6598
rect 2056 6458 2084 6831
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2056 6254 2084 6394
rect 2424 6390 2452 6870
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2412 6384 2464 6390
rect 2318 6352 2374 6361
rect 2412 6326 2464 6332
rect 2318 6287 2374 6296
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 1674 6080 1730 6089
rect 1674 6015 1730 6024
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 1032 5364 1084 5370
rect 1032 5306 1084 5312
rect 1780 5234 1808 5510
rect 2042 5264 2098 5273
rect 1768 5228 1820 5234
rect 2042 5199 2098 5208
rect 1768 5170 1820 5176
rect 2056 5166 2084 5199
rect 2148 5166 2176 5510
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 110 4040 166 4049
rect 110 3975 166 3984
rect 124 3602 152 3975
rect 112 3596 164 3602
rect 112 3538 164 3544
rect 1872 2990 1900 4626
rect 2148 4282 2176 5102
rect 2240 4826 2268 5646
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1964 3466 1992 3878
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 1964 2922 1992 3402
rect 1952 2916 2004 2922
rect 1952 2858 2004 2864
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 1688 82 1716 2042
rect 2332 785 2360 6287
rect 2424 5846 2452 6326
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 2424 5370 2452 5782
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2516 3942 2544 6598
rect 2608 6254 2636 6666
rect 2976 6361 3004 8230
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3160 7274 3188 7686
rect 3344 7449 3372 8230
rect 3330 7440 3386 7449
rect 3240 7404 3292 7410
rect 3330 7375 3386 7384
rect 3240 7346 3292 7352
rect 3252 7274 3280 7346
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3252 6458 3280 7210
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 2962 6352 3018 6361
rect 2962 6287 3018 6296
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2608 5030 2636 6190
rect 3436 6186 3464 8298
rect 4080 8265 4108 8366
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4066 8256 4122 8265
rect 4066 8191 4122 8200
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4172 7478 4200 7958
rect 4356 7886 4384 8298
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4356 7546 4384 7822
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 5166 3096 5510
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2964 4752 3016 4758
rect 3068 4740 3096 5102
rect 3016 4712 3096 4740
rect 2964 4694 3016 4700
rect 3068 4078 3096 4712
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3252 4078 3280 4558
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 3252 3670 3280 4014
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2608 2854 2636 3538
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2976 2990 3004 3402
rect 3436 2990 3464 5102
rect 3528 4758 3556 7142
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 3620 4690 3648 7414
rect 4528 7268 4580 7274
rect 4580 7228 4660 7256
rect 4528 7210 4580 7216
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3804 5574 3832 6734
rect 4080 6662 4108 7142
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6458 4108 6598
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4080 6118 4108 6394
rect 4264 6390 4292 6870
rect 4632 6798 4660 7228
rect 4816 6934 4844 8230
rect 5000 8090 5028 8774
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 4988 8084 5040 8090
rect 4908 8044 4988 8072
rect 4908 7478 4936 8044
rect 4988 8026 5040 8032
rect 5092 7993 5120 8230
rect 5828 8090 5856 15506
rect 6656 15475 6684 15506
rect 19996 15475 20024 15506
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 16762 10024 16818 10033
rect 16762 9959 16818 9968
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5078 7984 5134 7993
rect 5078 7919 5134 7928
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 5000 7410 5028 7822
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4264 5914 4292 6326
rect 4356 6322 4384 6598
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4448 5914 4476 6394
rect 4632 6322 4660 6734
rect 5000 6730 5028 7346
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 4988 6724 5040 6730
rect 4988 6666 5040 6672
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 3528 3602 3556 3946
rect 3804 3738 3832 5510
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4080 4554 4108 5102
rect 4448 5030 4476 5850
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4540 4826 4568 5646
rect 4528 4820 4580 4826
rect 4172 4780 4528 4808
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 4080 4078 4108 4490
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3528 3505 3556 3538
rect 3514 3496 3570 3505
rect 3514 3431 3570 3440
rect 3528 3126 3556 3431
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2608 2417 2636 2790
rect 2976 2650 3004 2926
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3436 2582 3464 2926
rect 3528 2650 3556 3062
rect 4080 2990 4108 4014
rect 4172 3058 4200 4780
rect 4528 4762 4580 4768
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 3942 4292 4558
rect 4632 4154 4660 6258
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 4356 4146 4660 4154
rect 4344 4140 4660 4146
rect 4396 4126 4660 4140
rect 4344 4082 4396 4088
rect 5000 4010 5028 5510
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5092 4826 5120 5102
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5184 4690 5212 5034
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5184 4282 5212 4626
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 3528 2514 3556 2586
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 2594 2408 2650 2417
rect 2594 2343 2650 2352
rect 2318 776 2374 785
rect 2318 711 2374 720
rect 1766 82 1822 480
rect 4264 377 4292 3878
rect 4632 3534 4660 3878
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4632 3194 4660 3470
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4816 2990 4844 3878
rect 5000 3738 5028 3946
rect 5092 3738 5120 4082
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5184 3602 5212 4218
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5184 3058 5212 3538
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 5368 2825 5396 7278
rect 5460 7206 5488 7890
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 13634 7848 13690 7857
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 9968 7206 9996 7822
rect 13634 7783 13690 7792
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 5460 4146 5488 7142
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 5736 6458 5764 6870
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5828 6390 5856 6870
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 6932 6322 6960 6734
rect 7208 6322 7236 7142
rect 9968 6905 9996 7142
rect 10336 6934 10364 7686
rect 13648 7342 13676 7783
rect 10692 7336 10744 7342
rect 13636 7336 13688 7342
rect 10692 7278 10744 7284
rect 12530 7304 12586 7313
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10324 6928 10376 6934
rect 9954 6896 10010 6905
rect 10324 6870 10376 6876
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 9954 6831 10010 6840
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 8588 6458 8616 6734
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6288 5098 6316 5850
rect 6564 5370 6592 6054
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 6656 5030 6684 5646
rect 7208 5642 7236 6258
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9140 5914 9168 6122
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7392 5370 7420 5646
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5736 4010 5764 4626
rect 6196 4282 6224 4626
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5736 3602 5764 3946
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 5448 2848 5500 2854
rect 5354 2816 5410 2825
rect 5448 2790 5500 2796
rect 5354 2751 5410 2760
rect 5460 2582 5488 2790
rect 6104 2650 6132 3538
rect 6196 3194 6224 4218
rect 6472 3942 6500 4626
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6472 3602 6500 3878
rect 6656 3738 6684 4966
rect 7484 4826 7512 5850
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 8128 5234 8156 5510
rect 9140 5370 9168 5850
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 8036 4214 8064 4558
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6472 3194 6500 3538
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 8036 3126 8064 3946
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 5448 2576 5500 2582
rect 7024 2553 7052 2926
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7576 2650 7604 2858
rect 7852 2650 7880 2994
rect 8128 2854 8156 5170
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 8220 4826 8248 5034
rect 9508 4826 9536 6122
rect 9968 5681 9996 6831
rect 10336 5914 10364 6870
rect 10428 6458 10456 6870
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10428 5846 10456 6394
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 9954 5672 10010 5681
rect 9954 5607 10010 5616
rect 10428 5370 10456 5782
rect 10520 5710 10548 7142
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10612 6322 10640 6666
rect 10704 6633 10732 7278
rect 14200 7313 14228 7890
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14476 7410 14504 7686
rect 16776 7546 16804 9959
rect 18602 9072 18658 9081
rect 18602 9007 18658 9016
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 13636 7278 13688 7284
rect 14186 7304 14242 7313
rect 12530 7239 12586 7248
rect 12544 6866 12572 7239
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 10690 6624 10746 6633
rect 10690 6559 10746 6568
rect 12544 6390 12572 6802
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10520 5234 10548 5646
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 12360 5166 12388 5510
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 9600 4826 9628 5102
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 8208 4820 8260 4826
rect 9496 4820 9548 4826
rect 8260 4780 8340 4808
rect 8208 4762 8260 4768
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8220 3942 8248 4082
rect 8312 4078 8340 4780
rect 9496 4762 9548 4768
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 10428 4690 10456 4966
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9508 4078 9536 4422
rect 9784 4282 9812 4626
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 8300 4072 8352 4078
rect 8576 4072 8628 4078
rect 8300 4014 8352 4020
rect 8496 4032 8576 4060
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8220 3058 8248 3878
rect 8496 3670 8524 4032
rect 8576 4014 8628 4020
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8496 2990 8524 3606
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8588 2990 8616 3470
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 5448 2518 5500 2524
rect 7010 2544 7066 2553
rect 4250 368 4306 377
rect 4250 303 4306 312
rect 1688 54 1822 82
rect 1766 0 1822 54
rect 5354 82 5410 480
rect 5460 82 5488 2518
rect 7944 2514 7972 2790
rect 8496 2650 8524 2926
rect 8680 2854 8708 3538
rect 8850 3360 8906 3369
rect 8850 3295 8906 3304
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 7010 2479 7066 2488
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8680 2378 8708 2790
rect 8864 2650 8892 3295
rect 9508 2990 9536 4014
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9600 3738 9628 3878
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9784 3534 9812 4218
rect 9876 3738 9904 4422
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 10428 3602 10456 4626
rect 10612 3942 10640 4626
rect 10980 4282 11008 4626
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3738 10640 3878
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 9772 3528 9824 3534
rect 10152 3505 10180 3538
rect 9772 3470 9824 3476
rect 10138 3496 10194 3505
rect 10138 3431 10194 3440
rect 10888 3058 10916 4150
rect 10980 4078 11008 4218
rect 11808 4078 11836 4966
rect 12360 4758 12388 5102
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11900 4486 11928 4626
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4078 11928 4422
rect 12360 4146 12388 4694
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11808 3942 11836 4014
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11518 3632 11574 3641
rect 11808 3602 11836 3878
rect 11518 3567 11574 3576
rect 11796 3596 11848 3602
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 11164 2990 11192 3402
rect 11532 3058 11560 3567
rect 11796 3538 11848 3544
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11808 2990 11836 3538
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11900 3194 11928 3470
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 12452 3058 12480 6190
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12636 5778 12664 6054
rect 13556 5846 13584 6122
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13280 5166 13308 5714
rect 13556 5370 13584 5782
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13280 4690 13308 5102
rect 13556 4826 13584 5102
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13556 4690 13584 4762
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 12808 4548 12860 4554
rect 12808 4490 12860 4496
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 10428 2514 10456 2790
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 10508 2508 10560 2514
rect 10508 2450 10560 2456
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 5354 54 5488 82
rect 8680 82 8708 2314
rect 10520 2310 10548 2450
rect 10980 2446 11008 2858
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10520 2106 10548 2246
rect 10508 2100 10560 2106
rect 10508 2042 10560 2048
rect 9034 82 9090 480
rect 8680 54 9090 82
rect 12360 82 12388 2926
rect 12452 2650 12480 2994
rect 12820 2650 12848 4490
rect 12912 4282 12940 4626
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12912 4078 12940 4218
rect 13280 4214 13308 4626
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 13004 3738 13032 4014
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 13648 1193 13676 7278
rect 14186 7239 14242 7248
rect 14832 7268 14884 7274
rect 14200 7206 14228 7239
rect 14832 7210 14884 7216
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14004 6928 14056 6934
rect 14004 6870 14056 6876
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 6254 13860 6598
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13740 4214 13768 5646
rect 13832 5302 13860 6190
rect 14016 5914 14044 6870
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14384 6390 14412 6734
rect 14844 6662 14872 7210
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14844 6186 14872 6598
rect 14936 6322 14964 7346
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15120 6322 15148 6598
rect 15212 6458 15240 7278
rect 15396 6798 15424 7414
rect 16394 7304 16450 7313
rect 16394 7239 16450 7248
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14752 5846 14780 6054
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 15212 5574 15240 6394
rect 15396 6118 15424 6734
rect 15488 6458 15516 6870
rect 15580 6798 15608 7142
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15580 5710 15608 6734
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 15028 5166 15056 5510
rect 15672 5370 15700 6122
rect 16408 5953 16436 7239
rect 18326 6896 18382 6905
rect 16764 6860 16816 6866
rect 18326 6831 18328 6840
rect 16764 6802 16816 6808
rect 18380 6831 18382 6840
rect 18328 6802 18380 6808
rect 16776 6118 16804 6802
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16394 5944 16450 5953
rect 16394 5879 16450 5888
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 13832 4826 13860 5102
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13728 4072 13780 4078
rect 13832 4060 13860 4626
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14660 4282 14688 4422
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 13780 4032 13860 4060
rect 13728 4014 13780 4020
rect 13740 3738 13768 4014
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13740 3126 13768 3538
rect 14200 3369 14228 4218
rect 14752 4214 14780 4762
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 14660 3534 14688 3878
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14186 3360 14242 3369
rect 14186 3295 14242 3304
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 13740 2514 13768 3062
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13820 2508 13872 2514
rect 13924 2496 13952 3062
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14016 2650 14044 2994
rect 14660 2990 14688 3470
rect 15212 3466 15240 3878
rect 15304 3602 15332 5034
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 15672 4758 15700 4966
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16132 4078 16160 4694
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16224 4146 16252 4626
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16224 3738 16252 4082
rect 16500 4078 16528 4218
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16408 3738 16436 4014
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14936 2922 14964 3334
rect 15304 3126 15332 3538
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15580 3126 15608 3334
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 14936 2650 14964 2858
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 13872 2468 13952 2496
rect 14278 2544 14334 2553
rect 14278 2479 14334 2488
rect 13820 2450 13872 2456
rect 13740 2258 13768 2450
rect 13832 2378 13860 2450
rect 14292 2446 14320 2479
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 14108 2258 14136 2382
rect 14936 2310 14964 2586
rect 15120 2514 15148 2858
rect 15304 2650 15332 3062
rect 15672 2650 15700 3674
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15948 3058 15976 3402
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 13740 2230 14136 2258
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 13634 1184 13690 1193
rect 13634 1119 13690 1128
rect 12622 82 12678 480
rect 12360 54 12678 82
rect 16224 82 16252 2926
rect 16316 2582 16344 3470
rect 16592 2990 16620 5102
rect 16776 3670 16804 6054
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16304 2576 16356 2582
rect 16304 2518 16356 2524
rect 16776 2446 16804 3470
rect 16868 2582 16896 5510
rect 16960 5030 16988 6598
rect 18340 6458 18368 6802
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18340 6361 18368 6394
rect 18326 6352 18382 6361
rect 18326 6287 18382 6296
rect 18616 6254 18644 9007
rect 20442 8936 20498 8945
rect 20442 8871 20498 8880
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 19154 7848 19210 7857
rect 19154 7783 19210 7792
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18788 6792 18840 6798
rect 18892 6769 18920 7278
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 18788 6734 18840 6740
rect 18878 6760 18934 6769
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 17500 6248 17552 6254
rect 17498 6216 17500 6225
rect 18604 6248 18656 6254
rect 17552 6216 17554 6225
rect 18604 6190 18656 6196
rect 17498 6151 17554 6160
rect 17512 6118 17540 6151
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17512 5817 17540 6054
rect 17498 5808 17554 5817
rect 17498 5743 17554 5752
rect 17788 5234 17816 6054
rect 18144 5840 18196 5846
rect 18144 5782 18196 5788
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16960 4554 16988 4966
rect 16948 4548 17000 4554
rect 16948 4490 17000 4496
rect 16960 4078 16988 4490
rect 17144 4146 17172 5170
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 17236 4214 17264 4626
rect 17224 4208 17276 4214
rect 17224 4150 17276 4156
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 17880 3942 17908 5510
rect 18156 5302 18184 5782
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 18156 5030 18184 5238
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18064 4078 18092 4626
rect 18156 4554 18184 4966
rect 18328 4752 18380 4758
rect 18328 4694 18380 4700
rect 18340 4554 18368 4694
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 18328 4548 18380 4554
rect 18328 4490 18380 4496
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17420 3738 17448 3878
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17972 3194 18000 3538
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18064 2990 18092 4014
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 18156 2650 18184 4490
rect 18340 4078 18368 4490
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18524 4010 18552 4218
rect 18616 4049 18644 6190
rect 18602 4040 18658 4049
rect 18512 4004 18564 4010
rect 18602 3975 18658 3984
rect 18512 3946 18564 3952
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3466 18276 3878
rect 18524 3602 18552 3946
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 18708 2854 18736 6598
rect 18800 6458 18828 6734
rect 18984 6730 19012 7142
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 18878 6695 18934 6704
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18984 6322 19012 6666
rect 19076 6662 19104 6870
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18972 6112 19024 6118
rect 19076 6100 19104 6598
rect 19168 6497 19196 7783
rect 19628 7206 19656 7890
rect 19984 7336 20036 7342
rect 20168 7336 20220 7342
rect 20036 7313 20116 7324
rect 20036 7304 20130 7313
rect 20036 7296 20074 7304
rect 19984 7278 20036 7284
rect 20168 7278 20220 7284
rect 20074 7239 20130 7248
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19154 6488 19210 6497
rect 19154 6423 19210 6432
rect 19024 6072 19104 6100
rect 18972 6054 19024 6060
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 18892 4622 18920 5510
rect 18984 5370 19012 6054
rect 19352 5846 19380 6598
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19352 4690 19380 4966
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 18880 4616 18932 4622
rect 18880 4558 18932 4564
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18800 3738 18828 4014
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18892 3602 18920 4558
rect 19352 4282 19380 4626
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 19076 2990 19104 4014
rect 19352 3126 19380 4218
rect 19628 3942 19656 7142
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19996 5778 20024 6666
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19812 4758 19840 5102
rect 19800 4752 19852 4758
rect 19800 4694 19852 4700
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 19720 4078 19748 4626
rect 20180 4154 20208 7278
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20364 6662 20392 7142
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20088 4126 20208 4154
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 18340 2514 18368 2790
rect 19352 2650 19380 3062
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16302 82 16358 480
rect 16224 54 16358 82
rect 19628 82 19656 3878
rect 19720 3602 19748 4014
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 19720 3398 19748 3538
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19720 3194 19748 3334
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 19720 2990 19748 3130
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 20088 1601 20116 4126
rect 20364 4078 20392 5510
rect 20456 4690 20484 8871
rect 20640 7002 20668 15506
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 29828 10464 29880 10470
rect 29828 10406 29880 10412
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 24214 7984 24270 7993
rect 24214 7919 24270 7928
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21362 7440 21418 7449
rect 21362 7375 21418 7384
rect 21272 7268 21324 7274
rect 21272 7210 21324 7216
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20720 6928 20772 6934
rect 20720 6870 20772 6876
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20548 5846 20576 6122
rect 20732 6118 20760 6870
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20824 6322 20852 6734
rect 20916 6730 20944 7142
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21284 6458 21312 7210
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20640 5098 20668 5646
rect 20732 5370 20760 6054
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20628 5092 20680 5098
rect 20628 5034 20680 5040
rect 20640 4826 20668 5034
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20824 4758 20852 6258
rect 21088 6180 21140 6186
rect 21284 6168 21312 6394
rect 21140 6140 21312 6168
rect 21088 6122 21140 6128
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 21284 5030 21312 5850
rect 21376 5409 21404 7375
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21560 6390 21588 6666
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21362 5400 21418 5409
rect 21362 5335 21418 5344
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 20812 4752 20864 4758
rect 20812 4694 20864 4700
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20364 3670 20392 4014
rect 21284 3670 21312 4762
rect 21376 4758 21404 5170
rect 21364 4752 21416 4758
rect 21364 4694 21416 4700
rect 21468 4154 21496 5646
rect 21560 5302 21588 6326
rect 21824 5568 21876 5574
rect 21824 5510 21876 5516
rect 21548 5296 21600 5302
rect 21548 5238 21600 5244
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 21640 4684 21692 4690
rect 21640 4626 21692 4632
rect 21376 4126 21496 4154
rect 20352 3664 20404 3670
rect 20352 3606 20404 3612
rect 21272 3664 21324 3670
rect 21272 3606 21324 3612
rect 21376 3534 21404 4126
rect 21652 3942 21680 4626
rect 21744 4282 21772 5034
rect 21836 4826 21864 5510
rect 22020 4826 22048 7686
rect 22374 7576 22430 7585
rect 22374 7511 22430 7520
rect 22388 6769 22416 7511
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22374 6760 22430 6769
rect 22374 6695 22430 6704
rect 22388 6322 22416 6695
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22572 5846 22600 6054
rect 22560 5840 22612 5846
rect 22560 5782 22612 5788
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 22284 5568 22336 5574
rect 22284 5510 22336 5516
rect 22112 5098 22140 5510
rect 22296 5234 22324 5510
rect 22284 5228 22336 5234
rect 22204 5188 22284 5216
rect 22100 5092 22152 5098
rect 22100 5034 22152 5040
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 21916 4752 21968 4758
rect 21916 4694 21968 4700
rect 21732 4276 21784 4282
rect 21732 4218 21784 4224
rect 21928 4154 21956 4694
rect 22020 4282 22048 4762
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 21836 4126 21956 4154
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 21456 3664 21508 3670
rect 21456 3606 21508 3612
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20640 2650 20668 3334
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 21008 2650 21036 2926
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 20640 2446 20668 2586
rect 21468 2514 21496 3606
rect 21652 2961 21680 3878
rect 21732 3392 21784 3398
rect 21732 3334 21784 3340
rect 21744 3194 21772 3334
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 21744 2990 21772 3130
rect 21836 2990 21864 4126
rect 22020 3602 22048 4218
rect 22112 4078 22140 4558
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 22112 3641 22140 4014
rect 22204 3670 22232 5188
rect 22284 5170 22336 5176
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22296 4078 22324 4966
rect 22756 4690 22784 7278
rect 23940 7268 23992 7274
rect 23940 7210 23992 7216
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23492 6458 23520 6802
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 22928 5840 22980 5846
rect 22928 5782 22980 5788
rect 22940 5370 22968 5782
rect 23492 5642 23520 6394
rect 23480 5636 23532 5642
rect 23480 5578 23532 5584
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 22836 5024 22888 5030
rect 22836 4966 22888 4972
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 22848 4690 22876 4966
rect 23492 4826 23520 4966
rect 23952 4826 23980 7210
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 24044 5710 24072 6054
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 24228 5302 24256 7919
rect 26146 7848 26202 7857
rect 26146 7783 26202 7792
rect 26160 7274 26188 7783
rect 26148 7268 26200 7274
rect 26148 7210 26200 7216
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24504 6458 24532 6802
rect 24584 6656 24636 6662
rect 24584 6598 24636 6604
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24400 6180 24452 6186
rect 24400 6122 24452 6128
rect 24306 5944 24362 5953
rect 24306 5879 24362 5888
rect 24216 5296 24268 5302
rect 24216 5238 24268 5244
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 23940 4820 23992 4826
rect 23940 4762 23992 4768
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 23112 4684 23164 4690
rect 23112 4626 23164 4632
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22756 4010 22784 4626
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 23032 4146 23060 4558
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 22744 4004 22796 4010
rect 22744 3946 22796 3952
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 22192 3664 22244 3670
rect 22098 3632 22154 3641
rect 22008 3596 22060 3602
rect 22192 3606 22244 3612
rect 22098 3567 22154 3576
rect 22008 3538 22060 3544
rect 22020 3058 22048 3538
rect 22296 3534 22324 3878
rect 22756 3738 22784 3946
rect 23032 3942 23060 4082
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 22204 3126 22232 3334
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 21732 2984 21784 2990
rect 21638 2952 21694 2961
rect 21732 2926 21784 2932
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21638 2887 21694 2896
rect 21744 2582 21772 2926
rect 21732 2576 21784 2582
rect 21732 2518 21784 2524
rect 22020 2514 22048 2994
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 22020 2310 22048 2450
rect 22296 2446 22324 3470
rect 23032 2650 23060 3878
rect 23124 3534 23152 4626
rect 23492 4146 23520 4762
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23204 4004 23256 4010
rect 23204 3946 23256 3952
rect 23216 3602 23244 3946
rect 23204 3596 23256 3602
rect 23388 3596 23440 3602
rect 23204 3538 23256 3544
rect 23308 3556 23388 3584
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23216 2854 23244 3538
rect 23308 2990 23336 3556
rect 23388 3538 23440 3544
rect 23664 3392 23716 3398
rect 23664 3334 23716 3340
rect 23676 2990 23704 3334
rect 23952 3194 23980 4762
rect 24320 4758 24348 5879
rect 24412 5370 24440 6122
rect 24596 5846 24624 6598
rect 24860 6452 24912 6458
rect 24860 6394 24912 6400
rect 24584 5840 24636 5846
rect 24584 5782 24636 5788
rect 24492 5704 24544 5710
rect 24492 5646 24544 5652
rect 24400 5364 24452 5370
rect 24400 5306 24452 5312
rect 24504 4826 24532 5646
rect 24596 5370 24624 5782
rect 24584 5364 24636 5370
rect 24584 5306 24636 5312
rect 24872 5098 24900 6394
rect 25148 6186 25176 6598
rect 25412 6316 25464 6322
rect 25412 6258 25464 6264
rect 25136 6180 25188 6186
rect 25136 6122 25188 6128
rect 25424 5914 25452 6258
rect 25504 6112 25556 6118
rect 25504 6054 25556 6060
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25320 5636 25372 5642
rect 25320 5578 25372 5584
rect 25332 5302 25360 5578
rect 25320 5296 25372 5302
rect 25320 5238 25372 5244
rect 25424 5234 25452 5850
rect 25516 5778 25544 6054
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 25504 5772 25556 5778
rect 25504 5714 25556 5720
rect 27252 5772 27304 5778
rect 27252 5714 27304 5720
rect 25228 5228 25280 5234
rect 25228 5170 25280 5176
rect 25412 5228 25464 5234
rect 25412 5170 25464 5176
rect 24860 5092 24912 5098
rect 24860 5034 24912 5040
rect 24492 4820 24544 4826
rect 24492 4762 24544 4768
rect 24308 4752 24360 4758
rect 24308 4694 24360 4700
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 24780 4010 24808 4558
rect 24872 4282 24900 5034
rect 24952 4820 25004 4826
rect 24952 4762 25004 4768
rect 24860 4276 24912 4282
rect 24860 4218 24912 4224
rect 24768 4004 24820 4010
rect 24768 3946 24820 3952
rect 24780 3670 24808 3946
rect 24964 3942 24992 4762
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 23940 3188 23992 3194
rect 23940 3130 23992 3136
rect 23952 2990 23980 3130
rect 24504 2990 24532 3470
rect 24688 2990 24716 3538
rect 25240 3534 25268 5170
rect 25516 4826 25544 5714
rect 26516 5704 26568 5710
rect 26516 5646 26568 5652
rect 25504 4820 25556 4826
rect 25504 4762 25556 4768
rect 25320 4752 25372 4758
rect 25320 4694 25372 4700
rect 25332 4146 25360 4694
rect 26424 4548 26476 4554
rect 26424 4490 26476 4496
rect 26332 4276 26384 4282
rect 26332 4218 26384 4224
rect 26344 4185 26372 4218
rect 26330 4176 26386 4185
rect 25320 4140 25372 4146
rect 25320 4082 25372 4088
rect 25964 4140 26016 4146
rect 26330 4111 26386 4120
rect 25964 4082 26016 4088
rect 25872 4072 25924 4078
rect 25872 4014 25924 4020
rect 25884 3738 25912 4014
rect 25976 3942 26004 4082
rect 26436 4078 26464 4490
rect 26424 4072 26476 4078
rect 26424 4014 26476 4020
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 25412 3664 25464 3670
rect 25412 3606 25464 3612
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25424 3194 25452 3606
rect 25412 3188 25464 3194
rect 25412 3130 25464 3136
rect 23296 2984 23348 2990
rect 23296 2926 23348 2932
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 23940 2984 23992 2990
rect 23940 2926 23992 2932
rect 24124 2984 24176 2990
rect 24124 2926 24176 2932
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 23032 2514 23060 2586
rect 23020 2508 23072 2514
rect 23020 2450 23072 2456
rect 22284 2440 22336 2446
rect 22190 2408 22246 2417
rect 22112 2378 22190 2394
rect 22100 2372 22190 2378
rect 22152 2366 22190 2372
rect 22284 2382 22336 2388
rect 22190 2343 22246 2352
rect 22100 2314 22152 2320
rect 22008 2304 22060 2310
rect 22008 2246 22060 2252
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 20074 1592 20130 1601
rect 20074 1527 20130 1536
rect 19890 82 19946 480
rect 19628 54 19946 82
rect 23400 82 23428 2790
rect 23676 2514 23704 2926
rect 24136 2650 24164 2926
rect 24952 2916 25004 2922
rect 24952 2858 25004 2864
rect 24124 2644 24176 2650
rect 24124 2586 24176 2592
rect 24136 2514 24164 2586
rect 24964 2514 24992 2858
rect 23664 2508 23716 2514
rect 23664 2450 23716 2456
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24952 2508 25004 2514
rect 24952 2450 25004 2456
rect 23676 2310 23704 2450
rect 24964 2378 24992 2450
rect 24952 2372 25004 2378
rect 24952 2314 25004 2320
rect 23664 2304 23716 2310
rect 23664 2246 23716 2252
rect 23570 82 23626 480
rect 25976 241 26004 3878
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26252 2990 26280 3334
rect 26436 3126 26464 4014
rect 26528 3670 26556 5646
rect 27264 5370 27292 5714
rect 27436 5568 27488 5574
rect 27436 5510 27488 5516
rect 27896 5568 27948 5574
rect 27896 5510 27948 5516
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 26792 5228 26844 5234
rect 26792 5170 26844 5176
rect 26804 4486 26832 5170
rect 26976 5160 27028 5166
rect 26974 5128 26976 5137
rect 27028 5128 27030 5137
rect 26974 5063 27030 5072
rect 27160 5092 27212 5098
rect 26988 5030 27016 5063
rect 27160 5034 27212 5040
rect 26976 5024 27028 5030
rect 26976 4966 27028 4972
rect 26884 4820 26936 4826
rect 26884 4762 26936 4768
rect 26896 4729 26924 4762
rect 26882 4720 26938 4729
rect 26882 4655 26938 4664
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26896 4282 26924 4655
rect 27172 4622 27200 5034
rect 27448 5030 27476 5510
rect 27908 5234 27936 5510
rect 27896 5228 27948 5234
rect 27896 5170 27948 5176
rect 28264 5092 28316 5098
rect 28264 5034 28316 5040
rect 27436 5024 27488 5030
rect 27436 4966 27488 4972
rect 27160 4616 27212 4622
rect 27160 4558 27212 4564
rect 27252 4480 27304 4486
rect 27252 4422 27304 4428
rect 26884 4276 26936 4282
rect 26884 4218 26936 4224
rect 27264 4010 27292 4422
rect 27252 4004 27304 4010
rect 27252 3946 27304 3952
rect 27264 3670 27292 3946
rect 27448 3738 27476 4966
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 28276 4758 28304 5034
rect 27712 4752 27764 4758
rect 27712 4694 27764 4700
rect 28264 4752 28316 4758
rect 28264 4694 28316 4700
rect 27724 4010 27752 4694
rect 28080 4616 28132 4622
rect 28080 4558 28132 4564
rect 28092 4282 28120 4558
rect 28080 4276 28132 4282
rect 28080 4218 28132 4224
rect 27712 4004 27764 4010
rect 27712 3946 27764 3952
rect 27988 3936 28040 3942
rect 27988 3878 28040 3884
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 27436 3732 27488 3738
rect 27436 3674 27488 3680
rect 26516 3664 26568 3670
rect 26516 3606 26568 3612
rect 27252 3664 27304 3670
rect 27252 3606 27304 3612
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26424 3120 26476 3126
rect 26424 3062 26476 3068
rect 26528 3058 26556 3470
rect 26516 3052 26568 3058
rect 26516 2994 26568 3000
rect 26240 2984 26292 2990
rect 26240 2926 26292 2932
rect 26148 2848 26200 2854
rect 26148 2790 26200 2796
rect 26160 2650 26188 2790
rect 26148 2644 26200 2650
rect 26148 2586 26200 2592
rect 26252 2582 26280 2926
rect 27264 2650 27292 3606
rect 27448 3126 27476 3674
rect 27436 3120 27488 3126
rect 27436 3062 27488 3068
rect 28000 3058 28028 3878
rect 28276 3738 28304 4694
rect 29184 4684 29236 4690
rect 29184 4626 29236 4632
rect 29196 4282 29224 4626
rect 29552 4480 29604 4486
rect 29552 4422 29604 4428
rect 28448 4276 28500 4282
rect 28448 4218 28500 4224
rect 29184 4276 29236 4282
rect 29184 4218 29236 4224
rect 28264 3732 28316 3738
rect 28264 3674 28316 3680
rect 28460 3670 28488 4218
rect 29184 4072 29236 4078
rect 29184 4014 29236 4020
rect 28448 3664 28500 3670
rect 28448 3606 28500 3612
rect 28460 3194 28488 3606
rect 29196 3369 29224 4014
rect 29276 3392 29328 3398
rect 29182 3360 29238 3369
rect 29276 3334 29328 3340
rect 29182 3295 29238 3304
rect 28448 3188 28500 3194
rect 28448 3130 28500 3136
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 27436 2848 27488 2854
rect 27436 2790 27488 2796
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 27252 2644 27304 2650
rect 27252 2586 27304 2592
rect 26240 2576 26292 2582
rect 26240 2518 26292 2524
rect 25962 232 26018 241
rect 25962 167 26018 176
rect 23400 54 23626 82
rect 5354 0 5410 54
rect 9034 0 9090 54
rect 12622 0 12678 54
rect 16302 0 16358 54
rect 19890 0 19946 54
rect 23570 0 23626 54
rect 27158 82 27214 480
rect 27264 82 27292 2586
rect 27448 2514 27476 2790
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 28092 2650 28120 2790
rect 28080 2644 28132 2650
rect 28080 2586 28132 2592
rect 27436 2508 27488 2514
rect 27436 2450 27488 2456
rect 29288 2446 29316 3334
rect 29564 2650 29592 4422
rect 29840 4282 29868 10406
rect 33428 10033 33456 15558
rect 35714 15056 35770 15065
rect 35714 14991 35770 15000
rect 35530 14240 35586 14249
rect 35530 14175 35586 14184
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 35452 10470 35480 11154
rect 35440 10464 35492 10470
rect 35440 10406 35492 10412
rect 35440 10124 35492 10130
rect 35440 10066 35492 10072
rect 33414 10024 33470 10033
rect 33414 9959 33470 9968
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 35452 9382 35480 10066
rect 35440 9376 35492 9382
rect 35440 9318 35492 9324
rect 35452 9081 35480 9318
rect 35438 9072 35494 9081
rect 35256 9036 35308 9042
rect 35438 9007 35494 9016
rect 35256 8978 35308 8984
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 34060 8424 34112 8430
rect 34060 8366 34112 8372
rect 34072 7721 34100 8366
rect 35268 8294 35296 8978
rect 35438 8392 35494 8401
rect 35438 8327 35494 8336
rect 34152 8288 34204 8294
rect 34152 8230 34204 8236
rect 35256 8288 35308 8294
rect 35256 8230 35308 8236
rect 34058 7712 34114 7721
rect 34058 7647 34114 7656
rect 34164 7585 34192 8230
rect 35452 7954 35480 8327
rect 35440 7948 35492 7954
rect 35440 7890 35492 7896
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34150 7576 34206 7585
rect 34289 7568 34585 7588
rect 35452 7546 35480 7890
rect 35544 7546 35572 14175
rect 35622 11520 35678 11529
rect 35622 11455 35678 11464
rect 35636 11354 35664 11455
rect 35624 11348 35676 11354
rect 35624 11290 35676 11296
rect 35622 10568 35678 10577
rect 35622 10503 35678 10512
rect 35636 10266 35664 10503
rect 35624 10260 35676 10266
rect 35624 10202 35676 10208
rect 35622 9752 35678 9761
rect 35622 9687 35678 9696
rect 35636 9178 35664 9687
rect 35624 9172 35676 9178
rect 35624 9114 35676 9120
rect 35622 8800 35678 8809
rect 35622 8735 35678 8744
rect 35636 8634 35664 8735
rect 35624 8628 35676 8634
rect 35624 8570 35676 8576
rect 35728 8090 35756 14991
rect 39578 13800 39634 13809
rect 39578 13735 39634 13744
rect 35806 12336 35862 12345
rect 35806 12271 35862 12280
rect 35716 8084 35768 8090
rect 35716 8026 35768 8032
rect 34150 7511 34206 7520
rect 35440 7540 35492 7546
rect 35440 7482 35492 7488
rect 35532 7540 35584 7546
rect 35532 7482 35584 7488
rect 35440 6860 35492 6866
rect 35440 6802 35492 6808
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 35452 6322 35480 6802
rect 35440 6316 35492 6322
rect 35440 6258 35492 6264
rect 35452 6225 35480 6258
rect 35438 6216 35494 6225
rect 35438 6151 35494 6160
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 30286 5400 30342 5409
rect 34289 5392 34585 5412
rect 35820 5370 35848 12271
rect 36726 7984 36782 7993
rect 36726 7919 36782 7928
rect 36740 7546 36768 7919
rect 36728 7540 36780 7546
rect 36728 7482 36780 7488
rect 35992 7404 36044 7410
rect 35992 7346 36044 7352
rect 36004 7313 36032 7346
rect 35990 7304 36046 7313
rect 35990 7239 36046 7248
rect 39592 7002 39620 13735
rect 39580 6996 39632 7002
rect 39580 6938 39632 6944
rect 30286 5335 30342 5344
rect 35808 5364 35860 5370
rect 30300 4758 30328 5335
rect 35808 5306 35860 5312
rect 35440 5160 35492 5166
rect 35440 5102 35492 5108
rect 30288 4752 30340 4758
rect 35452 4729 35480 5102
rect 30288 4694 30340 4700
rect 35438 4720 35494 4729
rect 31392 4684 31444 4690
rect 35438 4655 35494 4664
rect 31392 4626 31444 4632
rect 30564 4480 30616 4486
rect 30564 4422 30616 4428
rect 29828 4276 29880 4282
rect 29828 4218 29880 4224
rect 29840 4078 29868 4218
rect 29828 4072 29880 4078
rect 29828 4014 29880 4020
rect 30380 4004 30432 4010
rect 30380 3946 30432 3952
rect 30392 3738 30420 3946
rect 30380 3732 30432 3738
rect 30380 3674 30432 3680
rect 30576 3670 30604 4422
rect 31404 4078 31432 4626
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 31392 4072 31444 4078
rect 31390 4040 31392 4049
rect 31444 4040 31446 4049
rect 31024 4004 31076 4010
rect 31390 3975 31446 3984
rect 31024 3946 31076 3952
rect 31404 3949 31432 3975
rect 30564 3664 30616 3670
rect 30564 3606 30616 3612
rect 30656 3664 30708 3670
rect 30656 3606 30708 3612
rect 30668 3194 30696 3606
rect 31036 3534 31064 3946
rect 32220 3936 32272 3942
rect 32220 3878 32272 3884
rect 32232 3602 32260 3878
rect 32220 3596 32272 3602
rect 32220 3538 32272 3544
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 30656 3188 30708 3194
rect 30656 3130 30708 3136
rect 30932 2916 30984 2922
rect 31036 2904 31064 3470
rect 32232 3194 32260 3538
rect 32496 3392 32548 3398
rect 32496 3334 32548 3340
rect 32220 3188 32272 3194
rect 32220 3130 32272 3136
rect 32036 3052 32088 3058
rect 32036 2994 32088 3000
rect 31116 2916 31168 2922
rect 31036 2876 31116 2904
rect 30932 2858 30984 2864
rect 31116 2858 31168 2864
rect 29552 2644 29604 2650
rect 29552 2586 29604 2592
rect 30944 2582 30972 2858
rect 31208 2848 31260 2854
rect 31208 2790 31260 2796
rect 30932 2576 30984 2582
rect 30932 2518 30984 2524
rect 31220 2446 31248 2790
rect 32048 2650 32076 2994
rect 32508 2922 32536 3334
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 32496 2916 32548 2922
rect 32496 2858 32548 2864
rect 32680 2916 32732 2922
rect 32680 2858 32732 2864
rect 32036 2644 32088 2650
rect 32036 2586 32088 2592
rect 31852 2576 31904 2582
rect 31852 2518 31904 2524
rect 32128 2576 32180 2582
rect 32128 2518 32180 2524
rect 29276 2440 29328 2446
rect 31208 2440 31260 2446
rect 29276 2382 29328 2388
rect 30562 2408 30618 2417
rect 31864 2428 31892 2518
rect 32140 2428 32168 2518
rect 32692 2514 32720 2858
rect 32680 2508 32732 2514
rect 32680 2450 32732 2456
rect 31864 2400 32168 2428
rect 31208 2382 31260 2388
rect 30562 2343 30618 2352
rect 34152 2372 34204 2378
rect 27158 54 27292 82
rect 30576 82 30604 2343
rect 34152 2314 34204 2320
rect 30748 2304 30800 2310
rect 30748 2246 30800 2252
rect 30760 1193 30788 2246
rect 30746 1184 30802 1193
rect 30746 1119 30802 1128
rect 30838 82 30894 480
rect 30576 54 30894 82
rect 34164 82 34192 2314
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 39578 1320 39634 1329
rect 39578 1255 39634 1264
rect 38198 1184 38254 1193
rect 38198 1119 38254 1128
rect 34426 82 34482 480
rect 34164 54 34482 82
rect 27158 0 27214 54
rect 30838 0 30894 54
rect 34426 0 34482 54
rect 38106 82 38162 480
rect 38212 82 38240 1119
rect 39592 241 39620 1255
rect 39578 232 39634 241
rect 39578 167 39634 176
rect 38106 54 38240 82
rect 38106 0 38162 54
<< via2 >>
rect 1214 15000 1270 15056
rect 18 13776 74 13832
rect 1030 12280 1086 12336
rect 1490 14184 1546 14240
rect 1582 11464 1638 11520
rect 1582 10512 1638 10568
rect 1582 9696 1638 9752
rect 1674 8880 1730 8936
rect 1582 8744 1638 8800
rect 2686 8064 2742 8120
rect 2134 7248 2190 7304
rect 2042 7112 2098 7168
rect 2042 6840 2098 6896
rect 2318 6296 2374 6352
rect 1674 6024 1730 6080
rect 2042 5208 2098 5264
rect 110 3984 166 4040
rect 3330 7384 3386 7440
rect 2962 6296 3018 6352
rect 4066 8200 4122 8256
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 16762 9968 16818 10024
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 5078 7928 5134 7984
rect 3514 3440 3570 3496
rect 2594 2352 2650 2408
rect 2318 720 2374 776
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 13634 7792 13690 7848
rect 9954 6840 10010 6896
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 5354 2760 5410 2816
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 9954 5616 10010 5672
rect 12530 7248 12586 7304
rect 18602 9016 18658 9072
rect 10690 6568 10746 6624
rect 4250 312 4306 368
rect 7010 2488 7066 2544
rect 8850 3304 8906 3360
rect 10138 3440 10194 3496
rect 11518 3576 11574 3632
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 14186 7248 14242 7304
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 16394 7248 16450 7304
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 18326 6860 18382 6896
rect 18326 6840 18328 6860
rect 18328 6840 18380 6860
rect 18380 6840 18382 6860
rect 16394 5888 16450 5944
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 14186 3304 14242 3360
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 14278 2488 14334 2544
rect 13634 1128 13690 1184
rect 18326 6296 18382 6352
rect 20442 8880 20498 8936
rect 19154 7792 19210 7848
rect 17498 6196 17500 6216
rect 17500 6196 17552 6216
rect 17552 6196 17554 6216
rect 17498 6160 17554 6196
rect 17498 5752 17554 5808
rect 18602 3984 18658 4040
rect 18878 6704 18934 6760
rect 20074 7248 20130 7304
rect 19154 6432 19210 6488
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 24214 7928 24270 7984
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 21362 7384 21418 7440
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 21362 5344 21418 5400
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 22374 7520 22430 7576
rect 22374 6704 22430 6760
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 26146 7792 26202 7848
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 24306 5888 24362 5944
rect 22098 3576 22154 3632
rect 21638 2896 21694 2952
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 26330 4120 26386 4176
rect 22190 2352 22246 2408
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 20074 1536 20130 1592
rect 26974 5108 26976 5128
rect 26976 5108 27028 5128
rect 27028 5108 27030 5128
rect 26974 5072 27030 5108
rect 26882 4664 26938 4720
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 29182 3304 29238 3360
rect 25962 176 26018 232
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 35714 15000 35770 15056
rect 35530 14184 35586 14240
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 33414 9968 33470 10024
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 35438 9016 35494 9072
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 35438 8336 35494 8392
rect 34058 7656 34114 7712
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 34150 7520 34206 7576
rect 35622 11464 35678 11520
rect 35622 10512 35678 10568
rect 35622 9696 35678 9752
rect 35622 8744 35678 8800
rect 39578 13744 39634 13800
rect 35806 12280 35862 12336
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 35438 6160 35494 6216
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 30286 5344 30342 5400
rect 36726 7928 36782 7984
rect 35990 7248 36046 7304
rect 35438 4664 35494 4720
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 31390 4020 31392 4040
rect 31392 4020 31444 4040
rect 31444 4020 31446 4040
rect 31390 3984 31446 4020
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 30562 2352 30618 2408
rect 30746 1128 30802 1184
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 39578 1264 39634 1320
rect 38198 1128 38254 1184
rect 39578 176 39634 232
<< metal3 >>
rect 0 15512 480 15632
rect 39520 15512 40000 15632
rect 62 15058 122 15512
rect 1209 15058 1275 15061
rect 62 15056 1275 15058
rect 62 15000 1214 15056
rect 1270 15000 1275 15056
rect 62 14998 1275 15000
rect 1209 14995 1275 14998
rect 35709 15058 35775 15061
rect 39622 15058 39682 15512
rect 35709 15056 39682 15058
rect 35709 15000 35714 15056
rect 35770 15000 39682 15056
rect 35709 14998 39682 15000
rect 35709 14995 35775 14998
rect 0 14560 480 14680
rect 39520 14560 40000 14680
rect 62 14242 122 14560
rect 1485 14242 1551 14245
rect 62 14240 1551 14242
rect 62 14184 1490 14240
rect 1546 14184 1551 14240
rect 62 14182 1551 14184
rect 1485 14179 1551 14182
rect 35525 14242 35591 14245
rect 39622 14242 39682 14560
rect 35525 14240 39682 14242
rect 35525 14184 35530 14240
rect 35586 14184 39682 14240
rect 35525 14182 39682 14184
rect 35525 14179 35591 14182
rect 0 13832 480 13864
rect 0 13776 18 13832
rect 74 13776 480 13832
rect 39520 13802 40000 13864
rect 0 13744 480 13776
rect 39492 13800 40000 13802
rect 39492 13744 39578 13800
rect 39634 13744 40000 13800
rect 39492 13742 39639 13744
rect 39573 13739 39639 13742
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 0 12792 480 12912
rect 39520 12792 40000 12912
rect 62 12338 122 12792
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 1025 12338 1091 12341
rect 62 12336 1091 12338
rect 62 12280 1030 12336
rect 1086 12280 1091 12336
rect 62 12278 1091 12280
rect 1025 12275 1091 12278
rect 35801 12338 35867 12341
rect 39622 12338 39682 12792
rect 35801 12336 39682 12338
rect 35801 12280 35806 12336
rect 35862 12280 39682 12336
rect 35801 12278 39682 12280
rect 35801 12275 35867 12278
rect 0 11976 480 12096
rect 7610 12000 7930 12001
rect 62 11522 122 11976
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 39520 11976 40000 12096
rect 34277 11935 34597 11936
rect 1577 11522 1643 11525
rect 62 11520 1643 11522
rect 62 11464 1582 11520
rect 1638 11464 1643 11520
rect 62 11462 1643 11464
rect 1577 11459 1643 11462
rect 35617 11522 35683 11525
rect 39622 11522 39682 11976
rect 35617 11520 39682 11522
rect 35617 11464 35622 11520
rect 35678 11464 39682 11520
rect 35617 11462 39682 11464
rect 35617 11459 35683 11462
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 0 11024 480 11144
rect 39520 11024 40000 11144
rect 62 10570 122 11024
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 1577 10570 1643 10573
rect 62 10568 1643 10570
rect 62 10512 1582 10568
rect 1638 10512 1643 10568
rect 62 10510 1643 10512
rect 1577 10507 1643 10510
rect 35617 10570 35683 10573
rect 39622 10570 39682 11024
rect 35617 10568 39682 10570
rect 35617 10512 35622 10568
rect 35678 10512 39682 10568
rect 35617 10510 39682 10512
rect 35617 10507 35683 10510
rect 14277 10368 14597 10369
rect 0 10208 480 10328
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 39520 10208 40000 10328
rect 62 9754 122 10208
rect 16757 10026 16823 10029
rect 33409 10026 33475 10029
rect 16757 10024 33475 10026
rect 16757 9968 16762 10024
rect 16818 9968 33414 10024
rect 33470 9968 33475 10024
rect 16757 9966 33475 9968
rect 16757 9963 16823 9966
rect 33409 9963 33475 9966
rect 7610 9824 7930 9825
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 1577 9754 1643 9757
rect 62 9752 1643 9754
rect 62 9696 1582 9752
rect 1638 9696 1643 9752
rect 62 9694 1643 9696
rect 1577 9691 1643 9694
rect 35617 9754 35683 9757
rect 39622 9754 39682 10208
rect 35617 9752 39682 9754
rect 35617 9696 35622 9752
rect 35678 9696 39682 9752
rect 35617 9694 39682 9696
rect 35617 9691 35683 9694
rect 0 9256 480 9376
rect 14277 9280 14597 9281
rect 62 8802 122 9256
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 39520 9256 40000 9376
rect 27610 9215 27930 9216
rect 18597 9074 18663 9077
rect 35433 9074 35499 9077
rect 18597 9072 35499 9074
rect 18597 9016 18602 9072
rect 18658 9016 35438 9072
rect 35494 9016 35499 9072
rect 18597 9014 35499 9016
rect 18597 9011 18663 9014
rect 35433 9011 35499 9014
rect 1669 8938 1735 8941
rect 20437 8938 20503 8941
rect 1669 8936 20503 8938
rect 1669 8880 1674 8936
rect 1730 8880 20442 8936
rect 20498 8880 20503 8936
rect 1669 8878 20503 8880
rect 1669 8875 1735 8878
rect 20437 8875 20503 8878
rect 1577 8802 1643 8805
rect 62 8800 1643 8802
rect 62 8744 1582 8800
rect 1638 8744 1643 8800
rect 62 8742 1643 8744
rect 1577 8739 1643 8742
rect 35617 8802 35683 8805
rect 39622 8802 39682 9256
rect 35617 8800 39682 8802
rect 35617 8744 35622 8800
rect 35678 8744 39682 8800
rect 35617 8742 39682 8744
rect 35617 8739 35683 8742
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 0 8440 480 8560
rect 39520 8440 40000 8560
rect 62 8122 122 8440
rect 35433 8394 35499 8397
rect 4110 8392 35499 8394
rect 4110 8336 35438 8392
rect 35494 8336 35499 8392
rect 4110 8334 35499 8336
rect 4110 8261 4170 8334
rect 35433 8331 35499 8334
rect 4061 8256 4170 8261
rect 4061 8200 4066 8256
rect 4122 8200 4170 8256
rect 4061 8195 4170 8200
rect 2681 8122 2747 8125
rect 62 8120 2747 8122
rect 62 8064 2686 8120
rect 2742 8064 2747 8120
rect 62 8062 2747 8064
rect 2681 8059 2747 8062
rect 4110 7986 4170 8195
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 17910 8062 27538 8122
rect 62 7926 4170 7986
rect 5073 7986 5139 7989
rect 17910 7986 17970 8062
rect 24209 7986 24275 7989
rect 27478 7986 27538 8062
rect 36721 7986 36787 7989
rect 39622 7986 39682 8440
rect 5073 7984 17970 7986
rect 5073 7928 5078 7984
rect 5134 7928 17970 7984
rect 5073 7926 17970 7928
rect 18600 7984 26388 7986
rect 18600 7928 24214 7984
rect 24270 7928 26388 7984
rect 18600 7926 26388 7928
rect 27478 7926 33150 7986
rect 62 7608 122 7926
rect 5073 7923 5139 7926
rect 13629 7850 13695 7853
rect 18600 7850 18660 7926
rect 24209 7923 24275 7926
rect 13629 7848 18660 7850
rect 13629 7792 13634 7848
rect 13690 7792 18660 7848
rect 13629 7790 18660 7792
rect 19149 7850 19215 7853
rect 26141 7850 26207 7853
rect 19149 7848 26207 7850
rect 19149 7792 19154 7848
rect 19210 7792 26146 7848
rect 26202 7792 26207 7848
rect 19149 7790 26207 7792
rect 13629 7787 13695 7790
rect 19149 7787 19215 7790
rect 26141 7787 26207 7790
rect 26328 7714 26388 7926
rect 33090 7850 33150 7926
rect 36721 7984 39682 7986
rect 36721 7928 36726 7984
rect 36782 7928 39682 7984
rect 36721 7926 39682 7928
rect 36721 7923 36787 7926
rect 33090 7790 39682 7850
rect 34053 7714 34119 7717
rect 26328 7712 34119 7714
rect 26328 7656 34058 7712
rect 34114 7656 34119 7712
rect 26328 7654 34119 7656
rect 34053 7651 34119 7654
rect 7610 7648 7930 7649
rect 0 7488 480 7608
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 39622 7608 39682 7790
rect 34277 7583 34597 7584
rect 22369 7578 22435 7581
rect 34145 7578 34211 7581
rect 22369 7576 34211 7578
rect 22369 7520 22374 7576
rect 22430 7520 34150 7576
rect 34206 7520 34211 7576
rect 22369 7518 34211 7520
rect 22369 7515 22435 7518
rect 34145 7515 34211 7518
rect 39520 7488 40000 7608
rect 3325 7442 3391 7445
rect 21357 7442 21423 7445
rect 3325 7440 21423 7442
rect 3325 7384 3330 7440
rect 3386 7384 21362 7440
rect 21418 7384 21423 7440
rect 3325 7382 21423 7384
rect 3325 7379 3391 7382
rect 21357 7379 21423 7382
rect 2129 7306 2195 7309
rect 12525 7306 12591 7309
rect 14181 7306 14247 7309
rect 16389 7306 16455 7309
rect 2129 7304 12591 7306
rect 2129 7248 2134 7304
rect 2190 7248 12530 7304
rect 12586 7248 12591 7304
rect 2129 7246 12591 7248
rect 2129 7243 2195 7246
rect 12525 7243 12591 7246
rect 13770 7304 16455 7306
rect 13770 7248 14186 7304
rect 14242 7248 16394 7304
rect 16450 7248 16455 7304
rect 13770 7246 16455 7248
rect 2037 7170 2103 7173
rect 13770 7170 13830 7246
rect 14181 7243 14247 7246
rect 16389 7243 16455 7246
rect 20069 7306 20135 7309
rect 35985 7306 36051 7309
rect 20069 7304 36051 7306
rect 20069 7248 20074 7304
rect 20130 7248 35990 7304
rect 36046 7248 36051 7304
rect 20069 7246 36051 7248
rect 20069 7243 20135 7246
rect 35985 7243 36051 7246
rect 2037 7168 13830 7170
rect 2037 7112 2042 7168
rect 2098 7112 13830 7168
rect 2037 7110 13830 7112
rect 2037 7107 2103 7110
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 54 6836 60 6900
rect 124 6898 130 6900
rect 2037 6898 2103 6901
rect 9949 6898 10015 6901
rect 124 6838 674 6898
rect 124 6836 130 6838
rect 614 6762 674 6838
rect 2037 6896 10015 6898
rect 2037 6840 2042 6896
rect 2098 6840 9954 6896
rect 10010 6840 10015 6896
rect 2037 6838 10015 6840
rect 2037 6835 2103 6838
rect 9949 6835 10015 6838
rect 18321 6898 18387 6901
rect 18321 6896 39682 6898
rect 18321 6840 18326 6896
rect 18382 6840 39682 6896
rect 18321 6838 39682 6840
rect 18321 6835 18387 6838
rect 18873 6762 18939 6765
rect 22369 6762 22435 6765
rect 614 6760 18939 6762
rect 614 6704 18878 6760
rect 18934 6704 18939 6760
rect 614 6702 18939 6704
rect 18873 6699 18939 6702
rect 20716 6760 22435 6762
rect 20716 6704 22374 6760
rect 22430 6704 22435 6760
rect 20716 6702 22435 6704
rect 0 6628 480 6656
rect 0 6564 60 6628
rect 124 6564 480 6628
rect 0 6536 480 6564
rect 10685 6626 10751 6629
rect 20716 6626 20776 6702
rect 22369 6699 22435 6702
rect 39622 6656 39682 6838
rect 10685 6624 20776 6626
rect 10685 6568 10690 6624
rect 10746 6568 20776 6624
rect 10685 6566 20776 6568
rect 10685 6563 10751 6566
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 39520 6536 40000 6656
rect 34277 6495 34597 6496
rect 19149 6490 19215 6493
rect 13770 6488 19215 6490
rect 13770 6432 19154 6488
rect 19210 6432 19215 6488
rect 13770 6430 19215 6432
rect 2313 6354 2379 6357
rect 2957 6354 3023 6357
rect 13770 6354 13830 6430
rect 19149 6427 19215 6430
rect 18321 6354 18387 6357
rect 2313 6352 13830 6354
rect 2313 6296 2318 6352
rect 2374 6296 2962 6352
rect 3018 6296 13830 6352
rect 2313 6294 13830 6296
rect 14736 6352 18387 6354
rect 14736 6296 18326 6352
rect 18382 6296 18387 6352
rect 14736 6294 18387 6296
rect 2313 6291 2379 6294
rect 2957 6291 3023 6294
rect 14736 6218 14796 6294
rect 18321 6291 18387 6294
rect 4110 6158 14796 6218
rect 17493 6218 17559 6221
rect 35433 6218 35499 6221
rect 17493 6216 35499 6218
rect 17493 6160 17498 6216
rect 17554 6160 35438 6216
rect 35494 6160 35499 6216
rect 17493 6158 35499 6160
rect 54 6020 60 6084
rect 124 6082 130 6084
rect 1669 6082 1735 6085
rect 4110 6082 4170 6158
rect 17493 6155 17559 6158
rect 35433 6155 35499 6158
rect 124 6022 674 6082
rect 124 6020 130 6022
rect 614 5946 674 6022
rect 1669 6080 4170 6082
rect 1669 6024 1674 6080
rect 1730 6024 4170 6080
rect 1669 6022 4170 6024
rect 1669 6019 1735 6022
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 16389 5946 16455 5949
rect 24301 5946 24367 5949
rect 614 5886 9690 5946
rect 0 5812 480 5840
rect 0 5748 60 5812
rect 124 5748 480 5812
rect 9630 5810 9690 5886
rect 16389 5944 24367 5946
rect 16389 5888 16394 5944
rect 16450 5888 24306 5944
rect 24362 5888 24367 5944
rect 16389 5886 24367 5888
rect 16389 5883 16455 5886
rect 24301 5883 24367 5886
rect 17493 5810 17559 5813
rect 39520 5812 40000 5840
rect 39520 5810 39620 5812
rect 9630 5808 17559 5810
rect 9630 5752 17498 5808
rect 17554 5752 17559 5808
rect 9630 5750 17559 5752
rect 39492 5750 39620 5810
rect 0 5720 480 5748
rect 17493 5747 17559 5750
rect 39520 5748 39620 5750
rect 39684 5748 40000 5812
rect 39520 5720 40000 5748
rect 9949 5674 10015 5677
rect 9949 5672 39314 5674
rect 9949 5616 9954 5672
rect 10010 5616 39314 5672
rect 9949 5614 39314 5616
rect 9949 5611 10015 5614
rect 39254 5538 39314 5614
rect 39614 5538 39620 5540
rect 39254 5478 39620 5538
rect 39614 5476 39620 5478
rect 39684 5476 39690 5540
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 21357 5402 21423 5405
rect 30281 5402 30347 5405
rect 21357 5400 30347 5402
rect 21357 5344 21362 5400
rect 21418 5344 30286 5400
rect 30342 5344 30347 5400
rect 21357 5342 30347 5344
rect 21357 5339 21423 5342
rect 30281 5339 30347 5342
rect 2037 5266 2103 5269
rect 2037 5264 23490 5266
rect 2037 5208 2042 5264
rect 2098 5208 23490 5264
rect 2037 5206 23490 5208
rect 2037 5203 2103 5206
rect 23430 5130 23490 5206
rect 26969 5130 27035 5133
rect 23430 5128 39682 5130
rect 23430 5072 26974 5128
rect 27030 5072 39682 5128
rect 23430 5070 39682 5072
rect 26969 5067 27035 5070
rect 14277 4928 14597 4929
rect 0 4768 480 4888
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 39622 4888 39682 5070
rect 27610 4863 27930 4864
rect 39520 4768 40000 4888
rect 62 4314 122 4768
rect 26877 4722 26943 4725
rect 35433 4722 35499 4725
rect 26877 4720 35499 4722
rect 26877 4664 26882 4720
rect 26938 4664 35438 4720
rect 35494 4664 35499 4720
rect 26877 4662 35499 4664
rect 26877 4659 26943 4662
rect 35433 4659 35499 4662
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 62 4254 674 4314
rect 614 4178 674 4254
rect 26325 4178 26391 4181
rect 614 4176 26391 4178
rect 614 4120 26330 4176
rect 26386 4120 26391 4176
rect 614 4118 26391 4120
rect 26325 4115 26391 4118
rect 0 4040 480 4072
rect 18597 4042 18663 4045
rect 0 3984 110 4040
rect 166 3984 480 4040
rect 0 3952 480 3984
rect 4110 4040 18663 4042
rect 4110 3984 18602 4040
rect 18658 3984 18663 4040
rect 4110 3982 18663 3984
rect 4110 3770 4170 3982
rect 18597 3979 18663 3982
rect 31385 4042 31451 4045
rect 39520 4042 40000 4072
rect 31385 4040 40000 4042
rect 31385 3984 31390 4040
rect 31446 3984 40000 4040
rect 31385 3982 40000 3984
rect 31385 3979 31451 3982
rect 39520 3952 40000 3982
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 62 3710 4170 3770
rect 62 3120 122 3710
rect 11513 3634 11579 3637
rect 22093 3634 22159 3637
rect 11513 3632 22159 3634
rect 11513 3576 11518 3632
rect 11574 3576 22098 3632
rect 22154 3576 22159 3632
rect 11513 3574 22159 3576
rect 11513 3571 11579 3574
rect 22093 3571 22159 3574
rect 3509 3498 3575 3501
rect 10133 3498 10199 3501
rect 3509 3496 10199 3498
rect 3509 3440 3514 3496
rect 3570 3440 10138 3496
rect 10194 3440 10199 3496
rect 3509 3438 10199 3440
rect 3509 3435 3575 3438
rect 10133 3435 10199 3438
rect 8845 3362 8911 3365
rect 14181 3362 14247 3365
rect 8845 3360 14247 3362
rect 8845 3304 8850 3360
rect 8906 3304 14186 3360
rect 14242 3304 14247 3360
rect 8845 3302 14247 3304
rect 8845 3299 8911 3302
rect 14181 3299 14247 3302
rect 23422 3300 23428 3364
rect 23492 3362 23498 3364
rect 29177 3362 29243 3365
rect 23492 3360 29243 3362
rect 23492 3304 29182 3360
rect 29238 3304 29243 3360
rect 23492 3302 29243 3304
rect 23492 3300 23498 3302
rect 29177 3299 29243 3302
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 0 3000 480 3120
rect 39520 3092 40000 3120
rect 39520 3090 39620 3092
rect 39492 3030 39620 3090
rect 39520 3028 39620 3030
rect 39684 3028 40000 3092
rect 39520 3000 40000 3028
rect 21633 2954 21699 2957
rect 21633 2952 29010 2954
rect 21633 2896 21638 2952
rect 21694 2896 29010 2952
rect 21633 2894 29010 2896
rect 21633 2891 21699 2894
rect 5349 2818 5415 2821
rect 62 2816 5415 2818
rect 62 2760 5354 2816
rect 5410 2760 5415 2816
rect 62 2758 5415 2760
rect 28950 2818 29010 2894
rect 39614 2818 39620 2820
rect 28950 2758 39620 2818
rect 62 2304 122 2758
rect 5349 2755 5415 2758
rect 39614 2756 39620 2758
rect 39684 2756 39690 2820
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 7005 2546 7071 2549
rect 14273 2546 14339 2549
rect 7005 2544 14339 2546
rect 7005 2488 7010 2544
rect 7066 2488 14278 2544
rect 14334 2488 14339 2544
rect 7005 2486 14339 2488
rect 7005 2483 7071 2486
rect 14273 2483 14339 2486
rect 2589 2410 2655 2413
rect 4102 2410 4108 2412
rect 2589 2408 4108 2410
rect 2589 2352 2594 2408
rect 2650 2352 4108 2408
rect 2589 2350 4108 2352
rect 2589 2347 2655 2350
rect 4102 2348 4108 2350
rect 4172 2348 4178 2412
rect 22185 2410 22251 2413
rect 30557 2410 30623 2413
rect 22185 2408 30623 2410
rect 22185 2352 22190 2408
rect 22246 2352 30562 2408
rect 30618 2352 30623 2408
rect 22185 2350 30623 2352
rect 22185 2347 22251 2350
rect 30557 2347 30623 2350
rect 0 2184 480 2304
rect 7610 2208 7930 2209
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 39520 2184 40000 2304
rect 34277 2143 34597 2144
rect 20069 1594 20135 1597
rect 39622 1594 39682 2184
rect 20069 1592 39682 1594
rect 20069 1536 20074 1592
rect 20130 1536 39682 1592
rect 20069 1534 39682 1536
rect 20069 1531 20135 1534
rect 0 1324 480 1352
rect 0 1260 60 1324
rect 124 1260 480 1324
rect 39520 1322 40000 1352
rect 39492 1320 40000 1322
rect 39492 1264 39578 1320
rect 39634 1264 40000 1320
rect 39492 1262 40000 1264
rect 0 1232 480 1260
rect 39520 1232 40000 1262
rect 13629 1186 13695 1189
rect 9630 1184 13695 1186
rect 9630 1128 13634 1184
rect 13690 1128 13695 1184
rect 9630 1126 13695 1128
rect 54 988 60 1052
rect 124 1050 130 1052
rect 9630 1050 9690 1126
rect 13629 1123 13695 1126
rect 30741 1186 30807 1189
rect 38193 1186 38259 1189
rect 30741 1184 38259 1186
rect 30741 1128 30746 1184
rect 30802 1128 38198 1184
rect 38254 1128 38259 1184
rect 30741 1126 38259 1128
rect 30741 1123 30807 1126
rect 38193 1123 38259 1126
rect 124 990 9690 1050
rect 124 988 130 990
rect 2313 778 2379 781
rect 62 776 2379 778
rect 62 720 2318 776
rect 2374 720 2379 776
rect 62 718 2379 720
rect 62 536 122 718
rect 2313 715 2379 718
rect 0 416 480 536
rect 39520 508 40000 536
rect 39520 506 39620 508
rect 39492 446 39620 506
rect 39520 444 39620 446
rect 39684 444 40000 508
rect 39520 416 40000 444
rect 4245 370 4311 373
rect 39246 370 39252 372
rect 4245 368 39252 370
rect 4245 312 4250 368
rect 4306 312 39252 368
rect 4245 310 39252 312
rect 4245 307 4311 310
rect 39246 308 39252 310
rect 39316 308 39322 372
rect 25957 234 26023 237
rect 39573 234 39639 237
rect 25957 232 39639 234
rect 25957 176 25962 232
rect 26018 176 39578 232
rect 39634 176 39639 232
rect 25957 174 39639 176
rect 25957 171 26023 174
rect 39573 171 39639 174
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 60 6836 124 6900
rect 60 6564 124 6628
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 60 6020 124 6084
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 60 5748 124 5812
rect 39620 5748 39684 5812
rect 39620 5476 39684 5540
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 23428 3300 23492 3364
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 39620 3028 39684 3092
rect 39620 2756 39684 2820
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 4108 2348 4172 2412
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
rect 60 1260 124 1324
rect 60 988 124 1052
rect 39620 444 39684 508
rect 39252 308 39316 372
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 59 6900 125 6901
rect 59 6836 60 6900
rect 124 6836 125 6900
rect 59 6835 125 6836
rect 62 6629 122 6835
rect 59 6628 125 6629
rect 59 6564 60 6628
rect 124 6564 125 6628
rect 59 6563 125 6564
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 59 6084 125 6085
rect 59 6020 60 6084
rect 124 6020 125 6084
rect 59 6019 125 6020
rect 62 5813 122 6019
rect 59 5812 125 5813
rect 59 5748 60 5812
rect 124 5748 125 5812
rect 59 5747 125 5748
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 23427 3364 23493 3365
rect 23427 3300 23428 3364
rect 23492 3300 23493 3364
rect 23427 3299 23493 3300
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 23430 2498 23490 3299
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 2128 27930 2688
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 39619 5812 39685 5813
rect 39619 5748 39620 5812
rect 39684 5748 39685 5812
rect 39619 5747 39685 5748
rect 39622 5541 39682 5747
rect 39619 5540 39685 5541
rect 39619 5476 39620 5540
rect 39684 5476 39685 5540
rect 39619 5475 39685 5476
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 39619 3092 39685 3093
rect 39619 3028 39620 3092
rect 39684 3028 39685 3092
rect 39619 3027 39685 3028
rect 39622 2821 39682 3027
rect 39619 2820 39685 2821
rect 39619 2756 39620 2820
rect 39684 2756 39685 2820
rect 39619 2755 39685 2756
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
rect 59 1324 125 1325
rect 59 1260 60 1324
rect 124 1260 125 1324
rect 59 1259 125 1260
rect 62 1053 122 1259
rect 59 1052 125 1053
rect 59 988 60 1052
rect 124 988 125 1052
rect 59 987 125 988
rect 39619 508 39685 509
rect 39619 444 39620 508
rect 39684 444 39685 508
rect 39619 443 39685 444
rect 39251 372 39317 373
rect 39251 308 39252 372
rect 39316 370 39317 372
rect 39622 370 39682 443
rect 39316 310 39682 370
rect 39316 308 39317 310
rect 39251 307 39317 308
<< via4 >>
rect 4022 2412 4258 2498
rect 4022 2348 4108 2412
rect 4108 2348 4172 2412
rect 4172 2348 4258 2412
rect 4022 2262 4258 2348
rect 23342 2262 23578 2498
<< metal5 >>
rect 3980 2498 23620 2540
rect 3980 2262 4022 2498
rect 4258 2262 23342 2498
rect 23578 2262 23620 2498
rect 3980 2220 23620 2262
use scs8hd_decap_3  FILLER_1_8 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_8 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__050__B tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_13 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_16 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__049__D
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__C
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_nor4_4  _049_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__B
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_19
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__044__D
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__044__B
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _045_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_53 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_49
timestamp 1586364061
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_45
timestamp 1586364061
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__044__C
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_47
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_59
timestamp 1586364061
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_67
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _043_
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__D
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _037_
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_78
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_74
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__037__A
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_nor4_4  _056_
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 1602 592
use scs8hd_decap_8  FILLER_1_96
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_92
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_104
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__041__A
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use scs8hd_or2_4  _076_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 682 592
use scs8hd_inv_8  _041_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_117
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__038__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__039__A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _039_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_128
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _064_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__C
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_or4_4  _042_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__B
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_159
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__D
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _055_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_or4_4  _054_
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_167
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_163
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__D
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_176
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 866 592
use scs8hd_nor4_4  _068_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_180
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_201
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_198
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_205
timestamp 1586364061
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_202
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__C
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_209
timestamp 1586364061
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__D
timestamp 1586364061
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_213
timestamp 1586364061
transform 1 0 20700 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__C
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__D
timestamp 1586364061
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use scs8hd_nor4_4  _083_
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 1602 592
use scs8hd_nor4_4  _084_
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__D
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__D
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__D
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__D
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_nor4_4  _085_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1602 592
use scs8hd_nor4_4  _082_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25392 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_266
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_262
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_266
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_270
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_270
timestamp 1586364061
transform 1 0 25944 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 25760 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 26128 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 26496 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_284
timestamp 1586364061
transform 1 0 27232 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_278
timestamp 1586364061
transform 1 0 26680 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 26220 0 1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_288
timestamp 1586364061
transform 1 0 27600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_292
timestamp 1586364061
transform 1 0 27968 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_291
timestamp 1586364061
transform 1 0 27876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27784 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 28060 0 -1 2720
box -38 -48 222 592
use scs8hd_conb_1  _097_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_296
timestamp 1586364061
transform 1 0 28336 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_295
timestamp 1586364061
transform 1 0 28244 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_300
timestamp 1586364061
transform 1 0 28704 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28520 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__C
timestamp 1586364061
transform 1 0 28428 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28612 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_302
timestamp 1586364061
transform 1 0 28888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_306
timestamp 1586364061
transform 1 0 29256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_321
timestamp 1586364061
transform 1 0 30636 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_315
timestamp 1586364061
transform 1 0 30084 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_320
timestamp 1586364061
transform 1 0 30544 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _091_
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_0_329
timestamp 1586364061
transform 1 0 31372 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_325
timestamp 1586364061
transform 1 0 31004 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31188 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_336
timestamp 1586364061
transform 1 0 32016 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_332
timestamp 1586364061
transform 1 0 31648 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_337
timestamp 1586364061
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_333
timestamp 1586364061
transform 1 0 31740 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 32108 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31464 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30820 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _088_
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33396 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_351
timestamp 1586364061
transform 1 0 33396 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_1_339
timestamp 1586364061
transform 1 0 32292 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_349
timestamp 1586364061
transform 1 0 33212 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_353
timestamp 1586364061
transform 1 0 33580 0 1 2720
box -38 -48 1142 592
use scs8hd_conb_1  _096_
timestamp 1586364061
transform 1 0 34132 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_362
timestamp 1586364061
transform 1 0 34408 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_370
timestamp 1586364061
transform 1 0 35144 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_365
timestamp 1586364061
transform 1 0 34684 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__050__D
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__C
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_8
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_12
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__052__C
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__B
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_22
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_26
timestamp 1586364061
transform 1 0 3496 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 590 592
use scs8hd_nor4_4  _044_
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_38
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_62
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_70
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__C
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__C
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_1  _060_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 10120 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_96
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_100
timestamp 1586364061
transform 1 0 10304 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_8  _038_
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__C
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_118
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_8  _053_
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__D
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__D
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_133
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 314 592
use scs8hd_or4_4  _066_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__054__D
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _070_
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_175
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_195
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_conb_1  _095_
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__D
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__C
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__D
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _079_
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_2_249
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_253
timestamp 1586364061
transform 1 0 24380 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_257
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_267
timestamp 1586364061
transform 1 0 25668 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_271
timestamp 1586364061
transform 1 0 26036 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28244 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_287
timestamp 1586364061
transform 1 0 27508 0 -1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30268 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29900 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29256 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_304
timestamp 1586364061
transform 1 0 29072 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_308
timestamp 1586364061
transform 1 0 29440 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_315
timestamp 1586364061
transform 1 0 30084 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_328
timestamp 1586364061
transform 1 0 31280 0 -1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33120 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_346
timestamp 1586364061
transform 1 0 32936 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_350
timestamp 1586364061
transform 1 0 33304 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_362
timestamp 1586364061
transform 1 0 34408 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_374
timestamp 1586364061
transform 1 0 35512 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_386
timestamp 1586364061
transform 1 0 36616 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_394
timestamp 1586364061
transform 1 0 37352 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_nor4_4  _052_
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 1602 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__D
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_10
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_35
timestamp 1586364061
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__B
timestamp 1586364061
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_48
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_52
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_56
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__D
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_60
timestamp 1586364061
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__046__C
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_67
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _057_
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__C
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__D
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_96
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_100
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_104
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _061_
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_nor4_4  _063_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_108
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_140
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 406 592
use scs8hd_nor4_4  _072_
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__C
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__C
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_146
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_150
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_154
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _073_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__C
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_201
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_224
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_231
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__D
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_256
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_260
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_267
timestamp 1586364061
transform 1 0 25668 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_271
timestamp 1586364061
transform 1 0 26036 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27692 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_287
timestamp 1586364061
transform 1 0 27508 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_291
timestamp 1586364061
transform 1 0 27876 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_295
timestamp 1586364061
transform 1 0 28244 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30268 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_309
timestamp 1586364061
transform 1 0 29532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_313
timestamp 1586364061
transform 1 0 29900 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31280 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_326
timestamp 1586364061
transform 1 0 31096 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_nor4_4  _050_
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 1602 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__051__D
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_35
timestamp 1586364061
transform 1 0 4324 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _046_
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_39
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_61
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_69
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__057__D
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use scs8hd_nor4_4  _059_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_nor4_4  _062_
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__058__D
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_115
timestamp 1586364061
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_140
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__D
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__C
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_160
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _071_
timestamp 1586364061
transform 1 0 16192 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__071__C
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _074_
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_181
timestamp 1586364061
transform 1 0 17756 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_185
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _078_
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 1602 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 21344 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_218
timestamp 1586364061
transform 1 0 21160 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_222
timestamp 1586364061
transform 1 0 21528 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_226
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_266
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 26956 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27324 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_279
timestamp 1586364061
transform 1 0 26772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_283
timestamp 1586364061
transform 1 0 27140 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27508 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_296
timestamp 1586364061
transform 1 0 28336 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 29072 0 -1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30636 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_313
timestamp 1586364061
transform 1 0 29900 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_nor4_4  _051_
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1602 592
use scs8hd_buf_2  _101_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_32
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _092_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_65
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_69
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_103
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_107
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _048_
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use scs8hd_nor4_4  _058_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_140
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_144
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_or2_4  _081_
timestamp 1586364061
transform 1 0 16468 0 1 4896
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__D
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_163
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__C
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_199
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_218
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__C
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_235
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_239
timestamp 1586364061
transform 1 0 23092 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_248
timestamp 1586364061
transform 1 0 23920 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_252
timestamp 1586364061
transform 1 0 24288 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_265
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26864 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 27232 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_5_278
timestamp 1586364061
transform 1 0 26680 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_282
timestamp 1586364061
transform 1 0 27048 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27416 0 1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_5_295
timestamp 1586364061
transform 1 0 28244 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_303
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_342
timestamp 1586364061
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 35420 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_377
timestamp 1586364061
transform 1 0 35788 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_381
timestamp 1586364061
transform 1 0 36156 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_393
timestamp 1586364061
transform 1 0 37260 0 1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_5_405
timestamp 1586364061
transform 1 0 38364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_8
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__051__C
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__B
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_30
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_43
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_51
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_47
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_63
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_101
timestamp 1586364061
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_115
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_112
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__058__C
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__040__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_buf_1  _040_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_130
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_126
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_168
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_164
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_175
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_171
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_189
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_191
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_193
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__D
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_212
timestamp 1586364061
transform 1 0 20608 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_226
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_230
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_225
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_229
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_6_247
timestamp 1586364061
transform 1 0 23828 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_243
timestamp 1586364061
transform 1 0 23460 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_conb_1  _093_
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_262
timestamp 1586364061
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_266
timestamp 1586364061
transform 1 0 25576 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_252
timestamp 1586364061
transform 1 0 24288 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_256
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _087_
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_285
timestamp 1586364061
transform 1 0 27324 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_281
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27508 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27876 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_289
timestamp 1586364061
transform 1 0 27692 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_293
timestamp 1586364061
transform 1 0 28060 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_293
timestamp 1586364061
transform 1 0 28060 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_305
timestamp 1586364061
transform 1 0 29164 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_317
timestamp 1586364061
transform 1 0 30268 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_329
timestamp 1586364061
transform 1 0 31372 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_335
timestamp 1586364061
transform 1 0 31924 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_330
timestamp 1586364061
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_349
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_354
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 35420 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_361
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_375
timestamp 1586364061
transform 1 0 35604 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_387
timestamp 1586364061
transform 1 0 36708 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_399
timestamp 1586364061
transform 1 0 37812 0 1 5984
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _094_
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_76
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_108
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_112
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_124
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_128
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_132
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_1  _067_
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_228
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_240
timestamp 1586364061
transform 1 0 23184 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_244
timestamp 1586364061
transform 1 0 23552 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_8  _086_
timestamp 1586364061
transform 1 0 24288 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_261
timestamp 1586364061
transform 1 0 25116 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_265
timestamp 1586364061
transform 1 0 25484 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_273
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_288
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_300
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_377
timestamp 1586364061
transform 1 0 35788 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_389
timestamp 1586364061
transform 1 0 36892 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_17
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_30
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_47
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_55
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_97
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_102
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_106
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_131
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_165
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_192
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_198
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_202
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_209
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_213
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_281
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_293
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_318
timestamp 1586364061
transform 1 0 30360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_330
timestamp 1586364061
transform 1 0 31464 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_342
timestamp 1586364061
transform 1 0 32568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_354
timestamp 1586364061
transform 1 0 33672 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 35420 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 35236 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 406 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 36524 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 37076 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 35972 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_377
timestamp 1586364061
transform 1 0 35788 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_381
timestamp 1586364061
transform 1 0 36156 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_389
timestamp 1586364061
transform 1 0 36892 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_393
timestamp 1586364061
transform 1 0 37260 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_405
timestamp 1586364061
transform 1 0 38364 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_52
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_98
timestamp 1586364061
transform 1 0 10120 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_122
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_134
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_199
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_288
timestamp 1586364061
transform 1 0 27600 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_300
timestamp 1586364061
transform 1 0 28704 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_312
timestamp 1586364061
transform 1 0 29808 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_349
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 35420 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_361
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_377
timestamp 1586364061
transform 1 0 35788 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_389
timestamp 1586364061
transform 1 0 36892 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_18
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_22
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_44
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_281
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_293
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_318
timestamp 1586364061
transform 1 0 30360 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_330
timestamp 1586364061
transform 1 0 31464 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_342
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_354
timestamp 1586364061
transform 1 0 33672 0 1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 35420 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 35236 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_367
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 35972 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_377
timestamp 1586364061
transform 1 0 35788 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_381
timestamp 1586364061
transform 1 0 36156 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_393
timestamp 1586364061
transform 1 0 37260 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_11_405
timestamp 1586364061
transform 1 0 38364 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_300
timestamp 1586364061
transform 1 0 28704 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_324
timestamp 1586364061
transform 1 0 30912 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_349
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_361
timestamp 1586364061
transform 1 0 34316 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_377
timestamp 1586364061
transform 1 0 35788 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_389
timestamp 1586364061
transform 1 0 36892 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_293
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_288
timestamp 1586364061
transform 1 0 27600 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_300
timestamp 1586364061
transform 1 0 28704 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_318
timestamp 1586364061
transform 1 0 30360 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_312
timestamp 1586364061
transform 1 0 29808 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_330
timestamp 1586364061
transform 1 0 31464 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_324
timestamp 1586364061
transform 1 0 30912 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_342
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_354
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 35420 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 35420 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_361
timestamp 1586364061
transform 1 0 34316 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_375
timestamp 1586364061
transform 1 0 35604 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_387
timestamp 1586364061
transform 1 0 36708 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_377
timestamp 1586364061
transform 1 0 35788 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_389
timestamp 1586364061
transform 1 0 36892 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_399
timestamp 1586364061
transform 1 0 37812 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_43
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_318
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_342
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_354
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 35420 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_15_375
timestamp 1586364061
transform 1 0 35604 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_387
timestamp 1586364061
transform 1 0 36708 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_399
timestamp 1586364061
transform 1 0 37812 0 1 10336
box -38 -48 774 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_288
timestamp 1586364061
transform 1 0 27600 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_300
timestamp 1586364061
transform 1 0 28704 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_312
timestamp 1586364061
transform 1 0 29808 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_324
timestamp 1586364061
transform 1 0 30912 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_349
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_361
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_377
timestamp 1586364061
transform 1 0 35788 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_389
timestamp 1586364061
transform 1 0 36892 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_281
timestamp 1586364061
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_293
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_342
timestamp 1586364061
transform 1 0 32568 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_379
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_391
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_403
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_373
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_385
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_293
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_354
timestamp 1586364061
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_379
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_391
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_403
timestamp 1586364061
transform 1 0 38180 0 1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 5354 0 5410 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 9034 0 9090 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 12622 0 12678 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 16302 0 16358 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 19890 0 19946 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 23570 0 23626 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 30838 0 30894 480 6 bottom_grid_pin_0_
port 6 nsew default tristate
rlabel metal2 s 34426 0 34482 480 6 bottom_grid_pin_4_
port 7 nsew default tristate
rlabel metal2 s 38106 0 38162 480 6 bottom_grid_pin_8_
port 8 nsew default tristate
rlabel metal3 s 0 416 480 536 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal3 s 0 1232 480 1352 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal3 s 0 2184 480 2304 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 0 10208 480 10328 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal3 s 39520 416 40000 536 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 39520 1232 40000 1352 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal3 s 39520 2184 40000 2304 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal3 s 39520 3000 40000 3120 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 39520 3952 40000 4072 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal3 s 39520 4768 40000 4888 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 39520 5720 40000 5840 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal3 s 39520 6536 40000 6656 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 39520 7488 40000 7608 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal3 s 39520 8440 40000 8560 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal3 s 39520 9256 40000 9376 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal3 s 39520 10208 40000 10328 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 39520 11024 40000 11144 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 39520 11976 40000 12096 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal3 s 39520 12792 40000 12912 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal3 s 39520 13744 40000 13864 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 39520 14560 40000 14680 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal3 s 39520 15512 40000 15632 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 27158 0 27214 480 6 data_in
port 45 nsew default input
rlabel metal2 s 1766 0 1822 480 6 enable
port 46 nsew default input
rlabel metal2 s 33322 15520 33378 16000 6 top_grid_pin_14_
port 47 nsew default tristate
rlabel metal2 s 6642 15520 6698 16000 6 top_grid_pin_2_
port 48 nsew default tristate
rlabel metal2 s 19982 15520 20038 16000 6 top_grid_pin_6_
port 49 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 50 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 51 nsew default input
<< end >>
