magic
tech sky130A
magscale 1 2
timestamp 1606225941
<< locali >>
rect 10333 18539 10367 18709
rect 12265 18471 12299 18777
rect 11989 16839 12023 17145
rect 12173 14119 12207 14357
rect 15025 12487 15059 12657
rect 15761 7727 15795 7829
<< viali >>
rect 5089 19865 5123 19899
rect 18797 19865 18831 19899
rect 19349 19865 19383 19899
rect 20085 19865 20119 19899
rect 20637 19865 20671 19899
rect 4997 19797 5031 19831
rect 8493 19729 8527 19763
rect 18613 19729 18647 19763
rect 19165 19729 19199 19763
rect 19901 19729 19935 19763
rect 20453 19729 20487 19763
rect 5181 19661 5215 19695
rect 8585 19661 8619 19695
rect 8677 19661 8711 19695
rect 17233 19661 17267 19695
rect 4629 19525 4663 19559
rect 8125 19525 8159 19559
rect 16865 19253 16899 19287
rect 8677 19185 8711 19219
rect 10425 19185 10459 19219
rect 11897 19185 11931 19219
rect 16497 19185 16531 19219
rect 17509 19185 17543 19219
rect 18153 19185 18187 19219
rect 20269 19185 20303 19219
rect 4077 19117 4111 19151
rect 4344 19117 4378 19151
rect 7021 19117 7055 19151
rect 10333 19117 10367 19151
rect 13093 19117 13127 19151
rect 16313 19117 16347 19151
rect 17233 19117 17267 19151
rect 17877 19117 17911 19151
rect 18797 19117 18831 19151
rect 19349 19117 19383 19151
rect 20085 19117 20119 19151
rect 7288 19049 7322 19083
rect 11805 19049 11839 19083
rect 13360 19049 13394 19083
rect 17325 19049 17359 19083
rect 19625 19049 19659 19083
rect 5457 18981 5491 19015
rect 8401 18981 8435 19015
rect 9873 18981 9907 19015
rect 10241 18981 10275 19015
rect 11345 18981 11379 19015
rect 11713 18981 11747 19015
rect 14473 18981 14507 19015
rect 15853 18981 15887 19015
rect 16221 18981 16255 19015
rect 18981 18981 19015 19015
rect 3801 18777 3835 18811
rect 5181 18777 5215 18811
rect 8217 18777 8251 18811
rect 11805 18777 11839 18811
rect 12265 18777 12299 18811
rect 13829 18777 13863 18811
rect 15945 18777 15979 18811
rect 20729 18777 20763 18811
rect 9014 18709 9048 18743
rect 10333 18709 10367 18743
rect 10670 18709 10704 18743
rect 2688 18641 2722 18675
rect 5089 18641 5123 18675
rect 5733 18641 5767 18675
rect 6837 18641 6871 18675
rect 7104 18641 7138 18675
rect 8769 18641 8803 18675
rect 2421 18573 2455 18607
rect 5365 18573 5399 18607
rect 10425 18573 10459 18607
rect 10149 18505 10183 18539
rect 10333 18505 10367 18539
rect 12694 18709 12728 18743
rect 14810 18709 14844 18743
rect 16488 18709 16522 18743
rect 19625 18709 19659 18743
rect 14565 18641 14599 18675
rect 16221 18641 16255 18675
rect 18245 18641 18279 18675
rect 18521 18641 18555 18675
rect 19349 18641 19383 18675
rect 20545 18641 20579 18675
rect 12449 18573 12483 18607
rect 14105 18573 14139 18607
rect 4721 18437 4755 18471
rect 12265 18437 12299 18471
rect 17601 18437 17635 18471
rect 7941 18233 7975 18267
rect 14197 18233 14231 18267
rect 12909 18165 12943 18199
rect 8493 18097 8527 18131
rect 11713 18097 11747 18131
rect 13369 18097 13403 18131
rect 13553 18097 13587 18131
rect 14749 18097 14783 18131
rect 5181 18029 5215 18063
rect 8401 18029 8435 18063
rect 14565 18029 14599 18063
rect 20269 18029 20303 18063
rect 5457 17961 5491 17995
rect 13277 17961 13311 17995
rect 14657 17961 14691 17995
rect 8309 17893 8343 17927
rect 20453 17893 20487 17927
rect 2973 17689 3007 17723
rect 19625 17689 19659 17723
rect 5356 17621 5390 17655
rect 1593 17553 1627 17587
rect 1860 17553 1894 17587
rect 19441 17553 19475 17587
rect 19993 17553 20027 17587
rect 20545 17553 20579 17587
rect 3341 17485 3375 17519
rect 5089 17485 5123 17519
rect 6469 17349 6503 17383
rect 20177 17349 20211 17383
rect 20729 17349 20763 17383
rect 9689 17145 9723 17179
rect 11989 17145 12023 17179
rect 17693 17145 17727 17179
rect 3525 17009 3559 17043
rect 4537 17009 4571 17043
rect 4629 17009 4663 17043
rect 7481 17009 7515 17043
rect 8677 17009 8711 17043
rect 10241 17009 10275 17043
rect 11713 17009 11747 17043
rect 3341 16941 3375 16975
rect 4445 16941 4479 16975
rect 7205 16941 7239 16975
rect 8585 16941 8619 16975
rect 11621 16941 11655 16975
rect 10149 16873 10183 16907
rect 12173 17077 12207 17111
rect 12725 17009 12759 17043
rect 14565 17009 14599 17043
rect 15945 17009 15979 17043
rect 18245 17009 18279 17043
rect 19625 17009 19659 17043
rect 20361 17009 20395 17043
rect 14473 16941 14507 16975
rect 16212 16941 16246 16975
rect 19349 16941 19383 16975
rect 20085 16941 20119 16975
rect 12633 16873 12667 16907
rect 18061 16873 18095 16907
rect 18705 16873 18739 16907
rect 2973 16805 3007 16839
rect 3433 16805 3467 16839
rect 4077 16805 4111 16839
rect 8125 16805 8159 16839
rect 8493 16805 8527 16839
rect 10057 16805 10091 16839
rect 11161 16805 11195 16839
rect 11529 16805 11563 16839
rect 11989 16805 12023 16839
rect 12541 16805 12575 16839
rect 14013 16805 14047 16839
rect 14381 16805 14415 16839
rect 17325 16805 17359 16839
rect 18153 16805 18187 16839
rect 6837 16601 6871 16635
rect 7297 16601 7331 16635
rect 9597 16601 9631 16635
rect 11253 16601 11287 16635
rect 11897 16601 11931 16635
rect 15025 16601 15059 16635
rect 20729 16601 20763 16635
rect 8484 16533 8518 16567
rect 10140 16533 10174 16567
rect 19625 16533 19659 16567
rect 3893 16465 3927 16499
rect 4169 16465 4203 16499
rect 6285 16465 6319 16499
rect 7205 16465 7239 16499
rect 12889 16465 12923 16499
rect 14933 16465 14967 16499
rect 15577 16465 15611 16499
rect 16313 16465 16347 16499
rect 16580 16465 16614 16499
rect 19349 16465 19383 16499
rect 20545 16465 20579 16499
rect 7389 16397 7423 16431
rect 8217 16397 8251 16431
rect 9873 16397 9907 16431
rect 12633 16397 12667 16431
rect 15117 16397 15151 16431
rect 14013 16329 14047 16363
rect 14565 16329 14599 16363
rect 17693 16261 17727 16295
rect 3157 16057 3191 16091
rect 7113 16057 7147 16091
rect 12541 16057 12575 16091
rect 16773 16057 16807 16091
rect 19901 16057 19935 16091
rect 6837 15989 6871 16023
rect 20453 15989 20487 16023
rect 5457 15921 5491 15955
rect 7665 15921 7699 15955
rect 9873 15921 9907 15955
rect 11161 15921 11195 15955
rect 13553 15921 13587 15955
rect 17325 15921 17359 15955
rect 1777 15853 1811 15887
rect 5724 15853 5758 15887
rect 7573 15853 7607 15887
rect 13820 15853 13854 15887
rect 17233 15853 17267 15887
rect 19717 15853 19751 15887
rect 20269 15853 20303 15887
rect 2044 15785 2078 15819
rect 11428 15785 11462 15819
rect 17141 15785 17175 15819
rect 7481 15717 7515 15751
rect 14933 15717 14967 15751
rect 2973 15513 3007 15547
rect 6285 15513 6319 15547
rect 20729 15513 20763 15547
rect 19165 15445 19199 15479
rect 19901 15445 19935 15479
rect 3341 15377 3375 15411
rect 3985 15377 4019 15411
rect 4905 15377 4939 15411
rect 5172 15377 5206 15411
rect 16589 15377 16623 15411
rect 18889 15377 18923 15411
rect 19625 15377 19659 15411
rect 20545 15377 20579 15411
rect 3433 15309 3467 15343
rect 3525 15309 3559 15343
rect 16681 15309 16715 15343
rect 16773 15309 16807 15343
rect 16221 15173 16255 15207
rect 2973 14969 3007 15003
rect 4077 14969 4111 15003
rect 9321 14969 9355 15003
rect 9689 14969 9723 15003
rect 16129 14969 16163 15003
rect 20453 14969 20487 15003
rect 12265 14901 12299 14935
rect 1593 14833 1627 14867
rect 4629 14833 4663 14867
rect 10241 14833 10275 14867
rect 12817 14833 12851 14867
rect 16589 14833 16623 14867
rect 16773 14833 16807 14867
rect 4537 14765 4571 14799
rect 7205 14765 7239 14799
rect 7941 14765 7975 14799
rect 13645 14765 13679 14799
rect 18889 14765 18923 14799
rect 20269 14765 20303 14799
rect 1860 14697 1894 14731
rect 4445 14697 4479 14731
rect 8208 14697 8242 14731
rect 19165 14697 19199 14731
rect 7021 14629 7055 14663
rect 10057 14629 10091 14663
rect 10149 14629 10183 14663
rect 12633 14629 12667 14663
rect 12725 14629 12759 14663
rect 13461 14629 13495 14663
rect 16497 14629 16531 14663
rect 6101 14425 6135 14459
rect 8677 14425 8711 14459
rect 9781 14425 9815 14459
rect 12081 14425 12115 14459
rect 12449 14425 12483 14459
rect 12817 14425 12851 14459
rect 15577 14425 15611 14459
rect 17233 14425 17267 14459
rect 18705 14425 18739 14459
rect 20729 14425 20763 14459
rect 4160 14357 4194 14391
rect 7564 14357 7598 14391
rect 12173 14357 12207 14391
rect 12909 14357 12943 14391
rect 14464 14357 14498 14391
rect 16120 14357 16154 14391
rect 19349 14357 19383 14391
rect 20085 14357 20119 14391
rect 3893 14289 3927 14323
rect 6009 14289 6043 14323
rect 10957 14289 10991 14323
rect 6193 14221 6227 14255
rect 7297 14221 7331 14255
rect 10701 14221 10735 14255
rect 5273 14153 5307 14187
rect 14197 14289 14231 14323
rect 15853 14289 15887 14323
rect 18521 14289 18555 14323
rect 19073 14289 19107 14323
rect 19819 14289 19853 14323
rect 20545 14289 20579 14323
rect 13001 14221 13035 14255
rect 13461 14221 13495 14255
rect 17509 14221 17543 14255
rect 5641 14085 5675 14119
rect 12173 14085 12207 14119
rect 3709 13881 3743 13915
rect 6193 13881 6227 13915
rect 6469 13881 6503 13915
rect 8033 13881 8067 13915
rect 11253 13881 11287 13915
rect 12725 13881 12759 13915
rect 16589 13881 16623 13915
rect 20453 13881 20487 13915
rect 19901 13813 19935 13847
rect 2329 13745 2363 13779
rect 6929 13745 6963 13779
rect 7021 13745 7055 13779
rect 8493 13745 8527 13779
rect 8677 13745 8711 13779
rect 13277 13745 13311 13779
rect 17141 13745 17175 13779
rect 18429 13745 18463 13779
rect 2596 13677 2630 13711
rect 4813 13677 4847 13711
rect 5080 13677 5114 13711
rect 9229 13677 9263 13711
rect 9873 13677 9907 13711
rect 13093 13677 13127 13711
rect 16957 13677 16991 13711
rect 18153 13677 18187 13711
rect 19717 13677 19751 13711
rect 20269 13677 20303 13711
rect 8401 13609 8435 13643
rect 10140 13609 10174 13643
rect 13185 13609 13219 13643
rect 17049 13609 17083 13643
rect 6837 13541 6871 13575
rect 9045 13541 9079 13575
rect 6101 13337 6135 13371
rect 11437 13337 11471 13371
rect 19717 13337 19751 13371
rect 20729 13337 20763 13371
rect 10149 13269 10183 13303
rect 14105 13201 14139 13235
rect 19533 13201 19567 13235
rect 20545 13201 20579 13235
rect 14197 13133 14231 13167
rect 14289 13133 14323 13167
rect 13737 12997 13771 13031
rect 13185 12793 13219 12827
rect 19901 12793 19935 12827
rect 20453 12793 20487 12827
rect 7665 12725 7699 12759
rect 9873 12725 9907 12759
rect 14197 12725 14231 12759
rect 7113 12657 7147 12691
rect 7297 12657 7331 12691
rect 8217 12657 8251 12691
rect 10333 12657 10367 12691
rect 10425 12657 10459 12691
rect 11161 12657 11195 12691
rect 13645 12657 13679 12691
rect 13737 12657 13771 12691
rect 14749 12657 14783 12691
rect 15025 12657 15059 12691
rect 15577 12657 15611 12691
rect 18981 12657 19015 12691
rect 7021 12589 7055 12623
rect 10885 12589 10919 12623
rect 12909 12589 12943 12623
rect 8125 12521 8159 12555
rect 15301 12589 15335 12623
rect 16129 12589 16163 12623
rect 18705 12589 18739 12623
rect 19717 12589 19751 12623
rect 20269 12589 20303 12623
rect 16396 12521 16430 12555
rect 6653 12453 6687 12487
rect 8033 12453 8067 12487
rect 10241 12453 10275 12487
rect 12725 12453 12759 12487
rect 13553 12453 13587 12487
rect 14565 12453 14599 12487
rect 14657 12453 14691 12487
rect 15025 12453 15059 12487
rect 17509 12453 17543 12487
rect 10425 12249 10459 12283
rect 14473 12249 14507 12283
rect 18061 12249 18095 12283
rect 20177 12249 20211 12283
rect 20729 12249 20763 12283
rect 10793 12181 10827 12215
rect 11437 12181 11471 12215
rect 12716 12181 12750 12215
rect 14841 12181 14875 12215
rect 18429 12181 18463 12215
rect 7104 12113 7138 12147
rect 8944 12113 8978 12147
rect 10885 12113 10919 12147
rect 16580 12113 16614 12147
rect 19993 12113 20027 12147
rect 20545 12113 20579 12147
rect 6837 12045 6871 12079
rect 8677 12045 8711 12079
rect 10977 12045 11011 12079
rect 12449 12045 12483 12079
rect 14933 12045 14967 12079
rect 15117 12045 15151 12079
rect 16313 12045 16347 12079
rect 18521 12045 18555 12079
rect 18613 12045 18647 12079
rect 8217 11977 8251 12011
rect 10057 11977 10091 12011
rect 17693 11977 17727 12011
rect 13829 11909 13863 11943
rect 7941 11705 7975 11739
rect 13829 11705 13863 11739
rect 14105 11705 14139 11739
rect 18613 11705 18647 11739
rect 20453 11705 20487 11739
rect 8493 11569 8527 11603
rect 14657 11569 14691 11603
rect 16589 11569 16623 11603
rect 16681 11569 16715 11603
rect 19165 11569 19199 11603
rect 8401 11501 8435 11535
rect 11069 11501 11103 11535
rect 14013 11501 14047 11535
rect 20269 11501 20303 11535
rect 8309 11433 8343 11467
rect 11345 11433 11379 11467
rect 14473 11433 14507 11467
rect 15301 11433 15335 11467
rect 16497 11433 16531 11467
rect 18981 11433 19015 11467
rect 19625 11433 19659 11467
rect 14565 11365 14599 11399
rect 16129 11365 16163 11399
rect 19073 11365 19107 11399
rect 16865 11161 16899 11195
rect 19165 11161 19199 11195
rect 20729 11161 20763 11195
rect 8585 11025 8619 11059
rect 16773 11025 16807 11059
rect 19533 11025 19567 11059
rect 20545 11025 20579 11059
rect 17049 10957 17083 10991
rect 19625 10957 19659 10991
rect 19809 10957 19843 10991
rect 8401 10889 8435 10923
rect 16405 10889 16439 10923
rect 8033 10617 8067 10651
rect 10333 10617 10367 10651
rect 14473 10617 14507 10651
rect 16497 10617 16531 10651
rect 18521 10617 18555 10651
rect 20453 10617 20487 10651
rect 10885 10481 10919 10515
rect 11805 10481 11839 10515
rect 11989 10481 12023 10515
rect 13093 10481 13127 10515
rect 17141 10481 17175 10515
rect 19165 10481 19199 10515
rect 6653 10413 6687 10447
rect 6920 10413 6954 10447
rect 13360 10413 13394 10447
rect 20269 10413 20303 10447
rect 11713 10345 11747 10379
rect 16865 10345 16899 10379
rect 10701 10277 10735 10311
rect 10793 10277 10827 10311
rect 11345 10277 11379 10311
rect 16957 10277 16991 10311
rect 18889 10277 18923 10311
rect 18981 10277 19015 10311
rect 11253 10073 11287 10107
rect 12909 10073 12943 10107
rect 15117 10073 15151 10107
rect 17417 10073 17451 10107
rect 18245 10073 18279 10107
rect 20085 10073 20119 10107
rect 20729 10073 20763 10107
rect 8484 10005 8518 10039
rect 16304 10005 16338 10039
rect 10140 9937 10174 9971
rect 12817 9937 12851 9971
rect 13737 9937 13771 9971
rect 14004 9937 14038 9971
rect 18705 9937 18739 9971
rect 18972 9937 19006 9971
rect 20545 9937 20579 9971
rect 8217 9869 8251 9903
rect 9873 9869 9907 9903
rect 11529 9869 11563 9903
rect 13001 9869 13035 9903
rect 16037 9869 16071 9903
rect 9597 9801 9631 9835
rect 12449 9801 12483 9835
rect 18429 9529 18463 9563
rect 11161 9461 11195 9495
rect 13737 9461 13771 9495
rect 15485 9461 15519 9495
rect 20453 9461 20487 9495
rect 11805 9393 11839 9427
rect 13093 9393 13127 9427
rect 19073 9393 19107 9427
rect 11621 9325 11655 9359
rect 12909 9325 12943 9359
rect 13553 9325 13587 9359
rect 15301 9325 15335 9359
rect 18797 9325 18831 9359
rect 20269 9325 20303 9359
rect 11529 9257 11563 9291
rect 12541 9189 12575 9223
rect 13001 9189 13035 9223
rect 18889 9189 18923 9223
rect 10977 8985 11011 9019
rect 11345 8985 11379 9019
rect 20729 8985 20763 9019
rect 11437 8917 11471 8951
rect 15577 8917 15611 8951
rect 15301 8849 15335 8883
rect 20545 8849 20579 8883
rect 11621 8781 11655 8815
rect 11437 8441 11471 8475
rect 16129 8441 16163 8475
rect 19625 8441 19659 8475
rect 20453 8373 20487 8407
rect 13461 8305 13495 8339
rect 16773 8305 16807 8339
rect 11253 8237 11287 8271
rect 13185 8237 13219 8271
rect 18245 8237 18279 8271
rect 20269 8237 20303 8271
rect 16497 8169 16531 8203
rect 17141 8169 17175 8203
rect 18512 8169 18546 8203
rect 13921 8101 13955 8135
rect 16589 8101 16623 8135
rect 13185 7897 13219 7931
rect 13553 7897 13587 7931
rect 19441 7897 19475 7931
rect 20729 7897 20763 7931
rect 10977 7829 11011 7863
rect 15761 7829 15795 7863
rect 18306 7829 18340 7863
rect 9312 7761 9346 7795
rect 10701 7761 10735 7795
rect 14453 7761 14487 7795
rect 16120 7761 16154 7795
rect 18061 7761 18095 7795
rect 19993 7761 20027 7795
rect 20545 7761 20579 7795
rect 9045 7693 9079 7727
rect 11437 7693 11471 7727
rect 13645 7693 13679 7727
rect 13829 7693 13863 7727
rect 14197 7693 14231 7727
rect 15761 7693 15795 7727
rect 15853 7693 15887 7727
rect 15577 7625 15611 7659
rect 17233 7625 17267 7659
rect 10425 7557 10459 7591
rect 20177 7557 20211 7591
rect 9965 7353 9999 7387
rect 14013 7353 14047 7387
rect 16589 7353 16623 7387
rect 10517 7217 10551 7251
rect 17141 7217 17175 7251
rect 10333 7149 10367 7183
rect 10977 7149 11011 7183
rect 12633 7149 12667 7183
rect 17049 7149 17083 7183
rect 11222 7081 11256 7115
rect 12900 7081 12934 7115
rect 16957 7081 16991 7115
rect 10425 7013 10459 7047
rect 12357 7013 12391 7047
rect 10517 6809 10551 6843
rect 13645 6809 13679 6843
rect 10885 6741 10919 6775
rect 14013 6741 14047 6775
rect 7737 6673 7771 6707
rect 10977 6673 11011 6707
rect 7481 6605 7515 6639
rect 11069 6605 11103 6639
rect 14105 6605 14139 6639
rect 14289 6605 14323 6639
rect 8861 6537 8895 6571
rect 14197 6265 14231 6299
rect 14013 6061 14047 6095
rect 13093 5721 13127 5755
rect 12909 5585 12943 5619
rect 20729 4633 20763 4667
rect 20545 4497 20579 4531
<< metal1 >>
rect 10318 20536 10324 20588
rect 10376 20576 10382 20588
rect 17954 20576 17960 20588
rect 10376 20548 17960 20576
rect 10376 20536 10382 20548
rect 17954 20536 17960 20548
rect 18012 20536 18018 20588
rect 1104 20010 21620 20032
rect 1104 19958 7846 20010
rect 7898 19958 7910 20010
rect 7962 19958 7974 20010
rect 8026 19958 8038 20010
rect 8090 19958 14710 20010
rect 14762 19958 14774 20010
rect 14826 19958 14838 20010
rect 14890 19958 14902 20010
rect 14954 19958 21620 20010
rect 1104 19936 21620 19958
rect 4706 19856 4712 19908
rect 4764 19896 4770 19908
rect 5077 19899 5135 19905
rect 5077 19896 5089 19899
rect 4764 19868 5089 19896
rect 4764 19856 4770 19868
rect 5077 19865 5089 19868
rect 5123 19865 5135 19899
rect 18782 19896 18788 19908
rect 18743 19868 18788 19896
rect 5077 19859 5135 19865
rect 18782 19856 18788 19868
rect 18840 19856 18846 19908
rect 19334 19896 19340 19908
rect 19295 19868 19340 19896
rect 19334 19856 19340 19868
rect 19392 19856 19398 19908
rect 20070 19896 20076 19908
rect 20031 19868 20076 19896
rect 20070 19856 20076 19868
rect 20128 19856 20134 19908
rect 20622 19896 20628 19908
rect 20583 19868 20628 19896
rect 20622 19856 20628 19868
rect 20680 19856 20686 19908
rect 4985 19831 5043 19837
rect 4985 19797 4997 19831
rect 5031 19828 5043 19831
rect 9950 19828 9956 19840
rect 5031 19800 9956 19828
rect 5031 19797 5043 19800
rect 4985 19791 5043 19797
rect 9950 19788 9956 19800
rect 10008 19788 10014 19840
rect 8478 19760 8484 19772
rect 8439 19732 8484 19760
rect 8478 19720 8484 19732
rect 8536 19720 8542 19772
rect 18598 19760 18604 19772
rect 18559 19732 18604 19760
rect 18598 19720 18604 19732
rect 18656 19720 18662 19772
rect 19150 19760 19156 19772
rect 19111 19732 19156 19760
rect 19150 19720 19156 19732
rect 19208 19720 19214 19772
rect 19889 19763 19947 19769
rect 19889 19729 19901 19763
rect 19935 19760 19947 19763
rect 20254 19760 20260 19772
rect 19935 19732 20260 19760
rect 19935 19729 19947 19732
rect 19889 19723 19947 19729
rect 20254 19720 20260 19732
rect 20312 19720 20318 19772
rect 20438 19760 20444 19772
rect 20399 19732 20444 19760
rect 20438 19720 20444 19732
rect 20496 19720 20502 19772
rect 4706 19652 4712 19704
rect 4764 19692 4770 19704
rect 5169 19695 5227 19701
rect 5169 19692 5181 19695
rect 4764 19664 5181 19692
rect 4764 19652 4770 19664
rect 5169 19661 5181 19664
rect 5215 19661 5227 19695
rect 5169 19655 5227 19661
rect 8294 19652 8300 19704
rect 8352 19692 8358 19704
rect 8573 19695 8631 19701
rect 8573 19692 8585 19695
rect 8352 19664 8585 19692
rect 8352 19652 8358 19664
rect 8573 19661 8585 19664
rect 8619 19661 8631 19695
rect 8573 19655 8631 19661
rect 8665 19695 8723 19701
rect 8665 19661 8677 19695
rect 8711 19661 8723 19695
rect 17218 19692 17224 19704
rect 17179 19664 17224 19692
rect 8665 19655 8723 19661
rect 8386 19584 8392 19636
rect 8444 19624 8450 19636
rect 8680 19624 8708 19655
rect 17218 19652 17224 19664
rect 17276 19652 17282 19704
rect 8444 19596 8708 19624
rect 8444 19584 8450 19596
rect 4617 19559 4675 19565
rect 4617 19525 4629 19559
rect 4663 19556 4675 19559
rect 5166 19556 5172 19568
rect 4663 19528 5172 19556
rect 4663 19525 4675 19528
rect 4617 19519 4675 19525
rect 5166 19516 5172 19528
rect 5224 19516 5230 19568
rect 8110 19556 8116 19568
rect 8071 19528 8116 19556
rect 8110 19516 8116 19528
rect 8168 19516 8174 19568
rect 1104 19466 21620 19488
rect 1104 19414 4414 19466
rect 4466 19414 4478 19466
rect 4530 19414 4542 19466
rect 4594 19414 4606 19466
rect 4658 19414 11278 19466
rect 11330 19414 11342 19466
rect 11394 19414 11406 19466
rect 11458 19414 11470 19466
rect 11522 19414 18142 19466
rect 18194 19414 18206 19466
rect 18258 19414 18270 19466
rect 18322 19414 18334 19466
rect 18386 19414 21620 19466
rect 1104 19392 21620 19414
rect 8110 19312 8116 19364
rect 8168 19352 8174 19364
rect 8168 19324 19380 19352
rect 8168 19312 8174 19324
rect 16853 19287 16911 19293
rect 16853 19253 16865 19287
rect 16899 19284 16911 19287
rect 16899 19256 17632 19284
rect 16899 19253 16911 19256
rect 16853 19247 16911 19253
rect 8478 19176 8484 19228
rect 8536 19216 8542 19228
rect 8665 19219 8723 19225
rect 8665 19216 8677 19219
rect 8536 19188 8677 19216
rect 8536 19176 8542 19188
rect 8665 19185 8677 19188
rect 8711 19185 8723 19219
rect 10410 19216 10416 19228
rect 10371 19188 10416 19216
rect 8665 19179 8723 19185
rect 10410 19176 10416 19188
rect 10468 19176 10474 19228
rect 11882 19216 11888 19228
rect 11843 19188 11888 19216
rect 11882 19176 11888 19188
rect 11940 19176 11946 19228
rect 16482 19216 16488 19228
rect 16443 19188 16488 19216
rect 16482 19176 16488 19188
rect 16540 19176 16546 19228
rect 17494 19216 17500 19228
rect 17455 19188 17500 19216
rect 17494 19176 17500 19188
rect 17552 19176 17558 19228
rect 2406 19108 2412 19160
rect 2464 19148 2470 19160
rect 4065 19151 4123 19157
rect 4065 19148 4077 19151
rect 2464 19120 4077 19148
rect 2464 19108 2470 19120
rect 4065 19117 4077 19120
rect 4111 19117 4123 19151
rect 4065 19111 4123 19117
rect 4332 19151 4390 19157
rect 4332 19117 4344 19151
rect 4378 19148 4390 19151
rect 4706 19148 4712 19160
rect 4378 19120 4712 19148
rect 4378 19117 4390 19120
rect 4332 19111 4390 19117
rect 4080 19080 4108 19111
rect 4706 19108 4712 19120
rect 4764 19108 4770 19160
rect 7006 19148 7012 19160
rect 6967 19120 7012 19148
rect 7006 19108 7012 19120
rect 7064 19108 7070 19160
rect 7107 19120 8340 19148
rect 5074 19080 5080 19092
rect 4080 19052 5080 19080
rect 5074 19040 5080 19052
rect 5132 19040 5138 19092
rect 6730 19040 6736 19092
rect 6788 19080 6794 19092
rect 7107 19080 7135 19120
rect 6788 19052 7135 19080
rect 7276 19083 7334 19089
rect 6788 19040 6794 19052
rect 7276 19049 7288 19083
rect 7322 19080 7334 19083
rect 8202 19080 8208 19092
rect 7322 19052 8208 19080
rect 7322 19049 7334 19052
rect 7276 19043 7334 19049
rect 8202 19040 8208 19052
rect 8260 19040 8266 19092
rect 8312 19080 8340 19120
rect 9122 19108 9128 19160
rect 9180 19148 9186 19160
rect 10321 19151 10379 19157
rect 10321 19148 10333 19151
rect 9180 19120 10333 19148
rect 9180 19108 9186 19120
rect 10321 19117 10333 19120
rect 10367 19117 10379 19151
rect 10321 19111 10379 19117
rect 12618 19108 12624 19160
rect 12676 19148 12682 19160
rect 13081 19151 13139 19157
rect 13081 19148 13093 19151
rect 12676 19120 13093 19148
rect 12676 19108 12682 19120
rect 13081 19117 13093 19120
rect 13127 19117 13139 19151
rect 13081 19111 13139 19117
rect 14366 19108 14372 19160
rect 14424 19148 14430 19160
rect 16301 19151 16359 19157
rect 16301 19148 16313 19151
rect 14424 19120 16313 19148
rect 14424 19108 14430 19120
rect 16301 19117 16313 19120
rect 16347 19117 16359 19151
rect 17218 19148 17224 19160
rect 17179 19120 17224 19148
rect 16301 19111 16359 19117
rect 17218 19108 17224 19120
rect 17276 19108 17282 19160
rect 17604 19148 17632 19256
rect 18141 19219 18199 19225
rect 18141 19185 18153 19219
rect 18187 19216 18199 19219
rect 18598 19216 18604 19228
rect 18187 19188 18604 19216
rect 18187 19185 18199 19188
rect 18141 19179 18199 19185
rect 18598 19176 18604 19188
rect 18656 19176 18662 19228
rect 17865 19151 17923 19157
rect 17865 19148 17877 19151
rect 17604 19120 17877 19148
rect 17865 19117 17877 19120
rect 17911 19117 17923 19151
rect 18782 19148 18788 19160
rect 18743 19120 18788 19148
rect 17865 19111 17923 19117
rect 18782 19108 18788 19120
rect 18840 19108 18846 19160
rect 19352 19157 19380 19324
rect 20254 19216 20260 19228
rect 20215 19188 20260 19216
rect 20254 19176 20260 19188
rect 20312 19176 20318 19228
rect 19337 19151 19395 19157
rect 19337 19117 19349 19151
rect 19383 19117 19395 19151
rect 20070 19148 20076 19160
rect 20031 19120 20076 19148
rect 19337 19111 19395 19117
rect 20070 19108 20076 19120
rect 20128 19108 20134 19160
rect 9766 19080 9772 19092
rect 8312 19052 9772 19080
rect 9766 19040 9772 19052
rect 9824 19040 9830 19092
rect 11793 19083 11851 19089
rect 11793 19080 11805 19083
rect 9876 19052 11805 19080
rect 5442 19012 5448 19024
rect 5403 18984 5448 19012
rect 5442 18972 5448 18984
rect 5500 18972 5506 19024
rect 8386 19012 8392 19024
rect 8347 18984 8392 19012
rect 8386 18972 8392 18984
rect 8444 18972 8450 19024
rect 9876 19021 9904 19052
rect 11793 19049 11805 19052
rect 11839 19049 11851 19083
rect 11793 19043 11851 19049
rect 13348 19083 13406 19089
rect 13348 19049 13360 19083
rect 13394 19080 13406 19083
rect 13814 19080 13820 19092
rect 13394 19052 13820 19080
rect 13394 19049 13406 19052
rect 13348 19043 13406 19049
rect 13814 19040 13820 19052
rect 13872 19040 13878 19092
rect 15378 19080 15384 19092
rect 13924 19052 15384 19080
rect 9861 19015 9919 19021
rect 9861 18981 9873 19015
rect 9907 18981 9919 19015
rect 9861 18975 9919 18981
rect 9950 18972 9956 19024
rect 10008 19012 10014 19024
rect 10229 19015 10287 19021
rect 10229 19012 10241 19015
rect 10008 18984 10241 19012
rect 10008 18972 10014 18984
rect 10229 18981 10241 18984
rect 10275 19012 10287 19015
rect 11238 19012 11244 19024
rect 10275 18984 11244 19012
rect 10275 18981 10287 18984
rect 10229 18975 10287 18981
rect 11238 18972 11244 18984
rect 11296 18972 11302 19024
rect 11333 19015 11391 19021
rect 11333 18981 11345 19015
rect 11379 19012 11391 19015
rect 11514 19012 11520 19024
rect 11379 18984 11520 19012
rect 11379 18981 11391 18984
rect 11333 18975 11391 18981
rect 11514 18972 11520 18984
rect 11572 18972 11578 19024
rect 11701 19015 11759 19021
rect 11701 18981 11713 19015
rect 11747 19012 11759 19015
rect 12158 19012 12164 19024
rect 11747 18984 12164 19012
rect 11747 18981 11759 18984
rect 11701 18975 11759 18981
rect 12158 18972 12164 18984
rect 12216 18972 12222 19024
rect 12434 18972 12440 19024
rect 12492 19012 12498 19024
rect 13924 19012 13952 19052
rect 15378 19040 15384 19052
rect 15436 19040 15442 19092
rect 17313 19083 17371 19089
rect 17313 19080 17325 19083
rect 15856 19052 17325 19080
rect 14458 19012 14464 19024
rect 12492 18984 13952 19012
rect 14419 18984 14464 19012
rect 12492 18972 12498 18984
rect 14458 18972 14464 18984
rect 14516 18972 14522 19024
rect 15856 19021 15884 19052
rect 17313 19049 17325 19052
rect 17359 19049 17371 19083
rect 17313 19043 17371 19049
rect 19613 19083 19671 19089
rect 19613 19049 19625 19083
rect 19659 19080 19671 19083
rect 20438 19080 20444 19092
rect 19659 19052 20444 19080
rect 19659 19049 19671 19052
rect 19613 19043 19671 19049
rect 20438 19040 20444 19052
rect 20496 19040 20502 19092
rect 15841 19015 15899 19021
rect 15841 18981 15853 19015
rect 15887 18981 15899 19015
rect 15841 18975 15899 18981
rect 16209 19015 16267 19021
rect 16209 18981 16221 19015
rect 16255 19012 16267 19015
rect 16298 19012 16304 19024
rect 16255 18984 16304 19012
rect 16255 18981 16267 18984
rect 16209 18975 16267 18981
rect 16298 18972 16304 18984
rect 16356 18972 16362 19024
rect 18966 19012 18972 19024
rect 18927 18984 18972 19012
rect 18966 18972 18972 18984
rect 19024 18972 19030 19024
rect 1104 18922 21620 18944
rect 1104 18870 7846 18922
rect 7898 18870 7910 18922
rect 7962 18870 7974 18922
rect 8026 18870 8038 18922
rect 8090 18870 14710 18922
rect 14762 18870 14774 18922
rect 14826 18870 14838 18922
rect 14890 18870 14902 18922
rect 14954 18870 21620 18922
rect 1104 18848 21620 18870
rect 3789 18811 3847 18817
rect 3789 18777 3801 18811
rect 3835 18808 3847 18811
rect 4706 18808 4712 18820
rect 3835 18780 4712 18808
rect 3835 18777 3847 18780
rect 3789 18771 3847 18777
rect 4706 18768 4712 18780
rect 4764 18768 4770 18820
rect 5166 18808 5172 18820
rect 5127 18780 5172 18808
rect 5166 18768 5172 18780
rect 5224 18768 5230 18820
rect 6362 18768 6368 18820
rect 6420 18808 6426 18820
rect 8202 18808 8208 18820
rect 6420 18780 8064 18808
rect 8163 18780 8208 18808
rect 6420 18768 6426 18780
rect 290 18700 296 18752
rect 348 18740 354 18752
rect 6730 18740 6736 18752
rect 348 18712 6736 18740
rect 348 18700 354 18712
rect 6730 18700 6736 18712
rect 6788 18700 6794 18752
rect 7006 18740 7012 18752
rect 6840 18712 7012 18740
rect 2676 18675 2734 18681
rect 2676 18641 2688 18675
rect 2722 18672 2734 18675
rect 2958 18672 2964 18684
rect 2722 18644 2964 18672
rect 2722 18641 2734 18644
rect 2676 18635 2734 18641
rect 2958 18632 2964 18644
rect 3016 18632 3022 18684
rect 6840 18681 6868 18712
rect 7006 18700 7012 18712
rect 7064 18740 7070 18752
rect 8036 18740 8064 18780
rect 8202 18768 8208 18780
rect 8260 18768 8266 18820
rect 11698 18808 11704 18820
rect 8312 18780 11704 18808
rect 8312 18740 8340 18780
rect 11698 18768 11704 18780
rect 11756 18768 11762 18820
rect 11793 18811 11851 18817
rect 11793 18777 11805 18811
rect 11839 18808 11851 18811
rect 11882 18808 11888 18820
rect 11839 18780 11888 18808
rect 11839 18777 11851 18780
rect 11793 18771 11851 18777
rect 11882 18768 11888 18780
rect 11940 18768 11946 18820
rect 12253 18811 12311 18817
rect 12253 18777 12265 18811
rect 12299 18808 12311 18811
rect 12434 18808 12440 18820
rect 12299 18780 12440 18808
rect 12299 18777 12311 18780
rect 12253 18771 12311 18777
rect 12434 18768 12440 18780
rect 12492 18768 12498 18820
rect 12526 18768 12532 18820
rect 12584 18808 12590 18820
rect 12986 18808 12992 18820
rect 12584 18780 12992 18808
rect 12584 18768 12590 18780
rect 12986 18768 12992 18780
rect 13044 18768 13050 18820
rect 13814 18808 13820 18820
rect 13775 18780 13820 18808
rect 13814 18768 13820 18780
rect 13872 18768 13878 18820
rect 14090 18768 14096 18820
rect 14148 18808 14154 18820
rect 14550 18808 14556 18820
rect 14148 18780 14556 18808
rect 14148 18768 14154 18780
rect 14550 18768 14556 18780
rect 14608 18768 14614 18820
rect 15933 18811 15991 18817
rect 15933 18777 15945 18811
rect 15979 18777 15991 18811
rect 15933 18771 15991 18777
rect 7064 18712 7512 18740
rect 8036 18712 8340 18740
rect 7064 18700 7070 18712
rect 5077 18675 5135 18681
rect 5077 18641 5089 18675
rect 5123 18672 5135 18675
rect 5721 18675 5779 18681
rect 5721 18672 5733 18675
rect 5123 18644 5733 18672
rect 5123 18641 5135 18644
rect 5077 18635 5135 18641
rect 5721 18641 5733 18644
rect 5767 18641 5779 18675
rect 6825 18675 6883 18681
rect 6825 18672 6837 18675
rect 5721 18635 5779 18641
rect 5828 18644 6837 18672
rect 1578 18564 1584 18616
rect 1636 18604 1642 18616
rect 2406 18604 2412 18616
rect 1636 18576 2412 18604
rect 1636 18564 1642 18576
rect 2406 18564 2412 18576
rect 2464 18564 2470 18616
rect 5353 18607 5411 18613
rect 5353 18573 5365 18607
rect 5399 18604 5411 18607
rect 5442 18604 5448 18616
rect 5399 18576 5448 18604
rect 5399 18573 5411 18576
rect 5353 18567 5411 18573
rect 5442 18564 5448 18576
rect 5500 18564 5506 18616
rect 5828 18604 5856 18644
rect 6825 18641 6837 18644
rect 6871 18641 6883 18675
rect 6825 18635 6883 18641
rect 7092 18675 7150 18681
rect 7092 18641 7104 18675
rect 7138 18672 7150 18675
rect 7374 18672 7380 18684
rect 7138 18644 7380 18672
rect 7138 18641 7150 18644
rect 7092 18635 7150 18641
rect 7374 18632 7380 18644
rect 7432 18632 7438 18684
rect 7484 18672 7512 18712
rect 8386 18700 8392 18752
rect 8444 18740 8450 18752
rect 9002 18743 9060 18749
rect 9002 18740 9014 18743
rect 8444 18712 9014 18740
rect 8444 18700 8450 18712
rect 9002 18709 9014 18712
rect 9048 18709 9060 18743
rect 9002 18703 9060 18709
rect 10321 18743 10379 18749
rect 10321 18709 10333 18743
rect 10367 18740 10379 18743
rect 10410 18740 10416 18752
rect 10367 18712 10416 18740
rect 10367 18709 10379 18712
rect 10321 18703 10379 18709
rect 10410 18700 10416 18712
rect 10468 18740 10474 18752
rect 10658 18743 10716 18749
rect 10658 18740 10670 18743
rect 10468 18712 10670 18740
rect 10468 18700 10474 18712
rect 10658 18709 10670 18712
rect 10704 18709 10716 18743
rect 11900 18740 11928 18768
rect 12682 18743 12740 18749
rect 12682 18740 12694 18743
rect 11900 18712 12694 18740
rect 10658 18703 10716 18709
rect 12682 18709 12694 18712
rect 12728 18709 12740 18743
rect 12682 18703 12740 18709
rect 14458 18700 14464 18752
rect 14516 18740 14522 18752
rect 14798 18743 14856 18749
rect 14798 18740 14810 18743
rect 14516 18712 14810 18740
rect 14516 18700 14522 18712
rect 14798 18709 14810 18712
rect 14844 18709 14856 18743
rect 15948 18740 15976 18771
rect 17954 18768 17960 18820
rect 18012 18808 18018 18820
rect 19426 18808 19432 18820
rect 18012 18780 19432 18808
rect 18012 18768 18018 18780
rect 19426 18768 19432 18780
rect 19484 18768 19490 18820
rect 20714 18808 20720 18820
rect 20675 18780 20720 18808
rect 20714 18768 20720 18780
rect 20772 18768 20778 18820
rect 16482 18749 16488 18752
rect 16476 18740 16488 18749
rect 15948 18712 16488 18740
rect 14798 18703 14856 18709
rect 16476 18703 16488 18712
rect 16482 18700 16488 18703
rect 16540 18700 16546 18752
rect 18782 18700 18788 18752
rect 18840 18740 18846 18752
rect 19613 18743 19671 18749
rect 19613 18740 19625 18743
rect 18840 18712 19625 18740
rect 18840 18700 18846 18712
rect 19613 18709 19625 18712
rect 19659 18709 19671 18743
rect 19613 18703 19671 18709
rect 8757 18675 8815 18681
rect 8757 18672 8769 18675
rect 7484 18644 8769 18672
rect 8757 18641 8769 18644
rect 8803 18672 8815 18675
rect 8803 18644 9812 18672
rect 8803 18641 8815 18644
rect 8757 18635 8815 18641
rect 9784 18604 9812 18644
rect 10226 18632 10232 18684
rect 10284 18672 10290 18684
rect 14366 18672 14372 18684
rect 10284 18644 14372 18672
rect 10284 18632 10290 18644
rect 14366 18632 14372 18644
rect 14424 18632 14430 18684
rect 14553 18675 14611 18681
rect 14553 18641 14565 18675
rect 14599 18672 14611 18675
rect 15930 18672 15936 18684
rect 14599 18644 15936 18672
rect 14599 18641 14611 18644
rect 14553 18635 14611 18641
rect 15930 18632 15936 18644
rect 15988 18672 15994 18684
rect 16209 18675 16267 18681
rect 16209 18672 16221 18675
rect 15988 18644 16221 18672
rect 15988 18632 15994 18644
rect 16209 18641 16221 18644
rect 16255 18641 16267 18675
rect 16209 18635 16267 18641
rect 17954 18632 17960 18684
rect 18012 18672 18018 18684
rect 18233 18675 18291 18681
rect 18233 18672 18245 18675
rect 18012 18644 18245 18672
rect 18012 18632 18018 18644
rect 18233 18641 18245 18644
rect 18279 18641 18291 18675
rect 18233 18635 18291 18641
rect 18509 18675 18567 18681
rect 18509 18641 18521 18675
rect 18555 18672 18567 18675
rect 19150 18672 19156 18684
rect 18555 18644 19156 18672
rect 18555 18641 18567 18644
rect 18509 18635 18567 18641
rect 19150 18632 19156 18644
rect 19208 18632 19214 18684
rect 19334 18672 19340 18684
rect 19295 18644 19340 18672
rect 19334 18632 19340 18644
rect 19392 18632 19398 18684
rect 19518 18632 19524 18684
rect 19576 18672 19582 18684
rect 20533 18675 20591 18681
rect 20533 18672 20545 18675
rect 19576 18644 20545 18672
rect 19576 18632 19582 18644
rect 20533 18641 20545 18644
rect 20579 18641 20591 18675
rect 20533 18635 20591 18641
rect 9858 18604 9864 18616
rect 5552 18576 5856 18604
rect 9771 18576 9864 18604
rect 5074 18496 5080 18548
rect 5132 18536 5138 18548
rect 5552 18536 5580 18576
rect 9858 18564 9864 18576
rect 9916 18604 9922 18616
rect 10413 18607 10471 18613
rect 10413 18604 10425 18607
rect 9916 18576 10425 18604
rect 9916 18564 9922 18576
rect 10413 18573 10425 18576
rect 10459 18573 10471 18607
rect 10413 18567 10471 18573
rect 11422 18564 11428 18616
rect 11480 18604 11486 18616
rect 11882 18604 11888 18616
rect 11480 18576 11888 18604
rect 11480 18564 11486 18576
rect 11882 18564 11888 18576
rect 11940 18564 11946 18616
rect 12437 18607 12495 18613
rect 12437 18573 12449 18607
rect 12483 18573 12495 18607
rect 14090 18604 14096 18616
rect 14051 18576 14096 18604
rect 12437 18567 12495 18573
rect 5132 18508 5580 18536
rect 10137 18539 10195 18545
rect 5132 18496 5138 18508
rect 10137 18505 10149 18539
rect 10183 18536 10195 18539
rect 10321 18539 10379 18545
rect 10321 18536 10333 18539
rect 10183 18508 10333 18536
rect 10183 18505 10195 18508
rect 10137 18499 10195 18505
rect 10321 18505 10333 18508
rect 10367 18505 10379 18539
rect 10321 18499 10379 18505
rect 4709 18471 4767 18477
rect 4709 18437 4721 18471
rect 4755 18468 4767 18471
rect 5166 18468 5172 18480
rect 4755 18440 5172 18468
rect 4755 18437 4767 18440
rect 4709 18431 4767 18437
rect 5166 18428 5172 18440
rect 5224 18428 5230 18480
rect 7006 18428 7012 18480
rect 7064 18468 7070 18480
rect 12253 18471 12311 18477
rect 12253 18468 12265 18471
rect 7064 18440 12265 18468
rect 7064 18428 7070 18440
rect 12253 18437 12265 18440
rect 12299 18437 12311 18471
rect 12452 18468 12480 18567
rect 14090 18564 14096 18576
rect 14148 18564 14154 18616
rect 17678 18564 17684 18616
rect 17736 18604 17742 18616
rect 21174 18604 21180 18616
rect 17736 18576 21180 18604
rect 17736 18564 17742 18576
rect 21174 18564 21180 18576
rect 21232 18564 21238 18616
rect 20070 18536 20076 18548
rect 17144 18508 20076 18536
rect 12618 18468 12624 18480
rect 12452 18440 12624 18468
rect 12253 18431 12311 18437
rect 12618 18428 12624 18440
rect 12676 18428 12682 18480
rect 12710 18428 12716 18480
rect 12768 18468 12774 18480
rect 17144 18468 17172 18508
rect 20070 18496 20076 18508
rect 20128 18496 20134 18548
rect 17586 18468 17592 18480
rect 12768 18440 17172 18468
rect 17547 18440 17592 18468
rect 12768 18428 12774 18440
rect 17586 18428 17592 18440
rect 17644 18428 17650 18480
rect 19058 18428 19064 18480
rect 19116 18468 19122 18480
rect 20622 18468 20628 18480
rect 19116 18440 20628 18468
rect 19116 18428 19122 18440
rect 20622 18428 20628 18440
rect 20680 18428 20686 18480
rect 1104 18378 21620 18400
rect 1104 18326 4414 18378
rect 4466 18326 4478 18378
rect 4530 18326 4542 18378
rect 4594 18326 4606 18378
rect 4658 18326 11278 18378
rect 11330 18326 11342 18378
rect 11394 18326 11406 18378
rect 11458 18326 11470 18378
rect 11522 18326 18142 18378
rect 18194 18326 18206 18378
rect 18258 18326 18270 18378
rect 18322 18326 18334 18378
rect 18386 18326 21620 18378
rect 1104 18304 21620 18326
rect 1946 18224 1952 18276
rect 2004 18264 2010 18276
rect 2004 18236 3004 18264
rect 2004 18224 2010 18236
rect 2976 18196 3004 18236
rect 3050 18224 3056 18276
rect 3108 18264 3114 18276
rect 5350 18264 5356 18276
rect 3108 18236 5356 18264
rect 3108 18224 3114 18236
rect 5350 18224 5356 18236
rect 5408 18224 5414 18276
rect 7929 18267 7987 18273
rect 7929 18233 7941 18267
rect 7975 18264 7987 18267
rect 8294 18264 8300 18276
rect 7975 18236 8300 18264
rect 7975 18233 7987 18236
rect 7929 18227 7987 18233
rect 8294 18224 8300 18236
rect 8352 18224 8358 18276
rect 9766 18224 9772 18276
rect 9824 18264 9830 18276
rect 10686 18264 10692 18276
rect 9824 18236 10692 18264
rect 9824 18224 9830 18236
rect 10686 18224 10692 18236
rect 10744 18224 10750 18276
rect 11606 18224 11612 18276
rect 11664 18264 11670 18276
rect 12710 18264 12716 18276
rect 11664 18236 12716 18264
rect 11664 18224 11670 18236
rect 12710 18224 12716 18236
rect 12768 18224 12774 18276
rect 14185 18267 14243 18273
rect 12820 18236 13400 18264
rect 5718 18196 5724 18208
rect 2976 18168 5724 18196
rect 5718 18156 5724 18168
rect 5776 18156 5782 18208
rect 5810 18156 5816 18208
rect 5868 18196 5874 18208
rect 11514 18196 11520 18208
rect 5868 18168 11520 18196
rect 5868 18156 5874 18168
rect 11514 18156 11520 18168
rect 11572 18156 11578 18208
rect 12066 18196 12072 18208
rect 11624 18168 12072 18196
rect 8202 18088 8208 18140
rect 8260 18128 8266 18140
rect 8481 18131 8539 18137
rect 8481 18128 8493 18131
rect 8260 18100 8493 18128
rect 8260 18088 8266 18100
rect 8481 18097 8493 18100
rect 8527 18097 8539 18131
rect 8481 18091 8539 18097
rect 9766 18088 9772 18140
rect 9824 18128 9830 18140
rect 11624 18128 11652 18168
rect 12066 18156 12072 18168
rect 12124 18156 12130 18208
rect 9824 18100 11652 18128
rect 11701 18131 11759 18137
rect 9824 18088 9830 18100
rect 11701 18097 11713 18131
rect 11747 18128 11759 18131
rect 12158 18128 12164 18140
rect 11747 18100 12164 18128
rect 11747 18097 11759 18100
rect 11701 18091 11759 18097
rect 12158 18088 12164 18100
rect 12216 18088 12222 18140
rect 3602 18020 3608 18072
rect 3660 18060 3666 18072
rect 4246 18060 4252 18072
rect 3660 18032 4252 18060
rect 3660 18020 3666 18032
rect 4246 18020 4252 18032
rect 4304 18020 4310 18072
rect 5166 18060 5172 18072
rect 5127 18032 5172 18060
rect 5166 18020 5172 18032
rect 5224 18020 5230 18072
rect 8389 18063 8447 18069
rect 8389 18029 8401 18063
rect 8435 18060 8447 18063
rect 8570 18060 8576 18072
rect 8435 18032 8576 18060
rect 8435 18029 8447 18032
rect 8389 18023 8447 18029
rect 8570 18020 8576 18032
rect 8628 18020 8634 18072
rect 9674 18020 9680 18072
rect 9732 18060 9738 18072
rect 12820 18060 12848 18236
rect 12897 18199 12955 18205
rect 12897 18165 12909 18199
rect 12943 18165 12955 18199
rect 12897 18159 12955 18165
rect 9732 18032 12848 18060
rect 12912 18060 12940 18159
rect 13372 18137 13400 18236
rect 14185 18233 14197 18267
rect 14231 18264 14243 18267
rect 19334 18264 19340 18276
rect 14231 18236 19340 18264
rect 14231 18233 14243 18236
rect 14185 18227 14243 18233
rect 19334 18224 19340 18236
rect 19392 18224 19398 18276
rect 13630 18156 13636 18208
rect 13688 18196 13694 18208
rect 14274 18196 14280 18208
rect 13688 18168 14280 18196
rect 13688 18156 13694 18168
rect 14274 18156 14280 18168
rect 14332 18156 14338 18208
rect 19886 18156 19892 18208
rect 19944 18196 19950 18208
rect 21358 18196 21364 18208
rect 19944 18168 21364 18196
rect 19944 18156 19950 18168
rect 21358 18156 21364 18168
rect 21416 18156 21422 18208
rect 13357 18131 13415 18137
rect 13357 18097 13369 18131
rect 13403 18097 13415 18131
rect 13357 18091 13415 18097
rect 13541 18131 13599 18137
rect 13541 18097 13553 18131
rect 13587 18128 13599 18131
rect 13814 18128 13820 18140
rect 13587 18100 13820 18128
rect 13587 18097 13599 18100
rect 13541 18091 13599 18097
rect 13814 18088 13820 18100
rect 13872 18088 13878 18140
rect 14458 18088 14464 18140
rect 14516 18128 14522 18140
rect 14737 18131 14795 18137
rect 14737 18128 14749 18131
rect 14516 18100 14749 18128
rect 14516 18088 14522 18100
rect 14737 18097 14749 18100
rect 14783 18097 14795 18131
rect 14737 18091 14795 18097
rect 19794 18088 19800 18140
rect 19852 18128 19858 18140
rect 21910 18128 21916 18140
rect 19852 18100 21916 18128
rect 19852 18088 19858 18100
rect 21910 18088 21916 18100
rect 21968 18088 21974 18140
rect 12912 18032 13860 18060
rect 9732 18020 9738 18032
rect 5258 17952 5264 18004
rect 5316 17992 5322 18004
rect 5445 17995 5503 18001
rect 5445 17992 5457 17995
rect 5316 17964 5457 17992
rect 5316 17952 5322 17964
rect 5445 17961 5457 17964
rect 5491 17961 5503 17995
rect 5445 17955 5503 17961
rect 7466 17952 7472 18004
rect 7524 17992 7530 18004
rect 8478 17992 8484 18004
rect 7524 17964 8484 17992
rect 7524 17952 7530 17964
rect 8478 17952 8484 17964
rect 8536 17952 8542 18004
rect 10778 17952 10784 18004
rect 10836 17992 10842 18004
rect 12710 17992 12716 18004
rect 10836 17964 12716 17992
rect 10836 17952 10842 17964
rect 12710 17952 12716 17964
rect 12768 17952 12774 18004
rect 13265 17995 13323 18001
rect 13265 17992 13277 17995
rect 12820 17964 13277 17992
rect 8297 17927 8355 17933
rect 8297 17893 8309 17927
rect 8343 17924 8355 17927
rect 8754 17924 8760 17936
rect 8343 17896 8760 17924
rect 8343 17893 8355 17896
rect 8297 17887 8355 17893
rect 8754 17884 8760 17896
rect 8812 17884 8818 17936
rect 11146 17884 11152 17936
rect 11204 17924 11210 17936
rect 11974 17924 11980 17936
rect 11204 17896 11980 17924
rect 11204 17884 11210 17896
rect 11974 17884 11980 17896
rect 12032 17884 12038 17936
rect 12066 17884 12072 17936
rect 12124 17924 12130 17936
rect 12820 17924 12848 17964
rect 13265 17961 13277 17964
rect 13311 17961 13323 17995
rect 13265 17955 13323 17961
rect 13354 17952 13360 18004
rect 13412 17992 13418 18004
rect 13832 17992 13860 18032
rect 14090 18020 14096 18072
rect 14148 18060 14154 18072
rect 14553 18063 14611 18069
rect 14553 18060 14565 18063
rect 14148 18032 14565 18060
rect 14148 18020 14154 18032
rect 14553 18029 14565 18032
rect 14599 18029 14611 18063
rect 20254 18060 20260 18072
rect 20215 18032 20260 18060
rect 14553 18023 14611 18029
rect 20254 18020 20260 18032
rect 20312 18020 20318 18072
rect 14645 17995 14703 18001
rect 14645 17992 14657 17995
rect 13412 17964 13768 17992
rect 13832 17964 14657 17992
rect 13412 17952 13418 17964
rect 12124 17896 12848 17924
rect 12124 17884 12130 17896
rect 13078 17884 13084 17936
rect 13136 17924 13142 17936
rect 13630 17924 13636 17936
rect 13136 17896 13636 17924
rect 13136 17884 13142 17896
rect 13630 17884 13636 17896
rect 13688 17884 13694 17936
rect 13740 17924 13768 17964
rect 14645 17961 14657 17964
rect 14691 17961 14703 17995
rect 14645 17955 14703 17961
rect 15838 17952 15844 18004
rect 15896 17992 15902 18004
rect 19334 17992 19340 18004
rect 15896 17964 19340 17992
rect 15896 17952 15902 17964
rect 19334 17952 19340 17964
rect 19392 17952 19398 18004
rect 19702 17952 19708 18004
rect 19760 17992 19766 18004
rect 20346 17992 20352 18004
rect 19760 17964 20352 17992
rect 19760 17952 19766 17964
rect 20346 17952 20352 17964
rect 20404 17952 20410 18004
rect 15194 17924 15200 17936
rect 13740 17896 15200 17924
rect 15194 17884 15200 17896
rect 15252 17884 15258 17936
rect 15286 17884 15292 17936
rect 15344 17924 15350 17936
rect 16482 17924 16488 17936
rect 15344 17896 16488 17924
rect 15344 17884 15350 17896
rect 16482 17884 16488 17896
rect 16540 17884 16546 17936
rect 16942 17884 16948 17936
rect 17000 17924 17006 17936
rect 20070 17924 20076 17936
rect 17000 17896 20076 17924
rect 17000 17884 17006 17896
rect 20070 17884 20076 17896
rect 20128 17884 20134 17936
rect 20438 17924 20444 17936
rect 20399 17896 20444 17924
rect 20438 17884 20444 17896
rect 20496 17884 20502 17936
rect 20990 17884 20996 17936
rect 21048 17924 21054 17936
rect 22462 17924 22468 17936
rect 21048 17896 22468 17924
rect 21048 17884 21054 17896
rect 22462 17884 22468 17896
rect 22520 17884 22526 17936
rect 1104 17834 21620 17856
rect 1104 17782 7846 17834
rect 7898 17782 7910 17834
rect 7962 17782 7974 17834
rect 8026 17782 8038 17834
rect 8090 17782 14710 17834
rect 14762 17782 14774 17834
rect 14826 17782 14838 17834
rect 14890 17782 14902 17834
rect 14954 17782 21620 17834
rect 1104 17760 21620 17782
rect 2958 17720 2964 17732
rect 2919 17692 2964 17720
rect 2958 17680 2964 17692
rect 3016 17680 3022 17732
rect 5258 17680 5264 17732
rect 5316 17680 5322 17732
rect 12158 17680 12164 17732
rect 12216 17720 12222 17732
rect 19334 17720 19340 17732
rect 12216 17692 19340 17720
rect 12216 17680 12222 17692
rect 19334 17680 19340 17692
rect 19392 17680 19398 17732
rect 19610 17720 19616 17732
rect 19571 17692 19616 17720
rect 19610 17680 19616 17692
rect 19668 17680 19674 17732
rect 19702 17680 19708 17732
rect 19760 17720 19766 17732
rect 20070 17720 20076 17732
rect 19760 17692 20076 17720
rect 19760 17680 19766 17692
rect 20070 17680 20076 17692
rect 20128 17680 20134 17732
rect 20438 17680 20444 17732
rect 20496 17720 20502 17732
rect 20806 17720 20812 17732
rect 20496 17692 20812 17720
rect 20496 17680 20502 17692
rect 20806 17680 20812 17692
rect 20864 17680 20870 17732
rect 1578 17584 1584 17596
rect 1539 17556 1584 17584
rect 1578 17544 1584 17556
rect 1636 17544 1642 17596
rect 1848 17587 1906 17593
rect 1848 17553 1860 17587
rect 1894 17584 1906 17587
rect 3142 17584 3148 17596
rect 1894 17556 3148 17584
rect 1894 17553 1906 17556
rect 1848 17547 1906 17553
rect 3142 17544 3148 17556
rect 3200 17544 3206 17596
rect 5276 17584 5304 17680
rect 5344 17655 5402 17661
rect 5344 17621 5356 17655
rect 5390 17652 5402 17655
rect 5442 17652 5448 17664
rect 5390 17624 5448 17652
rect 5390 17621 5402 17624
rect 5344 17615 5402 17621
rect 5442 17612 5448 17624
rect 5500 17612 5506 17664
rect 5626 17612 5632 17664
rect 5684 17652 5690 17664
rect 16114 17652 16120 17664
rect 5684 17624 16120 17652
rect 5684 17612 5690 17624
rect 16114 17612 16120 17624
rect 16172 17612 16178 17664
rect 16224 17624 20024 17652
rect 16224 17584 16252 17624
rect 5276 17556 16252 17584
rect 16298 17544 16304 17596
rect 16356 17584 16362 17596
rect 17218 17584 17224 17596
rect 16356 17556 17224 17584
rect 16356 17544 16362 17556
rect 17218 17544 17224 17556
rect 17276 17544 17282 17596
rect 19996 17593 20024 17624
rect 19429 17587 19487 17593
rect 19429 17553 19441 17587
rect 19475 17584 19487 17587
rect 19981 17587 20039 17593
rect 19475 17556 19932 17584
rect 19475 17553 19487 17556
rect 19429 17547 19487 17553
rect 3326 17516 3332 17528
rect 3287 17488 3332 17516
rect 3326 17476 3332 17488
rect 3384 17476 3390 17528
rect 5074 17516 5080 17528
rect 5035 17488 5080 17516
rect 5074 17476 5080 17488
rect 5132 17476 5138 17528
rect 7466 17476 7472 17528
rect 7524 17516 7530 17528
rect 19518 17516 19524 17528
rect 7524 17488 19524 17516
rect 7524 17476 7530 17488
rect 19518 17476 19524 17488
rect 19576 17476 19582 17528
rect 19904 17516 19932 17556
rect 19981 17553 19993 17587
rect 20027 17553 20039 17587
rect 19981 17547 20039 17553
rect 20070 17544 20076 17596
rect 20128 17584 20134 17596
rect 20533 17587 20591 17593
rect 20533 17584 20545 17587
rect 20128 17556 20545 17584
rect 20128 17544 20134 17556
rect 20533 17553 20545 17556
rect 20579 17553 20591 17587
rect 20533 17547 20591 17553
rect 20806 17516 20812 17528
rect 19904 17488 20812 17516
rect 20806 17476 20812 17488
rect 20864 17476 20870 17528
rect 9674 17408 9680 17460
rect 9732 17448 9738 17460
rect 17402 17448 17408 17460
rect 9732 17420 17408 17448
rect 9732 17408 9738 17420
rect 17402 17408 17408 17420
rect 17460 17408 17466 17460
rect 6457 17383 6515 17389
rect 6457 17349 6469 17383
rect 6503 17380 6515 17383
rect 8662 17380 8668 17392
rect 6503 17352 8668 17380
rect 6503 17349 6515 17352
rect 6457 17343 6515 17349
rect 8662 17340 8668 17352
rect 8720 17340 8726 17392
rect 11698 17340 11704 17392
rect 11756 17380 11762 17392
rect 12342 17380 12348 17392
rect 11756 17352 12348 17380
rect 11756 17340 11762 17352
rect 12342 17340 12348 17352
rect 12400 17340 12406 17392
rect 16114 17340 16120 17392
rect 16172 17380 16178 17392
rect 18506 17380 18512 17392
rect 16172 17352 18512 17380
rect 16172 17340 16178 17352
rect 18506 17340 18512 17352
rect 18564 17340 18570 17392
rect 20162 17380 20168 17392
rect 20123 17352 20168 17380
rect 20162 17340 20168 17352
rect 20220 17340 20226 17392
rect 20714 17380 20720 17392
rect 20675 17352 20720 17380
rect 20714 17340 20720 17352
rect 20772 17340 20778 17392
rect 1104 17290 21620 17312
rect 1104 17238 4414 17290
rect 4466 17238 4478 17290
rect 4530 17238 4542 17290
rect 4594 17238 4606 17290
rect 4658 17238 11278 17290
rect 11330 17238 11342 17290
rect 11394 17238 11406 17290
rect 11458 17238 11470 17290
rect 11522 17238 18142 17290
rect 18194 17238 18206 17290
rect 18258 17238 18270 17290
rect 18322 17238 18334 17290
rect 18386 17238 21620 17290
rect 1104 17216 21620 17238
rect 9674 17176 9680 17188
rect 9635 17148 9680 17176
rect 9674 17136 9680 17148
rect 9732 17136 9738 17188
rect 11977 17179 12035 17185
rect 11977 17145 11989 17179
rect 12023 17176 12035 17179
rect 17218 17176 17224 17188
rect 12023 17148 17224 17176
rect 12023 17145 12035 17148
rect 11977 17139 12035 17145
rect 17218 17136 17224 17148
rect 17276 17136 17282 17188
rect 17681 17179 17739 17185
rect 17681 17145 17693 17179
rect 17727 17176 17739 17179
rect 17954 17176 17960 17188
rect 17727 17148 17960 17176
rect 17727 17145 17739 17148
rect 17681 17139 17739 17145
rect 17954 17136 17960 17148
rect 18012 17136 18018 17188
rect 3142 17068 3148 17120
rect 3200 17108 3206 17120
rect 8754 17108 8760 17120
rect 3200 17080 4660 17108
rect 3200 17068 3206 17080
rect 2958 17000 2964 17052
rect 3016 17040 3022 17052
rect 3513 17043 3571 17049
rect 3513 17040 3525 17043
rect 3016 17012 3525 17040
rect 3016 17000 3022 17012
rect 3513 17009 3525 17012
rect 3559 17009 3571 17043
rect 3513 17003 3571 17009
rect 4154 17000 4160 17052
rect 4212 17040 4218 17052
rect 4632 17049 4660 17080
rect 5460 17080 8760 17108
rect 4525 17043 4583 17049
rect 4525 17040 4537 17043
rect 4212 17012 4537 17040
rect 4212 17000 4218 17012
rect 4525 17009 4537 17012
rect 4571 17009 4583 17043
rect 4525 17003 4583 17009
rect 4617 17043 4675 17049
rect 4617 17009 4629 17043
rect 4663 17009 4675 17043
rect 4617 17003 4675 17009
rect 3326 16972 3332 16984
rect 3287 16944 3332 16972
rect 3326 16932 3332 16944
rect 3384 16932 3390 16984
rect 4433 16975 4491 16981
rect 4433 16941 4445 16975
rect 4479 16972 4491 16975
rect 5460 16972 5488 17080
rect 8754 17068 8760 17080
rect 8812 17068 8818 17120
rect 12158 17108 12164 17120
rect 12119 17080 12164 17108
rect 12158 17068 12164 17080
rect 12216 17068 12222 17120
rect 12342 17068 12348 17120
rect 12400 17108 12406 17120
rect 12400 17080 13584 17108
rect 12400 17068 12406 17080
rect 5534 17000 5540 17052
rect 5592 17040 5598 17052
rect 7466 17040 7472 17052
rect 5592 17012 7328 17040
rect 7427 17012 7472 17040
rect 5592 17000 5598 17012
rect 4479 16944 5488 16972
rect 4479 16941 4491 16944
rect 4433 16935 4491 16941
rect 6822 16932 6828 16984
rect 6880 16972 6886 16984
rect 7193 16975 7251 16981
rect 7193 16972 7205 16975
rect 6880 16944 7205 16972
rect 6880 16932 6886 16944
rect 7193 16941 7205 16944
rect 7239 16941 7251 16975
rect 7300 16972 7328 17012
rect 7466 17000 7472 17012
rect 7524 17000 7530 17052
rect 8662 17040 8668 17052
rect 8623 17012 8668 17040
rect 8662 17000 8668 17012
rect 8720 17000 8726 17052
rect 10226 17040 10232 17052
rect 10187 17012 10232 17040
rect 10226 17000 10232 17012
rect 10284 17000 10290 17052
rect 11698 17040 11704 17052
rect 11659 17012 11704 17040
rect 11698 17000 11704 17012
rect 11756 17000 11762 17052
rect 12710 17040 12716 17052
rect 12671 17012 12716 17040
rect 12710 17000 12716 17012
rect 12768 17000 12774 17052
rect 8573 16975 8631 16981
rect 8573 16972 8585 16975
rect 7300 16944 8585 16972
rect 7193 16935 7251 16941
rect 8573 16941 8585 16944
rect 8619 16941 8631 16975
rect 11606 16972 11612 16984
rect 11567 16944 11612 16972
rect 8573 16935 8631 16941
rect 11606 16932 11612 16944
rect 11664 16932 11670 16984
rect 13556 16972 13584 17080
rect 14090 17000 14096 17052
rect 14148 17040 14154 17052
rect 14553 17043 14611 17049
rect 14553 17040 14565 17043
rect 14148 17012 14565 17040
rect 14148 17000 14154 17012
rect 14553 17009 14565 17012
rect 14599 17009 14611 17043
rect 15930 17040 15936 17052
rect 15891 17012 15936 17040
rect 14553 17003 14611 17009
rect 15930 17000 15936 17012
rect 15988 17000 15994 17052
rect 17678 17000 17684 17052
rect 17736 17040 17742 17052
rect 18233 17043 18291 17049
rect 18233 17040 18245 17043
rect 17736 17012 18245 17040
rect 17736 17000 17742 17012
rect 18233 17009 18245 17012
rect 18279 17009 18291 17043
rect 18233 17003 18291 17009
rect 19613 17043 19671 17049
rect 19613 17009 19625 17043
rect 19659 17040 19671 17043
rect 20254 17040 20260 17052
rect 19659 17012 20260 17040
rect 19659 17009 19671 17012
rect 19613 17003 19671 17009
rect 20254 17000 20260 17012
rect 20312 17000 20318 17052
rect 20349 17043 20407 17049
rect 20349 17009 20361 17043
rect 20395 17040 20407 17043
rect 20806 17040 20812 17052
rect 20395 17012 20812 17040
rect 20395 17009 20407 17012
rect 20349 17003 20407 17009
rect 20806 17000 20812 17012
rect 20864 17000 20870 17052
rect 14461 16975 14519 16981
rect 14461 16972 14473 16975
rect 13556 16944 14473 16972
rect 14461 16941 14473 16944
rect 14507 16941 14519 16975
rect 14461 16935 14519 16941
rect 16200 16975 16258 16981
rect 16200 16941 16212 16975
rect 16246 16972 16258 16975
rect 17586 16972 17592 16984
rect 16246 16944 17592 16972
rect 16246 16941 16258 16944
rect 16200 16935 16258 16941
rect 17586 16932 17592 16944
rect 17644 16932 17650 16984
rect 19334 16972 19340 16984
rect 19295 16944 19340 16972
rect 19334 16932 19340 16944
rect 19392 16932 19398 16984
rect 19426 16932 19432 16984
rect 19484 16972 19490 16984
rect 20073 16975 20131 16981
rect 20073 16972 20085 16975
rect 19484 16944 20085 16972
rect 19484 16932 19490 16944
rect 20073 16941 20085 16944
rect 20119 16941 20131 16975
rect 20073 16935 20131 16941
rect 10137 16907 10195 16913
rect 10137 16904 10149 16907
rect 8128 16876 10149 16904
rect 2958 16836 2964 16848
rect 2919 16808 2964 16836
rect 2958 16796 2964 16808
rect 3016 16796 3022 16848
rect 8128 16845 8156 16876
rect 10137 16873 10149 16876
rect 10183 16873 10195 16907
rect 12621 16907 12679 16913
rect 12621 16904 12633 16907
rect 10137 16867 10195 16873
rect 11164 16876 12633 16904
rect 3421 16839 3479 16845
rect 3421 16805 3433 16839
rect 3467 16836 3479 16839
rect 4065 16839 4123 16845
rect 4065 16836 4077 16839
rect 3467 16808 4077 16836
rect 3467 16805 3479 16808
rect 3421 16799 3479 16805
rect 4065 16805 4077 16808
rect 4111 16805 4123 16839
rect 4065 16799 4123 16805
rect 8113 16839 8171 16845
rect 8113 16805 8125 16839
rect 8159 16805 8171 16839
rect 8113 16799 8171 16805
rect 8481 16839 8539 16845
rect 8481 16805 8493 16839
rect 8527 16836 8539 16839
rect 9766 16836 9772 16848
rect 8527 16808 9772 16836
rect 8527 16805 8539 16808
rect 8481 16799 8539 16805
rect 9766 16796 9772 16808
rect 9824 16796 9830 16848
rect 10042 16836 10048 16848
rect 10003 16808 10048 16836
rect 10042 16796 10048 16808
rect 10100 16796 10106 16848
rect 11164 16845 11192 16876
rect 12621 16873 12633 16876
rect 12667 16873 12679 16907
rect 12621 16867 12679 16873
rect 18049 16907 18107 16913
rect 18049 16873 18061 16907
rect 18095 16904 18107 16907
rect 18693 16907 18751 16913
rect 18693 16904 18705 16907
rect 18095 16876 18705 16904
rect 18095 16873 18107 16876
rect 18049 16867 18107 16873
rect 18693 16873 18705 16876
rect 18739 16873 18751 16907
rect 18693 16867 18751 16873
rect 11149 16839 11207 16845
rect 11149 16805 11161 16839
rect 11195 16805 11207 16839
rect 11149 16799 11207 16805
rect 11517 16839 11575 16845
rect 11517 16805 11529 16839
rect 11563 16836 11575 16839
rect 11977 16839 12035 16845
rect 11977 16836 11989 16839
rect 11563 16808 11989 16836
rect 11563 16805 11575 16808
rect 11517 16799 11575 16805
rect 11977 16805 11989 16808
rect 12023 16805 12035 16839
rect 12526 16836 12532 16848
rect 12487 16808 12532 16836
rect 11977 16799 12035 16805
rect 12526 16796 12532 16808
rect 12584 16796 12590 16848
rect 13998 16836 14004 16848
rect 13959 16808 14004 16836
rect 13998 16796 14004 16808
rect 14056 16796 14062 16848
rect 14366 16836 14372 16848
rect 14327 16808 14372 16836
rect 14366 16796 14372 16808
rect 14424 16796 14430 16848
rect 17310 16836 17316 16848
rect 17271 16808 17316 16836
rect 17310 16796 17316 16808
rect 17368 16796 17374 16848
rect 17954 16796 17960 16848
rect 18012 16836 18018 16848
rect 18141 16839 18199 16845
rect 18141 16836 18153 16839
rect 18012 16808 18153 16836
rect 18012 16796 18018 16808
rect 18141 16805 18153 16808
rect 18187 16805 18199 16839
rect 18141 16799 18199 16805
rect 1104 16746 21620 16768
rect 1104 16694 7846 16746
rect 7898 16694 7910 16746
rect 7962 16694 7974 16746
rect 8026 16694 8038 16746
rect 8090 16694 14710 16746
rect 14762 16694 14774 16746
rect 14826 16694 14838 16746
rect 14890 16694 14902 16746
rect 14954 16694 21620 16746
rect 1104 16672 21620 16694
rect 6822 16632 6828 16644
rect 6783 16604 6828 16632
rect 6822 16592 6828 16604
rect 6880 16592 6886 16644
rect 7282 16632 7288 16644
rect 7243 16604 7288 16632
rect 7282 16592 7288 16604
rect 7340 16592 7346 16644
rect 9585 16635 9643 16641
rect 9585 16601 9597 16635
rect 9631 16601 9643 16635
rect 9585 16595 9643 16601
rect 11241 16635 11299 16641
rect 11241 16601 11253 16635
rect 11287 16632 11299 16635
rect 11698 16632 11704 16644
rect 11287 16604 11704 16632
rect 11287 16601 11299 16604
rect 11241 16595 11299 16601
rect 8472 16567 8530 16573
rect 8472 16533 8484 16567
rect 8518 16564 8530 16567
rect 8662 16564 8668 16576
rect 8518 16536 8668 16564
rect 8518 16533 8530 16536
rect 8472 16527 8530 16533
rect 8662 16524 8668 16536
rect 8720 16524 8726 16576
rect 9600 16564 9628 16595
rect 11698 16592 11704 16604
rect 11756 16592 11762 16644
rect 11885 16635 11943 16641
rect 11885 16601 11897 16635
rect 11931 16632 11943 16635
rect 12526 16632 12532 16644
rect 11931 16604 12532 16632
rect 11931 16601 11943 16604
rect 11885 16595 11943 16601
rect 12526 16592 12532 16604
rect 12584 16592 12590 16644
rect 13998 16592 14004 16644
rect 14056 16632 14062 16644
rect 15013 16635 15071 16641
rect 15013 16632 15025 16635
rect 14056 16604 15025 16632
rect 14056 16592 14062 16604
rect 15013 16601 15025 16604
rect 15059 16601 15071 16635
rect 15013 16595 15071 16601
rect 18506 16592 18512 16644
rect 18564 16632 18570 16644
rect 18564 16604 19564 16632
rect 18564 16592 18570 16604
rect 10128 16567 10186 16573
rect 10128 16564 10140 16567
rect 9600 16536 10140 16564
rect 10128 16533 10140 16536
rect 10174 16564 10186 16567
rect 10226 16564 10232 16576
rect 10174 16536 10232 16564
rect 10174 16533 10186 16536
rect 10128 16527 10186 16533
rect 10226 16524 10232 16536
rect 10284 16524 10290 16576
rect 19426 16564 19432 16576
rect 14844 16536 19432 16564
rect 2958 16456 2964 16508
rect 3016 16496 3022 16508
rect 3881 16499 3939 16505
rect 3881 16496 3893 16499
rect 3016 16468 3893 16496
rect 3016 16456 3022 16468
rect 3881 16465 3893 16468
rect 3927 16465 3939 16499
rect 3881 16459 3939 16465
rect 4157 16499 4215 16505
rect 4157 16465 4169 16499
rect 4203 16496 4215 16499
rect 5626 16496 5632 16508
rect 4203 16468 5632 16496
rect 4203 16465 4215 16468
rect 4157 16459 4215 16465
rect 5626 16456 5632 16468
rect 5684 16456 5690 16508
rect 6273 16499 6331 16505
rect 6273 16465 6285 16499
rect 6319 16496 6331 16499
rect 7193 16499 7251 16505
rect 7193 16496 7205 16499
rect 6319 16468 7205 16496
rect 6319 16465 6331 16468
rect 6273 16459 6331 16465
rect 7193 16465 7205 16468
rect 7239 16465 7251 16499
rect 7193 16459 7251 16465
rect 9600 16468 12388 16496
rect 9600 16440 9628 16468
rect 7374 16428 7380 16440
rect 7335 16400 7380 16428
rect 7374 16388 7380 16400
rect 7432 16388 7438 16440
rect 8202 16428 8208 16440
rect 8163 16400 8208 16428
rect 8202 16388 8208 16400
rect 8260 16388 8266 16440
rect 9582 16388 9588 16440
rect 9640 16388 9646 16440
rect 9858 16428 9864 16440
rect 9819 16400 9864 16428
rect 9858 16388 9864 16400
rect 9916 16388 9922 16440
rect 12360 16292 12388 16468
rect 12526 16456 12532 16508
rect 12584 16496 12590 16508
rect 12710 16496 12716 16508
rect 12584 16468 12716 16496
rect 12584 16456 12590 16468
rect 12710 16456 12716 16468
rect 12768 16496 12774 16508
rect 12877 16499 12935 16505
rect 12877 16496 12889 16499
rect 12768 16468 12889 16496
rect 12768 16456 12774 16468
rect 12877 16465 12889 16468
rect 12923 16465 12935 16499
rect 14844 16496 14872 16536
rect 19426 16524 19432 16536
rect 19484 16524 19490 16576
rect 12877 16459 12935 16465
rect 14568 16468 14872 16496
rect 14921 16499 14979 16505
rect 12618 16428 12624 16440
rect 12579 16400 12624 16428
rect 12618 16388 12624 16400
rect 12676 16388 12682 16440
rect 14001 16363 14059 16369
rect 14001 16329 14013 16363
rect 14047 16360 14059 16363
rect 14090 16360 14096 16372
rect 14047 16332 14096 16360
rect 14047 16329 14059 16332
rect 14001 16323 14059 16329
rect 14090 16320 14096 16332
rect 14148 16320 14154 16372
rect 14568 16369 14596 16468
rect 14921 16465 14933 16499
rect 14967 16496 14979 16499
rect 15565 16499 15623 16505
rect 15565 16496 15577 16499
rect 14967 16468 15577 16496
rect 14967 16465 14979 16468
rect 14921 16459 14979 16465
rect 15565 16465 15577 16468
rect 15611 16465 15623 16499
rect 15565 16459 15623 16465
rect 15930 16456 15936 16508
rect 15988 16496 15994 16508
rect 16301 16499 16359 16505
rect 16301 16496 16313 16499
rect 15988 16468 16313 16496
rect 15988 16456 15994 16468
rect 16301 16465 16313 16468
rect 16347 16465 16359 16499
rect 16301 16459 16359 16465
rect 16568 16499 16626 16505
rect 16568 16465 16580 16499
rect 16614 16496 16626 16499
rect 17310 16496 17316 16508
rect 16614 16468 17316 16496
rect 16614 16465 16626 16468
rect 16568 16459 16626 16465
rect 17310 16456 17316 16468
rect 17368 16456 17374 16508
rect 17402 16456 17408 16508
rect 17460 16496 17466 16508
rect 19337 16499 19395 16505
rect 19337 16496 19349 16499
rect 17460 16468 19349 16496
rect 17460 16456 17466 16468
rect 19337 16465 19349 16468
rect 19383 16465 19395 16499
rect 19536 16496 19564 16604
rect 19702 16592 19708 16644
rect 19760 16632 19766 16644
rect 20254 16632 20260 16644
rect 19760 16604 20260 16632
rect 19760 16592 19766 16604
rect 20254 16592 20260 16604
rect 20312 16592 20318 16644
rect 20622 16592 20628 16644
rect 20680 16632 20686 16644
rect 20717 16635 20775 16641
rect 20717 16632 20729 16635
rect 20680 16604 20729 16632
rect 20680 16592 20686 16604
rect 20717 16601 20729 16604
rect 20763 16601 20775 16635
rect 20717 16595 20775 16601
rect 19613 16567 19671 16573
rect 19613 16533 19625 16567
rect 19659 16564 19671 16567
rect 20070 16564 20076 16576
rect 19659 16536 20076 16564
rect 19659 16533 19671 16536
rect 19613 16527 19671 16533
rect 20070 16524 20076 16536
rect 20128 16524 20134 16576
rect 20533 16499 20591 16505
rect 20533 16496 20545 16499
rect 19536 16468 20545 16496
rect 19337 16459 19395 16465
rect 20533 16465 20545 16468
rect 20579 16465 20591 16499
rect 20533 16459 20591 16465
rect 15102 16428 15108 16440
rect 15063 16400 15108 16428
rect 15102 16388 15108 16400
rect 15160 16388 15166 16440
rect 14553 16363 14611 16369
rect 14553 16329 14565 16363
rect 14599 16329 14611 16363
rect 14553 16323 14611 16329
rect 17678 16292 17684 16304
rect 12360 16264 17684 16292
rect 17678 16252 17684 16264
rect 17736 16252 17742 16304
rect 19610 16252 19616 16304
rect 19668 16292 19674 16304
rect 19886 16292 19892 16304
rect 19668 16264 19892 16292
rect 19668 16252 19674 16264
rect 19886 16252 19892 16264
rect 19944 16252 19950 16304
rect 1104 16202 21620 16224
rect 1104 16150 4414 16202
rect 4466 16150 4478 16202
rect 4530 16150 4542 16202
rect 4594 16150 4606 16202
rect 4658 16150 11278 16202
rect 11330 16150 11342 16202
rect 11394 16150 11406 16202
rect 11458 16150 11470 16202
rect 11522 16150 18142 16202
rect 18194 16150 18206 16202
rect 18258 16150 18270 16202
rect 18322 16150 18334 16202
rect 18386 16150 21620 16202
rect 1104 16128 21620 16150
rect 3142 16088 3148 16100
rect 3103 16060 3148 16088
rect 3142 16048 3148 16060
rect 3200 16048 3206 16100
rect 7101 16091 7159 16097
rect 7101 16057 7113 16091
rect 7147 16088 7159 16091
rect 7282 16088 7288 16100
rect 7147 16060 7288 16088
rect 7147 16057 7159 16060
rect 7101 16051 7159 16057
rect 7282 16048 7288 16060
rect 7340 16048 7346 16100
rect 12526 16088 12532 16100
rect 11164 16060 12112 16088
rect 12487 16060 12532 16088
rect 6825 16023 6883 16029
rect 6825 15989 6837 16023
rect 6871 16020 6883 16023
rect 7374 16020 7380 16032
rect 6871 15992 7380 16020
rect 6871 15989 6883 15992
rect 6825 15983 6883 15989
rect 7374 15980 7380 15992
rect 7432 15980 7438 16032
rect 5074 15912 5080 15964
rect 5132 15952 5138 15964
rect 5445 15955 5503 15961
rect 5445 15952 5457 15955
rect 5132 15924 5457 15952
rect 5132 15912 5138 15924
rect 5445 15921 5457 15924
rect 5491 15921 5503 15955
rect 7650 15952 7656 15964
rect 5445 15915 5503 15921
rect 6564 15924 7656 15952
rect 1578 15844 1584 15896
rect 1636 15884 1642 15896
rect 1765 15887 1823 15893
rect 1765 15884 1777 15887
rect 1636 15856 1777 15884
rect 1636 15844 1642 15856
rect 1765 15853 1777 15856
rect 1811 15853 1823 15887
rect 1765 15847 1823 15853
rect 5712 15887 5770 15893
rect 5712 15853 5724 15887
rect 5758 15884 5770 15887
rect 6564 15884 6592 15924
rect 7650 15912 7656 15924
rect 7708 15912 7714 15964
rect 9861 15955 9919 15961
rect 9861 15921 9873 15955
rect 9907 15952 9919 15955
rect 10042 15952 10048 15964
rect 9907 15924 10048 15952
rect 9907 15921 9919 15924
rect 9861 15915 9919 15921
rect 10042 15912 10048 15924
rect 10100 15912 10106 15964
rect 11164 15961 11192 16060
rect 12084 16020 12112 16060
rect 12526 16048 12532 16060
rect 12584 16048 12590 16100
rect 12618 16048 12624 16100
rect 12676 16088 12682 16100
rect 15930 16088 15936 16100
rect 12676 16060 15936 16088
rect 12676 16048 12682 16060
rect 12636 16020 12664 16048
rect 12084 15992 12664 16020
rect 11149 15955 11207 15961
rect 11149 15921 11161 15955
rect 11195 15921 11207 15955
rect 11149 15915 11207 15921
rect 13446 15912 13452 15964
rect 13504 15952 13510 15964
rect 13556 15961 13584 16060
rect 15930 16048 15936 16060
rect 15988 16048 15994 16100
rect 16761 16091 16819 16097
rect 16761 16057 16773 16091
rect 16807 16088 16819 16091
rect 17954 16088 17960 16100
rect 16807 16060 17960 16088
rect 16807 16057 16819 16060
rect 16761 16051 16819 16057
rect 17954 16048 17960 16060
rect 18012 16048 18018 16100
rect 18874 16048 18880 16100
rect 18932 16088 18938 16100
rect 19889 16091 19947 16097
rect 19889 16088 19901 16091
rect 18932 16060 19901 16088
rect 18932 16048 18938 16060
rect 19889 16057 19901 16060
rect 19935 16057 19947 16091
rect 19889 16051 19947 16057
rect 20438 16020 20444 16032
rect 20399 15992 20444 16020
rect 20438 15980 20444 15992
rect 20496 15980 20502 16032
rect 13541 15955 13599 15961
rect 13541 15952 13553 15955
rect 13504 15924 13553 15952
rect 13504 15912 13510 15924
rect 13541 15921 13553 15924
rect 13587 15921 13599 15955
rect 17310 15952 17316 15964
rect 17271 15924 17316 15952
rect 13541 15915 13599 15921
rect 17310 15912 17316 15924
rect 17368 15912 17374 15964
rect 5758 15856 6592 15884
rect 7561 15887 7619 15893
rect 5758 15853 5770 15856
rect 5712 15847 5770 15853
rect 7561 15853 7573 15887
rect 7607 15884 7619 15887
rect 7742 15884 7748 15896
rect 7607 15856 7748 15884
rect 7607 15853 7619 15856
rect 7561 15847 7619 15853
rect 7742 15844 7748 15856
rect 7800 15844 7806 15896
rect 13808 15887 13866 15893
rect 13808 15853 13820 15887
rect 13854 15884 13866 15887
rect 14090 15884 14096 15896
rect 13854 15856 14096 15884
rect 13854 15853 13866 15856
rect 13808 15847 13866 15853
rect 14090 15844 14096 15856
rect 14148 15844 14154 15896
rect 15194 15844 15200 15896
rect 15252 15884 15258 15896
rect 17221 15887 17279 15893
rect 17221 15884 17233 15887
rect 15252 15856 17233 15884
rect 15252 15844 15258 15856
rect 17221 15853 17233 15856
rect 17267 15853 17279 15887
rect 17221 15847 17279 15853
rect 19150 15844 19156 15896
rect 19208 15884 19214 15896
rect 19705 15887 19763 15893
rect 19705 15884 19717 15887
rect 19208 15856 19717 15884
rect 19208 15844 19214 15856
rect 19705 15853 19717 15856
rect 19751 15853 19763 15887
rect 19705 15847 19763 15853
rect 19886 15844 19892 15896
rect 19944 15884 19950 15896
rect 20257 15887 20315 15893
rect 20257 15884 20269 15887
rect 19944 15856 20269 15884
rect 19944 15844 19950 15856
rect 20257 15853 20269 15856
rect 20303 15853 20315 15887
rect 20257 15847 20315 15853
rect 2032 15819 2090 15825
rect 2032 15785 2044 15819
rect 2078 15816 2090 15819
rect 2958 15816 2964 15828
rect 2078 15788 2964 15816
rect 2078 15785 2090 15788
rect 2032 15779 2090 15785
rect 2958 15776 2964 15788
rect 3016 15776 3022 15828
rect 11416 15819 11474 15825
rect 11416 15785 11428 15819
rect 11462 15816 11474 15819
rect 11698 15816 11704 15828
rect 11462 15788 11704 15816
rect 11462 15785 11474 15788
rect 11416 15779 11474 15785
rect 11698 15776 11704 15788
rect 11756 15776 11762 15828
rect 14366 15776 14372 15828
rect 14424 15816 14430 15828
rect 17129 15819 17187 15825
rect 17129 15816 17141 15819
rect 14424 15788 17141 15816
rect 14424 15776 14430 15788
rect 15212 15760 15240 15788
rect 17129 15785 17141 15788
rect 17175 15785 17187 15819
rect 17129 15779 17187 15785
rect 7469 15751 7527 15757
rect 7469 15717 7481 15751
rect 7515 15748 7527 15751
rect 7742 15748 7748 15760
rect 7515 15720 7748 15748
rect 7515 15717 7527 15720
rect 7469 15711 7527 15717
rect 7742 15708 7748 15720
rect 7800 15708 7806 15760
rect 14550 15708 14556 15760
rect 14608 15748 14614 15760
rect 14921 15751 14979 15757
rect 14921 15748 14933 15751
rect 14608 15720 14933 15748
rect 14608 15708 14614 15720
rect 14921 15717 14933 15720
rect 14967 15748 14979 15751
rect 15102 15748 15108 15760
rect 14967 15720 15108 15748
rect 14967 15717 14979 15720
rect 14921 15711 14979 15717
rect 15102 15708 15108 15720
rect 15160 15708 15166 15760
rect 15194 15708 15200 15760
rect 15252 15708 15258 15760
rect 1104 15658 21620 15680
rect 1104 15606 7846 15658
rect 7898 15606 7910 15658
rect 7962 15606 7974 15658
rect 8026 15606 8038 15658
rect 8090 15606 14710 15658
rect 14762 15606 14774 15658
rect 14826 15606 14838 15658
rect 14890 15606 14902 15658
rect 14954 15606 21620 15658
rect 1104 15584 21620 15606
rect 2961 15547 3019 15553
rect 2961 15513 2973 15547
rect 3007 15513 3019 15547
rect 2961 15507 3019 15513
rect 6273 15547 6331 15553
rect 6273 15513 6285 15547
rect 6319 15544 6331 15547
rect 7650 15544 7656 15556
rect 6319 15516 7656 15544
rect 6319 15513 6331 15516
rect 6273 15507 6331 15513
rect 2976 15476 3004 15507
rect 7650 15504 7656 15516
rect 7708 15504 7714 15556
rect 20714 15544 20720 15556
rect 20675 15516 20720 15544
rect 20714 15504 20720 15516
rect 20772 15504 20778 15556
rect 19150 15476 19156 15488
rect 2976 15448 19012 15476
rect 19111 15448 19156 15476
rect 3329 15411 3387 15417
rect 3329 15377 3341 15411
rect 3375 15408 3387 15411
rect 3973 15411 4031 15417
rect 3973 15408 3985 15411
rect 3375 15380 3985 15408
rect 3375 15377 3387 15380
rect 3329 15371 3387 15377
rect 3973 15377 3985 15380
rect 4019 15377 4031 15411
rect 3973 15371 4031 15377
rect 4893 15411 4951 15417
rect 4893 15377 4905 15411
rect 4939 15408 4951 15411
rect 4982 15408 4988 15420
rect 4939 15380 4988 15408
rect 4939 15377 4951 15380
rect 4893 15371 4951 15377
rect 4982 15368 4988 15380
rect 5040 15368 5046 15420
rect 5160 15411 5218 15417
rect 5160 15377 5172 15411
rect 5206 15408 5218 15411
rect 6822 15408 6828 15420
rect 5206 15380 6828 15408
rect 5206 15377 5218 15380
rect 5160 15371 5218 15377
rect 6822 15368 6828 15380
rect 6880 15368 6886 15420
rect 16574 15408 16580 15420
rect 16535 15380 16580 15408
rect 16574 15368 16580 15380
rect 16632 15368 16638 15420
rect 18877 15411 18935 15417
rect 18877 15377 18889 15411
rect 18923 15377 18935 15411
rect 18984 15408 19012 15448
rect 19150 15436 19156 15448
rect 19208 15436 19214 15488
rect 19886 15476 19892 15488
rect 19847 15448 19892 15476
rect 19886 15436 19892 15448
rect 19944 15436 19950 15488
rect 19613 15411 19671 15417
rect 19613 15408 19625 15411
rect 18984 15380 19625 15408
rect 18877 15371 18935 15377
rect 19613 15377 19625 15380
rect 19659 15377 19671 15411
rect 19613 15371 19671 15377
rect 2958 15300 2964 15352
rect 3016 15300 3022 15352
rect 3418 15340 3424 15352
rect 3379 15312 3424 15340
rect 3418 15300 3424 15312
rect 3476 15300 3482 15352
rect 3513 15343 3571 15349
rect 3513 15309 3525 15343
rect 3559 15309 3571 15343
rect 16666 15340 16672 15352
rect 16627 15312 16672 15340
rect 3513 15303 3571 15309
rect 2976 15272 3004 15300
rect 3528 15272 3556 15303
rect 16666 15300 16672 15312
rect 16724 15300 16730 15352
rect 16758 15300 16764 15352
rect 16816 15340 16822 15352
rect 16816 15312 16861 15340
rect 16816 15300 16822 15312
rect 2976 15244 3556 15272
rect 15102 15232 15108 15284
rect 15160 15272 15166 15284
rect 18892 15272 18920 15371
rect 20070 15368 20076 15420
rect 20128 15408 20134 15420
rect 20533 15411 20591 15417
rect 20533 15408 20545 15411
rect 20128 15380 20545 15408
rect 20128 15368 20134 15380
rect 20533 15377 20545 15380
rect 20579 15377 20591 15411
rect 20533 15371 20591 15377
rect 15160 15244 18920 15272
rect 15160 15232 15166 15244
rect 16209 15207 16267 15213
rect 16209 15173 16221 15207
rect 16255 15204 16267 15207
rect 17862 15204 17868 15216
rect 16255 15176 17868 15204
rect 16255 15173 16267 15176
rect 16209 15167 16267 15173
rect 17862 15164 17868 15176
rect 17920 15164 17926 15216
rect 1104 15114 21620 15136
rect 1104 15062 4414 15114
rect 4466 15062 4478 15114
rect 4530 15062 4542 15114
rect 4594 15062 4606 15114
rect 4658 15062 11278 15114
rect 11330 15062 11342 15114
rect 11394 15062 11406 15114
rect 11458 15062 11470 15114
rect 11522 15062 18142 15114
rect 18194 15062 18206 15114
rect 18258 15062 18270 15114
rect 18322 15062 18334 15114
rect 18386 15062 21620 15114
rect 1104 15040 21620 15062
rect 2498 14960 2504 15012
rect 2556 14960 2562 15012
rect 2958 15000 2964 15012
rect 2919 14972 2964 15000
rect 2958 14960 2964 14972
rect 3016 14960 3022 15012
rect 3418 14960 3424 15012
rect 3476 15000 3482 15012
rect 4065 15003 4123 15009
rect 4065 15000 4077 15003
rect 3476 14972 4077 15000
rect 3476 14960 3482 14972
rect 4065 14969 4077 14972
rect 4111 14969 4123 15003
rect 4065 14963 4123 14969
rect 6822 14960 6828 15012
rect 6880 15000 6886 15012
rect 9309 15003 9367 15009
rect 9309 15000 9321 15003
rect 6880 14972 9321 15000
rect 6880 14960 6886 14972
rect 9309 14969 9321 14972
rect 9355 14969 9367 15003
rect 9309 14963 9367 14969
rect 9677 15003 9735 15009
rect 9677 14969 9689 15003
rect 9723 15000 9735 15003
rect 15102 15000 15108 15012
rect 9723 14972 15108 15000
rect 9723 14969 9735 14972
rect 9677 14963 9735 14969
rect 2516 14932 2544 14960
rect 2516 14904 7604 14932
rect 1578 14864 1584 14876
rect 1539 14836 1584 14864
rect 1578 14824 1584 14836
rect 1636 14824 1642 14876
rect 3694 14824 3700 14876
rect 3752 14864 3758 14876
rect 4617 14867 4675 14873
rect 4617 14864 4629 14867
rect 3752 14836 4629 14864
rect 3752 14824 3758 14836
rect 4617 14833 4629 14836
rect 4663 14833 4675 14867
rect 7466 14864 7472 14876
rect 4617 14827 4675 14833
rect 7116 14836 7472 14864
rect 4246 14756 4252 14808
rect 4304 14796 4310 14808
rect 4525 14799 4583 14805
rect 4525 14796 4537 14799
rect 4304 14768 4537 14796
rect 4304 14756 4310 14768
rect 4525 14765 4537 14768
rect 4571 14765 4583 14799
rect 4525 14759 4583 14765
rect 1848 14731 1906 14737
rect 1848 14697 1860 14731
rect 1894 14728 1906 14731
rect 3694 14728 3700 14740
rect 1894 14700 3700 14728
rect 1894 14697 1906 14700
rect 1848 14691 1906 14697
rect 3694 14688 3700 14700
rect 3752 14688 3758 14740
rect 4433 14731 4491 14737
rect 4433 14697 4445 14731
rect 4479 14728 4491 14731
rect 7116 14728 7144 14836
rect 7466 14824 7472 14836
rect 7524 14824 7530 14876
rect 7576 14864 7604 14904
rect 9324 14864 9352 14963
rect 15102 14960 15108 14972
rect 15160 14960 15166 15012
rect 16117 15003 16175 15009
rect 16117 14969 16129 15003
rect 16163 15000 16175 15003
rect 16666 15000 16672 15012
rect 16163 14972 16672 15000
rect 16163 14969 16175 14972
rect 16117 14963 16175 14969
rect 16666 14960 16672 14972
rect 16724 14960 16730 15012
rect 20438 15000 20444 15012
rect 20399 14972 20444 15000
rect 20438 14960 20444 14972
rect 20496 14960 20502 15012
rect 9398 14892 9404 14944
rect 9456 14932 9462 14944
rect 12158 14932 12164 14944
rect 9456 14904 12164 14932
rect 9456 14892 9462 14904
rect 12158 14892 12164 14904
rect 12216 14892 12222 14944
rect 12253 14935 12311 14941
rect 12253 14901 12265 14935
rect 12299 14901 12311 14935
rect 12253 14895 12311 14901
rect 10229 14867 10287 14873
rect 10229 14864 10241 14867
rect 7576 14836 8064 14864
rect 9324 14836 10241 14864
rect 7193 14799 7251 14805
rect 7193 14765 7205 14799
rect 7239 14796 7251 14799
rect 7239 14768 7604 14796
rect 7239 14765 7251 14768
rect 7193 14759 7251 14765
rect 4479 14700 7144 14728
rect 4479 14697 4491 14700
rect 4433 14691 4491 14697
rect 5074 14620 5080 14672
rect 5132 14660 5138 14672
rect 7009 14663 7067 14669
rect 7009 14660 7021 14663
rect 5132 14632 7021 14660
rect 5132 14620 5138 14632
rect 7009 14629 7021 14632
rect 7055 14629 7067 14663
rect 7576 14660 7604 14768
rect 7650 14756 7656 14808
rect 7708 14796 7714 14808
rect 7926 14796 7932 14808
rect 7708 14768 7932 14796
rect 7708 14756 7714 14768
rect 7926 14756 7932 14768
rect 7984 14756 7990 14808
rect 8036 14796 8064 14836
rect 10229 14833 10241 14836
rect 10275 14833 10287 14867
rect 12268 14864 12296 14895
rect 12802 14864 12808 14876
rect 12268 14836 12725 14864
rect 12763 14836 12808 14864
rect 10229 14827 10287 14833
rect 12250 14796 12256 14808
rect 8036 14768 12256 14796
rect 12250 14756 12256 14768
rect 12308 14756 12314 14808
rect 12697 14796 12725 14836
rect 12802 14824 12808 14836
rect 12860 14824 12866 14876
rect 13556 14836 15332 14864
rect 13556 14796 13584 14836
rect 12697 14768 13584 14796
rect 13633 14799 13691 14805
rect 13633 14765 13645 14799
rect 13679 14796 13691 14799
rect 13906 14796 13912 14808
rect 13679 14768 13912 14796
rect 13679 14765 13691 14768
rect 13633 14759 13691 14765
rect 13906 14756 13912 14768
rect 13964 14756 13970 14808
rect 15304 14796 15332 14836
rect 15378 14824 15384 14876
rect 15436 14864 15442 14876
rect 16577 14867 16635 14873
rect 16577 14864 16589 14867
rect 15436 14836 16589 14864
rect 15436 14824 15442 14836
rect 16577 14833 16589 14836
rect 16623 14833 16635 14867
rect 16758 14864 16764 14876
rect 16719 14836 16764 14864
rect 16577 14827 16635 14833
rect 16758 14824 16764 14836
rect 16816 14824 16822 14876
rect 17770 14796 17776 14808
rect 15304 14768 17776 14796
rect 17770 14756 17776 14768
rect 17828 14756 17834 14808
rect 17862 14756 17868 14808
rect 17920 14796 17926 14808
rect 18877 14799 18935 14805
rect 18877 14796 18889 14799
rect 17920 14768 18889 14796
rect 17920 14756 17926 14768
rect 18877 14765 18889 14768
rect 18923 14765 18935 14799
rect 18877 14759 18935 14765
rect 19334 14756 19340 14808
rect 19392 14796 19398 14808
rect 20257 14799 20315 14805
rect 20257 14796 20269 14799
rect 19392 14768 20269 14796
rect 19392 14756 19398 14768
rect 20257 14765 20269 14768
rect 20303 14765 20315 14799
rect 20257 14759 20315 14765
rect 8196 14731 8254 14737
rect 8196 14697 8208 14731
rect 8242 14728 8254 14731
rect 8662 14728 8668 14740
rect 8242 14700 8668 14728
rect 8242 14697 8254 14700
rect 8196 14691 8254 14697
rect 8662 14688 8668 14700
rect 8720 14688 8726 14740
rect 19153 14731 19211 14737
rect 19153 14697 19165 14731
rect 19199 14728 19211 14731
rect 20530 14728 20536 14740
rect 19199 14700 20536 14728
rect 19199 14697 19211 14700
rect 19153 14691 19211 14697
rect 20530 14688 20536 14700
rect 20588 14688 20594 14740
rect 9030 14660 9036 14672
rect 7576 14632 9036 14660
rect 7009 14623 7067 14629
rect 9030 14620 9036 14632
rect 9088 14620 9094 14672
rect 9766 14620 9772 14672
rect 9824 14660 9830 14672
rect 10045 14663 10103 14669
rect 10045 14660 10057 14663
rect 9824 14632 10057 14660
rect 9824 14620 9830 14632
rect 10045 14629 10057 14632
rect 10091 14629 10103 14663
rect 10045 14623 10103 14629
rect 10134 14620 10140 14672
rect 10192 14660 10198 14672
rect 12618 14660 12624 14672
rect 10192 14632 10237 14660
rect 12579 14632 12624 14660
rect 10192 14620 10198 14632
rect 12618 14620 12624 14632
rect 12676 14620 12682 14672
rect 12710 14620 12716 14672
rect 12768 14660 12774 14672
rect 13446 14660 13452 14672
rect 12768 14632 12813 14660
rect 13407 14632 13452 14660
rect 12768 14620 12774 14632
rect 13446 14620 13452 14632
rect 13504 14620 13510 14672
rect 15470 14620 15476 14672
rect 15528 14660 15534 14672
rect 16298 14660 16304 14672
rect 15528 14632 16304 14660
rect 15528 14620 15534 14632
rect 16298 14620 16304 14632
rect 16356 14660 16362 14672
rect 16485 14663 16543 14669
rect 16485 14660 16497 14663
rect 16356 14632 16497 14660
rect 16356 14620 16362 14632
rect 16485 14629 16497 14632
rect 16531 14629 16543 14663
rect 16485 14623 16543 14629
rect 1104 14570 21620 14592
rect 1104 14518 7846 14570
rect 7898 14518 7910 14570
rect 7962 14518 7974 14570
rect 8026 14518 8038 14570
rect 8090 14518 14710 14570
rect 14762 14518 14774 14570
rect 14826 14518 14838 14570
rect 14890 14518 14902 14570
rect 14954 14518 21620 14570
rect 1104 14496 21620 14518
rect 5350 14416 5356 14468
rect 5408 14456 5414 14468
rect 6089 14459 6147 14465
rect 6089 14456 6101 14459
rect 5408 14428 6101 14456
rect 5408 14416 5414 14428
rect 6089 14425 6101 14428
rect 6135 14425 6147 14459
rect 8662 14456 8668 14468
rect 8623 14428 8668 14456
rect 6089 14419 6147 14425
rect 8662 14416 8668 14428
rect 8720 14416 8726 14468
rect 9766 14456 9772 14468
rect 9727 14428 9772 14456
rect 9766 14416 9772 14428
rect 9824 14416 9830 14468
rect 12069 14459 12127 14465
rect 12069 14425 12081 14459
rect 12115 14425 12127 14459
rect 12069 14419 12127 14425
rect 12437 14459 12495 14465
rect 12437 14425 12449 14459
rect 12483 14456 12495 14459
rect 12710 14456 12716 14468
rect 12483 14428 12716 14456
rect 12483 14425 12495 14428
rect 12437 14419 12495 14425
rect 4148 14391 4206 14397
rect 4148 14357 4160 14391
rect 4194 14388 4206 14391
rect 7552 14391 7610 14397
rect 4194 14360 7512 14388
rect 4194 14357 4206 14360
rect 4148 14351 4206 14357
rect 1578 14280 1584 14332
rect 1636 14320 1642 14332
rect 2314 14320 2320 14332
rect 1636 14292 2320 14320
rect 1636 14280 1642 14292
rect 2314 14280 2320 14292
rect 2372 14320 2378 14332
rect 3881 14323 3939 14329
rect 3881 14320 3893 14323
rect 2372 14292 3893 14320
rect 2372 14280 2378 14292
rect 3881 14289 3893 14292
rect 3927 14320 3939 14323
rect 4890 14320 4896 14332
rect 3927 14292 4896 14320
rect 3927 14289 3939 14292
rect 3881 14283 3939 14289
rect 4890 14280 4896 14292
rect 4948 14320 4954 14332
rect 5074 14320 5080 14332
rect 4948 14292 5080 14320
rect 4948 14280 4954 14292
rect 5074 14280 5080 14292
rect 5132 14280 5138 14332
rect 5997 14323 6055 14329
rect 5997 14289 6009 14323
rect 6043 14320 6055 14323
rect 7006 14320 7012 14332
rect 6043 14292 7012 14320
rect 6043 14289 6055 14292
rect 5997 14283 6055 14289
rect 7006 14280 7012 14292
rect 7064 14280 7070 14332
rect 7484 14320 7512 14360
rect 7552 14357 7564 14391
rect 7598 14388 7610 14391
rect 9398 14388 9404 14400
rect 7598 14360 9404 14388
rect 7598 14357 7610 14360
rect 7552 14351 7610 14357
rect 9398 14348 9404 14360
rect 9456 14348 9462 14400
rect 12084 14388 12112 14419
rect 12710 14416 12716 14428
rect 12768 14416 12774 14468
rect 12805 14459 12863 14465
rect 12805 14425 12817 14459
rect 12851 14456 12863 14459
rect 15470 14456 15476 14468
rect 12851 14428 15476 14456
rect 12851 14425 12863 14428
rect 12805 14419 12863 14425
rect 15470 14416 15476 14428
rect 15528 14416 15534 14468
rect 15565 14459 15623 14465
rect 15565 14425 15577 14459
rect 15611 14425 15623 14459
rect 15565 14419 15623 14425
rect 12161 14391 12219 14397
rect 12161 14388 12173 14391
rect 9508 14360 12173 14388
rect 9508 14320 9536 14360
rect 12161 14357 12173 14360
rect 12207 14357 12219 14391
rect 12161 14351 12219 14357
rect 12250 14348 12256 14400
rect 12308 14388 12314 14400
rect 12897 14391 12955 14397
rect 12897 14388 12909 14391
rect 12308 14360 12909 14388
rect 12308 14348 12314 14360
rect 12897 14357 12909 14360
rect 12943 14357 12955 14391
rect 12897 14351 12955 14357
rect 13446 14348 13452 14400
rect 13504 14388 13510 14400
rect 14452 14391 14510 14397
rect 13504 14360 14228 14388
rect 13504 14348 13510 14360
rect 10962 14329 10968 14332
rect 7484 14292 9536 14320
rect 10945 14323 10968 14329
rect 10945 14289 10957 14323
rect 10945 14283 10968 14289
rect 10962 14280 10968 14283
rect 11020 14280 11026 14332
rect 14200 14329 14228 14360
rect 14452 14357 14464 14391
rect 14498 14388 14510 14391
rect 14550 14388 14556 14400
rect 14498 14360 14556 14388
rect 14498 14357 14510 14360
rect 14452 14351 14510 14357
rect 14550 14348 14556 14360
rect 14608 14348 14614 14400
rect 15580 14388 15608 14419
rect 16850 14416 16856 14468
rect 16908 14456 16914 14468
rect 17221 14459 17279 14465
rect 17221 14456 17233 14459
rect 16908 14428 17233 14456
rect 16908 14416 16914 14428
rect 17221 14425 17233 14428
rect 17267 14425 17279 14459
rect 18690 14456 18696 14468
rect 18651 14428 18696 14456
rect 17221 14419 17279 14425
rect 18690 14416 18696 14428
rect 18748 14416 18754 14468
rect 20622 14416 20628 14468
rect 20680 14456 20686 14468
rect 20717 14459 20775 14465
rect 20717 14456 20729 14459
rect 20680 14428 20729 14456
rect 20680 14416 20686 14428
rect 20717 14425 20729 14428
rect 20763 14425 20775 14459
rect 20717 14419 20775 14425
rect 16108 14391 16166 14397
rect 16108 14388 16120 14391
rect 15580 14360 16120 14388
rect 16108 14357 16120 14360
rect 16154 14388 16166 14391
rect 16758 14388 16764 14400
rect 16154 14360 16764 14388
rect 16154 14357 16166 14360
rect 16108 14351 16166 14357
rect 16758 14348 16764 14360
rect 16816 14348 16822 14400
rect 17770 14348 17776 14400
rect 17828 14388 17834 14400
rect 19334 14388 19340 14400
rect 17828 14360 19104 14388
rect 19295 14360 19340 14388
rect 17828 14348 17834 14360
rect 14185 14323 14243 14329
rect 14185 14289 14197 14323
rect 14231 14320 14243 14323
rect 15841 14323 15899 14329
rect 15841 14320 15853 14323
rect 14231 14292 15853 14320
rect 14231 14289 14243 14292
rect 14185 14283 14243 14289
rect 15841 14289 15853 14292
rect 15887 14289 15899 14323
rect 18506 14320 18512 14332
rect 18467 14292 18512 14320
rect 15841 14283 15899 14289
rect 18506 14280 18512 14292
rect 18564 14280 18570 14332
rect 19076 14329 19104 14360
rect 19334 14348 19340 14360
rect 19392 14348 19398 14400
rect 20070 14388 20076 14400
rect 20031 14360 20076 14388
rect 20070 14348 20076 14360
rect 20128 14348 20134 14400
rect 19061 14323 19119 14329
rect 19061 14289 19073 14323
rect 19107 14289 19119 14323
rect 19061 14283 19119 14289
rect 19794 14280 19800 14332
rect 19852 14329 19858 14332
rect 19852 14323 19865 14329
rect 19853 14320 19865 14323
rect 20530 14320 20536 14332
rect 19853 14292 19897 14320
rect 20491 14292 20536 14320
rect 19853 14289 19865 14292
rect 19852 14283 19865 14289
rect 19852 14280 19858 14283
rect 20530 14280 20536 14292
rect 20588 14280 20594 14332
rect 6181 14255 6239 14261
rect 6181 14221 6193 14255
rect 6227 14221 6239 14255
rect 6181 14215 6239 14221
rect 7285 14255 7343 14261
rect 7285 14221 7297 14255
rect 7331 14221 7343 14255
rect 7285 14215 7343 14221
rect 10689 14255 10747 14261
rect 10689 14221 10701 14255
rect 10735 14221 10747 14255
rect 10689 14215 10747 14221
rect 12989 14255 13047 14261
rect 12989 14221 13001 14255
rect 13035 14221 13047 14255
rect 13446 14252 13452 14264
rect 13407 14224 13452 14252
rect 12989 14215 13047 14221
rect 5074 14144 5080 14196
rect 5132 14184 5138 14196
rect 5261 14187 5319 14193
rect 5261 14184 5273 14187
rect 5132 14156 5273 14184
rect 5132 14144 5138 14156
rect 5261 14153 5273 14156
rect 5307 14184 5319 14187
rect 6196 14184 6224 14215
rect 5307 14156 6224 14184
rect 5307 14153 5319 14156
rect 5261 14147 5319 14153
rect 5629 14119 5687 14125
rect 5629 14085 5641 14119
rect 5675 14116 5687 14119
rect 6914 14116 6920 14128
rect 5675 14088 6920 14116
rect 5675 14085 5687 14088
rect 5629 14079 5687 14085
rect 6914 14076 6920 14088
rect 6972 14076 6978 14128
rect 7300 14116 7328 14215
rect 8294 14144 8300 14196
rect 8352 14184 8358 14196
rect 9950 14184 9956 14196
rect 8352 14156 9956 14184
rect 8352 14144 8358 14156
rect 9950 14144 9956 14156
rect 10008 14184 10014 14196
rect 10704 14184 10732 14215
rect 10008 14156 10732 14184
rect 10008 14144 10014 14156
rect 12526 14144 12532 14196
rect 12584 14184 12590 14196
rect 13004 14184 13032 14215
rect 13446 14212 13452 14224
rect 13504 14212 13510 14264
rect 17494 14252 17500 14264
rect 17455 14224 17500 14252
rect 17494 14212 17500 14224
rect 17552 14212 17558 14264
rect 12584 14156 13032 14184
rect 12584 14144 12590 14156
rect 7650 14116 7656 14128
rect 7300 14088 7656 14116
rect 7650 14076 7656 14088
rect 7708 14076 7714 14128
rect 7926 14076 7932 14128
rect 7984 14116 7990 14128
rect 12066 14116 12072 14128
rect 7984 14088 12072 14116
rect 7984 14076 7990 14088
rect 12066 14076 12072 14088
rect 12124 14076 12130 14128
rect 12161 14119 12219 14125
rect 12161 14085 12173 14119
rect 12207 14116 12219 14119
rect 12802 14116 12808 14128
rect 12207 14088 12808 14116
rect 12207 14085 12219 14088
rect 12161 14079 12219 14085
rect 12802 14076 12808 14088
rect 12860 14076 12866 14128
rect 1104 14026 21620 14048
rect 1104 13974 4414 14026
rect 4466 13974 4478 14026
rect 4530 13974 4542 14026
rect 4594 13974 4606 14026
rect 4658 13974 11278 14026
rect 11330 13974 11342 14026
rect 11394 13974 11406 14026
rect 11458 13974 11470 14026
rect 11522 13974 18142 14026
rect 18194 13974 18206 14026
rect 18258 13974 18270 14026
rect 18322 13974 18334 14026
rect 18386 13974 21620 14026
rect 1104 13952 21620 13974
rect 3694 13912 3700 13924
rect 3655 13884 3700 13912
rect 3694 13872 3700 13884
rect 3752 13872 3758 13924
rect 6181 13915 6239 13921
rect 6181 13912 6193 13915
rect 4724 13884 6193 13912
rect 2314 13776 2320 13788
rect 2275 13748 2320 13776
rect 2314 13736 2320 13748
rect 2372 13736 2378 13788
rect 2584 13711 2642 13717
rect 2584 13677 2596 13711
rect 2630 13708 2642 13711
rect 4724 13708 4752 13884
rect 6181 13881 6193 13884
rect 6227 13881 6239 13915
rect 6181 13875 6239 13881
rect 6457 13915 6515 13921
rect 6457 13881 6469 13915
rect 6503 13912 6515 13915
rect 8021 13915 8079 13921
rect 6503 13884 7972 13912
rect 6503 13881 6515 13884
rect 6457 13875 6515 13881
rect 6196 13844 6224 13875
rect 7944 13844 7972 13884
rect 8021 13881 8033 13915
rect 8067 13912 8079 13915
rect 10134 13912 10140 13924
rect 8067 13884 10140 13912
rect 8067 13881 8079 13884
rect 8021 13875 8079 13881
rect 10134 13872 10140 13884
rect 10192 13872 10198 13924
rect 10962 13872 10968 13924
rect 11020 13912 11026 13924
rect 11241 13915 11299 13921
rect 11241 13912 11253 13915
rect 11020 13884 11253 13912
rect 11020 13872 11026 13884
rect 11241 13881 11253 13884
rect 11287 13912 11299 13915
rect 12526 13912 12532 13924
rect 11287 13884 12532 13912
rect 11287 13881 11299 13884
rect 11241 13875 11299 13881
rect 12526 13872 12532 13884
rect 12584 13872 12590 13924
rect 12618 13872 12624 13924
rect 12676 13912 12682 13924
rect 12713 13915 12771 13921
rect 12713 13912 12725 13915
rect 12676 13884 12725 13912
rect 12676 13872 12682 13884
rect 12713 13881 12725 13884
rect 12759 13881 12771 13915
rect 16574 13912 16580 13924
rect 16535 13884 16580 13912
rect 12713 13875 12771 13881
rect 16574 13872 16580 13884
rect 16632 13872 16638 13924
rect 16666 13872 16672 13924
rect 16724 13912 16730 13924
rect 20438 13912 20444 13924
rect 16724 13884 20300 13912
rect 20399 13884 20444 13912
rect 16724 13872 16730 13884
rect 9858 13844 9864 13856
rect 6196 13816 7052 13844
rect 7944 13816 9864 13844
rect 6914 13776 6920 13788
rect 6875 13748 6920 13776
rect 6914 13736 6920 13748
rect 6972 13736 6978 13788
rect 7024 13785 7052 13816
rect 9858 13804 9864 13816
rect 9916 13804 9922 13856
rect 19886 13804 19892 13856
rect 19944 13844 19950 13856
rect 19944 13816 19989 13844
rect 19944 13804 19950 13816
rect 7009 13779 7067 13785
rect 7009 13745 7021 13779
rect 7055 13745 7067 13779
rect 8478 13776 8484 13788
rect 8439 13748 8484 13776
rect 7009 13739 7067 13745
rect 8478 13736 8484 13748
rect 8536 13736 8542 13788
rect 8662 13776 8668 13788
rect 8623 13748 8668 13776
rect 8662 13736 8668 13748
rect 8720 13736 8726 13788
rect 12526 13736 12532 13788
rect 12584 13776 12590 13788
rect 13265 13779 13323 13785
rect 13265 13776 13277 13779
rect 12584 13748 13277 13776
rect 12584 13736 12590 13748
rect 13265 13745 13277 13748
rect 13311 13745 13323 13779
rect 13265 13739 13323 13745
rect 16758 13736 16764 13788
rect 16816 13776 16822 13788
rect 17129 13779 17187 13785
rect 17129 13776 17141 13779
rect 16816 13748 17141 13776
rect 16816 13736 16822 13748
rect 17129 13745 17141 13748
rect 17175 13745 17187 13779
rect 17129 13739 17187 13745
rect 18417 13779 18475 13785
rect 18417 13745 18429 13779
rect 18463 13776 18475 13779
rect 18506 13776 18512 13788
rect 18463 13748 18512 13776
rect 18463 13745 18475 13748
rect 18417 13739 18475 13745
rect 18506 13736 18512 13748
rect 18564 13736 18570 13788
rect 2630 13680 4752 13708
rect 4801 13711 4859 13717
rect 2630 13677 2642 13680
rect 2584 13671 2642 13677
rect 4801 13677 4813 13711
rect 4847 13708 4859 13711
rect 4890 13708 4896 13720
rect 4847 13680 4896 13708
rect 4847 13677 4859 13680
rect 4801 13671 4859 13677
rect 4890 13668 4896 13680
rect 4948 13668 4954 13720
rect 5074 13717 5080 13720
rect 5068 13708 5080 13717
rect 5035 13680 5080 13708
rect 5068 13671 5080 13680
rect 5074 13668 5080 13671
rect 5132 13668 5138 13720
rect 9217 13711 9275 13717
rect 9217 13677 9229 13711
rect 9263 13708 9275 13711
rect 9766 13708 9772 13720
rect 9263 13680 9772 13708
rect 9263 13677 9275 13680
rect 9217 13671 9275 13677
rect 9766 13668 9772 13680
rect 9824 13668 9830 13720
rect 9861 13711 9919 13717
rect 9861 13677 9873 13711
rect 9907 13677 9919 13711
rect 9861 13671 9919 13677
rect 13081 13711 13139 13717
rect 13081 13677 13093 13711
rect 13127 13708 13139 13711
rect 13446 13708 13452 13720
rect 13127 13680 13452 13708
rect 13127 13677 13139 13680
rect 13081 13671 13139 13677
rect 7006 13600 7012 13652
rect 7064 13640 7070 13652
rect 8389 13643 8447 13649
rect 8389 13640 8401 13643
rect 7064 13612 8401 13640
rect 7064 13600 7070 13612
rect 8389 13609 8401 13612
rect 8435 13640 8447 13643
rect 9876 13640 9904 13671
rect 13446 13668 13452 13680
rect 13504 13668 13510 13720
rect 16945 13711 17003 13717
rect 13556 13680 16896 13708
rect 9950 13640 9956 13652
rect 8435 13612 9168 13640
rect 9876 13612 9956 13640
rect 8435 13609 8447 13612
rect 8389 13603 8447 13609
rect 6822 13572 6828 13584
rect 6783 13544 6828 13572
rect 6822 13532 6828 13544
rect 6880 13532 6886 13584
rect 9030 13572 9036 13584
rect 8991 13544 9036 13572
rect 9030 13532 9036 13544
rect 9088 13532 9094 13584
rect 9140 13572 9168 13612
rect 9950 13600 9956 13612
rect 10008 13600 10014 13652
rect 10128 13643 10186 13649
rect 10128 13609 10140 13643
rect 10174 13640 10186 13643
rect 10410 13640 10416 13652
rect 10174 13612 10416 13640
rect 10174 13609 10186 13612
rect 10128 13603 10186 13609
rect 10410 13600 10416 13612
rect 10468 13600 10474 13652
rect 13173 13643 13231 13649
rect 13173 13609 13185 13643
rect 13219 13640 13231 13643
rect 13556 13640 13584 13680
rect 13219 13612 13584 13640
rect 16868 13640 16896 13680
rect 16945 13677 16957 13711
rect 16991 13708 17003 13711
rect 17494 13708 17500 13720
rect 16991 13680 17500 13708
rect 16991 13677 17003 13680
rect 16945 13671 17003 13677
rect 17494 13668 17500 13680
rect 17552 13668 17558 13720
rect 18141 13711 18199 13717
rect 18141 13677 18153 13711
rect 18187 13708 18199 13711
rect 19705 13711 19763 13717
rect 18187 13680 18552 13708
rect 18187 13677 18199 13680
rect 18141 13671 18199 13677
rect 18524 13652 18552 13680
rect 19705 13677 19717 13711
rect 19751 13708 19763 13711
rect 19794 13708 19800 13720
rect 19751 13680 19800 13708
rect 19751 13677 19763 13680
rect 19705 13671 19763 13677
rect 19794 13668 19800 13680
rect 19852 13668 19858 13720
rect 20272 13717 20300 13884
rect 20438 13872 20444 13884
rect 20496 13872 20502 13924
rect 20257 13711 20315 13717
rect 20257 13677 20269 13711
rect 20303 13677 20315 13711
rect 20257 13671 20315 13677
rect 17037 13643 17095 13649
rect 17037 13640 17049 13643
rect 16868 13612 17049 13640
rect 13219 13609 13231 13612
rect 13173 13603 13231 13609
rect 17037 13609 17049 13612
rect 17083 13640 17095 13643
rect 17402 13640 17408 13652
rect 17083 13612 17408 13640
rect 17083 13609 17095 13612
rect 17037 13603 17095 13609
rect 17402 13600 17408 13612
rect 17460 13600 17466 13652
rect 18506 13600 18512 13652
rect 18564 13600 18570 13652
rect 14366 13572 14372 13584
rect 9140 13544 14372 13572
rect 14366 13532 14372 13544
rect 14424 13532 14430 13584
rect 1104 13482 21620 13504
rect 1104 13430 7846 13482
rect 7898 13430 7910 13482
rect 7962 13430 7974 13482
rect 8026 13430 8038 13482
rect 8090 13430 14710 13482
rect 14762 13430 14774 13482
rect 14826 13430 14838 13482
rect 14890 13430 14902 13482
rect 14954 13430 21620 13482
rect 1104 13408 21620 13430
rect 6089 13371 6147 13377
rect 6089 13337 6101 13371
rect 6135 13368 6147 13371
rect 6822 13368 6828 13380
rect 6135 13340 6828 13368
rect 6135 13337 6147 13340
rect 6089 13331 6147 13337
rect 6822 13328 6828 13340
rect 6880 13328 6886 13380
rect 9766 13328 9772 13380
rect 9824 13368 9830 13380
rect 10962 13368 10968 13380
rect 9824 13340 10968 13368
rect 9824 13328 9830 13340
rect 10962 13328 10968 13340
rect 11020 13368 11026 13380
rect 11425 13371 11483 13377
rect 11425 13368 11437 13371
rect 11020 13340 11437 13368
rect 11020 13328 11026 13340
rect 11425 13337 11437 13340
rect 11471 13337 11483 13371
rect 19702 13368 19708 13380
rect 19663 13340 19708 13368
rect 11425 13331 11483 13337
rect 19702 13328 19708 13340
rect 19760 13328 19766 13380
rect 20714 13368 20720 13380
rect 20675 13340 20720 13368
rect 20714 13328 20720 13340
rect 20772 13328 20778 13380
rect 10137 13303 10195 13309
rect 10137 13269 10149 13303
rect 10183 13300 10195 13303
rect 10318 13300 10324 13312
rect 10183 13272 10324 13300
rect 10183 13269 10195 13272
rect 10137 13263 10195 13269
rect 10318 13260 10324 13272
rect 10376 13260 10382 13312
rect 14090 13232 14096 13244
rect 14051 13204 14096 13232
rect 14090 13192 14096 13204
rect 14148 13192 14154 13244
rect 18966 13192 18972 13244
rect 19024 13232 19030 13244
rect 19521 13235 19579 13241
rect 19521 13232 19533 13235
rect 19024 13204 19533 13232
rect 19024 13192 19030 13204
rect 19521 13201 19533 13204
rect 19567 13201 19579 13235
rect 19521 13195 19579 13201
rect 20533 13235 20591 13241
rect 20533 13201 20545 13235
rect 20579 13201 20591 13235
rect 20533 13195 20591 13201
rect 13170 13124 13176 13176
rect 13228 13164 13234 13176
rect 14185 13167 14243 13173
rect 14185 13164 14197 13167
rect 13228 13136 14197 13164
rect 13228 13124 13234 13136
rect 14185 13133 14197 13136
rect 14231 13133 14243 13167
rect 14185 13127 14243 13133
rect 14277 13167 14335 13173
rect 14277 13133 14289 13167
rect 14323 13133 14335 13167
rect 14277 13127 14335 13133
rect 13814 13056 13820 13108
rect 13872 13096 13878 13108
rect 14292 13096 14320 13127
rect 15562 13124 15568 13176
rect 15620 13164 15626 13176
rect 20548 13164 20576 13195
rect 15620 13136 20576 13164
rect 15620 13124 15626 13136
rect 13872 13068 14320 13096
rect 13872 13056 13878 13068
rect 13725 13031 13783 13037
rect 13725 12997 13737 13031
rect 13771 13028 13783 13031
rect 14826 13028 14832 13040
rect 13771 13000 14832 13028
rect 13771 12997 13783 13000
rect 13725 12991 13783 12997
rect 14826 12988 14832 13000
rect 14884 12988 14890 13040
rect 1104 12938 21620 12960
rect 1104 12886 4414 12938
rect 4466 12886 4478 12938
rect 4530 12886 4542 12938
rect 4594 12886 4606 12938
rect 4658 12886 11278 12938
rect 11330 12886 11342 12938
rect 11394 12886 11406 12938
rect 11458 12886 11470 12938
rect 11522 12886 18142 12938
rect 18194 12886 18206 12938
rect 18258 12886 18270 12938
rect 18322 12886 18334 12938
rect 18386 12886 21620 12938
rect 1104 12864 21620 12886
rect 13170 12824 13176 12836
rect 2884 12796 11008 12824
rect 13131 12796 13176 12824
rect 842 12648 848 12700
rect 900 12688 906 12700
rect 2884 12688 2912 12796
rect 7653 12759 7711 12765
rect 7653 12725 7665 12759
rect 7699 12756 7711 12759
rect 9861 12759 9919 12765
rect 7699 12728 9076 12756
rect 7699 12725 7711 12728
rect 7653 12719 7711 12725
rect 900 12660 2912 12688
rect 900 12648 906 12660
rect 5718 12648 5724 12700
rect 5776 12688 5782 12700
rect 7101 12691 7159 12697
rect 7101 12688 7113 12691
rect 5776 12660 7113 12688
rect 5776 12648 5782 12660
rect 7101 12657 7113 12660
rect 7147 12657 7159 12691
rect 7101 12651 7159 12657
rect 7285 12691 7343 12697
rect 7285 12657 7297 12691
rect 7331 12688 7343 12691
rect 7374 12688 7380 12700
rect 7331 12660 7380 12688
rect 7331 12657 7343 12660
rect 7285 12651 7343 12657
rect 7374 12648 7380 12660
rect 7432 12648 7438 12700
rect 8202 12688 8208 12700
rect 8163 12660 8208 12688
rect 8202 12648 8208 12660
rect 8260 12648 8266 12700
rect 9048 12688 9076 12728
rect 9861 12725 9873 12759
rect 9907 12756 9919 12759
rect 10980 12756 11008 12796
rect 13170 12784 13176 12796
rect 13228 12784 13234 12836
rect 13538 12784 13544 12836
rect 13596 12824 13602 12836
rect 16482 12824 16488 12836
rect 13596 12796 16488 12824
rect 13596 12784 13602 12796
rect 16482 12784 16488 12796
rect 16540 12784 16546 12836
rect 19610 12784 19616 12836
rect 19668 12824 19674 12836
rect 19889 12827 19947 12833
rect 19889 12824 19901 12827
rect 19668 12796 19901 12824
rect 19668 12784 19674 12796
rect 19889 12793 19901 12796
rect 19935 12793 19947 12827
rect 19889 12787 19947 12793
rect 20346 12784 20352 12836
rect 20404 12824 20410 12836
rect 20441 12827 20499 12833
rect 20441 12824 20453 12827
rect 20404 12796 20453 12824
rect 20404 12784 20410 12796
rect 20441 12793 20453 12796
rect 20487 12793 20499 12827
rect 20441 12787 20499 12793
rect 14185 12759 14243 12765
rect 9907 12728 10916 12756
rect 10980 12728 13676 12756
rect 9907 12725 9919 12728
rect 9861 12719 9919 12725
rect 10321 12691 10379 12697
rect 10321 12688 10333 12691
rect 9048 12660 10333 12688
rect 10321 12657 10333 12660
rect 10367 12657 10379 12691
rect 10321 12651 10379 12657
rect 10410 12648 10416 12700
rect 10468 12688 10474 12700
rect 10468 12660 10513 12688
rect 10468 12648 10474 12660
rect 7006 12620 7012 12632
rect 6967 12592 7012 12620
rect 7006 12580 7012 12592
rect 7064 12580 7070 12632
rect 10888 12629 10916 12728
rect 11149 12691 11207 12697
rect 11149 12657 11161 12691
rect 11195 12688 11207 12691
rect 13538 12688 13544 12700
rect 11195 12660 13544 12688
rect 11195 12657 11207 12660
rect 11149 12651 11207 12657
rect 13538 12648 13544 12660
rect 13596 12648 13602 12700
rect 13648 12697 13676 12728
rect 14185 12725 14197 12759
rect 14231 12725 14243 12759
rect 14185 12719 14243 12725
rect 13633 12691 13691 12697
rect 13633 12657 13645 12691
rect 13679 12657 13691 12691
rect 13633 12651 13691 12657
rect 13722 12648 13728 12700
rect 13780 12688 13786 12700
rect 13780 12660 14136 12688
rect 13780 12648 13786 12660
rect 10873 12623 10931 12629
rect 10873 12589 10885 12623
rect 10919 12589 10931 12623
rect 10873 12583 10931 12589
rect 10962 12580 10968 12632
rect 11020 12620 11026 12632
rect 12897 12623 12955 12629
rect 12897 12620 12909 12623
rect 11020 12592 12909 12620
rect 11020 12580 11026 12592
rect 12897 12589 12909 12592
rect 12943 12589 12955 12623
rect 12897 12583 12955 12589
rect 8113 12555 8171 12561
rect 8113 12552 8125 12555
rect 6656 12524 8125 12552
rect 6656 12493 6684 12524
rect 8113 12521 8125 12524
rect 8159 12521 8171 12555
rect 13906 12552 13912 12564
rect 8113 12515 8171 12521
rect 12728 12524 13912 12552
rect 6641 12487 6699 12493
rect 6641 12453 6653 12487
rect 6687 12453 6699 12487
rect 6641 12447 6699 12453
rect 7742 12444 7748 12496
rect 7800 12484 7806 12496
rect 8021 12487 8079 12493
rect 8021 12484 8033 12487
rect 7800 12456 8033 12484
rect 7800 12444 7806 12456
rect 8021 12453 8033 12456
rect 8067 12453 8079 12487
rect 10226 12484 10232 12496
rect 10187 12456 10232 12484
rect 8021 12447 8079 12453
rect 10226 12444 10232 12456
rect 10284 12444 10290 12496
rect 12728 12493 12756 12524
rect 13906 12512 13912 12524
rect 13964 12512 13970 12564
rect 14108 12552 14136 12660
rect 14200 12620 14228 12719
rect 14366 12716 14372 12768
rect 14424 12756 14430 12768
rect 14424 12728 15700 12756
rect 14424 12716 14430 12728
rect 14734 12688 14740 12700
rect 14695 12660 14740 12688
rect 14734 12648 14740 12660
rect 14792 12648 14798 12700
rect 14826 12648 14832 12700
rect 14884 12688 14890 12700
rect 15013 12691 15071 12697
rect 15013 12688 15025 12691
rect 14884 12660 15025 12688
rect 14884 12648 14890 12660
rect 15013 12657 15025 12660
rect 15059 12657 15071 12691
rect 15562 12688 15568 12700
rect 15523 12660 15568 12688
rect 15013 12651 15071 12657
rect 15562 12648 15568 12660
rect 15620 12648 15626 12700
rect 15672 12688 15700 12728
rect 18966 12688 18972 12700
rect 15672 12660 16252 12688
rect 18927 12660 18972 12688
rect 15289 12623 15347 12629
rect 15289 12620 15301 12623
rect 14200 12592 15301 12620
rect 15289 12589 15301 12592
rect 15335 12589 15347 12623
rect 15289 12583 15347 12589
rect 16022 12580 16028 12632
rect 16080 12620 16086 12632
rect 16117 12623 16175 12629
rect 16117 12620 16129 12623
rect 16080 12592 16129 12620
rect 16080 12580 16086 12592
rect 16117 12589 16129 12592
rect 16163 12589 16175 12623
rect 16224 12620 16252 12660
rect 18966 12648 18972 12660
rect 19024 12648 19030 12700
rect 17310 12620 17316 12632
rect 16224 12592 17316 12620
rect 16117 12583 16175 12589
rect 17310 12580 17316 12592
rect 17368 12580 17374 12632
rect 18690 12620 18696 12632
rect 18651 12592 18696 12620
rect 18690 12580 18696 12592
rect 18748 12580 18754 12632
rect 19702 12620 19708 12632
rect 19663 12592 19708 12620
rect 19702 12580 19708 12592
rect 19760 12580 19766 12632
rect 20254 12620 20260 12632
rect 20215 12592 20260 12620
rect 20254 12580 20260 12592
rect 20312 12580 20318 12632
rect 16384 12555 16442 12561
rect 14108 12524 15148 12552
rect 15120 12496 15148 12524
rect 16384 12521 16396 12555
rect 16430 12552 16442 12555
rect 17678 12552 17684 12564
rect 16430 12524 17684 12552
rect 16430 12521 16442 12524
rect 16384 12515 16442 12521
rect 17678 12512 17684 12524
rect 17736 12512 17742 12564
rect 12713 12487 12771 12493
rect 12713 12453 12725 12487
rect 12759 12453 12771 12487
rect 12713 12447 12771 12453
rect 13541 12487 13599 12493
rect 13541 12453 13553 12487
rect 13587 12484 13599 12487
rect 14366 12484 14372 12496
rect 13587 12456 14372 12484
rect 13587 12453 13599 12456
rect 13541 12447 13599 12453
rect 14366 12444 14372 12456
rect 14424 12444 14430 12496
rect 14550 12484 14556 12496
rect 14511 12456 14556 12484
rect 14550 12444 14556 12456
rect 14608 12444 14614 12496
rect 14645 12487 14703 12493
rect 14645 12453 14657 12487
rect 14691 12484 14703 12487
rect 15013 12487 15071 12493
rect 15013 12484 15025 12487
rect 14691 12456 15025 12484
rect 14691 12453 14703 12456
rect 14645 12447 14703 12453
rect 15013 12453 15025 12456
rect 15059 12453 15071 12487
rect 15013 12447 15071 12453
rect 15102 12444 15108 12496
rect 15160 12484 15166 12496
rect 17497 12487 17555 12493
rect 17497 12484 17509 12487
rect 15160 12456 17509 12484
rect 15160 12444 15166 12456
rect 17497 12453 17509 12456
rect 17543 12453 17555 12487
rect 17497 12447 17555 12453
rect 1104 12394 21620 12416
rect 1104 12342 7846 12394
rect 7898 12342 7910 12394
rect 7962 12342 7974 12394
rect 8026 12342 8038 12394
rect 8090 12342 14710 12394
rect 14762 12342 14774 12394
rect 14826 12342 14838 12394
rect 14890 12342 14902 12394
rect 14954 12342 21620 12394
rect 1104 12320 21620 12342
rect 10226 12240 10232 12292
rect 10284 12280 10290 12292
rect 10413 12283 10471 12289
rect 10413 12280 10425 12283
rect 10284 12252 10425 12280
rect 10284 12240 10290 12252
rect 10413 12249 10425 12252
rect 10459 12249 10471 12283
rect 10413 12243 10471 12249
rect 10520 12252 14044 12280
rect 7650 12172 7656 12224
rect 7708 12212 7714 12224
rect 8294 12212 8300 12224
rect 7708 12184 8300 12212
rect 7708 12172 7714 12184
rect 8294 12172 8300 12184
rect 8352 12172 8358 12224
rect 9674 12172 9680 12224
rect 9732 12212 9738 12224
rect 10520 12212 10548 12252
rect 9732 12184 10548 12212
rect 10781 12215 10839 12221
rect 9732 12172 9738 12184
rect 10781 12181 10793 12215
rect 10827 12212 10839 12215
rect 11425 12215 11483 12221
rect 11425 12212 11437 12215
rect 10827 12184 11437 12212
rect 10827 12181 10839 12184
rect 10781 12175 10839 12181
rect 11425 12181 11437 12184
rect 11471 12181 11483 12215
rect 11425 12175 11483 12181
rect 12704 12215 12762 12221
rect 12704 12181 12716 12215
rect 12750 12212 12762 12215
rect 13722 12212 13728 12224
rect 12750 12184 13728 12212
rect 12750 12181 12762 12184
rect 12704 12175 12762 12181
rect 13722 12172 13728 12184
rect 13780 12172 13786 12224
rect 14016 12212 14044 12252
rect 14090 12240 14096 12292
rect 14148 12280 14154 12292
rect 14461 12283 14519 12289
rect 14461 12280 14473 12283
rect 14148 12252 14473 12280
rect 14148 12240 14154 12252
rect 14461 12249 14473 12252
rect 14507 12249 14519 12283
rect 14461 12243 14519 12249
rect 17402 12240 17408 12292
rect 17460 12280 17466 12292
rect 17770 12280 17776 12292
rect 17460 12252 17776 12280
rect 17460 12240 17466 12252
rect 17770 12240 17776 12252
rect 17828 12240 17834 12292
rect 18049 12283 18107 12289
rect 18049 12249 18061 12283
rect 18095 12280 18107 12283
rect 18690 12280 18696 12292
rect 18095 12252 18696 12280
rect 18095 12249 18107 12252
rect 18049 12243 18107 12249
rect 18690 12240 18696 12252
rect 18748 12240 18754 12292
rect 19978 12240 19984 12292
rect 20036 12280 20042 12292
rect 20165 12283 20223 12289
rect 20165 12280 20177 12283
rect 20036 12252 20177 12280
rect 20036 12240 20042 12252
rect 20165 12249 20177 12252
rect 20211 12249 20223 12283
rect 20165 12243 20223 12249
rect 20717 12283 20775 12289
rect 20717 12249 20729 12283
rect 20763 12280 20775 12283
rect 21082 12280 21088 12292
rect 20763 12252 21088 12280
rect 20763 12249 20775 12252
rect 20717 12243 20775 12249
rect 21082 12240 21088 12252
rect 21140 12240 21146 12292
rect 14829 12215 14887 12221
rect 14829 12212 14841 12215
rect 14016 12184 14841 12212
rect 14829 12181 14841 12184
rect 14875 12212 14887 12215
rect 17954 12212 17960 12224
rect 14875 12184 17960 12212
rect 14875 12181 14887 12184
rect 14829 12175 14887 12181
rect 17954 12172 17960 12184
rect 18012 12172 18018 12224
rect 18417 12215 18475 12221
rect 18417 12181 18429 12215
rect 18463 12212 18475 12215
rect 18598 12212 18604 12224
rect 18463 12184 18604 12212
rect 18463 12181 18475 12184
rect 18417 12175 18475 12181
rect 18598 12172 18604 12184
rect 18656 12172 18662 12224
rect 7092 12147 7150 12153
rect 7092 12113 7104 12147
rect 7138 12144 7150 12147
rect 7374 12144 7380 12156
rect 7138 12116 7380 12144
rect 7138 12113 7150 12116
rect 7092 12107 7150 12113
rect 7374 12104 7380 12116
rect 7432 12104 7438 12156
rect 8202 12144 8208 12156
rect 8115 12116 8208 12144
rect 8202 12104 8208 12116
rect 8260 12144 8266 12156
rect 8932 12147 8990 12153
rect 8932 12144 8944 12147
rect 8260 12116 8944 12144
rect 8260 12104 8266 12116
rect 8932 12113 8944 12116
rect 8978 12144 8990 12147
rect 10873 12147 10931 12153
rect 8978 12116 10364 12144
rect 8978 12113 8990 12116
rect 8932 12107 8990 12113
rect 6822 12076 6828 12088
rect 6783 12048 6828 12076
rect 6822 12036 6828 12048
rect 6880 12036 6886 12088
rect 8220 12017 8248 12104
rect 8294 12036 8300 12088
rect 8352 12076 8358 12088
rect 8665 12079 8723 12085
rect 8665 12076 8677 12079
rect 8352 12048 8677 12076
rect 8352 12036 8358 12048
rect 8665 12045 8677 12048
rect 8711 12045 8723 12079
rect 10336 12076 10364 12116
rect 10873 12113 10885 12147
rect 10919 12144 10931 12147
rect 15194 12144 15200 12156
rect 10919 12116 15200 12144
rect 10919 12113 10931 12116
rect 10873 12107 10931 12113
rect 15194 12104 15200 12116
rect 15252 12104 15258 12156
rect 16568 12147 16626 12153
rect 16568 12113 16580 12147
rect 16614 12144 16626 12147
rect 17034 12144 17040 12156
rect 16614 12116 17040 12144
rect 16614 12113 16626 12116
rect 16568 12107 16626 12113
rect 17034 12104 17040 12116
rect 17092 12104 17098 12156
rect 19978 12144 19984 12156
rect 19939 12116 19984 12144
rect 19978 12104 19984 12116
rect 20036 12104 20042 12156
rect 20070 12104 20076 12156
rect 20128 12144 20134 12156
rect 20533 12147 20591 12153
rect 20533 12144 20545 12147
rect 20128 12116 20545 12144
rect 20128 12104 20134 12116
rect 20533 12113 20545 12116
rect 20579 12113 20591 12147
rect 20533 12107 20591 12113
rect 10965 12079 11023 12085
rect 10965 12076 10977 12079
rect 10336 12048 10977 12076
rect 8665 12039 8723 12045
rect 10965 12045 10977 12048
rect 11011 12045 11023 12079
rect 10965 12039 11023 12045
rect 12434 12036 12440 12088
rect 12492 12076 12498 12088
rect 14921 12079 14979 12085
rect 12492 12048 12537 12076
rect 12492 12036 12498 12048
rect 14921 12045 14933 12079
rect 14967 12045 14979 12079
rect 15102 12076 15108 12088
rect 15063 12048 15108 12076
rect 14921 12039 14979 12045
rect 8205 12011 8263 12017
rect 8205 11977 8217 12011
rect 8251 11977 8263 12011
rect 8205 11971 8263 11977
rect 10045 12011 10103 12017
rect 10045 11977 10057 12011
rect 10091 12008 10103 12011
rect 10410 12008 10416 12020
rect 10091 11980 10416 12008
rect 10091 11977 10103 11980
rect 10045 11971 10103 11977
rect 10410 11968 10416 11980
rect 10468 11968 10474 12020
rect 14936 12008 14964 12039
rect 15102 12036 15108 12048
rect 15160 12036 15166 12088
rect 15838 12036 15844 12088
rect 15896 12076 15902 12088
rect 16301 12079 16359 12085
rect 16301 12076 16313 12079
rect 15896 12048 16313 12076
rect 15896 12036 15902 12048
rect 16301 12045 16313 12048
rect 16347 12045 16359 12079
rect 16301 12039 16359 12045
rect 17402 12036 17408 12088
rect 17460 12076 17466 12088
rect 18509 12079 18567 12085
rect 18509 12076 18521 12079
rect 17460 12048 18521 12076
rect 17460 12036 17466 12048
rect 18509 12045 18521 12048
rect 18555 12045 18567 12079
rect 18509 12039 18567 12045
rect 18601 12079 18659 12085
rect 18601 12045 18613 12079
rect 18647 12045 18659 12079
rect 18601 12039 18659 12045
rect 17678 12008 17684 12020
rect 13648 11980 14964 12008
rect 17591 11980 17684 12008
rect 8662 11900 8668 11952
rect 8720 11940 8726 11952
rect 13648 11940 13676 11980
rect 13814 11940 13820 11952
rect 8720 11912 13676 11940
rect 13775 11912 13820 11940
rect 8720 11900 8726 11912
rect 13814 11900 13820 11912
rect 13872 11900 13878 11952
rect 14936 11940 14964 11980
rect 17678 11968 17684 11980
rect 17736 12008 17742 12020
rect 18616 12008 18644 12039
rect 17736 11980 18644 12008
rect 17736 11968 17742 11980
rect 18690 11940 18696 11952
rect 14936 11912 18696 11940
rect 18690 11900 18696 11912
rect 18748 11900 18754 11952
rect 1104 11850 21620 11872
rect 1104 11798 4414 11850
rect 4466 11798 4478 11850
rect 4530 11798 4542 11850
rect 4594 11798 4606 11850
rect 4658 11798 11278 11850
rect 11330 11798 11342 11850
rect 11394 11798 11406 11850
rect 11458 11798 11470 11850
rect 11522 11798 18142 11850
rect 18194 11798 18206 11850
rect 18258 11798 18270 11850
rect 18322 11798 18334 11850
rect 18386 11798 21620 11850
rect 1104 11776 21620 11798
rect 7742 11696 7748 11748
rect 7800 11736 7806 11748
rect 7929 11739 7987 11745
rect 7929 11736 7941 11739
rect 7800 11708 7941 11736
rect 7800 11696 7806 11708
rect 7929 11705 7941 11708
rect 7975 11705 7987 11739
rect 7929 11699 7987 11705
rect 12434 11696 12440 11748
rect 12492 11736 12498 11748
rect 13078 11736 13084 11748
rect 12492 11708 13084 11736
rect 12492 11696 12498 11708
rect 13078 11696 13084 11708
rect 13136 11736 13142 11748
rect 13817 11739 13875 11745
rect 13817 11736 13829 11739
rect 13136 11708 13829 11736
rect 13136 11696 13142 11708
rect 13817 11705 13829 11708
rect 13863 11705 13875 11739
rect 13817 11699 13875 11705
rect 14093 11739 14151 11745
rect 14093 11705 14105 11739
rect 14139 11736 14151 11739
rect 14550 11736 14556 11748
rect 14139 11708 14556 11736
rect 14139 11705 14151 11708
rect 14093 11699 14151 11705
rect 14550 11696 14556 11708
rect 14608 11696 14614 11748
rect 18598 11736 18604 11748
rect 18559 11708 18604 11736
rect 18598 11696 18604 11708
rect 18656 11696 18662 11748
rect 20162 11696 20168 11748
rect 20220 11736 20226 11748
rect 20441 11739 20499 11745
rect 20441 11736 20453 11739
rect 20220 11708 20453 11736
rect 20220 11696 20226 11708
rect 20441 11705 20453 11708
rect 20487 11705 20499 11739
rect 20441 11699 20499 11705
rect 11054 11628 11060 11680
rect 11112 11668 11118 11680
rect 11112 11640 14780 11668
rect 11112 11628 11118 11640
rect 7374 11560 7380 11612
rect 7432 11600 7438 11612
rect 8202 11600 8208 11612
rect 7432 11572 8208 11600
rect 7432 11560 7438 11572
rect 8202 11560 8208 11572
rect 8260 11600 8266 11612
rect 8481 11603 8539 11609
rect 8481 11600 8493 11603
rect 8260 11572 8493 11600
rect 8260 11560 8266 11572
rect 8481 11569 8493 11572
rect 8527 11569 8539 11603
rect 8481 11563 8539 11569
rect 13814 11560 13820 11612
rect 13872 11600 13878 11612
rect 14645 11603 14703 11609
rect 14645 11600 14657 11603
rect 13872 11572 14657 11600
rect 13872 11560 13878 11572
rect 14645 11569 14657 11572
rect 14691 11569 14703 11603
rect 14752 11600 14780 11640
rect 16298 11628 16304 11680
rect 16356 11668 16362 11680
rect 16356 11640 16712 11668
rect 16356 11628 16362 11640
rect 16684 11609 16712 11640
rect 16577 11603 16635 11609
rect 16577 11600 16589 11603
rect 14752 11572 16589 11600
rect 14645 11563 14703 11569
rect 16577 11569 16589 11572
rect 16623 11569 16635 11603
rect 16577 11563 16635 11569
rect 16669 11603 16727 11609
rect 16669 11569 16681 11603
rect 16715 11569 16727 11603
rect 16669 11563 16727 11569
rect 17034 11560 17040 11612
rect 17092 11600 17098 11612
rect 19153 11603 19211 11609
rect 19153 11600 19165 11603
rect 17092 11572 19165 11600
rect 17092 11560 17098 11572
rect 19153 11569 19165 11572
rect 19199 11569 19211 11603
rect 19153 11563 19211 11569
rect 8389 11535 8447 11541
rect 8389 11501 8401 11535
rect 8435 11532 8447 11535
rect 8662 11532 8668 11544
rect 8435 11504 8668 11532
rect 8435 11501 8447 11504
rect 8389 11495 8447 11501
rect 8662 11492 8668 11504
rect 8720 11492 8726 11544
rect 11054 11532 11060 11544
rect 11015 11504 11060 11532
rect 11054 11492 11060 11504
rect 11112 11492 11118 11544
rect 13906 11492 13912 11544
rect 13964 11532 13970 11544
rect 14001 11535 14059 11541
rect 14001 11532 14013 11535
rect 13964 11504 14013 11532
rect 13964 11492 13970 11504
rect 14001 11501 14013 11504
rect 14047 11501 14059 11535
rect 20070 11532 20076 11544
rect 14001 11495 14059 11501
rect 14384 11504 20076 11532
rect 8297 11467 8355 11473
rect 8297 11433 8309 11467
rect 8343 11464 8355 11467
rect 9674 11464 9680 11476
rect 8343 11436 9680 11464
rect 8343 11433 8355 11436
rect 8297 11427 8355 11433
rect 9674 11424 9680 11436
rect 9732 11424 9738 11476
rect 11333 11467 11391 11473
rect 11333 11433 11345 11467
rect 11379 11464 11391 11467
rect 14384 11464 14412 11504
rect 20070 11492 20076 11504
rect 20128 11492 20134 11544
rect 20254 11532 20260 11544
rect 20215 11504 20260 11532
rect 20254 11492 20260 11504
rect 20312 11492 20318 11544
rect 11379 11436 14412 11464
rect 14461 11467 14519 11473
rect 11379 11433 11391 11436
rect 11333 11427 11391 11433
rect 14461 11433 14473 11467
rect 14507 11464 14519 11467
rect 15289 11467 15347 11473
rect 15289 11464 15301 11467
rect 14507 11436 15301 11464
rect 14507 11433 14519 11436
rect 14461 11427 14519 11433
rect 15289 11433 15301 11436
rect 15335 11433 15347 11467
rect 15289 11427 15347 11433
rect 16022 11424 16028 11476
rect 16080 11464 16086 11476
rect 16390 11464 16396 11476
rect 16080 11436 16396 11464
rect 16080 11424 16086 11436
rect 16390 11424 16396 11436
rect 16448 11464 16454 11476
rect 16485 11467 16543 11473
rect 16485 11464 16497 11467
rect 16448 11436 16497 11464
rect 16448 11424 16454 11436
rect 16485 11433 16497 11436
rect 16531 11433 16543 11467
rect 16485 11427 16543 11433
rect 18969 11467 19027 11473
rect 18969 11433 18981 11467
rect 19015 11464 19027 11467
rect 19613 11467 19671 11473
rect 19613 11464 19625 11467
rect 19015 11436 19625 11464
rect 19015 11433 19027 11436
rect 18969 11427 19027 11433
rect 19613 11433 19625 11436
rect 19659 11433 19671 11467
rect 19613 11427 19671 11433
rect 14550 11396 14556 11408
rect 14463 11368 14556 11396
rect 14550 11356 14556 11368
rect 14608 11396 14614 11408
rect 15194 11396 15200 11408
rect 14608 11368 15200 11396
rect 14608 11356 14614 11368
rect 15194 11356 15200 11368
rect 15252 11356 15258 11408
rect 16114 11396 16120 11408
rect 16075 11368 16120 11396
rect 16114 11356 16120 11368
rect 16172 11356 16178 11408
rect 19061 11399 19119 11405
rect 19061 11365 19073 11399
rect 19107 11396 19119 11399
rect 19150 11396 19156 11408
rect 19107 11368 19156 11396
rect 19107 11365 19119 11368
rect 19061 11359 19119 11365
rect 19150 11356 19156 11368
rect 19208 11356 19214 11408
rect 1104 11306 21620 11328
rect 1104 11254 7846 11306
rect 7898 11254 7910 11306
rect 7962 11254 7974 11306
rect 8026 11254 8038 11306
rect 8090 11254 14710 11306
rect 14762 11254 14774 11306
rect 14826 11254 14838 11306
rect 14890 11254 14902 11306
rect 14954 11254 21620 11306
rect 1104 11232 21620 11254
rect 16114 11152 16120 11204
rect 16172 11192 16178 11204
rect 16853 11195 16911 11201
rect 16853 11192 16865 11195
rect 16172 11164 16865 11192
rect 16172 11152 16178 11164
rect 16853 11161 16865 11164
rect 16899 11161 16911 11195
rect 19150 11192 19156 11204
rect 19111 11164 19156 11192
rect 16853 11155 16911 11161
rect 19150 11152 19156 11164
rect 19208 11152 19214 11204
rect 20622 11152 20628 11204
rect 20680 11192 20686 11204
rect 20717 11195 20775 11201
rect 20717 11192 20729 11195
rect 20680 11164 20729 11192
rect 20680 11152 20686 11164
rect 20717 11161 20729 11164
rect 20763 11161 20775 11195
rect 20717 11155 20775 11161
rect 8573 11059 8631 11065
rect 8573 11025 8585 11059
rect 8619 11056 8631 11059
rect 9030 11056 9036 11068
rect 8619 11028 9036 11056
rect 8619 11025 8631 11028
rect 8573 11019 8631 11025
rect 9030 11016 9036 11028
rect 9088 11016 9094 11068
rect 16758 11056 16764 11068
rect 16719 11028 16764 11056
rect 16758 11016 16764 11028
rect 16816 11016 16822 11068
rect 17770 11016 17776 11068
rect 17828 11056 17834 11068
rect 19521 11059 19579 11065
rect 19521 11056 19533 11059
rect 17828 11028 19533 11056
rect 17828 11016 17834 11028
rect 19521 11025 19533 11028
rect 19567 11025 19579 11059
rect 20530 11056 20536 11068
rect 20491 11028 20536 11056
rect 19521 11019 19579 11025
rect 20530 11016 20536 11028
rect 20588 11016 20594 11068
rect 17034 10988 17040 11000
rect 16995 10960 17040 10988
rect 17034 10948 17040 10960
rect 17092 10948 17098 11000
rect 17218 10948 17224 11000
rect 17276 10988 17282 11000
rect 17862 10988 17868 11000
rect 17276 10960 17868 10988
rect 17276 10948 17282 10960
rect 17862 10948 17868 10960
rect 17920 10988 17926 11000
rect 19613 10991 19671 10997
rect 19613 10988 19625 10991
rect 17920 10960 19625 10988
rect 17920 10948 17926 10960
rect 19613 10957 19625 10960
rect 19659 10957 19671 10991
rect 19794 10988 19800 11000
rect 19755 10960 19800 10988
rect 19613 10951 19671 10957
rect 19794 10948 19800 10960
rect 19852 10948 19858 11000
rect 8294 10880 8300 10932
rect 8352 10920 8358 10932
rect 8389 10923 8447 10929
rect 8389 10920 8401 10923
rect 8352 10892 8401 10920
rect 8352 10880 8358 10892
rect 8389 10889 8401 10892
rect 8435 10889 8447 10923
rect 8389 10883 8447 10889
rect 16393 10923 16451 10929
rect 16393 10889 16405 10923
rect 16439 10920 16451 10923
rect 17402 10920 17408 10932
rect 16439 10892 17408 10920
rect 16439 10889 16451 10892
rect 16393 10883 16451 10889
rect 17402 10880 17408 10892
rect 17460 10880 17466 10932
rect 1104 10762 21620 10784
rect 1104 10710 4414 10762
rect 4466 10710 4478 10762
rect 4530 10710 4542 10762
rect 4594 10710 4606 10762
rect 4658 10710 11278 10762
rect 11330 10710 11342 10762
rect 11394 10710 11406 10762
rect 11458 10710 11470 10762
rect 11522 10710 18142 10762
rect 18194 10710 18206 10762
rect 18258 10710 18270 10762
rect 18322 10710 18334 10762
rect 18386 10710 21620 10762
rect 1104 10688 21620 10710
rect 1670 10608 1676 10660
rect 1728 10648 1734 10660
rect 8021 10651 8079 10657
rect 1728 10620 7604 10648
rect 1728 10608 1734 10620
rect 7576 10580 7604 10620
rect 8021 10617 8033 10651
rect 8067 10648 8079 10651
rect 8202 10648 8208 10660
rect 8067 10620 8208 10648
rect 8067 10617 8079 10620
rect 8021 10611 8079 10617
rect 8202 10608 8208 10620
rect 8260 10608 8266 10660
rect 10321 10651 10379 10657
rect 10321 10617 10333 10651
rect 10367 10648 10379 10651
rect 11054 10648 11060 10660
rect 10367 10620 11060 10648
rect 10367 10617 10379 10620
rect 10321 10611 10379 10617
rect 11054 10608 11060 10620
rect 11112 10608 11118 10660
rect 14458 10648 14464 10660
rect 14419 10620 14464 10648
rect 14458 10608 14464 10620
rect 14516 10608 14522 10660
rect 16485 10651 16543 10657
rect 16485 10617 16497 10651
rect 16531 10648 16543 10651
rect 16758 10648 16764 10660
rect 16531 10620 16764 10648
rect 16531 10617 16543 10620
rect 16485 10611 16543 10617
rect 16758 10608 16764 10620
rect 16816 10608 16822 10660
rect 18506 10648 18512 10660
rect 18467 10620 18512 10648
rect 18506 10608 18512 10620
rect 18564 10608 18570 10660
rect 19610 10608 19616 10660
rect 19668 10648 19674 10660
rect 20441 10651 20499 10657
rect 20441 10648 20453 10651
rect 19668 10620 20453 10648
rect 19668 10608 19674 10620
rect 20441 10617 20453 10620
rect 20487 10617 20499 10651
rect 20441 10611 20499 10617
rect 7576 10552 11836 10580
rect 11808 10521 11836 10552
rect 10873 10515 10931 10521
rect 10873 10481 10885 10515
rect 10919 10481 10931 10515
rect 10873 10475 10931 10481
rect 11793 10515 11851 10521
rect 11793 10481 11805 10515
rect 11839 10481 11851 10515
rect 11974 10512 11980 10524
rect 11935 10484 11980 10512
rect 11793 10475 11851 10481
rect 6641 10447 6699 10453
rect 6641 10413 6653 10447
rect 6687 10413 6699 10447
rect 6641 10407 6699 10413
rect 6908 10447 6966 10453
rect 6908 10413 6920 10447
rect 6954 10444 6966 10447
rect 10888 10444 10916 10475
rect 11974 10472 11980 10484
rect 12032 10472 12038 10524
rect 13078 10512 13084 10524
rect 13039 10484 13084 10512
rect 13078 10472 13084 10484
rect 13136 10472 13142 10524
rect 17129 10515 17187 10521
rect 17129 10481 17141 10515
rect 17175 10481 17187 10515
rect 17129 10475 17187 10481
rect 19153 10515 19211 10521
rect 19153 10481 19165 10515
rect 19199 10512 19211 10515
rect 19334 10512 19340 10524
rect 19199 10484 19340 10512
rect 19199 10481 19211 10484
rect 19153 10475 19211 10481
rect 11238 10444 11244 10456
rect 6954 10416 11244 10444
rect 6954 10413 6966 10416
rect 6908 10407 6966 10413
rect 6656 10376 6684 10407
rect 11238 10404 11244 10416
rect 11296 10404 11302 10456
rect 13348 10447 13406 10453
rect 13348 10413 13360 10447
rect 13394 10444 13406 10447
rect 13814 10444 13820 10456
rect 13394 10416 13820 10444
rect 13394 10413 13406 10416
rect 13348 10407 13406 10413
rect 13814 10404 13820 10416
rect 13872 10404 13878 10456
rect 16298 10404 16304 10456
rect 16356 10444 16362 10456
rect 17144 10444 17172 10475
rect 19334 10472 19340 10484
rect 19392 10472 19398 10524
rect 19794 10444 19800 10456
rect 16356 10416 19800 10444
rect 16356 10404 16362 10416
rect 19794 10404 19800 10416
rect 19852 10404 19858 10456
rect 20254 10444 20260 10456
rect 20215 10416 20260 10444
rect 20254 10404 20260 10416
rect 20312 10404 20318 10456
rect 6822 10376 6828 10388
rect 6656 10348 6828 10376
rect 6822 10336 6828 10348
rect 6880 10376 6886 10388
rect 8202 10376 8208 10388
rect 6880 10348 8208 10376
rect 6880 10336 6886 10348
rect 8202 10336 8208 10348
rect 8260 10336 8266 10388
rect 11701 10379 11759 10385
rect 11701 10345 11713 10379
rect 11747 10376 11759 10379
rect 16022 10376 16028 10388
rect 11747 10348 16028 10376
rect 11747 10345 11759 10348
rect 11701 10339 11759 10345
rect 16022 10336 16028 10348
rect 16080 10336 16086 10388
rect 16850 10376 16856 10388
rect 16811 10348 16856 10376
rect 16850 10336 16856 10348
rect 16908 10336 16914 10388
rect 10686 10308 10692 10320
rect 10647 10280 10692 10308
rect 10686 10268 10692 10280
rect 10744 10268 10750 10320
rect 10781 10311 10839 10317
rect 10781 10277 10793 10311
rect 10827 10308 10839 10311
rect 11146 10308 11152 10320
rect 10827 10280 11152 10308
rect 10827 10277 10839 10280
rect 10781 10271 10839 10277
rect 11146 10268 11152 10280
rect 11204 10268 11210 10320
rect 11330 10308 11336 10320
rect 11291 10280 11336 10308
rect 11330 10268 11336 10280
rect 11388 10268 11394 10320
rect 16942 10308 16948 10320
rect 16903 10280 16948 10308
rect 16942 10268 16948 10280
rect 17000 10268 17006 10320
rect 18230 10268 18236 10320
rect 18288 10308 18294 10320
rect 18877 10311 18935 10317
rect 18877 10308 18889 10311
rect 18288 10280 18889 10308
rect 18288 10268 18294 10280
rect 18877 10277 18889 10280
rect 18923 10277 18935 10311
rect 18877 10271 18935 10277
rect 18966 10268 18972 10320
rect 19024 10308 19030 10320
rect 19024 10280 19069 10308
rect 19024 10268 19030 10280
rect 1104 10218 21620 10240
rect 1104 10166 7846 10218
rect 7898 10166 7910 10218
rect 7962 10166 7974 10218
rect 8026 10166 8038 10218
rect 8090 10166 14710 10218
rect 14762 10166 14774 10218
rect 14826 10166 14838 10218
rect 14890 10166 14902 10218
rect 14954 10166 21620 10218
rect 1104 10144 21620 10166
rect 11238 10104 11244 10116
rect 11199 10076 11244 10104
rect 11238 10064 11244 10076
rect 11296 10064 11302 10116
rect 11330 10064 11336 10116
rect 11388 10104 11394 10116
rect 12897 10107 12955 10113
rect 12897 10104 12909 10107
rect 11388 10076 12909 10104
rect 11388 10064 11394 10076
rect 12897 10073 12909 10076
rect 12943 10073 12955 10107
rect 12897 10067 12955 10073
rect 15105 10107 15163 10113
rect 15105 10073 15117 10107
rect 15151 10073 15163 10107
rect 15105 10067 15163 10073
rect 8472 10039 8530 10045
rect 8472 10005 8484 10039
rect 8518 10036 8530 10039
rect 11790 10036 11796 10048
rect 8518 10008 11796 10036
rect 8518 10005 8530 10008
rect 8472 9999 8530 10005
rect 11790 9996 11796 10008
rect 11848 10036 11854 10048
rect 11974 10036 11980 10048
rect 11848 10008 11980 10036
rect 11848 9996 11854 10008
rect 11974 9996 11980 10008
rect 12032 10036 12038 10048
rect 15120 10036 15148 10067
rect 17034 10064 17040 10116
rect 17092 10104 17098 10116
rect 17405 10107 17463 10113
rect 17405 10104 17417 10107
rect 17092 10076 17417 10104
rect 17092 10064 17098 10076
rect 17405 10073 17417 10076
rect 17451 10073 17463 10107
rect 18230 10104 18236 10116
rect 18191 10076 18236 10104
rect 17405 10067 17463 10073
rect 18230 10064 18236 10076
rect 18288 10064 18294 10116
rect 19794 10064 19800 10116
rect 19852 10104 19858 10116
rect 20073 10107 20131 10113
rect 20073 10104 20085 10107
rect 19852 10076 20085 10104
rect 19852 10064 19858 10076
rect 20073 10073 20085 10076
rect 20119 10073 20131 10107
rect 20073 10067 20131 10073
rect 20717 10107 20775 10113
rect 20717 10073 20729 10107
rect 20763 10104 20775 10107
rect 21174 10104 21180 10116
rect 20763 10076 21180 10104
rect 20763 10073 20775 10076
rect 20717 10067 20775 10073
rect 21174 10064 21180 10076
rect 21232 10064 21238 10116
rect 16298 10045 16304 10048
rect 16292 10036 16304 10045
rect 12032 10008 15148 10036
rect 16259 10008 16304 10036
rect 12032 9996 12038 10008
rect 16292 9999 16304 10008
rect 16298 9996 16304 9999
rect 16356 9996 16362 10048
rect 10128 9971 10186 9977
rect 10128 9968 10140 9971
rect 9600 9940 10140 9968
rect 8202 9900 8208 9912
rect 8163 9872 8208 9900
rect 8202 9860 8208 9872
rect 8260 9860 8266 9912
rect 9600 9841 9628 9940
rect 10128 9937 10140 9940
rect 10174 9968 10186 9971
rect 12802 9968 12808 9980
rect 10174 9940 11744 9968
rect 12763 9940 12808 9968
rect 10174 9937 10186 9940
rect 10128 9931 10186 9937
rect 11716 9912 11744 9940
rect 12802 9928 12808 9940
rect 12860 9928 12866 9980
rect 13078 9928 13084 9980
rect 13136 9968 13142 9980
rect 13725 9971 13783 9977
rect 13725 9968 13737 9971
rect 13136 9940 13737 9968
rect 13136 9928 13142 9940
rect 13725 9937 13737 9940
rect 13771 9937 13783 9971
rect 13725 9931 13783 9937
rect 13992 9971 14050 9977
rect 13992 9937 14004 9971
rect 14038 9968 14050 9971
rect 14458 9968 14464 9980
rect 14038 9940 14464 9968
rect 14038 9937 14050 9940
rect 13992 9931 14050 9937
rect 9861 9903 9919 9909
rect 9861 9900 9873 9903
rect 9692 9872 9873 9900
rect 9585 9835 9643 9841
rect 9585 9801 9597 9835
rect 9631 9801 9643 9835
rect 9585 9795 9643 9801
rect 8202 9724 8208 9776
rect 8260 9764 8266 9776
rect 9692 9764 9720 9872
rect 9861 9869 9873 9872
rect 9907 9869 9919 9903
rect 9861 9863 9919 9869
rect 11517 9903 11575 9909
rect 11517 9869 11529 9903
rect 11563 9900 11575 9903
rect 11606 9900 11612 9912
rect 11563 9872 11612 9900
rect 11563 9869 11575 9872
rect 11517 9863 11575 9869
rect 11606 9860 11612 9872
rect 11664 9860 11670 9912
rect 11698 9860 11704 9912
rect 11756 9900 11762 9912
rect 12989 9903 13047 9909
rect 11756 9872 12756 9900
rect 11756 9860 11762 9872
rect 11146 9792 11152 9844
rect 11204 9832 11210 9844
rect 12437 9835 12495 9841
rect 12437 9832 12449 9835
rect 11204 9804 12449 9832
rect 11204 9792 11210 9804
rect 12437 9801 12449 9804
rect 12483 9801 12495 9835
rect 12728 9832 12756 9872
rect 12989 9869 13001 9903
rect 13035 9869 13047 9903
rect 12989 9863 13047 9869
rect 13004 9832 13032 9863
rect 12728 9804 13032 9832
rect 12437 9795 12495 9801
rect 8260 9736 9720 9764
rect 13740 9764 13768 9931
rect 14458 9928 14464 9940
rect 14516 9928 14522 9980
rect 18693 9971 18751 9977
rect 18693 9968 18705 9971
rect 16040 9940 18705 9968
rect 15838 9900 15844 9912
rect 15212 9872 15844 9900
rect 14090 9764 14096 9776
rect 13740 9736 14096 9764
rect 8260 9724 8266 9736
rect 14090 9724 14096 9736
rect 14148 9764 14154 9776
rect 15212 9764 15240 9872
rect 15838 9860 15844 9872
rect 15896 9900 15902 9912
rect 16040 9909 16068 9940
rect 18693 9937 18705 9940
rect 18739 9937 18751 9971
rect 18693 9931 18751 9937
rect 18960 9971 19018 9977
rect 18960 9937 18972 9971
rect 19006 9968 19018 9971
rect 19334 9968 19340 9980
rect 19006 9940 19340 9968
rect 19006 9937 19018 9940
rect 18960 9931 19018 9937
rect 19334 9928 19340 9940
rect 19392 9928 19398 9980
rect 20530 9968 20536 9980
rect 20491 9940 20536 9968
rect 20530 9928 20536 9940
rect 20588 9928 20594 9980
rect 16025 9903 16083 9909
rect 16025 9900 16037 9903
rect 15896 9872 16037 9900
rect 15896 9860 15902 9872
rect 16025 9869 16037 9872
rect 16071 9869 16083 9903
rect 16025 9863 16083 9869
rect 14148 9736 15240 9764
rect 14148 9724 14154 9736
rect 1104 9674 21620 9696
rect 1104 9622 4414 9674
rect 4466 9622 4478 9674
rect 4530 9622 4542 9674
rect 4594 9622 4606 9674
rect 4658 9622 11278 9674
rect 11330 9622 11342 9674
rect 11394 9622 11406 9674
rect 11458 9622 11470 9674
rect 11522 9622 18142 9674
rect 18194 9622 18206 9674
rect 18258 9622 18270 9674
rect 18322 9622 18334 9674
rect 18386 9622 21620 9674
rect 1104 9600 21620 9622
rect 18417 9563 18475 9569
rect 18417 9529 18429 9563
rect 18463 9560 18475 9563
rect 18966 9560 18972 9572
rect 18463 9532 18972 9560
rect 18463 9529 18475 9532
rect 18417 9523 18475 9529
rect 18966 9520 18972 9532
rect 19024 9520 19030 9572
rect 11149 9495 11207 9501
rect 11149 9461 11161 9495
rect 11195 9492 11207 9495
rect 12802 9492 12808 9504
rect 11195 9464 12808 9492
rect 11195 9461 11207 9464
rect 11149 9455 11207 9461
rect 12802 9452 12808 9464
rect 12860 9452 12866 9504
rect 13630 9452 13636 9504
rect 13688 9492 13694 9504
rect 13725 9495 13783 9501
rect 13725 9492 13737 9495
rect 13688 9464 13737 9492
rect 13688 9452 13694 9464
rect 13725 9461 13737 9464
rect 13771 9461 13783 9495
rect 13725 9455 13783 9461
rect 15010 9452 15016 9504
rect 15068 9492 15074 9504
rect 15473 9495 15531 9501
rect 15473 9492 15485 9495
rect 15068 9464 15485 9492
rect 15068 9452 15074 9464
rect 15473 9461 15485 9464
rect 15519 9461 15531 9495
rect 15473 9455 15531 9461
rect 20346 9452 20352 9504
rect 20404 9492 20410 9504
rect 20441 9495 20499 9501
rect 20441 9492 20453 9495
rect 20404 9464 20453 9492
rect 20404 9452 20410 9464
rect 20441 9461 20453 9464
rect 20487 9461 20499 9495
rect 20441 9455 20499 9461
rect 11790 9424 11796 9436
rect 11751 9396 11796 9424
rect 11790 9384 11796 9396
rect 11848 9424 11854 9436
rect 13081 9427 13139 9433
rect 13081 9424 13093 9427
rect 11848 9396 13093 9424
rect 11848 9384 11854 9396
rect 13081 9393 13093 9396
rect 13127 9393 13139 9427
rect 17770 9424 17776 9436
rect 13081 9387 13139 9393
rect 13372 9396 17776 9424
rect 11609 9359 11667 9365
rect 11609 9325 11621 9359
rect 11655 9356 11667 9359
rect 12066 9356 12072 9368
rect 11655 9328 12072 9356
rect 11655 9325 11667 9328
rect 11609 9319 11667 9325
rect 12066 9316 12072 9328
rect 12124 9316 12130 9368
rect 12897 9359 12955 9365
rect 12897 9325 12909 9359
rect 12943 9356 12955 9359
rect 13372 9356 13400 9396
rect 17770 9384 17776 9396
rect 17828 9384 17834 9436
rect 19061 9427 19119 9433
rect 19061 9393 19073 9427
rect 19107 9424 19119 9427
rect 19426 9424 19432 9436
rect 19107 9396 19432 9424
rect 19107 9393 19119 9396
rect 19061 9387 19119 9393
rect 19426 9384 19432 9396
rect 19484 9384 19490 9436
rect 12943 9328 13400 9356
rect 12943 9325 12955 9328
rect 12897 9319 12955 9325
rect 13446 9316 13452 9368
rect 13504 9356 13510 9368
rect 13541 9359 13599 9365
rect 13541 9356 13553 9359
rect 13504 9328 13553 9356
rect 13504 9316 13510 9328
rect 13541 9325 13553 9328
rect 13587 9325 13599 9359
rect 13541 9319 13599 9325
rect 15289 9359 15347 9365
rect 15289 9325 15301 9359
rect 15335 9356 15347 9359
rect 15562 9356 15568 9368
rect 15335 9328 15568 9356
rect 15335 9325 15347 9328
rect 15289 9319 15347 9325
rect 15562 9316 15568 9328
rect 15620 9316 15626 9368
rect 18782 9356 18788 9368
rect 18743 9328 18788 9356
rect 18782 9316 18788 9328
rect 18840 9316 18846 9368
rect 20254 9356 20260 9368
rect 20215 9328 20260 9356
rect 20254 9316 20260 9328
rect 20312 9316 20318 9368
rect 11517 9291 11575 9297
rect 11517 9257 11529 9291
rect 11563 9288 11575 9291
rect 11882 9288 11888 9300
rect 11563 9260 11888 9288
rect 11563 9257 11575 9260
rect 11517 9251 11575 9257
rect 11882 9248 11888 9260
rect 11940 9288 11946 9300
rect 16850 9288 16856 9300
rect 11940 9260 16856 9288
rect 11940 9248 11946 9260
rect 16850 9248 16856 9260
rect 16908 9248 16914 9300
rect 16942 9248 16948 9300
rect 17000 9288 17006 9300
rect 19058 9288 19064 9300
rect 17000 9260 19064 9288
rect 17000 9248 17006 9260
rect 19058 9248 19064 9260
rect 19116 9248 19122 9300
rect 12526 9220 12532 9232
rect 12487 9192 12532 9220
rect 12526 9180 12532 9192
rect 12584 9180 12590 9232
rect 12989 9223 13047 9229
rect 12989 9189 13001 9223
rect 13035 9220 13047 9223
rect 17862 9220 17868 9232
rect 13035 9192 17868 9220
rect 13035 9189 13047 9192
rect 12989 9183 13047 9189
rect 17862 9180 17868 9192
rect 17920 9180 17926 9232
rect 18874 9220 18880 9232
rect 18835 9192 18880 9220
rect 18874 9180 18880 9192
rect 18932 9180 18938 9232
rect 1104 9130 21620 9152
rect 1104 9078 7846 9130
rect 7898 9078 7910 9130
rect 7962 9078 7974 9130
rect 8026 9078 8038 9130
rect 8090 9078 14710 9130
rect 14762 9078 14774 9130
rect 14826 9078 14838 9130
rect 14890 9078 14902 9130
rect 14954 9078 21620 9130
rect 1104 9056 21620 9078
rect 10686 8976 10692 9028
rect 10744 9016 10750 9028
rect 10965 9019 11023 9025
rect 10965 9016 10977 9019
rect 10744 8988 10977 9016
rect 10744 8976 10750 8988
rect 10965 8985 10977 8988
rect 11011 8985 11023 9019
rect 10965 8979 11023 8985
rect 11333 9019 11391 9025
rect 11333 8985 11345 9019
rect 11379 9016 11391 9019
rect 11606 9016 11612 9028
rect 11379 8988 11612 9016
rect 11379 8985 11391 8988
rect 11333 8979 11391 8985
rect 11606 8976 11612 8988
rect 11664 8976 11670 9028
rect 12066 8976 12072 9028
rect 12124 9016 12130 9028
rect 12124 8988 16160 9016
rect 12124 8976 12130 8988
rect 11425 8951 11483 8957
rect 11425 8917 11437 8951
rect 11471 8948 11483 8951
rect 12526 8948 12532 8960
rect 11471 8920 12532 8948
rect 11471 8917 11483 8920
rect 11425 8911 11483 8917
rect 12526 8908 12532 8920
rect 12584 8908 12590 8960
rect 15562 8948 15568 8960
rect 15523 8920 15568 8948
rect 15562 8908 15568 8920
rect 15620 8908 15626 8960
rect 16132 8948 16160 8988
rect 16206 8976 16212 9028
rect 16264 9016 16270 9028
rect 20717 9019 20775 9025
rect 20717 9016 20729 9019
rect 16264 8988 20729 9016
rect 16264 8976 16270 8988
rect 20717 8985 20729 8988
rect 20763 8985 20775 9019
rect 20717 8979 20775 8985
rect 16132 8920 16252 8948
rect 15289 8883 15347 8889
rect 15289 8849 15301 8883
rect 15335 8880 15347 8883
rect 16114 8880 16120 8892
rect 15335 8852 16120 8880
rect 15335 8849 15347 8852
rect 15289 8843 15347 8849
rect 16114 8840 16120 8852
rect 16172 8840 16178 8892
rect 16224 8880 16252 8920
rect 16850 8908 16856 8960
rect 16908 8948 16914 8960
rect 18782 8948 18788 8960
rect 16908 8920 18788 8948
rect 16908 8908 16914 8920
rect 18782 8908 18788 8920
rect 18840 8908 18846 8960
rect 16942 8880 16948 8892
rect 16224 8852 16948 8880
rect 16942 8840 16948 8852
rect 17000 8840 17006 8892
rect 20530 8880 20536 8892
rect 20491 8852 20536 8880
rect 20530 8840 20536 8852
rect 20588 8840 20594 8892
rect 11609 8815 11667 8821
rect 11609 8781 11621 8815
rect 11655 8812 11667 8815
rect 11698 8812 11704 8824
rect 11655 8784 11704 8812
rect 11655 8781 11667 8784
rect 11609 8775 11667 8781
rect 11698 8772 11704 8784
rect 11756 8772 11762 8824
rect 1104 8586 21620 8608
rect 1104 8534 4414 8586
rect 4466 8534 4478 8586
rect 4530 8534 4542 8586
rect 4594 8534 4606 8586
rect 4658 8534 11278 8586
rect 11330 8534 11342 8586
rect 11394 8534 11406 8586
rect 11458 8534 11470 8586
rect 11522 8534 18142 8586
rect 18194 8534 18206 8586
rect 18258 8534 18270 8586
rect 18322 8534 18334 8586
rect 18386 8534 21620 8586
rect 1104 8512 21620 8534
rect 11054 8432 11060 8484
rect 11112 8472 11118 8484
rect 11425 8475 11483 8481
rect 11425 8472 11437 8475
rect 11112 8444 11437 8472
rect 11112 8432 11118 8444
rect 11425 8441 11437 8444
rect 11471 8441 11483 8475
rect 16114 8472 16120 8484
rect 16075 8444 16120 8472
rect 11425 8435 11483 8441
rect 16114 8432 16120 8444
rect 16172 8432 16178 8484
rect 19334 8432 19340 8484
rect 19392 8472 19398 8484
rect 19613 8475 19671 8481
rect 19613 8472 19625 8475
rect 19392 8444 19625 8472
rect 19392 8432 19398 8444
rect 19613 8441 19625 8444
rect 19659 8441 19671 8475
rect 19613 8435 19671 8441
rect 19518 8364 19524 8416
rect 19576 8404 19582 8416
rect 20441 8407 20499 8413
rect 20441 8404 20453 8407
rect 19576 8376 20453 8404
rect 19576 8364 19582 8376
rect 20441 8373 20453 8376
rect 20487 8373 20499 8407
rect 20441 8367 20499 8373
rect 13446 8336 13452 8348
rect 13407 8308 13452 8336
rect 13446 8296 13452 8308
rect 13504 8296 13510 8348
rect 16761 8339 16819 8345
rect 16761 8305 16773 8339
rect 16807 8336 16819 8339
rect 17218 8336 17224 8348
rect 16807 8308 17224 8336
rect 16807 8305 16819 8308
rect 16761 8299 16819 8305
rect 17218 8296 17224 8308
rect 17276 8296 17282 8348
rect 11238 8268 11244 8280
rect 11199 8240 11244 8268
rect 11238 8228 11244 8240
rect 11296 8228 11302 8280
rect 13170 8268 13176 8280
rect 13131 8240 13176 8268
rect 13170 8228 13176 8240
rect 13228 8228 13234 8280
rect 18046 8228 18052 8280
rect 18104 8268 18110 8280
rect 18233 8271 18291 8277
rect 18233 8268 18245 8271
rect 18104 8240 18245 8268
rect 18104 8228 18110 8240
rect 18233 8237 18245 8240
rect 18279 8237 18291 8271
rect 20254 8268 20260 8280
rect 20215 8240 20260 8268
rect 18233 8231 18291 8237
rect 20254 8228 20260 8240
rect 20312 8228 20318 8280
rect 16485 8203 16543 8209
rect 16485 8169 16497 8203
rect 16531 8200 16543 8203
rect 17129 8203 17187 8209
rect 17129 8200 17141 8203
rect 16531 8172 17141 8200
rect 16531 8169 16543 8172
rect 16485 8163 16543 8169
rect 17129 8169 17141 8172
rect 17175 8169 17187 8203
rect 17129 8163 17187 8169
rect 18500 8203 18558 8209
rect 18500 8169 18512 8203
rect 18546 8200 18558 8203
rect 19426 8200 19432 8212
rect 18546 8172 19432 8200
rect 18546 8169 18558 8172
rect 18500 8163 18558 8169
rect 19426 8160 19432 8172
rect 19484 8160 19490 8212
rect 13906 8132 13912 8144
rect 13867 8104 13912 8132
rect 13906 8092 13912 8104
rect 13964 8092 13970 8144
rect 16574 8092 16580 8144
rect 16632 8132 16638 8144
rect 16632 8104 16677 8132
rect 16632 8092 16638 8104
rect 1104 8042 21620 8064
rect 1104 7990 7846 8042
rect 7898 7990 7910 8042
rect 7962 7990 7974 8042
rect 8026 7990 8038 8042
rect 8090 7990 14710 8042
rect 14762 7990 14774 8042
rect 14826 7990 14838 8042
rect 14890 7990 14902 8042
rect 14954 7990 21620 8042
rect 1104 7968 21620 7990
rect 13170 7928 13176 7940
rect 13131 7900 13176 7928
rect 13170 7888 13176 7900
rect 13228 7888 13234 7940
rect 13541 7931 13599 7937
rect 13541 7897 13553 7931
rect 13587 7928 13599 7931
rect 13906 7928 13912 7940
rect 13587 7900 13912 7928
rect 13587 7897 13599 7900
rect 13541 7891 13599 7897
rect 13906 7888 13912 7900
rect 13964 7888 13970 7940
rect 14182 7888 14188 7940
rect 14240 7928 14246 7940
rect 19426 7928 19432 7940
rect 14240 7900 18460 7928
rect 19387 7900 19432 7928
rect 14240 7888 14246 7900
rect 10965 7863 11023 7869
rect 10965 7829 10977 7863
rect 11011 7860 11023 7863
rect 11238 7860 11244 7872
rect 11011 7832 11244 7860
rect 11011 7829 11023 7832
rect 10965 7823 11023 7829
rect 11238 7820 11244 7832
rect 11296 7820 11302 7872
rect 15749 7863 15807 7869
rect 15749 7829 15761 7863
rect 15795 7860 15807 7863
rect 15795 7832 16252 7860
rect 15795 7829 15807 7832
rect 15749 7823 15807 7829
rect 9306 7801 9312 7804
rect 9300 7792 9312 7801
rect 9267 7764 9312 7792
rect 9300 7755 9312 7764
rect 9306 7752 9312 7755
rect 9364 7752 9370 7804
rect 10686 7792 10692 7804
rect 10647 7764 10692 7792
rect 10686 7752 10692 7764
rect 10744 7752 10750 7804
rect 13998 7792 14004 7804
rect 13832 7764 14004 7792
rect 7466 7684 7472 7736
rect 7524 7724 7530 7736
rect 8202 7724 8208 7736
rect 7524 7696 8208 7724
rect 7524 7684 7530 7696
rect 8202 7684 8208 7696
rect 8260 7724 8266 7736
rect 9033 7727 9091 7733
rect 9033 7724 9045 7727
rect 8260 7696 9045 7724
rect 8260 7684 8266 7696
rect 9033 7693 9045 7696
rect 9079 7693 9091 7727
rect 9033 7687 9091 7693
rect 10318 7684 10324 7736
rect 10376 7724 10382 7736
rect 11425 7727 11483 7733
rect 11425 7724 11437 7727
rect 10376 7696 11437 7724
rect 10376 7684 10382 7696
rect 11425 7693 11437 7696
rect 11471 7693 11483 7727
rect 13630 7724 13636 7736
rect 13591 7696 13636 7724
rect 11425 7687 11483 7693
rect 13630 7684 13636 7696
rect 13688 7684 13694 7736
rect 13832 7733 13860 7764
rect 13998 7752 14004 7764
rect 14056 7792 14062 7804
rect 16114 7801 16120 7804
rect 14441 7795 14499 7801
rect 14441 7792 14453 7795
rect 14056 7764 14453 7792
rect 14056 7752 14062 7764
rect 14441 7761 14453 7764
rect 14487 7761 14499 7795
rect 16108 7792 16120 7801
rect 14441 7755 14499 7761
rect 15672 7764 16120 7792
rect 13817 7727 13875 7733
rect 13817 7693 13829 7727
rect 13863 7693 13875 7727
rect 13817 7687 13875 7693
rect 14090 7684 14096 7736
rect 14148 7724 14154 7736
rect 14185 7727 14243 7733
rect 14185 7724 14197 7727
rect 14148 7696 14197 7724
rect 14148 7684 14154 7696
rect 14185 7693 14197 7696
rect 14231 7693 14243 7727
rect 14185 7687 14243 7693
rect 10413 7591 10471 7597
rect 10413 7557 10425 7591
rect 10459 7588 10471 7591
rect 10502 7588 10508 7600
rect 10459 7560 10508 7588
rect 10459 7557 10471 7560
rect 10413 7551 10471 7557
rect 10502 7548 10508 7560
rect 10560 7548 10566 7600
rect 14200 7588 14228 7687
rect 15565 7659 15623 7665
rect 15565 7625 15577 7659
rect 15611 7656 15623 7659
rect 15672 7656 15700 7764
rect 16108 7755 16120 7764
rect 16114 7752 16120 7755
rect 16172 7752 16178 7804
rect 16224 7792 16252 7832
rect 17218 7820 17224 7872
rect 17276 7860 17282 7872
rect 18294 7863 18352 7869
rect 18294 7860 18306 7863
rect 17276 7832 18306 7860
rect 17276 7820 17282 7832
rect 18294 7829 18306 7832
rect 18340 7829 18352 7863
rect 18432 7860 18460 7900
rect 19426 7888 19432 7900
rect 19484 7888 19490 7940
rect 20717 7931 20775 7937
rect 20717 7897 20729 7931
rect 20763 7897 20775 7931
rect 20717 7891 20775 7897
rect 20732 7860 20760 7891
rect 18432 7832 20760 7860
rect 18294 7823 18352 7829
rect 18046 7792 18052 7804
rect 16224 7764 18052 7792
rect 18046 7752 18052 7764
rect 18104 7752 18110 7804
rect 19978 7792 19984 7804
rect 19939 7764 19984 7792
rect 19978 7752 19984 7764
rect 20036 7752 20042 7804
rect 20530 7792 20536 7804
rect 20491 7764 20536 7792
rect 20530 7752 20536 7764
rect 20588 7752 20594 7804
rect 15749 7727 15807 7733
rect 15749 7693 15761 7727
rect 15795 7724 15807 7727
rect 15841 7727 15899 7733
rect 15841 7724 15853 7727
rect 15795 7696 15853 7724
rect 15795 7693 15807 7696
rect 15749 7687 15807 7693
rect 15841 7693 15853 7696
rect 15887 7693 15899 7727
rect 15841 7687 15899 7693
rect 15611 7628 15700 7656
rect 15611 7625 15623 7628
rect 15565 7619 15623 7625
rect 15856 7588 15884 7687
rect 17218 7656 17224 7668
rect 17179 7628 17224 7656
rect 17218 7616 17224 7628
rect 17276 7616 17282 7668
rect 14200 7560 15884 7588
rect 16482 7548 16488 7600
rect 16540 7588 16546 7600
rect 20165 7591 20223 7597
rect 20165 7588 20177 7591
rect 16540 7560 20177 7588
rect 16540 7548 16546 7560
rect 20165 7557 20177 7560
rect 20211 7557 20223 7591
rect 20165 7551 20223 7557
rect 1104 7498 21620 7520
rect 1104 7446 4414 7498
rect 4466 7446 4478 7498
rect 4530 7446 4542 7498
rect 4594 7446 4606 7498
rect 4658 7446 11278 7498
rect 11330 7446 11342 7498
rect 11394 7446 11406 7498
rect 11458 7446 11470 7498
rect 11522 7446 18142 7498
rect 18194 7446 18206 7498
rect 18258 7446 18270 7498
rect 18322 7446 18334 7498
rect 18386 7446 21620 7498
rect 1104 7424 21620 7446
rect 9953 7387 10011 7393
rect 9953 7353 9965 7387
rect 9999 7384 10011 7387
rect 10686 7384 10692 7396
rect 9999 7356 10692 7384
rect 9999 7353 10011 7356
rect 9953 7347 10011 7353
rect 10686 7344 10692 7356
rect 10744 7344 10750 7396
rect 13998 7384 14004 7396
rect 13959 7356 14004 7384
rect 13998 7344 14004 7356
rect 14056 7344 14062 7396
rect 16574 7384 16580 7396
rect 16535 7356 16580 7384
rect 16574 7344 16580 7356
rect 16632 7344 16638 7396
rect 10502 7248 10508 7260
rect 10463 7220 10508 7248
rect 10502 7208 10508 7220
rect 10560 7208 10566 7260
rect 16114 7208 16120 7260
rect 16172 7248 16178 7260
rect 17129 7251 17187 7257
rect 17129 7248 17141 7251
rect 16172 7220 17141 7248
rect 16172 7208 16178 7220
rect 17129 7217 17141 7220
rect 17175 7217 17187 7251
rect 17129 7211 17187 7217
rect 10318 7180 10324 7192
rect 10279 7152 10324 7180
rect 10318 7140 10324 7152
rect 10376 7140 10382 7192
rect 10520 7112 10548 7208
rect 10965 7183 11023 7189
rect 10965 7149 10977 7183
rect 11011 7180 11023 7183
rect 12621 7183 12679 7189
rect 12621 7180 12633 7183
rect 11011 7152 12633 7180
rect 11011 7149 11023 7152
rect 10965 7143 11023 7149
rect 12621 7149 12633 7152
rect 12667 7180 12679 7183
rect 14090 7180 14096 7192
rect 12667 7152 14096 7180
rect 12667 7149 12679 7152
rect 12621 7143 12679 7149
rect 14090 7140 14096 7152
rect 14148 7140 14154 7192
rect 14182 7140 14188 7192
rect 14240 7180 14246 7192
rect 17037 7183 17095 7189
rect 17037 7180 17049 7183
rect 14240 7152 17049 7180
rect 14240 7140 14246 7152
rect 17037 7149 17049 7152
rect 17083 7180 17095 7183
rect 18874 7180 18880 7192
rect 17083 7152 18880 7180
rect 17083 7149 17095 7152
rect 17037 7143 17095 7149
rect 18874 7140 18880 7152
rect 18932 7140 18938 7192
rect 11210 7115 11268 7121
rect 11210 7112 11222 7115
rect 10520 7084 11222 7112
rect 11210 7081 11222 7084
rect 11256 7081 11268 7115
rect 12888 7115 12946 7121
rect 12888 7112 12900 7115
rect 11210 7075 11268 7081
rect 12360 7084 12900 7112
rect 10410 7004 10416 7056
rect 10468 7044 10474 7056
rect 12360 7053 12388 7084
rect 12888 7081 12900 7084
rect 12934 7112 12946 7115
rect 14366 7112 14372 7124
rect 12934 7084 14372 7112
rect 12934 7081 12946 7084
rect 12888 7075 12946 7081
rect 14366 7072 14372 7084
rect 14424 7072 14430 7124
rect 16945 7115 17003 7121
rect 16945 7081 16957 7115
rect 16991 7112 17003 7115
rect 18598 7112 18604 7124
rect 16991 7084 18604 7112
rect 16991 7081 17003 7084
rect 16945 7075 17003 7081
rect 18598 7072 18604 7084
rect 18656 7072 18662 7124
rect 12345 7047 12403 7053
rect 10468 7016 10513 7044
rect 10468 7004 10474 7016
rect 12345 7013 12357 7047
rect 12391 7013 12403 7047
rect 12345 7007 12403 7013
rect 17954 7004 17960 7056
rect 18012 7044 18018 7056
rect 18874 7044 18880 7056
rect 18012 7016 18880 7044
rect 18012 7004 18018 7016
rect 18874 7004 18880 7016
rect 18932 7004 18938 7056
rect 1104 6954 21620 6976
rect 1104 6902 7846 6954
rect 7898 6902 7910 6954
rect 7962 6902 7974 6954
rect 8026 6902 8038 6954
rect 8090 6902 14710 6954
rect 14762 6902 14774 6954
rect 14826 6902 14838 6954
rect 14890 6902 14902 6954
rect 14954 6902 21620 6954
rect 1104 6880 21620 6902
rect 10410 6800 10416 6852
rect 10468 6840 10474 6852
rect 10505 6843 10563 6849
rect 10505 6840 10517 6843
rect 10468 6812 10517 6840
rect 10468 6800 10474 6812
rect 10505 6809 10517 6812
rect 10551 6809 10563 6843
rect 13630 6840 13636 6852
rect 13591 6812 13636 6840
rect 10505 6803 10563 6809
rect 13630 6800 13636 6812
rect 13688 6800 13694 6852
rect 16482 6840 16488 6852
rect 13924 6812 16488 6840
rect 10873 6775 10931 6781
rect 10873 6741 10885 6775
rect 10919 6772 10931 6775
rect 13924 6772 13952 6812
rect 16482 6800 16488 6812
rect 16540 6800 16546 6852
rect 10919 6744 13952 6772
rect 14001 6775 14059 6781
rect 10919 6741 10931 6744
rect 10873 6735 10931 6741
rect 14001 6741 14013 6775
rect 14047 6772 14059 6775
rect 14047 6744 16528 6772
rect 14047 6741 14059 6744
rect 14001 6735 14059 6741
rect 3602 6664 3608 6716
rect 3660 6704 3666 6716
rect 7725 6707 7783 6713
rect 7725 6704 7737 6707
rect 3660 6676 7737 6704
rect 3660 6664 3666 6676
rect 7725 6673 7737 6676
rect 7771 6673 7783 6707
rect 7725 6667 7783 6673
rect 10778 6664 10784 6716
rect 10836 6704 10842 6716
rect 10965 6707 11023 6713
rect 10965 6704 10977 6707
rect 10836 6676 10977 6704
rect 10836 6664 10842 6676
rect 10965 6673 10977 6676
rect 11011 6704 11023 6707
rect 16500 6704 16528 6744
rect 18506 6704 18512 6716
rect 11011 6676 11836 6704
rect 16500 6676 18512 6704
rect 11011 6673 11023 6676
rect 10965 6667 11023 6673
rect 7466 6636 7472 6648
rect 7427 6608 7472 6636
rect 7466 6596 7472 6608
rect 7524 6596 7530 6648
rect 11057 6639 11115 6645
rect 11057 6605 11069 6639
rect 11103 6605 11115 6639
rect 11808 6636 11836 6676
rect 18506 6664 18512 6676
rect 18564 6664 18570 6716
rect 14090 6636 14096 6648
rect 11808 6608 14096 6636
rect 11057 6599 11115 6605
rect 8849 6571 8907 6577
rect 8849 6537 8861 6571
rect 8895 6568 8907 6571
rect 9306 6568 9312 6580
rect 8895 6540 9312 6568
rect 8895 6537 8907 6540
rect 8849 6531 8907 6537
rect 9306 6528 9312 6540
rect 9364 6568 9370 6580
rect 11072 6568 11100 6599
rect 14090 6596 14096 6608
rect 14148 6596 14154 6648
rect 14277 6639 14335 6645
rect 14277 6605 14289 6639
rect 14323 6636 14335 6639
rect 14366 6636 14372 6648
rect 14323 6608 14372 6636
rect 14323 6605 14335 6608
rect 14277 6599 14335 6605
rect 14366 6596 14372 6608
rect 14424 6596 14430 6648
rect 9364 6540 11100 6568
rect 9364 6528 9370 6540
rect 1104 6410 21620 6432
rect 1104 6358 4414 6410
rect 4466 6358 4478 6410
rect 4530 6358 4542 6410
rect 4594 6358 4606 6410
rect 4658 6358 11278 6410
rect 11330 6358 11342 6410
rect 11394 6358 11406 6410
rect 11458 6358 11470 6410
rect 11522 6358 18142 6410
rect 18194 6358 18206 6410
rect 18258 6358 18270 6410
rect 18322 6358 18334 6410
rect 18386 6358 21620 6410
rect 1104 6336 21620 6358
rect 14185 6299 14243 6305
rect 14185 6265 14197 6299
rect 14231 6296 14243 6299
rect 14274 6296 14280 6308
rect 14231 6268 14280 6296
rect 14231 6265 14243 6268
rect 14185 6259 14243 6265
rect 14274 6256 14280 6268
rect 14332 6256 14338 6308
rect 14001 6095 14059 6101
rect 14001 6061 14013 6095
rect 14047 6092 14059 6095
rect 17954 6092 17960 6104
rect 14047 6064 17960 6092
rect 14047 6061 14059 6064
rect 14001 6055 14059 6061
rect 17954 6052 17960 6064
rect 18012 6052 18018 6104
rect 1104 5866 21620 5888
rect 1104 5814 7846 5866
rect 7898 5814 7910 5866
rect 7962 5814 7974 5866
rect 8026 5814 8038 5866
rect 8090 5814 14710 5866
rect 14762 5814 14774 5866
rect 14826 5814 14838 5866
rect 14890 5814 14902 5866
rect 14954 5814 21620 5866
rect 1104 5792 21620 5814
rect 12986 5712 12992 5764
rect 13044 5752 13050 5764
rect 13081 5755 13139 5761
rect 13081 5752 13093 5755
rect 13044 5724 13093 5752
rect 13044 5712 13050 5724
rect 13081 5721 13093 5724
rect 13127 5721 13139 5755
rect 13081 5715 13139 5721
rect 12897 5619 12955 5625
rect 12897 5585 12909 5619
rect 12943 5616 12955 5619
rect 13814 5616 13820 5628
rect 12943 5588 13820 5616
rect 12943 5585 12955 5588
rect 12897 5579 12955 5585
rect 13814 5576 13820 5588
rect 13872 5576 13878 5628
rect 1104 5322 21620 5344
rect 1104 5270 4414 5322
rect 4466 5270 4478 5322
rect 4530 5270 4542 5322
rect 4594 5270 4606 5322
rect 4658 5270 11278 5322
rect 11330 5270 11342 5322
rect 11394 5270 11406 5322
rect 11458 5270 11470 5322
rect 11522 5270 18142 5322
rect 18194 5270 18206 5322
rect 18258 5270 18270 5322
rect 18322 5270 18334 5322
rect 18386 5270 21620 5322
rect 1104 5248 21620 5270
rect 13814 5168 13820 5220
rect 13872 5208 13878 5220
rect 17954 5208 17960 5220
rect 13872 5180 17960 5208
rect 13872 5168 13878 5180
rect 17954 5168 17960 5180
rect 18012 5168 18018 5220
rect 16482 5100 16488 5152
rect 16540 5140 16546 5152
rect 18046 5140 18052 5152
rect 16540 5112 18052 5140
rect 16540 5100 16546 5112
rect 18046 5100 18052 5112
rect 18104 5100 18110 5152
rect 1104 4778 21620 4800
rect 1104 4726 7846 4778
rect 7898 4726 7910 4778
rect 7962 4726 7974 4778
rect 8026 4726 8038 4778
rect 8090 4726 14710 4778
rect 14762 4726 14774 4778
rect 14826 4726 14838 4778
rect 14890 4726 14902 4778
rect 14954 4726 21620 4778
rect 1104 4704 21620 4726
rect 20717 4667 20775 4673
rect 20717 4633 20729 4667
rect 20763 4664 20775 4667
rect 20990 4664 20996 4676
rect 20763 4636 20996 4664
rect 20763 4633 20775 4636
rect 20717 4627 20775 4633
rect 20990 4624 20996 4636
rect 21048 4624 21054 4676
rect 20530 4528 20536 4540
rect 20491 4500 20536 4528
rect 20530 4488 20536 4500
rect 20588 4488 20594 4540
rect 1104 4234 21620 4256
rect 1104 4182 4414 4234
rect 4466 4182 4478 4234
rect 4530 4182 4542 4234
rect 4594 4182 4606 4234
rect 4658 4182 11278 4234
rect 11330 4182 11342 4234
rect 11394 4182 11406 4234
rect 11458 4182 11470 4234
rect 11522 4182 18142 4234
rect 18194 4182 18206 4234
rect 18258 4182 18270 4234
rect 18322 4182 18334 4234
rect 18386 4182 21620 4234
rect 1104 4160 21620 4182
rect 14550 3944 14556 3996
rect 14608 3984 14614 3996
rect 18506 3984 18512 3996
rect 14608 3956 18512 3984
rect 14608 3944 14614 3956
rect 18506 3944 18512 3956
rect 18564 3944 18570 3996
rect 1104 3690 21620 3712
rect 1104 3638 7846 3690
rect 7898 3638 7910 3690
rect 7962 3638 7974 3690
rect 8026 3638 8038 3690
rect 8090 3638 14710 3690
rect 14762 3638 14774 3690
rect 14826 3638 14838 3690
rect 14890 3638 14902 3690
rect 14954 3638 21620 3690
rect 1104 3616 21620 3638
rect 1104 3146 21620 3168
rect 1104 3094 4414 3146
rect 4466 3094 4478 3146
rect 4530 3094 4542 3146
rect 4594 3094 4606 3146
rect 4658 3094 11278 3146
rect 11330 3094 11342 3146
rect 11394 3094 11406 3146
rect 11458 3094 11470 3146
rect 11522 3094 18142 3146
rect 18194 3094 18206 3146
rect 18258 3094 18270 3146
rect 18322 3094 18334 3146
rect 18386 3094 21620 3146
rect 1104 3072 21620 3094
rect 1104 2602 21620 2624
rect 1104 2550 7846 2602
rect 7898 2550 7910 2602
rect 7962 2550 7974 2602
rect 8026 2550 8038 2602
rect 8090 2550 14710 2602
rect 14762 2550 14774 2602
rect 14826 2550 14838 2602
rect 14890 2550 14902 2602
rect 14954 2550 21620 2602
rect 1104 2528 21620 2550
rect 1104 2058 21620 2080
rect 1104 2006 4414 2058
rect 4466 2006 4478 2058
rect 4530 2006 4542 2058
rect 4594 2006 4606 2058
rect 4658 2006 11278 2058
rect 11330 2006 11342 2058
rect 11394 2006 11406 2058
rect 11458 2006 11470 2058
rect 11522 2006 18142 2058
rect 18194 2006 18206 2058
rect 18258 2006 18270 2058
rect 18322 2006 18334 2058
rect 18386 2006 21620 2058
rect 1104 1984 21620 2006
rect 16022 1156 16028 1208
rect 16080 1196 16086 1208
rect 18138 1196 18144 1208
rect 16080 1168 18144 1196
rect 16080 1156 16086 1168
rect 18138 1156 18144 1168
rect 18196 1156 18202 1208
<< via1 >>
rect 10324 20536 10376 20588
rect 17960 20536 18012 20588
rect 7846 19958 7898 20010
rect 7910 19958 7962 20010
rect 7974 19958 8026 20010
rect 8038 19958 8090 20010
rect 14710 19958 14762 20010
rect 14774 19958 14826 20010
rect 14838 19958 14890 20010
rect 14902 19958 14954 20010
rect 4712 19856 4764 19908
rect 18788 19899 18840 19908
rect 18788 19865 18797 19899
rect 18797 19865 18831 19899
rect 18831 19865 18840 19899
rect 18788 19856 18840 19865
rect 19340 19899 19392 19908
rect 19340 19865 19349 19899
rect 19349 19865 19383 19899
rect 19383 19865 19392 19899
rect 19340 19856 19392 19865
rect 20076 19899 20128 19908
rect 20076 19865 20085 19899
rect 20085 19865 20119 19899
rect 20119 19865 20128 19899
rect 20076 19856 20128 19865
rect 20628 19899 20680 19908
rect 20628 19865 20637 19899
rect 20637 19865 20671 19899
rect 20671 19865 20680 19899
rect 20628 19856 20680 19865
rect 9956 19788 10008 19840
rect 8484 19763 8536 19772
rect 8484 19729 8493 19763
rect 8493 19729 8527 19763
rect 8527 19729 8536 19763
rect 8484 19720 8536 19729
rect 18604 19763 18656 19772
rect 18604 19729 18613 19763
rect 18613 19729 18647 19763
rect 18647 19729 18656 19763
rect 18604 19720 18656 19729
rect 19156 19763 19208 19772
rect 19156 19729 19165 19763
rect 19165 19729 19199 19763
rect 19199 19729 19208 19763
rect 19156 19720 19208 19729
rect 20260 19720 20312 19772
rect 20444 19763 20496 19772
rect 20444 19729 20453 19763
rect 20453 19729 20487 19763
rect 20487 19729 20496 19763
rect 20444 19720 20496 19729
rect 4712 19652 4764 19704
rect 8300 19652 8352 19704
rect 17224 19695 17276 19704
rect 8392 19584 8444 19636
rect 17224 19661 17233 19695
rect 17233 19661 17267 19695
rect 17267 19661 17276 19695
rect 17224 19652 17276 19661
rect 5172 19516 5224 19568
rect 8116 19559 8168 19568
rect 8116 19525 8125 19559
rect 8125 19525 8159 19559
rect 8159 19525 8168 19559
rect 8116 19516 8168 19525
rect 4414 19414 4466 19466
rect 4478 19414 4530 19466
rect 4542 19414 4594 19466
rect 4606 19414 4658 19466
rect 11278 19414 11330 19466
rect 11342 19414 11394 19466
rect 11406 19414 11458 19466
rect 11470 19414 11522 19466
rect 18142 19414 18194 19466
rect 18206 19414 18258 19466
rect 18270 19414 18322 19466
rect 18334 19414 18386 19466
rect 8116 19312 8168 19364
rect 8484 19176 8536 19228
rect 10416 19219 10468 19228
rect 10416 19185 10425 19219
rect 10425 19185 10459 19219
rect 10459 19185 10468 19219
rect 10416 19176 10468 19185
rect 11888 19219 11940 19228
rect 11888 19185 11897 19219
rect 11897 19185 11931 19219
rect 11931 19185 11940 19219
rect 11888 19176 11940 19185
rect 16488 19219 16540 19228
rect 16488 19185 16497 19219
rect 16497 19185 16531 19219
rect 16531 19185 16540 19219
rect 16488 19176 16540 19185
rect 17500 19219 17552 19228
rect 17500 19185 17509 19219
rect 17509 19185 17543 19219
rect 17543 19185 17552 19219
rect 17500 19176 17552 19185
rect 2412 19108 2464 19160
rect 4712 19108 4764 19160
rect 7012 19151 7064 19160
rect 7012 19117 7021 19151
rect 7021 19117 7055 19151
rect 7055 19117 7064 19151
rect 7012 19108 7064 19117
rect 5080 19040 5132 19092
rect 6736 19040 6788 19092
rect 8208 19040 8260 19092
rect 9128 19108 9180 19160
rect 12624 19108 12676 19160
rect 14372 19108 14424 19160
rect 17224 19151 17276 19160
rect 17224 19117 17233 19151
rect 17233 19117 17267 19151
rect 17267 19117 17276 19151
rect 17224 19108 17276 19117
rect 18604 19176 18656 19228
rect 18788 19151 18840 19160
rect 18788 19117 18797 19151
rect 18797 19117 18831 19151
rect 18831 19117 18840 19151
rect 18788 19108 18840 19117
rect 20260 19219 20312 19228
rect 20260 19185 20269 19219
rect 20269 19185 20303 19219
rect 20303 19185 20312 19219
rect 20260 19176 20312 19185
rect 20076 19151 20128 19160
rect 20076 19117 20085 19151
rect 20085 19117 20119 19151
rect 20119 19117 20128 19151
rect 20076 19108 20128 19117
rect 9772 19040 9824 19092
rect 5448 19015 5500 19024
rect 5448 18981 5457 19015
rect 5457 18981 5491 19015
rect 5491 18981 5500 19015
rect 5448 18972 5500 18981
rect 8392 19015 8444 19024
rect 8392 18981 8401 19015
rect 8401 18981 8435 19015
rect 8435 18981 8444 19015
rect 8392 18972 8444 18981
rect 13820 19040 13872 19092
rect 9956 18972 10008 19024
rect 11244 18972 11296 19024
rect 11520 18972 11572 19024
rect 12164 18972 12216 19024
rect 12440 18972 12492 19024
rect 15384 19040 15436 19092
rect 14464 19015 14516 19024
rect 14464 18981 14473 19015
rect 14473 18981 14507 19015
rect 14507 18981 14516 19015
rect 14464 18972 14516 18981
rect 20444 19040 20496 19092
rect 16304 18972 16356 19024
rect 18972 19015 19024 19024
rect 18972 18981 18981 19015
rect 18981 18981 19015 19015
rect 19015 18981 19024 19015
rect 18972 18972 19024 18981
rect 7846 18870 7898 18922
rect 7910 18870 7962 18922
rect 7974 18870 8026 18922
rect 8038 18870 8090 18922
rect 14710 18870 14762 18922
rect 14774 18870 14826 18922
rect 14838 18870 14890 18922
rect 14902 18870 14954 18922
rect 4712 18768 4764 18820
rect 5172 18811 5224 18820
rect 5172 18777 5181 18811
rect 5181 18777 5215 18811
rect 5215 18777 5224 18811
rect 5172 18768 5224 18777
rect 6368 18768 6420 18820
rect 8208 18811 8260 18820
rect 296 18700 348 18752
rect 6736 18700 6788 18752
rect 2964 18632 3016 18684
rect 7012 18700 7064 18752
rect 8208 18777 8217 18811
rect 8217 18777 8251 18811
rect 8251 18777 8260 18811
rect 8208 18768 8260 18777
rect 11704 18768 11756 18820
rect 11888 18768 11940 18820
rect 12440 18768 12492 18820
rect 12532 18768 12584 18820
rect 12992 18768 13044 18820
rect 13820 18811 13872 18820
rect 13820 18777 13829 18811
rect 13829 18777 13863 18811
rect 13863 18777 13872 18811
rect 13820 18768 13872 18777
rect 14096 18768 14148 18820
rect 14556 18768 14608 18820
rect 1584 18564 1636 18616
rect 2412 18607 2464 18616
rect 2412 18573 2421 18607
rect 2421 18573 2455 18607
rect 2455 18573 2464 18607
rect 2412 18564 2464 18573
rect 5448 18564 5500 18616
rect 7380 18632 7432 18684
rect 8392 18700 8444 18752
rect 10416 18700 10468 18752
rect 14464 18700 14516 18752
rect 17960 18768 18012 18820
rect 19432 18768 19484 18820
rect 20720 18811 20772 18820
rect 20720 18777 20729 18811
rect 20729 18777 20763 18811
rect 20763 18777 20772 18811
rect 20720 18768 20772 18777
rect 16488 18743 16540 18752
rect 16488 18709 16522 18743
rect 16522 18709 16540 18743
rect 16488 18700 16540 18709
rect 18788 18700 18840 18752
rect 10232 18632 10284 18684
rect 14372 18632 14424 18684
rect 15936 18632 15988 18684
rect 17960 18632 18012 18684
rect 19156 18632 19208 18684
rect 19340 18675 19392 18684
rect 19340 18641 19349 18675
rect 19349 18641 19383 18675
rect 19383 18641 19392 18675
rect 19340 18632 19392 18641
rect 19524 18632 19576 18684
rect 5080 18496 5132 18548
rect 9864 18564 9916 18616
rect 11428 18564 11480 18616
rect 11888 18564 11940 18616
rect 14096 18607 14148 18616
rect 5172 18428 5224 18480
rect 7012 18428 7064 18480
rect 14096 18573 14105 18607
rect 14105 18573 14139 18607
rect 14139 18573 14148 18607
rect 14096 18564 14148 18573
rect 17684 18564 17736 18616
rect 21180 18564 21232 18616
rect 12624 18428 12676 18480
rect 12716 18428 12768 18480
rect 20076 18496 20128 18548
rect 17592 18471 17644 18480
rect 17592 18437 17601 18471
rect 17601 18437 17635 18471
rect 17635 18437 17644 18471
rect 17592 18428 17644 18437
rect 19064 18428 19116 18480
rect 20628 18428 20680 18480
rect 4414 18326 4466 18378
rect 4478 18326 4530 18378
rect 4542 18326 4594 18378
rect 4606 18326 4658 18378
rect 11278 18326 11330 18378
rect 11342 18326 11394 18378
rect 11406 18326 11458 18378
rect 11470 18326 11522 18378
rect 18142 18326 18194 18378
rect 18206 18326 18258 18378
rect 18270 18326 18322 18378
rect 18334 18326 18386 18378
rect 1952 18224 2004 18276
rect 3056 18224 3108 18276
rect 5356 18224 5408 18276
rect 8300 18224 8352 18276
rect 9772 18224 9824 18276
rect 10692 18224 10744 18276
rect 11612 18224 11664 18276
rect 12716 18224 12768 18276
rect 5724 18156 5776 18208
rect 5816 18156 5868 18208
rect 11520 18156 11572 18208
rect 8208 18088 8260 18140
rect 9772 18088 9824 18140
rect 12072 18156 12124 18208
rect 12164 18088 12216 18140
rect 3608 18020 3660 18072
rect 4252 18020 4304 18072
rect 5172 18063 5224 18072
rect 5172 18029 5181 18063
rect 5181 18029 5215 18063
rect 5215 18029 5224 18063
rect 5172 18020 5224 18029
rect 8576 18020 8628 18072
rect 9680 18020 9732 18072
rect 19340 18224 19392 18276
rect 13636 18156 13688 18208
rect 14280 18156 14332 18208
rect 19892 18156 19944 18208
rect 21364 18156 21416 18208
rect 13820 18088 13872 18140
rect 14464 18088 14516 18140
rect 19800 18088 19852 18140
rect 21916 18088 21968 18140
rect 5264 17952 5316 18004
rect 7472 17952 7524 18004
rect 8484 17952 8536 18004
rect 10784 17952 10836 18004
rect 12716 17952 12768 18004
rect 8760 17884 8812 17936
rect 11152 17884 11204 17936
rect 11980 17884 12032 17936
rect 12072 17884 12124 17936
rect 13360 17952 13412 18004
rect 14096 18020 14148 18072
rect 20260 18063 20312 18072
rect 20260 18029 20269 18063
rect 20269 18029 20303 18063
rect 20303 18029 20312 18063
rect 20260 18020 20312 18029
rect 13084 17884 13136 17936
rect 13636 17884 13688 17936
rect 15844 17952 15896 18004
rect 19340 17952 19392 18004
rect 19708 17952 19760 18004
rect 20352 17952 20404 18004
rect 15200 17884 15252 17936
rect 15292 17884 15344 17936
rect 16488 17884 16540 17936
rect 16948 17884 17000 17936
rect 20076 17884 20128 17936
rect 20444 17927 20496 17936
rect 20444 17893 20453 17927
rect 20453 17893 20487 17927
rect 20487 17893 20496 17927
rect 20444 17884 20496 17893
rect 20996 17884 21048 17936
rect 22468 17884 22520 17936
rect 7846 17782 7898 17834
rect 7910 17782 7962 17834
rect 7974 17782 8026 17834
rect 8038 17782 8090 17834
rect 14710 17782 14762 17834
rect 14774 17782 14826 17834
rect 14838 17782 14890 17834
rect 14902 17782 14954 17834
rect 2964 17723 3016 17732
rect 2964 17689 2973 17723
rect 2973 17689 3007 17723
rect 3007 17689 3016 17723
rect 2964 17680 3016 17689
rect 5264 17680 5316 17732
rect 12164 17680 12216 17732
rect 19340 17680 19392 17732
rect 19616 17723 19668 17732
rect 19616 17689 19625 17723
rect 19625 17689 19659 17723
rect 19659 17689 19668 17723
rect 19616 17680 19668 17689
rect 19708 17680 19760 17732
rect 20076 17680 20128 17732
rect 20444 17680 20496 17732
rect 20812 17680 20864 17732
rect 1584 17587 1636 17596
rect 1584 17553 1593 17587
rect 1593 17553 1627 17587
rect 1627 17553 1636 17587
rect 1584 17544 1636 17553
rect 3148 17544 3200 17596
rect 5448 17612 5500 17664
rect 5632 17612 5684 17664
rect 16120 17612 16172 17664
rect 16304 17544 16356 17596
rect 17224 17544 17276 17596
rect 3332 17519 3384 17528
rect 3332 17485 3341 17519
rect 3341 17485 3375 17519
rect 3375 17485 3384 17519
rect 3332 17476 3384 17485
rect 5080 17519 5132 17528
rect 5080 17485 5089 17519
rect 5089 17485 5123 17519
rect 5123 17485 5132 17519
rect 5080 17476 5132 17485
rect 7472 17476 7524 17528
rect 19524 17476 19576 17528
rect 20076 17544 20128 17596
rect 20812 17476 20864 17528
rect 9680 17408 9732 17460
rect 17408 17408 17460 17460
rect 8668 17340 8720 17392
rect 11704 17340 11756 17392
rect 12348 17340 12400 17392
rect 16120 17340 16172 17392
rect 18512 17340 18564 17392
rect 20168 17383 20220 17392
rect 20168 17349 20177 17383
rect 20177 17349 20211 17383
rect 20211 17349 20220 17383
rect 20168 17340 20220 17349
rect 20720 17383 20772 17392
rect 20720 17349 20729 17383
rect 20729 17349 20763 17383
rect 20763 17349 20772 17383
rect 20720 17340 20772 17349
rect 4414 17238 4466 17290
rect 4478 17238 4530 17290
rect 4542 17238 4594 17290
rect 4606 17238 4658 17290
rect 11278 17238 11330 17290
rect 11342 17238 11394 17290
rect 11406 17238 11458 17290
rect 11470 17238 11522 17290
rect 18142 17238 18194 17290
rect 18206 17238 18258 17290
rect 18270 17238 18322 17290
rect 18334 17238 18386 17290
rect 9680 17179 9732 17188
rect 9680 17145 9689 17179
rect 9689 17145 9723 17179
rect 9723 17145 9732 17179
rect 9680 17136 9732 17145
rect 17224 17136 17276 17188
rect 17960 17136 18012 17188
rect 3148 17068 3200 17120
rect 2964 17000 3016 17052
rect 4160 17000 4212 17052
rect 3332 16975 3384 16984
rect 3332 16941 3341 16975
rect 3341 16941 3375 16975
rect 3375 16941 3384 16975
rect 3332 16932 3384 16941
rect 8760 17068 8812 17120
rect 12164 17111 12216 17120
rect 12164 17077 12173 17111
rect 12173 17077 12207 17111
rect 12207 17077 12216 17111
rect 12164 17068 12216 17077
rect 12348 17068 12400 17120
rect 5540 17000 5592 17052
rect 7472 17043 7524 17052
rect 6828 16932 6880 16984
rect 7472 17009 7481 17043
rect 7481 17009 7515 17043
rect 7515 17009 7524 17043
rect 7472 17000 7524 17009
rect 8668 17043 8720 17052
rect 8668 17009 8677 17043
rect 8677 17009 8711 17043
rect 8711 17009 8720 17043
rect 8668 17000 8720 17009
rect 10232 17043 10284 17052
rect 10232 17009 10241 17043
rect 10241 17009 10275 17043
rect 10275 17009 10284 17043
rect 10232 17000 10284 17009
rect 11704 17043 11756 17052
rect 11704 17009 11713 17043
rect 11713 17009 11747 17043
rect 11747 17009 11756 17043
rect 11704 17000 11756 17009
rect 12716 17043 12768 17052
rect 12716 17009 12725 17043
rect 12725 17009 12759 17043
rect 12759 17009 12768 17043
rect 12716 17000 12768 17009
rect 11612 16975 11664 16984
rect 11612 16941 11621 16975
rect 11621 16941 11655 16975
rect 11655 16941 11664 16975
rect 11612 16932 11664 16941
rect 14096 17000 14148 17052
rect 15936 17043 15988 17052
rect 15936 17009 15945 17043
rect 15945 17009 15979 17043
rect 15979 17009 15988 17043
rect 15936 17000 15988 17009
rect 17684 17000 17736 17052
rect 20260 17000 20312 17052
rect 20812 17000 20864 17052
rect 17592 16932 17644 16984
rect 19340 16975 19392 16984
rect 19340 16941 19349 16975
rect 19349 16941 19383 16975
rect 19383 16941 19392 16975
rect 19340 16932 19392 16941
rect 19432 16932 19484 16984
rect 2964 16839 3016 16848
rect 2964 16805 2973 16839
rect 2973 16805 3007 16839
rect 3007 16805 3016 16839
rect 2964 16796 3016 16805
rect 9772 16796 9824 16848
rect 10048 16839 10100 16848
rect 10048 16805 10057 16839
rect 10057 16805 10091 16839
rect 10091 16805 10100 16839
rect 10048 16796 10100 16805
rect 12532 16839 12584 16848
rect 12532 16805 12541 16839
rect 12541 16805 12575 16839
rect 12575 16805 12584 16839
rect 12532 16796 12584 16805
rect 14004 16839 14056 16848
rect 14004 16805 14013 16839
rect 14013 16805 14047 16839
rect 14047 16805 14056 16839
rect 14004 16796 14056 16805
rect 14372 16839 14424 16848
rect 14372 16805 14381 16839
rect 14381 16805 14415 16839
rect 14415 16805 14424 16839
rect 14372 16796 14424 16805
rect 17316 16839 17368 16848
rect 17316 16805 17325 16839
rect 17325 16805 17359 16839
rect 17359 16805 17368 16839
rect 17316 16796 17368 16805
rect 17960 16796 18012 16848
rect 7846 16694 7898 16746
rect 7910 16694 7962 16746
rect 7974 16694 8026 16746
rect 8038 16694 8090 16746
rect 14710 16694 14762 16746
rect 14774 16694 14826 16746
rect 14838 16694 14890 16746
rect 14902 16694 14954 16746
rect 6828 16635 6880 16644
rect 6828 16601 6837 16635
rect 6837 16601 6871 16635
rect 6871 16601 6880 16635
rect 6828 16592 6880 16601
rect 7288 16635 7340 16644
rect 7288 16601 7297 16635
rect 7297 16601 7331 16635
rect 7331 16601 7340 16635
rect 7288 16592 7340 16601
rect 8668 16524 8720 16576
rect 11704 16592 11756 16644
rect 12532 16592 12584 16644
rect 14004 16592 14056 16644
rect 18512 16592 18564 16644
rect 10232 16524 10284 16576
rect 2964 16456 3016 16508
rect 5632 16456 5684 16508
rect 7380 16431 7432 16440
rect 7380 16397 7389 16431
rect 7389 16397 7423 16431
rect 7423 16397 7432 16431
rect 7380 16388 7432 16397
rect 8208 16431 8260 16440
rect 8208 16397 8217 16431
rect 8217 16397 8251 16431
rect 8251 16397 8260 16431
rect 8208 16388 8260 16397
rect 9588 16388 9640 16440
rect 9864 16431 9916 16440
rect 9864 16397 9873 16431
rect 9873 16397 9907 16431
rect 9907 16397 9916 16431
rect 9864 16388 9916 16397
rect 12532 16456 12584 16508
rect 12716 16456 12768 16508
rect 19432 16524 19484 16576
rect 12624 16431 12676 16440
rect 12624 16397 12633 16431
rect 12633 16397 12667 16431
rect 12667 16397 12676 16431
rect 12624 16388 12676 16397
rect 14096 16320 14148 16372
rect 15936 16456 15988 16508
rect 17316 16456 17368 16508
rect 17408 16456 17460 16508
rect 19708 16592 19760 16644
rect 20260 16592 20312 16644
rect 20628 16592 20680 16644
rect 20076 16524 20128 16576
rect 15108 16431 15160 16440
rect 15108 16397 15117 16431
rect 15117 16397 15151 16431
rect 15151 16397 15160 16431
rect 15108 16388 15160 16397
rect 17684 16295 17736 16304
rect 17684 16261 17693 16295
rect 17693 16261 17727 16295
rect 17727 16261 17736 16295
rect 17684 16252 17736 16261
rect 19616 16252 19668 16304
rect 19892 16252 19944 16304
rect 4414 16150 4466 16202
rect 4478 16150 4530 16202
rect 4542 16150 4594 16202
rect 4606 16150 4658 16202
rect 11278 16150 11330 16202
rect 11342 16150 11394 16202
rect 11406 16150 11458 16202
rect 11470 16150 11522 16202
rect 18142 16150 18194 16202
rect 18206 16150 18258 16202
rect 18270 16150 18322 16202
rect 18334 16150 18386 16202
rect 3148 16091 3200 16100
rect 3148 16057 3157 16091
rect 3157 16057 3191 16091
rect 3191 16057 3200 16091
rect 3148 16048 3200 16057
rect 7288 16048 7340 16100
rect 12532 16091 12584 16100
rect 7380 15980 7432 16032
rect 5080 15912 5132 15964
rect 7656 15955 7708 15964
rect 1584 15844 1636 15896
rect 7656 15921 7665 15955
rect 7665 15921 7699 15955
rect 7699 15921 7708 15955
rect 7656 15912 7708 15921
rect 10048 15912 10100 15964
rect 12532 16057 12541 16091
rect 12541 16057 12575 16091
rect 12575 16057 12584 16091
rect 12532 16048 12584 16057
rect 12624 16048 12676 16100
rect 13452 15912 13504 15964
rect 15936 16048 15988 16100
rect 17960 16048 18012 16100
rect 18880 16048 18932 16100
rect 20444 16023 20496 16032
rect 20444 15989 20453 16023
rect 20453 15989 20487 16023
rect 20487 15989 20496 16023
rect 20444 15980 20496 15989
rect 17316 15955 17368 15964
rect 17316 15921 17325 15955
rect 17325 15921 17359 15955
rect 17359 15921 17368 15955
rect 17316 15912 17368 15921
rect 7748 15844 7800 15896
rect 14096 15844 14148 15896
rect 15200 15844 15252 15896
rect 19156 15844 19208 15896
rect 19892 15844 19944 15896
rect 2964 15776 3016 15828
rect 11704 15776 11756 15828
rect 14372 15776 14424 15828
rect 7748 15708 7800 15760
rect 14556 15708 14608 15760
rect 15108 15708 15160 15760
rect 15200 15708 15252 15760
rect 7846 15606 7898 15658
rect 7910 15606 7962 15658
rect 7974 15606 8026 15658
rect 8038 15606 8090 15658
rect 14710 15606 14762 15658
rect 14774 15606 14826 15658
rect 14838 15606 14890 15658
rect 14902 15606 14954 15658
rect 7656 15504 7708 15556
rect 20720 15547 20772 15556
rect 20720 15513 20729 15547
rect 20729 15513 20763 15547
rect 20763 15513 20772 15547
rect 20720 15504 20772 15513
rect 19156 15479 19208 15488
rect 4988 15368 5040 15420
rect 6828 15368 6880 15420
rect 16580 15411 16632 15420
rect 16580 15377 16589 15411
rect 16589 15377 16623 15411
rect 16623 15377 16632 15411
rect 16580 15368 16632 15377
rect 19156 15445 19165 15479
rect 19165 15445 19199 15479
rect 19199 15445 19208 15479
rect 19156 15436 19208 15445
rect 19892 15479 19944 15488
rect 19892 15445 19901 15479
rect 19901 15445 19935 15479
rect 19935 15445 19944 15479
rect 19892 15436 19944 15445
rect 2964 15300 3016 15352
rect 3424 15343 3476 15352
rect 3424 15309 3433 15343
rect 3433 15309 3467 15343
rect 3467 15309 3476 15343
rect 3424 15300 3476 15309
rect 16672 15343 16724 15352
rect 16672 15309 16681 15343
rect 16681 15309 16715 15343
rect 16715 15309 16724 15343
rect 16672 15300 16724 15309
rect 16764 15343 16816 15352
rect 16764 15309 16773 15343
rect 16773 15309 16807 15343
rect 16807 15309 16816 15343
rect 16764 15300 16816 15309
rect 15108 15232 15160 15284
rect 20076 15368 20128 15420
rect 17868 15164 17920 15216
rect 4414 15062 4466 15114
rect 4478 15062 4530 15114
rect 4542 15062 4594 15114
rect 4606 15062 4658 15114
rect 11278 15062 11330 15114
rect 11342 15062 11394 15114
rect 11406 15062 11458 15114
rect 11470 15062 11522 15114
rect 18142 15062 18194 15114
rect 18206 15062 18258 15114
rect 18270 15062 18322 15114
rect 18334 15062 18386 15114
rect 2504 14960 2556 15012
rect 2964 15003 3016 15012
rect 2964 14969 2973 15003
rect 2973 14969 3007 15003
rect 3007 14969 3016 15003
rect 2964 14960 3016 14969
rect 3424 14960 3476 15012
rect 6828 14960 6880 15012
rect 1584 14867 1636 14876
rect 1584 14833 1593 14867
rect 1593 14833 1627 14867
rect 1627 14833 1636 14867
rect 1584 14824 1636 14833
rect 3700 14824 3752 14876
rect 4252 14756 4304 14808
rect 3700 14688 3752 14740
rect 7472 14824 7524 14876
rect 15108 14960 15160 15012
rect 16672 14960 16724 15012
rect 20444 15003 20496 15012
rect 20444 14969 20453 15003
rect 20453 14969 20487 15003
rect 20487 14969 20496 15003
rect 20444 14960 20496 14969
rect 9404 14892 9456 14944
rect 12164 14892 12216 14944
rect 5080 14620 5132 14672
rect 7656 14756 7708 14808
rect 7932 14799 7984 14808
rect 7932 14765 7941 14799
rect 7941 14765 7975 14799
rect 7975 14765 7984 14799
rect 7932 14756 7984 14765
rect 12808 14867 12860 14876
rect 12256 14756 12308 14808
rect 12808 14833 12817 14867
rect 12817 14833 12851 14867
rect 12851 14833 12860 14867
rect 12808 14824 12860 14833
rect 13912 14756 13964 14808
rect 15384 14824 15436 14876
rect 16764 14867 16816 14876
rect 16764 14833 16773 14867
rect 16773 14833 16807 14867
rect 16807 14833 16816 14867
rect 16764 14824 16816 14833
rect 17776 14756 17828 14808
rect 17868 14756 17920 14808
rect 19340 14756 19392 14808
rect 8668 14688 8720 14740
rect 20536 14688 20588 14740
rect 9036 14620 9088 14672
rect 9772 14620 9824 14672
rect 10140 14663 10192 14672
rect 10140 14629 10149 14663
rect 10149 14629 10183 14663
rect 10183 14629 10192 14663
rect 12624 14663 12676 14672
rect 10140 14620 10192 14629
rect 12624 14629 12633 14663
rect 12633 14629 12667 14663
rect 12667 14629 12676 14663
rect 12624 14620 12676 14629
rect 12716 14663 12768 14672
rect 12716 14629 12725 14663
rect 12725 14629 12759 14663
rect 12759 14629 12768 14663
rect 13452 14663 13504 14672
rect 12716 14620 12768 14629
rect 13452 14629 13461 14663
rect 13461 14629 13495 14663
rect 13495 14629 13504 14663
rect 13452 14620 13504 14629
rect 15476 14620 15528 14672
rect 16304 14620 16356 14672
rect 7846 14518 7898 14570
rect 7910 14518 7962 14570
rect 7974 14518 8026 14570
rect 8038 14518 8090 14570
rect 14710 14518 14762 14570
rect 14774 14518 14826 14570
rect 14838 14518 14890 14570
rect 14902 14518 14954 14570
rect 5356 14416 5408 14468
rect 8668 14459 8720 14468
rect 8668 14425 8677 14459
rect 8677 14425 8711 14459
rect 8711 14425 8720 14459
rect 8668 14416 8720 14425
rect 9772 14459 9824 14468
rect 9772 14425 9781 14459
rect 9781 14425 9815 14459
rect 9815 14425 9824 14459
rect 9772 14416 9824 14425
rect 1584 14280 1636 14332
rect 2320 14280 2372 14332
rect 4896 14280 4948 14332
rect 5080 14280 5132 14332
rect 7012 14280 7064 14332
rect 9404 14348 9456 14400
rect 12716 14416 12768 14468
rect 15476 14416 15528 14468
rect 12256 14348 12308 14400
rect 13452 14348 13504 14400
rect 10968 14323 11020 14332
rect 10968 14289 10991 14323
rect 10991 14289 11020 14323
rect 10968 14280 11020 14289
rect 14556 14348 14608 14400
rect 16856 14416 16908 14468
rect 18696 14459 18748 14468
rect 18696 14425 18705 14459
rect 18705 14425 18739 14459
rect 18739 14425 18748 14459
rect 18696 14416 18748 14425
rect 20628 14416 20680 14468
rect 16764 14348 16816 14400
rect 17776 14348 17828 14400
rect 19340 14391 19392 14400
rect 18512 14323 18564 14332
rect 18512 14289 18521 14323
rect 18521 14289 18555 14323
rect 18555 14289 18564 14323
rect 18512 14280 18564 14289
rect 19340 14357 19349 14391
rect 19349 14357 19383 14391
rect 19383 14357 19392 14391
rect 19340 14348 19392 14357
rect 20076 14391 20128 14400
rect 20076 14357 20085 14391
rect 20085 14357 20119 14391
rect 20119 14357 20128 14391
rect 20076 14348 20128 14357
rect 19800 14323 19852 14332
rect 19800 14289 19819 14323
rect 19819 14289 19852 14323
rect 20536 14323 20588 14332
rect 19800 14280 19852 14289
rect 20536 14289 20545 14323
rect 20545 14289 20579 14323
rect 20579 14289 20588 14323
rect 20536 14280 20588 14289
rect 13452 14255 13504 14264
rect 5080 14144 5132 14196
rect 6920 14076 6972 14128
rect 8300 14144 8352 14196
rect 9956 14144 10008 14196
rect 12532 14144 12584 14196
rect 13452 14221 13461 14255
rect 13461 14221 13495 14255
rect 13495 14221 13504 14255
rect 13452 14212 13504 14221
rect 17500 14255 17552 14264
rect 17500 14221 17509 14255
rect 17509 14221 17543 14255
rect 17543 14221 17552 14255
rect 17500 14212 17552 14221
rect 7656 14076 7708 14128
rect 7932 14076 7984 14128
rect 12072 14076 12124 14128
rect 12808 14076 12860 14128
rect 4414 13974 4466 14026
rect 4478 13974 4530 14026
rect 4542 13974 4594 14026
rect 4606 13974 4658 14026
rect 11278 13974 11330 14026
rect 11342 13974 11394 14026
rect 11406 13974 11458 14026
rect 11470 13974 11522 14026
rect 18142 13974 18194 14026
rect 18206 13974 18258 14026
rect 18270 13974 18322 14026
rect 18334 13974 18386 14026
rect 3700 13915 3752 13924
rect 3700 13881 3709 13915
rect 3709 13881 3743 13915
rect 3743 13881 3752 13915
rect 3700 13872 3752 13881
rect 2320 13779 2372 13788
rect 2320 13745 2329 13779
rect 2329 13745 2363 13779
rect 2363 13745 2372 13779
rect 2320 13736 2372 13745
rect 10140 13872 10192 13924
rect 10968 13872 11020 13924
rect 12532 13872 12584 13924
rect 12624 13872 12676 13924
rect 16580 13915 16632 13924
rect 16580 13881 16589 13915
rect 16589 13881 16623 13915
rect 16623 13881 16632 13915
rect 16580 13872 16632 13881
rect 16672 13872 16724 13924
rect 20444 13915 20496 13924
rect 6920 13779 6972 13788
rect 6920 13745 6929 13779
rect 6929 13745 6963 13779
rect 6963 13745 6972 13779
rect 6920 13736 6972 13745
rect 9864 13804 9916 13856
rect 19892 13847 19944 13856
rect 19892 13813 19901 13847
rect 19901 13813 19935 13847
rect 19935 13813 19944 13847
rect 19892 13804 19944 13813
rect 8484 13779 8536 13788
rect 8484 13745 8493 13779
rect 8493 13745 8527 13779
rect 8527 13745 8536 13779
rect 8484 13736 8536 13745
rect 8668 13779 8720 13788
rect 8668 13745 8677 13779
rect 8677 13745 8711 13779
rect 8711 13745 8720 13779
rect 8668 13736 8720 13745
rect 12532 13736 12584 13788
rect 16764 13736 16816 13788
rect 18512 13736 18564 13788
rect 4896 13668 4948 13720
rect 5080 13711 5132 13720
rect 5080 13677 5114 13711
rect 5114 13677 5132 13711
rect 5080 13668 5132 13677
rect 9772 13668 9824 13720
rect 7012 13600 7064 13652
rect 13452 13668 13504 13720
rect 6828 13575 6880 13584
rect 6828 13541 6837 13575
rect 6837 13541 6871 13575
rect 6871 13541 6880 13575
rect 6828 13532 6880 13541
rect 9036 13575 9088 13584
rect 9036 13541 9045 13575
rect 9045 13541 9079 13575
rect 9079 13541 9088 13575
rect 9036 13532 9088 13541
rect 9956 13600 10008 13652
rect 10416 13600 10468 13652
rect 17500 13668 17552 13720
rect 19800 13668 19852 13720
rect 20444 13881 20453 13915
rect 20453 13881 20487 13915
rect 20487 13881 20496 13915
rect 20444 13872 20496 13881
rect 17408 13600 17460 13652
rect 18512 13600 18564 13652
rect 14372 13532 14424 13584
rect 7846 13430 7898 13482
rect 7910 13430 7962 13482
rect 7974 13430 8026 13482
rect 8038 13430 8090 13482
rect 14710 13430 14762 13482
rect 14774 13430 14826 13482
rect 14838 13430 14890 13482
rect 14902 13430 14954 13482
rect 6828 13328 6880 13380
rect 9772 13328 9824 13380
rect 10968 13328 11020 13380
rect 19708 13371 19760 13380
rect 19708 13337 19717 13371
rect 19717 13337 19751 13371
rect 19751 13337 19760 13371
rect 19708 13328 19760 13337
rect 20720 13371 20772 13380
rect 20720 13337 20729 13371
rect 20729 13337 20763 13371
rect 20763 13337 20772 13371
rect 20720 13328 20772 13337
rect 10324 13260 10376 13312
rect 14096 13235 14148 13244
rect 14096 13201 14105 13235
rect 14105 13201 14139 13235
rect 14139 13201 14148 13235
rect 14096 13192 14148 13201
rect 18972 13192 19024 13244
rect 13176 13124 13228 13176
rect 13820 13056 13872 13108
rect 15568 13124 15620 13176
rect 14832 12988 14884 13040
rect 4414 12886 4466 12938
rect 4478 12886 4530 12938
rect 4542 12886 4594 12938
rect 4606 12886 4658 12938
rect 11278 12886 11330 12938
rect 11342 12886 11394 12938
rect 11406 12886 11458 12938
rect 11470 12886 11522 12938
rect 18142 12886 18194 12938
rect 18206 12886 18258 12938
rect 18270 12886 18322 12938
rect 18334 12886 18386 12938
rect 13176 12827 13228 12836
rect 848 12648 900 12700
rect 5724 12648 5776 12700
rect 7380 12648 7432 12700
rect 8208 12691 8260 12700
rect 8208 12657 8217 12691
rect 8217 12657 8251 12691
rect 8251 12657 8260 12691
rect 8208 12648 8260 12657
rect 13176 12793 13185 12827
rect 13185 12793 13219 12827
rect 13219 12793 13228 12827
rect 13176 12784 13228 12793
rect 13544 12784 13596 12836
rect 16488 12784 16540 12836
rect 19616 12784 19668 12836
rect 20352 12784 20404 12836
rect 10416 12691 10468 12700
rect 10416 12657 10425 12691
rect 10425 12657 10459 12691
rect 10459 12657 10468 12691
rect 10416 12648 10468 12657
rect 7012 12623 7064 12632
rect 7012 12589 7021 12623
rect 7021 12589 7055 12623
rect 7055 12589 7064 12623
rect 7012 12580 7064 12589
rect 13544 12648 13596 12700
rect 13728 12691 13780 12700
rect 13728 12657 13737 12691
rect 13737 12657 13771 12691
rect 13771 12657 13780 12691
rect 13728 12648 13780 12657
rect 10968 12580 11020 12632
rect 7748 12444 7800 12496
rect 10232 12487 10284 12496
rect 10232 12453 10241 12487
rect 10241 12453 10275 12487
rect 10275 12453 10284 12487
rect 10232 12444 10284 12453
rect 13912 12512 13964 12564
rect 14372 12716 14424 12768
rect 14740 12691 14792 12700
rect 14740 12657 14749 12691
rect 14749 12657 14783 12691
rect 14783 12657 14792 12691
rect 14740 12648 14792 12657
rect 14832 12648 14884 12700
rect 15568 12691 15620 12700
rect 15568 12657 15577 12691
rect 15577 12657 15611 12691
rect 15611 12657 15620 12691
rect 15568 12648 15620 12657
rect 18972 12691 19024 12700
rect 16028 12580 16080 12632
rect 18972 12657 18981 12691
rect 18981 12657 19015 12691
rect 19015 12657 19024 12691
rect 18972 12648 19024 12657
rect 17316 12580 17368 12632
rect 18696 12623 18748 12632
rect 18696 12589 18705 12623
rect 18705 12589 18739 12623
rect 18739 12589 18748 12623
rect 18696 12580 18748 12589
rect 19708 12623 19760 12632
rect 19708 12589 19717 12623
rect 19717 12589 19751 12623
rect 19751 12589 19760 12623
rect 19708 12580 19760 12589
rect 20260 12623 20312 12632
rect 20260 12589 20269 12623
rect 20269 12589 20303 12623
rect 20303 12589 20312 12623
rect 20260 12580 20312 12589
rect 17684 12512 17736 12564
rect 14372 12444 14424 12496
rect 14556 12487 14608 12496
rect 14556 12453 14565 12487
rect 14565 12453 14599 12487
rect 14599 12453 14608 12487
rect 14556 12444 14608 12453
rect 15108 12444 15160 12496
rect 7846 12342 7898 12394
rect 7910 12342 7962 12394
rect 7974 12342 8026 12394
rect 8038 12342 8090 12394
rect 14710 12342 14762 12394
rect 14774 12342 14826 12394
rect 14838 12342 14890 12394
rect 14902 12342 14954 12394
rect 10232 12240 10284 12292
rect 7656 12172 7708 12224
rect 8300 12172 8352 12224
rect 9680 12172 9732 12224
rect 13728 12172 13780 12224
rect 14096 12240 14148 12292
rect 17408 12240 17460 12292
rect 17776 12240 17828 12292
rect 18696 12240 18748 12292
rect 19984 12240 20036 12292
rect 21088 12240 21140 12292
rect 17960 12172 18012 12224
rect 18604 12172 18656 12224
rect 7380 12104 7432 12156
rect 8208 12104 8260 12156
rect 6828 12079 6880 12088
rect 6828 12045 6837 12079
rect 6837 12045 6871 12079
rect 6871 12045 6880 12079
rect 6828 12036 6880 12045
rect 8300 12036 8352 12088
rect 15200 12104 15252 12156
rect 17040 12104 17092 12156
rect 19984 12147 20036 12156
rect 19984 12113 19993 12147
rect 19993 12113 20027 12147
rect 20027 12113 20036 12147
rect 19984 12104 20036 12113
rect 20076 12104 20128 12156
rect 12440 12079 12492 12088
rect 12440 12045 12449 12079
rect 12449 12045 12483 12079
rect 12483 12045 12492 12079
rect 12440 12036 12492 12045
rect 15108 12079 15160 12088
rect 10416 11968 10468 12020
rect 15108 12045 15117 12079
rect 15117 12045 15151 12079
rect 15151 12045 15160 12079
rect 15108 12036 15160 12045
rect 15844 12036 15896 12088
rect 17408 12036 17460 12088
rect 17684 12011 17736 12020
rect 8668 11900 8720 11952
rect 13820 11943 13872 11952
rect 13820 11909 13829 11943
rect 13829 11909 13863 11943
rect 13863 11909 13872 11943
rect 13820 11900 13872 11909
rect 17684 11977 17693 12011
rect 17693 11977 17727 12011
rect 17727 11977 17736 12011
rect 17684 11968 17736 11977
rect 18696 11900 18748 11952
rect 4414 11798 4466 11850
rect 4478 11798 4530 11850
rect 4542 11798 4594 11850
rect 4606 11798 4658 11850
rect 11278 11798 11330 11850
rect 11342 11798 11394 11850
rect 11406 11798 11458 11850
rect 11470 11798 11522 11850
rect 18142 11798 18194 11850
rect 18206 11798 18258 11850
rect 18270 11798 18322 11850
rect 18334 11798 18386 11850
rect 7748 11696 7800 11748
rect 12440 11696 12492 11748
rect 13084 11696 13136 11748
rect 14556 11696 14608 11748
rect 18604 11739 18656 11748
rect 18604 11705 18613 11739
rect 18613 11705 18647 11739
rect 18647 11705 18656 11739
rect 18604 11696 18656 11705
rect 20168 11696 20220 11748
rect 11060 11628 11112 11680
rect 7380 11560 7432 11612
rect 8208 11560 8260 11612
rect 13820 11560 13872 11612
rect 16304 11628 16356 11680
rect 17040 11560 17092 11612
rect 8668 11492 8720 11544
rect 11060 11535 11112 11544
rect 11060 11501 11069 11535
rect 11069 11501 11103 11535
rect 11103 11501 11112 11535
rect 11060 11492 11112 11501
rect 13912 11492 13964 11544
rect 9680 11424 9732 11476
rect 20076 11492 20128 11544
rect 20260 11535 20312 11544
rect 20260 11501 20269 11535
rect 20269 11501 20303 11535
rect 20303 11501 20312 11535
rect 20260 11492 20312 11501
rect 16028 11424 16080 11476
rect 16396 11424 16448 11476
rect 14556 11399 14608 11408
rect 14556 11365 14565 11399
rect 14565 11365 14599 11399
rect 14599 11365 14608 11399
rect 14556 11356 14608 11365
rect 15200 11356 15252 11408
rect 16120 11399 16172 11408
rect 16120 11365 16129 11399
rect 16129 11365 16163 11399
rect 16163 11365 16172 11399
rect 16120 11356 16172 11365
rect 19156 11356 19208 11408
rect 7846 11254 7898 11306
rect 7910 11254 7962 11306
rect 7974 11254 8026 11306
rect 8038 11254 8090 11306
rect 14710 11254 14762 11306
rect 14774 11254 14826 11306
rect 14838 11254 14890 11306
rect 14902 11254 14954 11306
rect 16120 11152 16172 11204
rect 19156 11195 19208 11204
rect 19156 11161 19165 11195
rect 19165 11161 19199 11195
rect 19199 11161 19208 11195
rect 19156 11152 19208 11161
rect 20628 11152 20680 11204
rect 9036 11016 9088 11068
rect 16764 11059 16816 11068
rect 16764 11025 16773 11059
rect 16773 11025 16807 11059
rect 16807 11025 16816 11059
rect 16764 11016 16816 11025
rect 17776 11016 17828 11068
rect 20536 11059 20588 11068
rect 20536 11025 20545 11059
rect 20545 11025 20579 11059
rect 20579 11025 20588 11059
rect 20536 11016 20588 11025
rect 17040 10991 17092 11000
rect 17040 10957 17049 10991
rect 17049 10957 17083 10991
rect 17083 10957 17092 10991
rect 17040 10948 17092 10957
rect 17224 10948 17276 11000
rect 17868 10948 17920 11000
rect 19800 10991 19852 11000
rect 19800 10957 19809 10991
rect 19809 10957 19843 10991
rect 19843 10957 19852 10991
rect 19800 10948 19852 10957
rect 8300 10880 8352 10932
rect 17408 10880 17460 10932
rect 4414 10710 4466 10762
rect 4478 10710 4530 10762
rect 4542 10710 4594 10762
rect 4606 10710 4658 10762
rect 11278 10710 11330 10762
rect 11342 10710 11394 10762
rect 11406 10710 11458 10762
rect 11470 10710 11522 10762
rect 18142 10710 18194 10762
rect 18206 10710 18258 10762
rect 18270 10710 18322 10762
rect 18334 10710 18386 10762
rect 1676 10608 1728 10660
rect 8208 10608 8260 10660
rect 11060 10608 11112 10660
rect 14464 10651 14516 10660
rect 14464 10617 14473 10651
rect 14473 10617 14507 10651
rect 14507 10617 14516 10651
rect 14464 10608 14516 10617
rect 16764 10608 16816 10660
rect 18512 10651 18564 10660
rect 18512 10617 18521 10651
rect 18521 10617 18555 10651
rect 18555 10617 18564 10651
rect 18512 10608 18564 10617
rect 19616 10608 19668 10660
rect 11980 10515 12032 10524
rect 11980 10481 11989 10515
rect 11989 10481 12023 10515
rect 12023 10481 12032 10515
rect 11980 10472 12032 10481
rect 13084 10515 13136 10524
rect 13084 10481 13093 10515
rect 13093 10481 13127 10515
rect 13127 10481 13136 10515
rect 13084 10472 13136 10481
rect 11244 10404 11296 10456
rect 13820 10404 13872 10456
rect 16304 10404 16356 10456
rect 19340 10472 19392 10524
rect 19800 10404 19852 10456
rect 20260 10447 20312 10456
rect 20260 10413 20269 10447
rect 20269 10413 20303 10447
rect 20303 10413 20312 10447
rect 20260 10404 20312 10413
rect 6828 10336 6880 10388
rect 8208 10336 8260 10388
rect 16028 10336 16080 10388
rect 16856 10379 16908 10388
rect 16856 10345 16865 10379
rect 16865 10345 16899 10379
rect 16899 10345 16908 10379
rect 16856 10336 16908 10345
rect 10692 10311 10744 10320
rect 10692 10277 10701 10311
rect 10701 10277 10735 10311
rect 10735 10277 10744 10311
rect 10692 10268 10744 10277
rect 11152 10268 11204 10320
rect 11336 10311 11388 10320
rect 11336 10277 11345 10311
rect 11345 10277 11379 10311
rect 11379 10277 11388 10311
rect 11336 10268 11388 10277
rect 16948 10311 17000 10320
rect 16948 10277 16957 10311
rect 16957 10277 16991 10311
rect 16991 10277 17000 10311
rect 16948 10268 17000 10277
rect 18236 10268 18288 10320
rect 18972 10311 19024 10320
rect 18972 10277 18981 10311
rect 18981 10277 19015 10311
rect 19015 10277 19024 10311
rect 18972 10268 19024 10277
rect 7846 10166 7898 10218
rect 7910 10166 7962 10218
rect 7974 10166 8026 10218
rect 8038 10166 8090 10218
rect 14710 10166 14762 10218
rect 14774 10166 14826 10218
rect 14838 10166 14890 10218
rect 14902 10166 14954 10218
rect 11244 10107 11296 10116
rect 11244 10073 11253 10107
rect 11253 10073 11287 10107
rect 11287 10073 11296 10107
rect 11244 10064 11296 10073
rect 11336 10064 11388 10116
rect 11796 9996 11848 10048
rect 11980 9996 12032 10048
rect 17040 10064 17092 10116
rect 18236 10107 18288 10116
rect 18236 10073 18245 10107
rect 18245 10073 18279 10107
rect 18279 10073 18288 10107
rect 18236 10064 18288 10073
rect 19800 10064 19852 10116
rect 21180 10064 21232 10116
rect 16304 10039 16356 10048
rect 16304 10005 16338 10039
rect 16338 10005 16356 10039
rect 16304 9996 16356 10005
rect 8208 9903 8260 9912
rect 8208 9869 8217 9903
rect 8217 9869 8251 9903
rect 8251 9869 8260 9903
rect 8208 9860 8260 9869
rect 12808 9971 12860 9980
rect 12808 9937 12817 9971
rect 12817 9937 12851 9971
rect 12851 9937 12860 9971
rect 12808 9928 12860 9937
rect 13084 9928 13136 9980
rect 8208 9724 8260 9776
rect 11612 9860 11664 9912
rect 11704 9860 11756 9912
rect 11152 9792 11204 9844
rect 14464 9928 14516 9980
rect 14096 9724 14148 9776
rect 15844 9860 15896 9912
rect 19340 9928 19392 9980
rect 20536 9971 20588 9980
rect 20536 9937 20545 9971
rect 20545 9937 20579 9971
rect 20579 9937 20588 9971
rect 20536 9928 20588 9937
rect 4414 9622 4466 9674
rect 4478 9622 4530 9674
rect 4542 9622 4594 9674
rect 4606 9622 4658 9674
rect 11278 9622 11330 9674
rect 11342 9622 11394 9674
rect 11406 9622 11458 9674
rect 11470 9622 11522 9674
rect 18142 9622 18194 9674
rect 18206 9622 18258 9674
rect 18270 9622 18322 9674
rect 18334 9622 18386 9674
rect 18972 9520 19024 9572
rect 12808 9452 12860 9504
rect 13636 9452 13688 9504
rect 15016 9452 15068 9504
rect 20352 9452 20404 9504
rect 11796 9427 11848 9436
rect 11796 9393 11805 9427
rect 11805 9393 11839 9427
rect 11839 9393 11848 9427
rect 11796 9384 11848 9393
rect 12072 9316 12124 9368
rect 17776 9384 17828 9436
rect 19432 9384 19484 9436
rect 13452 9316 13504 9368
rect 15568 9316 15620 9368
rect 18788 9359 18840 9368
rect 18788 9325 18797 9359
rect 18797 9325 18831 9359
rect 18831 9325 18840 9359
rect 18788 9316 18840 9325
rect 20260 9359 20312 9368
rect 20260 9325 20269 9359
rect 20269 9325 20303 9359
rect 20303 9325 20312 9359
rect 20260 9316 20312 9325
rect 11888 9248 11940 9300
rect 16856 9248 16908 9300
rect 16948 9248 17000 9300
rect 19064 9248 19116 9300
rect 12532 9223 12584 9232
rect 12532 9189 12541 9223
rect 12541 9189 12575 9223
rect 12575 9189 12584 9223
rect 12532 9180 12584 9189
rect 17868 9180 17920 9232
rect 18880 9223 18932 9232
rect 18880 9189 18889 9223
rect 18889 9189 18923 9223
rect 18923 9189 18932 9223
rect 18880 9180 18932 9189
rect 7846 9078 7898 9130
rect 7910 9078 7962 9130
rect 7974 9078 8026 9130
rect 8038 9078 8090 9130
rect 14710 9078 14762 9130
rect 14774 9078 14826 9130
rect 14838 9078 14890 9130
rect 14902 9078 14954 9130
rect 10692 8976 10744 9028
rect 11612 8976 11664 9028
rect 12072 8976 12124 9028
rect 12532 8908 12584 8960
rect 15568 8951 15620 8960
rect 15568 8917 15577 8951
rect 15577 8917 15611 8951
rect 15611 8917 15620 8951
rect 15568 8908 15620 8917
rect 16212 8976 16264 9028
rect 16120 8840 16172 8892
rect 16856 8908 16908 8960
rect 18788 8908 18840 8960
rect 16948 8840 17000 8892
rect 20536 8883 20588 8892
rect 20536 8849 20545 8883
rect 20545 8849 20579 8883
rect 20579 8849 20588 8883
rect 20536 8840 20588 8849
rect 11704 8772 11756 8824
rect 4414 8534 4466 8586
rect 4478 8534 4530 8586
rect 4542 8534 4594 8586
rect 4606 8534 4658 8586
rect 11278 8534 11330 8586
rect 11342 8534 11394 8586
rect 11406 8534 11458 8586
rect 11470 8534 11522 8586
rect 18142 8534 18194 8586
rect 18206 8534 18258 8586
rect 18270 8534 18322 8586
rect 18334 8534 18386 8586
rect 11060 8432 11112 8484
rect 16120 8475 16172 8484
rect 16120 8441 16129 8475
rect 16129 8441 16163 8475
rect 16163 8441 16172 8475
rect 16120 8432 16172 8441
rect 19340 8432 19392 8484
rect 19524 8364 19576 8416
rect 13452 8339 13504 8348
rect 13452 8305 13461 8339
rect 13461 8305 13495 8339
rect 13495 8305 13504 8339
rect 13452 8296 13504 8305
rect 17224 8296 17276 8348
rect 11244 8271 11296 8280
rect 11244 8237 11253 8271
rect 11253 8237 11287 8271
rect 11287 8237 11296 8271
rect 11244 8228 11296 8237
rect 13176 8271 13228 8280
rect 13176 8237 13185 8271
rect 13185 8237 13219 8271
rect 13219 8237 13228 8271
rect 13176 8228 13228 8237
rect 18052 8228 18104 8280
rect 20260 8271 20312 8280
rect 20260 8237 20269 8271
rect 20269 8237 20303 8271
rect 20303 8237 20312 8271
rect 20260 8228 20312 8237
rect 19432 8160 19484 8212
rect 13912 8135 13964 8144
rect 13912 8101 13921 8135
rect 13921 8101 13955 8135
rect 13955 8101 13964 8135
rect 13912 8092 13964 8101
rect 16580 8135 16632 8144
rect 16580 8101 16589 8135
rect 16589 8101 16623 8135
rect 16623 8101 16632 8135
rect 16580 8092 16632 8101
rect 7846 7990 7898 8042
rect 7910 7990 7962 8042
rect 7974 7990 8026 8042
rect 8038 7990 8090 8042
rect 14710 7990 14762 8042
rect 14774 7990 14826 8042
rect 14838 7990 14890 8042
rect 14902 7990 14954 8042
rect 13176 7931 13228 7940
rect 13176 7897 13185 7931
rect 13185 7897 13219 7931
rect 13219 7897 13228 7931
rect 13176 7888 13228 7897
rect 13912 7888 13964 7940
rect 14188 7888 14240 7940
rect 19432 7931 19484 7940
rect 11244 7820 11296 7872
rect 9312 7795 9364 7804
rect 9312 7761 9346 7795
rect 9346 7761 9364 7795
rect 9312 7752 9364 7761
rect 10692 7795 10744 7804
rect 10692 7761 10701 7795
rect 10701 7761 10735 7795
rect 10735 7761 10744 7795
rect 10692 7752 10744 7761
rect 7472 7684 7524 7736
rect 8208 7684 8260 7736
rect 10324 7684 10376 7736
rect 13636 7727 13688 7736
rect 13636 7693 13645 7727
rect 13645 7693 13679 7727
rect 13679 7693 13688 7727
rect 13636 7684 13688 7693
rect 14004 7752 14056 7804
rect 16120 7795 16172 7804
rect 14096 7684 14148 7736
rect 10508 7548 10560 7600
rect 16120 7761 16154 7795
rect 16154 7761 16172 7795
rect 16120 7752 16172 7761
rect 17224 7820 17276 7872
rect 19432 7897 19441 7931
rect 19441 7897 19475 7931
rect 19475 7897 19484 7931
rect 19432 7888 19484 7897
rect 18052 7795 18104 7804
rect 18052 7761 18061 7795
rect 18061 7761 18095 7795
rect 18095 7761 18104 7795
rect 18052 7752 18104 7761
rect 19984 7795 20036 7804
rect 19984 7761 19993 7795
rect 19993 7761 20027 7795
rect 20027 7761 20036 7795
rect 19984 7752 20036 7761
rect 20536 7795 20588 7804
rect 20536 7761 20545 7795
rect 20545 7761 20579 7795
rect 20579 7761 20588 7795
rect 20536 7752 20588 7761
rect 17224 7659 17276 7668
rect 17224 7625 17233 7659
rect 17233 7625 17267 7659
rect 17267 7625 17276 7659
rect 17224 7616 17276 7625
rect 16488 7548 16540 7600
rect 4414 7446 4466 7498
rect 4478 7446 4530 7498
rect 4542 7446 4594 7498
rect 4606 7446 4658 7498
rect 11278 7446 11330 7498
rect 11342 7446 11394 7498
rect 11406 7446 11458 7498
rect 11470 7446 11522 7498
rect 18142 7446 18194 7498
rect 18206 7446 18258 7498
rect 18270 7446 18322 7498
rect 18334 7446 18386 7498
rect 10692 7344 10744 7396
rect 14004 7387 14056 7396
rect 14004 7353 14013 7387
rect 14013 7353 14047 7387
rect 14047 7353 14056 7387
rect 14004 7344 14056 7353
rect 16580 7387 16632 7396
rect 16580 7353 16589 7387
rect 16589 7353 16623 7387
rect 16623 7353 16632 7387
rect 16580 7344 16632 7353
rect 10508 7251 10560 7260
rect 10508 7217 10517 7251
rect 10517 7217 10551 7251
rect 10551 7217 10560 7251
rect 10508 7208 10560 7217
rect 16120 7208 16172 7260
rect 10324 7183 10376 7192
rect 10324 7149 10333 7183
rect 10333 7149 10367 7183
rect 10367 7149 10376 7183
rect 10324 7140 10376 7149
rect 14096 7140 14148 7192
rect 14188 7140 14240 7192
rect 18880 7140 18932 7192
rect 10416 7047 10468 7056
rect 10416 7013 10425 7047
rect 10425 7013 10459 7047
rect 10459 7013 10468 7047
rect 14372 7072 14424 7124
rect 18604 7072 18656 7124
rect 10416 7004 10468 7013
rect 17960 7004 18012 7056
rect 18880 7004 18932 7056
rect 7846 6902 7898 6954
rect 7910 6902 7962 6954
rect 7974 6902 8026 6954
rect 8038 6902 8090 6954
rect 14710 6902 14762 6954
rect 14774 6902 14826 6954
rect 14838 6902 14890 6954
rect 14902 6902 14954 6954
rect 10416 6800 10468 6852
rect 13636 6843 13688 6852
rect 13636 6809 13645 6843
rect 13645 6809 13679 6843
rect 13679 6809 13688 6843
rect 13636 6800 13688 6809
rect 16488 6800 16540 6852
rect 3608 6664 3660 6716
rect 10784 6664 10836 6716
rect 7472 6639 7524 6648
rect 7472 6605 7481 6639
rect 7481 6605 7515 6639
rect 7515 6605 7524 6639
rect 7472 6596 7524 6605
rect 18512 6664 18564 6716
rect 14096 6639 14148 6648
rect 9312 6528 9364 6580
rect 14096 6605 14105 6639
rect 14105 6605 14139 6639
rect 14139 6605 14148 6639
rect 14096 6596 14148 6605
rect 14372 6596 14424 6648
rect 4414 6358 4466 6410
rect 4478 6358 4530 6410
rect 4542 6358 4594 6410
rect 4606 6358 4658 6410
rect 11278 6358 11330 6410
rect 11342 6358 11394 6410
rect 11406 6358 11458 6410
rect 11470 6358 11522 6410
rect 18142 6358 18194 6410
rect 18206 6358 18258 6410
rect 18270 6358 18322 6410
rect 18334 6358 18386 6410
rect 14280 6256 14332 6308
rect 17960 6052 18012 6104
rect 7846 5814 7898 5866
rect 7910 5814 7962 5866
rect 7974 5814 8026 5866
rect 8038 5814 8090 5866
rect 14710 5814 14762 5866
rect 14774 5814 14826 5866
rect 14838 5814 14890 5866
rect 14902 5814 14954 5866
rect 12992 5712 13044 5764
rect 13820 5576 13872 5628
rect 4414 5270 4466 5322
rect 4478 5270 4530 5322
rect 4542 5270 4594 5322
rect 4606 5270 4658 5322
rect 11278 5270 11330 5322
rect 11342 5270 11394 5322
rect 11406 5270 11458 5322
rect 11470 5270 11522 5322
rect 18142 5270 18194 5322
rect 18206 5270 18258 5322
rect 18270 5270 18322 5322
rect 18334 5270 18386 5322
rect 13820 5168 13872 5220
rect 17960 5168 18012 5220
rect 16488 5100 16540 5152
rect 18052 5100 18104 5152
rect 7846 4726 7898 4778
rect 7910 4726 7962 4778
rect 7974 4726 8026 4778
rect 8038 4726 8090 4778
rect 14710 4726 14762 4778
rect 14774 4726 14826 4778
rect 14838 4726 14890 4778
rect 14902 4726 14954 4778
rect 20996 4624 21048 4676
rect 20536 4531 20588 4540
rect 20536 4497 20545 4531
rect 20545 4497 20579 4531
rect 20579 4497 20588 4531
rect 20536 4488 20588 4497
rect 4414 4182 4466 4234
rect 4478 4182 4530 4234
rect 4542 4182 4594 4234
rect 4606 4182 4658 4234
rect 11278 4182 11330 4234
rect 11342 4182 11394 4234
rect 11406 4182 11458 4234
rect 11470 4182 11522 4234
rect 18142 4182 18194 4234
rect 18206 4182 18258 4234
rect 18270 4182 18322 4234
rect 18334 4182 18386 4234
rect 14556 3944 14608 3996
rect 18512 3944 18564 3996
rect 7846 3638 7898 3690
rect 7910 3638 7962 3690
rect 7974 3638 8026 3690
rect 8038 3638 8090 3690
rect 14710 3638 14762 3690
rect 14774 3638 14826 3690
rect 14838 3638 14890 3690
rect 14902 3638 14954 3690
rect 4414 3094 4466 3146
rect 4478 3094 4530 3146
rect 4542 3094 4594 3146
rect 4606 3094 4658 3146
rect 11278 3094 11330 3146
rect 11342 3094 11394 3146
rect 11406 3094 11458 3146
rect 11470 3094 11522 3146
rect 18142 3094 18194 3146
rect 18206 3094 18258 3146
rect 18270 3094 18322 3146
rect 18334 3094 18386 3146
rect 7846 2550 7898 2602
rect 7910 2550 7962 2602
rect 7974 2550 8026 2602
rect 8038 2550 8090 2602
rect 14710 2550 14762 2602
rect 14774 2550 14826 2602
rect 14838 2550 14890 2602
rect 14902 2550 14954 2602
rect 4414 2006 4466 2058
rect 4478 2006 4530 2058
rect 4542 2006 4594 2058
rect 4606 2006 4658 2058
rect 11278 2006 11330 2058
rect 11342 2006 11394 2058
rect 11406 2006 11458 2058
rect 11470 2006 11522 2058
rect 18142 2006 18194 2058
rect 18206 2006 18258 2058
rect 18270 2006 18322 2058
rect 18334 2006 18386 2058
rect 16028 1156 16080 1208
rect 18144 1156 18196 1208
<< metal2 >>
rect 294 22176 350 22656
rect 846 22176 902 22656
rect 1398 22176 1454 22656
rect 1950 22176 2006 22656
rect 2502 22176 2558 22656
rect 3054 22176 3110 22656
rect 3606 22176 3662 22656
rect 4158 22176 4214 22656
rect 4710 22176 4766 22656
rect 5262 22176 5318 22656
rect 5814 22176 5870 22656
rect 6366 22176 6422 22656
rect 6918 22176 6974 22656
rect 7470 22176 7526 22656
rect 8022 22176 8078 22656
rect 8574 22176 8630 22656
rect 9126 22176 9182 22656
rect 9678 22176 9734 22656
rect 10230 22176 10286 22656
rect 10782 22176 10838 22656
rect 11334 22176 11390 22656
rect 11978 22176 12034 22656
rect 12530 22176 12586 22656
rect 13082 22176 13138 22656
rect 13634 22176 13690 22656
rect 14186 22176 14242 22656
rect 14738 22176 14794 22656
rect 15290 22176 15346 22656
rect 15842 22176 15898 22656
rect 16394 22176 16450 22656
rect 16946 22176 17002 22656
rect 17498 22176 17554 22656
rect 17958 22392 18014 22401
rect 17958 22327 18014 22336
rect 308 18758 336 22176
rect 296 18752 348 18758
rect 296 18694 348 18700
rect 860 12706 888 22176
rect 1412 17210 1440 22176
rect 1584 18616 1636 18622
rect 1584 18558 1636 18564
rect 1596 17602 1624 18558
rect 1964 18282 1992 22176
rect 2412 19160 2464 19166
rect 2412 19102 2464 19108
rect 2424 18622 2452 19102
rect 2412 18616 2464 18622
rect 2412 18558 2464 18564
rect 1952 18276 2004 18282
rect 1952 18218 2004 18224
rect 1584 17596 1636 17602
rect 1584 17538 1636 17544
rect 1412 17182 1716 17210
rect 1584 15896 1636 15902
rect 1584 15838 1636 15844
rect 1596 14882 1624 15838
rect 1584 14876 1636 14882
rect 1584 14818 1636 14824
rect 1596 14338 1624 14818
rect 1584 14332 1636 14338
rect 1584 14274 1636 14280
rect 848 12700 900 12706
rect 848 12642 900 12648
rect 1688 10666 1716 17182
rect 2516 15018 2544 22176
rect 2964 18684 3016 18690
rect 2964 18626 3016 18632
rect 2976 17738 3004 18626
rect 3068 18282 3096 22176
rect 3056 18276 3108 18282
rect 3056 18218 3108 18224
rect 3620 18078 3648 22176
rect 3608 18072 3660 18078
rect 3608 18014 3660 18020
rect 2964 17732 3016 17738
rect 2964 17674 3016 17680
rect 2976 17058 3004 17674
rect 3148 17596 3200 17602
rect 3148 17538 3200 17544
rect 3160 17126 3188 17538
rect 3332 17528 3384 17534
rect 3332 17470 3384 17476
rect 3148 17120 3200 17126
rect 3148 17062 3200 17068
rect 2964 17052 3016 17058
rect 2964 16994 3016 17000
rect 2964 16848 3016 16854
rect 2964 16790 3016 16796
rect 2976 16514 3004 16790
rect 2964 16508 3016 16514
rect 2964 16450 3016 16456
rect 3160 16106 3188 17062
rect 3344 16990 3372 17470
rect 4172 17058 4200 22176
rect 4724 19914 4752 22176
rect 4712 19908 4764 19914
rect 4712 19850 4764 19856
rect 4712 19704 4764 19710
rect 4712 19646 4764 19652
rect 4388 19468 4684 19488
rect 4444 19466 4468 19468
rect 4524 19466 4548 19468
rect 4604 19466 4628 19468
rect 4466 19414 4468 19466
rect 4530 19414 4542 19466
rect 4604 19414 4606 19466
rect 4444 19412 4468 19414
rect 4524 19412 4548 19414
rect 4604 19412 4628 19414
rect 4388 19392 4684 19412
rect 4724 19166 4752 19646
rect 5172 19568 5224 19574
rect 5172 19510 5224 19516
rect 4712 19160 4764 19166
rect 4712 19102 4764 19108
rect 4724 18826 4752 19102
rect 5080 19092 5132 19098
rect 5080 19034 5132 19040
rect 4712 18820 4764 18826
rect 4712 18762 4764 18768
rect 5092 18554 5120 19034
rect 5184 18826 5212 19510
rect 5276 19114 5304 22176
rect 5276 19086 5580 19114
rect 5448 19024 5500 19030
rect 5448 18966 5500 18972
rect 5172 18820 5224 18826
rect 5172 18762 5224 18768
rect 5460 18622 5488 18966
rect 5448 18616 5500 18622
rect 5448 18558 5500 18564
rect 5080 18548 5132 18554
rect 5080 18490 5132 18496
rect 4388 18380 4684 18400
rect 4444 18378 4468 18380
rect 4524 18378 4548 18380
rect 4604 18378 4628 18380
rect 4466 18326 4468 18378
rect 4530 18326 4542 18378
rect 4604 18326 4606 18378
rect 4444 18324 4468 18326
rect 4524 18324 4548 18326
rect 4604 18324 4628 18326
rect 4388 18304 4684 18324
rect 4252 18072 4304 18078
rect 4252 18014 4304 18020
rect 4160 17052 4212 17058
rect 4160 16994 4212 17000
rect 3332 16984 3384 16990
rect 3332 16926 3384 16932
rect 3148 16100 3200 16106
rect 3148 16042 3200 16048
rect 2964 15828 3016 15834
rect 2964 15770 3016 15776
rect 2976 15358 3004 15770
rect 2964 15352 3016 15358
rect 2964 15294 3016 15300
rect 3424 15352 3476 15358
rect 3424 15294 3476 15300
rect 2976 15018 3004 15294
rect 3436 15018 3464 15294
rect 2504 15012 2556 15018
rect 2504 14954 2556 14960
rect 2964 15012 3016 15018
rect 2964 14954 3016 14960
rect 3424 15012 3476 15018
rect 3424 14954 3476 14960
rect 3700 14876 3752 14882
rect 3700 14818 3752 14824
rect 3712 14746 3740 14818
rect 4264 14814 4292 18014
rect 5092 17534 5120 18490
rect 5172 18480 5224 18486
rect 5172 18422 5224 18428
rect 5184 18078 5212 18422
rect 5356 18276 5408 18282
rect 5356 18218 5408 18224
rect 5172 18072 5224 18078
rect 5172 18014 5224 18020
rect 5264 18004 5316 18010
rect 5264 17946 5316 17952
rect 5276 17738 5304 17946
rect 5264 17732 5316 17738
rect 5264 17674 5316 17680
rect 5080 17528 5132 17534
rect 5080 17470 5132 17476
rect 4388 17292 4684 17312
rect 4444 17290 4468 17292
rect 4524 17290 4548 17292
rect 4604 17290 4628 17292
rect 4466 17238 4468 17290
rect 4530 17238 4542 17290
rect 4604 17238 4606 17290
rect 4444 17236 4468 17238
rect 4524 17236 4548 17238
rect 4604 17236 4628 17238
rect 4388 17216 4684 17236
rect 4388 16204 4684 16224
rect 4444 16202 4468 16204
rect 4524 16202 4548 16204
rect 4604 16202 4628 16204
rect 4466 16150 4468 16202
rect 4530 16150 4542 16202
rect 4604 16150 4606 16202
rect 4444 16148 4468 16150
rect 4524 16148 4548 16150
rect 4604 16148 4628 16150
rect 4388 16128 4684 16148
rect 5092 15970 5120 17470
rect 5080 15964 5132 15970
rect 5080 15906 5132 15912
rect 5092 15442 5120 15906
rect 5000 15426 5120 15442
rect 4988 15420 5120 15426
rect 5040 15414 5120 15420
rect 4988 15362 5040 15368
rect 4388 15116 4684 15136
rect 4444 15114 4468 15116
rect 4524 15114 4548 15116
rect 4604 15114 4628 15116
rect 4466 15062 4468 15114
rect 4530 15062 4542 15114
rect 4604 15062 4606 15114
rect 4444 15060 4468 15062
rect 4524 15060 4548 15062
rect 4604 15060 4628 15062
rect 4388 15040 4684 15060
rect 4252 14808 4304 14814
rect 4252 14750 4304 14756
rect 3700 14740 3752 14746
rect 3700 14682 3752 14688
rect 2320 14332 2372 14338
rect 2320 14274 2372 14280
rect 2332 13794 2360 14274
rect 3712 13930 3740 14682
rect 5092 14678 5120 15414
rect 5080 14672 5132 14678
rect 5080 14614 5132 14620
rect 5092 14338 5120 14614
rect 5368 14474 5396 18218
rect 5460 17670 5488 18558
rect 5448 17664 5500 17670
rect 5448 17606 5500 17612
rect 5552 17058 5580 19086
rect 5828 18214 5856 22176
rect 6380 18826 6408 22176
rect 6736 19092 6788 19098
rect 6736 19034 6788 19040
rect 6368 18820 6420 18826
rect 6368 18762 6420 18768
rect 6748 18758 6776 19034
rect 6736 18752 6788 18758
rect 6736 18694 6788 18700
rect 6932 18468 6960 22176
rect 7012 19160 7064 19166
rect 7012 19102 7064 19108
rect 7024 18758 7052 19102
rect 7012 18752 7064 18758
rect 7012 18694 7064 18700
rect 7380 18684 7432 18690
rect 7380 18626 7432 18632
rect 7012 18480 7064 18486
rect 6932 18440 7012 18468
rect 7012 18422 7064 18428
rect 5724 18208 5776 18214
rect 5724 18150 5776 18156
rect 5816 18208 5868 18214
rect 5816 18150 5868 18156
rect 5632 17664 5684 17670
rect 5632 17606 5684 17612
rect 5540 17052 5592 17058
rect 5540 16994 5592 17000
rect 5644 16514 5672 17606
rect 5632 16508 5684 16514
rect 5632 16450 5684 16456
rect 5356 14468 5408 14474
rect 5356 14410 5408 14416
rect 4896 14332 4948 14338
rect 4896 14274 4948 14280
rect 5080 14332 5132 14338
rect 5080 14274 5132 14280
rect 4388 14028 4684 14048
rect 4444 14026 4468 14028
rect 4524 14026 4548 14028
rect 4604 14026 4628 14028
rect 4466 13974 4468 14026
rect 4530 13974 4542 14026
rect 4604 13974 4606 14026
rect 4444 13972 4468 13974
rect 4524 13972 4548 13974
rect 4604 13972 4628 13974
rect 4388 13952 4684 13972
rect 3700 13924 3752 13930
rect 3700 13866 3752 13872
rect 2320 13788 2372 13794
rect 2320 13730 2372 13736
rect 4908 13726 4936 14274
rect 5080 14196 5132 14202
rect 5080 14138 5132 14144
rect 5092 13726 5120 14138
rect 4896 13720 4948 13726
rect 4896 13662 4948 13668
rect 5080 13720 5132 13726
rect 5080 13662 5132 13668
rect 4388 12940 4684 12960
rect 4444 12938 4468 12940
rect 4524 12938 4548 12940
rect 4604 12938 4628 12940
rect 4466 12886 4468 12938
rect 4530 12886 4542 12938
rect 4604 12886 4606 12938
rect 4444 12884 4468 12886
rect 4524 12884 4548 12886
rect 4604 12884 4628 12886
rect 4388 12864 4684 12884
rect 5736 12706 5764 18150
rect 6828 16984 6880 16990
rect 6828 16926 6880 16932
rect 6840 16650 6868 16926
rect 6828 16644 6880 16650
rect 6828 16586 6880 16592
rect 7288 16644 7340 16650
rect 7288 16586 7340 16592
rect 7300 16106 7328 16586
rect 7392 16446 7420 18626
rect 7484 18010 7512 22176
rect 8036 20202 8064 22176
rect 7760 20174 8064 20202
rect 7472 18004 7524 18010
rect 7472 17946 7524 17952
rect 7472 17528 7524 17534
rect 7472 17470 7524 17476
rect 7484 17058 7512 17470
rect 7472 17052 7524 17058
rect 7472 16994 7524 17000
rect 7380 16440 7432 16446
rect 7380 16382 7432 16388
rect 7288 16100 7340 16106
rect 7288 16042 7340 16048
rect 7392 16038 7420 16382
rect 7380 16032 7432 16038
rect 7380 15974 7432 15980
rect 7656 15964 7708 15970
rect 7656 15906 7708 15912
rect 7668 15562 7696 15906
rect 7760 15902 7788 20174
rect 7820 20012 8116 20032
rect 7876 20010 7900 20012
rect 7956 20010 7980 20012
rect 8036 20010 8060 20012
rect 7898 19958 7900 20010
rect 7962 19958 7974 20010
rect 8036 19958 8038 20010
rect 7876 19956 7900 19958
rect 7956 19956 7980 19958
rect 8036 19956 8060 19958
rect 7820 19936 8116 19956
rect 8484 19772 8536 19778
rect 8484 19714 8536 19720
rect 8300 19704 8352 19710
rect 8300 19646 8352 19652
rect 8116 19568 8168 19574
rect 8116 19510 8168 19516
rect 8128 19370 8156 19510
rect 8116 19364 8168 19370
rect 8116 19306 8168 19312
rect 8208 19092 8260 19098
rect 8208 19034 8260 19040
rect 7820 18924 8116 18944
rect 7876 18922 7900 18924
rect 7956 18922 7980 18924
rect 8036 18922 8060 18924
rect 7898 18870 7900 18922
rect 7962 18870 7974 18922
rect 8036 18870 8038 18922
rect 7876 18868 7900 18870
rect 7956 18868 7980 18870
rect 8036 18868 8060 18870
rect 7820 18848 8116 18868
rect 8220 18826 8248 19034
rect 8208 18820 8260 18826
rect 8208 18762 8260 18768
rect 8220 18146 8248 18762
rect 8312 18282 8340 19646
rect 8392 19636 8444 19642
rect 8392 19578 8444 19584
rect 8404 19030 8432 19578
rect 8496 19234 8524 19714
rect 8484 19228 8536 19234
rect 8484 19170 8536 19176
rect 8392 19024 8444 19030
rect 8392 18966 8444 18972
rect 8404 18758 8432 18966
rect 8392 18752 8444 18758
rect 8392 18694 8444 18700
rect 8300 18276 8352 18282
rect 8300 18218 8352 18224
rect 8208 18140 8260 18146
rect 8208 18082 8260 18088
rect 8588 18078 8616 22176
rect 9140 19166 9168 22176
rect 9128 19160 9180 19166
rect 9128 19102 9180 19108
rect 9692 18078 9720 22176
rect 9956 19840 10008 19846
rect 9956 19782 10008 19788
rect 9772 19092 9824 19098
rect 9772 19034 9824 19040
rect 9784 18282 9812 19034
rect 9968 19030 9996 19782
rect 9956 19024 10008 19030
rect 9956 18966 10008 18972
rect 10244 18690 10272 22176
rect 10324 20588 10376 20594
rect 10324 20530 10376 20536
rect 10232 18684 10284 18690
rect 10232 18626 10284 18632
rect 9864 18616 9916 18622
rect 9864 18558 9916 18564
rect 9772 18276 9824 18282
rect 9772 18218 9824 18224
rect 9772 18140 9824 18146
rect 9772 18082 9824 18088
rect 8576 18072 8628 18078
rect 8576 18014 8628 18020
rect 9680 18072 9732 18078
rect 9680 18014 9732 18020
rect 8484 18004 8536 18010
rect 8484 17946 8536 17952
rect 7820 17836 8116 17856
rect 7876 17834 7900 17836
rect 7956 17834 7980 17836
rect 8036 17834 8060 17836
rect 7898 17782 7900 17834
rect 7962 17782 7974 17834
rect 8036 17782 8038 17834
rect 7876 17780 7900 17782
rect 7956 17780 7980 17782
rect 8036 17780 8060 17782
rect 7820 17760 8116 17780
rect 7820 16748 8116 16768
rect 7876 16746 7900 16748
rect 7956 16746 7980 16748
rect 8036 16746 8060 16748
rect 7898 16694 7900 16746
rect 7962 16694 7974 16746
rect 8036 16694 8038 16746
rect 7876 16692 7900 16694
rect 7956 16692 7980 16694
rect 8036 16692 8060 16694
rect 7820 16672 8116 16692
rect 8208 16440 8260 16446
rect 8208 16382 8260 16388
rect 7748 15896 7800 15902
rect 7748 15838 7800 15844
rect 7748 15760 7800 15766
rect 7748 15702 7800 15708
rect 7656 15556 7708 15562
rect 7656 15498 7708 15504
rect 6828 15420 6880 15426
rect 6828 15362 6880 15368
rect 6840 15018 6868 15362
rect 6828 15012 6880 15018
rect 6828 14954 6880 14960
rect 7760 14898 7788 15702
rect 7820 15660 8116 15680
rect 7876 15658 7900 15660
rect 7956 15658 7980 15660
rect 8036 15658 8060 15660
rect 7898 15606 7900 15658
rect 7962 15606 7974 15658
rect 8036 15606 8038 15658
rect 7876 15604 7900 15606
rect 7956 15604 7980 15606
rect 8036 15604 8060 15606
rect 7820 15584 8116 15604
rect 8220 14898 8248 16382
rect 7484 14882 7788 14898
rect 7472 14876 7788 14882
rect 7524 14870 7788 14876
rect 7472 14818 7524 14824
rect 7656 14808 7708 14814
rect 7656 14750 7708 14756
rect 7012 14332 7064 14338
rect 7012 14274 7064 14280
rect 6920 14128 6972 14134
rect 6920 14070 6972 14076
rect 6932 13794 6960 14070
rect 6920 13788 6972 13794
rect 6920 13730 6972 13736
rect 7024 13658 7052 14274
rect 7668 14134 7696 14750
rect 7760 14456 7788 14870
rect 7944 14870 8248 14898
rect 7944 14814 7972 14870
rect 7932 14808 7984 14814
rect 7932 14750 7984 14756
rect 7820 14572 8116 14592
rect 7876 14570 7900 14572
rect 7956 14570 7980 14572
rect 8036 14570 8060 14572
rect 7898 14518 7900 14570
rect 7962 14518 7974 14570
rect 8036 14518 8038 14570
rect 7876 14516 7900 14518
rect 7956 14516 7980 14518
rect 8036 14516 8060 14518
rect 7820 14496 8116 14516
rect 7760 14428 7972 14456
rect 7944 14134 7972 14428
rect 8220 14218 8248 14870
rect 8220 14202 8340 14218
rect 8220 14196 8352 14202
rect 8220 14190 8300 14196
rect 8300 14138 8352 14144
rect 7656 14128 7708 14134
rect 7656 14070 7708 14076
rect 7932 14128 7984 14134
rect 7932 14070 7984 14076
rect 7012 13652 7064 13658
rect 7012 13594 7064 13600
rect 6828 13584 6880 13590
rect 6828 13526 6880 13532
rect 6840 13386 6868 13526
rect 6828 13380 6880 13386
rect 6828 13322 6880 13328
rect 5724 12700 5776 12706
rect 5724 12642 5776 12648
rect 7024 12638 7052 13594
rect 7380 12700 7432 12706
rect 7380 12642 7432 12648
rect 7012 12632 7064 12638
rect 7012 12574 7064 12580
rect 7392 12162 7420 12642
rect 7668 12230 7696 14070
rect 8496 13794 8524 17946
rect 8760 17936 8812 17942
rect 8760 17878 8812 17884
rect 8668 17392 8720 17398
rect 8668 17334 8720 17340
rect 8680 17058 8708 17334
rect 8772 17126 8800 17878
rect 9680 17460 9732 17466
rect 9680 17402 9732 17408
rect 9692 17194 9720 17402
rect 9680 17188 9732 17194
rect 9680 17130 9732 17136
rect 8760 17120 8812 17126
rect 8760 17062 8812 17068
rect 9586 17088 9642 17097
rect 8668 17052 8720 17058
rect 8668 16994 8720 17000
rect 8680 16582 8708 16994
rect 8668 16576 8720 16582
rect 8668 16518 8720 16524
rect 8668 14740 8720 14746
rect 8668 14682 8720 14688
rect 8680 14474 8708 14682
rect 8668 14468 8720 14474
rect 8668 14410 8720 14416
rect 8680 13794 8708 14410
rect 8484 13788 8536 13794
rect 8484 13730 8536 13736
rect 8668 13788 8720 13794
rect 8668 13730 8720 13736
rect 7820 13484 8116 13504
rect 7876 13482 7900 13484
rect 7956 13482 7980 13484
rect 8036 13482 8060 13484
rect 7898 13430 7900 13482
rect 7962 13430 7974 13482
rect 8036 13430 8038 13482
rect 7876 13428 7900 13430
rect 7956 13428 7980 13430
rect 8036 13428 8060 13430
rect 7820 13408 8116 13428
rect 8208 12700 8260 12706
rect 8208 12642 8260 12648
rect 7748 12496 7800 12502
rect 7748 12438 7800 12444
rect 7656 12224 7708 12230
rect 7656 12166 7708 12172
rect 7380 12156 7432 12162
rect 7380 12098 7432 12104
rect 6828 12088 6880 12094
rect 6828 12030 6880 12036
rect 4388 11852 4684 11872
rect 4444 11850 4468 11852
rect 4524 11850 4548 11852
rect 4604 11850 4628 11852
rect 4466 11798 4468 11850
rect 4530 11798 4542 11850
rect 4604 11798 4606 11850
rect 4444 11796 4468 11798
rect 4524 11796 4548 11798
rect 4604 11796 4628 11798
rect 4388 11776 4684 11796
rect 4388 10764 4684 10784
rect 4444 10762 4468 10764
rect 4524 10762 4548 10764
rect 4604 10762 4628 10764
rect 4466 10710 4468 10762
rect 4530 10710 4542 10762
rect 4604 10710 4606 10762
rect 4444 10708 4468 10710
rect 4524 10708 4548 10710
rect 4604 10708 4628 10710
rect 4388 10688 4684 10708
rect 1676 10660 1728 10666
rect 1676 10602 1728 10608
rect 6840 10394 6868 12030
rect 7392 11618 7420 12098
rect 7760 11754 7788 12438
rect 7820 12396 8116 12416
rect 7876 12394 7900 12396
rect 7956 12394 7980 12396
rect 8036 12394 8060 12396
rect 7898 12342 7900 12394
rect 7962 12342 7974 12394
rect 8036 12342 8038 12394
rect 7876 12340 7900 12342
rect 7956 12340 7980 12342
rect 8036 12340 8060 12342
rect 7820 12320 8116 12340
rect 8220 12162 8248 12642
rect 8300 12224 8352 12230
rect 8300 12166 8352 12172
rect 8208 12156 8260 12162
rect 8208 12098 8260 12104
rect 8312 12094 8340 12166
rect 8300 12088 8352 12094
rect 8772 12042 8800 17062
rect 9586 17023 9642 17032
rect 9600 16446 9628 17023
rect 9784 16854 9812 18082
rect 9772 16848 9824 16854
rect 9692 16808 9772 16836
rect 9588 16440 9640 16446
rect 9588 16382 9640 16388
rect 9404 14944 9456 14950
rect 9404 14886 9456 14892
rect 9036 14672 9088 14678
rect 9036 14614 9088 14620
rect 9048 13590 9076 14614
rect 9416 14406 9444 14886
rect 9404 14400 9456 14406
rect 9404 14342 9456 14348
rect 9036 13584 9088 13590
rect 9036 13526 9088 13532
rect 8300 12030 8352 12036
rect 7748 11748 7800 11754
rect 7748 11690 7800 11696
rect 7380 11612 7432 11618
rect 7380 11554 7432 11560
rect 8208 11612 8260 11618
rect 8208 11554 8260 11560
rect 7820 11308 8116 11328
rect 7876 11306 7900 11308
rect 7956 11306 7980 11308
rect 8036 11306 8060 11308
rect 7898 11254 7900 11306
rect 7962 11254 7974 11306
rect 8036 11254 8038 11306
rect 7876 11252 7900 11254
rect 7956 11252 7980 11254
rect 8036 11252 8060 11254
rect 7820 11232 8116 11252
rect 8220 10666 8248 11554
rect 8312 10938 8340 12030
rect 8680 12014 8800 12042
rect 8680 11958 8708 12014
rect 8668 11952 8720 11958
rect 8668 11894 8720 11900
rect 8680 11550 8708 11894
rect 8668 11544 8720 11550
rect 8668 11486 8720 11492
rect 9048 11074 9076 13526
rect 9692 12230 9720 16808
rect 9772 16790 9824 16796
rect 9876 16446 9904 18558
rect 10232 17052 10284 17058
rect 10232 16994 10284 17000
rect 10048 16848 10100 16854
rect 10048 16790 10100 16796
rect 9864 16440 9916 16446
rect 9864 16382 9916 16388
rect 10060 15970 10088 16790
rect 10244 16582 10272 16994
rect 10232 16576 10284 16582
rect 10232 16518 10284 16524
rect 10048 15964 10100 15970
rect 10048 15906 10100 15912
rect 9772 14672 9824 14678
rect 9772 14614 9824 14620
rect 10140 14672 10192 14678
rect 10140 14614 10192 14620
rect 9784 14474 9812 14614
rect 9772 14468 9824 14474
rect 9772 14410 9824 14416
rect 9956 14196 10008 14202
rect 9956 14138 10008 14144
rect 9864 13856 9916 13862
rect 9862 13824 9864 13833
rect 9916 13824 9918 13833
rect 9862 13759 9918 13768
rect 9772 13720 9824 13726
rect 9772 13662 9824 13668
rect 9784 13386 9812 13662
rect 9968 13658 9996 14138
rect 10152 13930 10180 14614
rect 10140 13924 10192 13930
rect 10140 13866 10192 13872
rect 9956 13652 10008 13658
rect 9956 13594 10008 13600
rect 9772 13380 9824 13386
rect 9772 13322 9824 13328
rect 10336 13318 10364 20530
rect 10416 19228 10468 19234
rect 10416 19170 10468 19176
rect 10428 18758 10456 19170
rect 10416 18752 10468 18758
rect 10416 18694 10468 18700
rect 10692 18276 10744 18282
rect 10692 18218 10744 18224
rect 10704 17890 10732 18218
rect 10796 18010 10824 22176
rect 11348 19658 11376 22176
rect 11072 19630 11376 19658
rect 10784 18004 10836 18010
rect 10784 17946 10836 17952
rect 10704 17862 10824 17890
rect 10416 13652 10468 13658
rect 10416 13594 10468 13600
rect 10324 13312 10376 13318
rect 10324 13254 10376 13260
rect 10428 12706 10456 13594
rect 10416 12700 10468 12706
rect 10416 12642 10468 12648
rect 10232 12496 10284 12502
rect 10232 12438 10284 12444
rect 10244 12298 10272 12438
rect 10232 12292 10284 12298
rect 10232 12234 10284 12240
rect 9680 12224 9732 12230
rect 9680 12166 9732 12172
rect 9692 11482 9720 12166
rect 10428 12026 10456 12642
rect 10416 12020 10468 12026
rect 10416 11962 10468 11968
rect 9680 11476 9732 11482
rect 9680 11418 9732 11424
rect 9036 11068 9088 11074
rect 9036 11010 9088 11016
rect 8300 10932 8352 10938
rect 8300 10874 8352 10880
rect 8208 10660 8260 10666
rect 8208 10602 8260 10608
rect 8312 10546 8340 10874
rect 8220 10518 8340 10546
rect 8220 10394 8248 10518
rect 6828 10388 6880 10394
rect 6828 10330 6880 10336
rect 8208 10388 8260 10394
rect 8208 10330 8260 10336
rect 7820 10220 8116 10240
rect 7876 10218 7900 10220
rect 7956 10218 7980 10220
rect 8036 10218 8060 10220
rect 7898 10166 7900 10218
rect 7962 10166 7974 10218
rect 8036 10166 8038 10218
rect 7876 10164 7900 10166
rect 7956 10164 7980 10166
rect 8036 10164 8060 10166
rect 7820 10144 8116 10164
rect 8220 9918 8248 10330
rect 10692 10320 10744 10326
rect 10692 10262 10744 10268
rect 8208 9912 8260 9918
rect 8208 9854 8260 9860
rect 8220 9782 8248 9854
rect 8208 9776 8260 9782
rect 8208 9718 8260 9724
rect 4388 9676 4684 9696
rect 4444 9674 4468 9676
rect 4524 9674 4548 9676
rect 4604 9674 4628 9676
rect 4466 9622 4468 9674
rect 4530 9622 4542 9674
rect 4604 9622 4606 9674
rect 4444 9620 4468 9622
rect 4524 9620 4548 9622
rect 4604 9620 4628 9622
rect 4388 9600 4684 9620
rect 7820 9132 8116 9152
rect 7876 9130 7900 9132
rect 7956 9130 7980 9132
rect 8036 9130 8060 9132
rect 7898 9078 7900 9130
rect 7962 9078 7974 9130
rect 8036 9078 8038 9130
rect 7876 9076 7900 9078
rect 7956 9076 7980 9078
rect 8036 9076 8060 9078
rect 7820 9056 8116 9076
rect 4388 8588 4684 8608
rect 4444 8586 4468 8588
rect 4524 8586 4548 8588
rect 4604 8586 4628 8588
rect 4466 8534 4468 8586
rect 4530 8534 4542 8586
rect 4604 8534 4606 8586
rect 4444 8532 4468 8534
rect 4524 8532 4548 8534
rect 4604 8532 4628 8534
rect 4388 8512 4684 8532
rect 7820 8044 8116 8064
rect 7876 8042 7900 8044
rect 7956 8042 7980 8044
rect 8036 8042 8060 8044
rect 7898 7990 7900 8042
rect 7962 7990 7974 8042
rect 8036 7990 8038 8042
rect 7876 7988 7900 7990
rect 7956 7988 7980 7990
rect 8036 7988 8060 7990
rect 7820 7968 8116 7988
rect 8220 7742 8248 9718
rect 10704 9034 10732 10262
rect 10692 9028 10744 9034
rect 10692 8970 10744 8976
rect 9312 7804 9364 7810
rect 9312 7746 9364 7752
rect 10692 7804 10744 7810
rect 10692 7746 10744 7752
rect 7472 7736 7524 7742
rect 7472 7678 7524 7684
rect 8208 7736 8260 7742
rect 8208 7678 8260 7684
rect 4388 7500 4684 7520
rect 4444 7498 4468 7500
rect 4524 7498 4548 7500
rect 4604 7498 4628 7500
rect 4466 7446 4468 7498
rect 4530 7446 4542 7498
rect 4604 7446 4606 7498
rect 4444 7444 4468 7446
rect 4524 7444 4548 7446
rect 4604 7444 4628 7446
rect 4388 7424 4684 7444
rect 3608 6716 3660 6722
rect 3608 6658 3660 6664
rect 3620 5673 3648 6658
rect 7484 6654 7512 7678
rect 7820 6956 8116 6976
rect 7876 6954 7900 6956
rect 7956 6954 7980 6956
rect 8036 6954 8060 6956
rect 7898 6902 7900 6954
rect 7962 6902 7974 6954
rect 8036 6902 8038 6954
rect 7876 6900 7900 6902
rect 7956 6900 7980 6902
rect 8036 6900 8060 6902
rect 7820 6880 8116 6900
rect 7472 6648 7524 6654
rect 7472 6590 7524 6596
rect 9324 6586 9352 7746
rect 10324 7736 10376 7742
rect 10324 7678 10376 7684
rect 10336 7198 10364 7678
rect 10508 7600 10560 7606
rect 10508 7542 10560 7548
rect 10520 7266 10548 7542
rect 10704 7402 10732 7746
rect 10692 7396 10744 7402
rect 10692 7338 10744 7344
rect 10508 7260 10560 7266
rect 10508 7202 10560 7208
rect 10324 7192 10376 7198
rect 10324 7134 10376 7140
rect 10416 7056 10468 7062
rect 10416 6998 10468 7004
rect 10428 6858 10456 6998
rect 10416 6852 10468 6858
rect 10416 6794 10468 6800
rect 10796 6722 10824 17862
rect 10968 14332 11020 14338
rect 10968 14274 11020 14280
rect 10980 13930 11008 14274
rect 10968 13924 11020 13930
rect 10968 13866 11020 13872
rect 10968 13380 11020 13386
rect 10968 13322 11020 13328
rect 10980 12638 11008 13322
rect 10968 12632 11020 12638
rect 10968 12574 11020 12580
rect 11072 11686 11100 19630
rect 11252 19468 11548 19488
rect 11308 19466 11332 19468
rect 11388 19466 11412 19468
rect 11468 19466 11492 19468
rect 11330 19414 11332 19466
rect 11394 19414 11406 19466
rect 11468 19414 11470 19466
rect 11308 19412 11332 19414
rect 11388 19412 11412 19414
rect 11468 19412 11492 19414
rect 11252 19392 11548 19412
rect 11888 19228 11940 19234
rect 11888 19170 11940 19176
rect 11244 19024 11296 19030
rect 11244 18966 11296 18972
rect 11520 19024 11572 19030
rect 11572 18984 11652 19012
rect 11520 18966 11572 18972
rect 11256 18604 11284 18966
rect 11428 18616 11480 18622
rect 11256 18576 11428 18604
rect 11428 18558 11480 18564
rect 11252 18380 11548 18400
rect 11308 18378 11332 18380
rect 11388 18378 11412 18380
rect 11468 18378 11492 18380
rect 11330 18326 11332 18378
rect 11394 18326 11406 18378
rect 11468 18326 11470 18378
rect 11308 18324 11332 18326
rect 11388 18324 11412 18326
rect 11468 18324 11492 18326
rect 11252 18304 11548 18324
rect 11624 18282 11652 18984
rect 11900 18826 11928 19170
rect 11704 18820 11756 18826
rect 11704 18762 11756 18768
rect 11888 18820 11940 18826
rect 11888 18762 11940 18768
rect 11612 18276 11664 18282
rect 11612 18218 11664 18224
rect 11520 18208 11572 18214
rect 11572 18156 11652 18162
rect 11520 18150 11652 18156
rect 11532 18134 11652 18150
rect 11152 17936 11204 17942
rect 11152 17878 11204 17884
rect 11060 11680 11112 11686
rect 11060 11622 11112 11628
rect 11060 11544 11112 11550
rect 11060 11486 11112 11492
rect 11072 10666 11100 11486
rect 11060 10660 11112 10666
rect 11060 10602 11112 10608
rect 11164 10410 11192 17878
rect 11252 17292 11548 17312
rect 11308 17290 11332 17292
rect 11388 17290 11412 17292
rect 11468 17290 11492 17292
rect 11330 17238 11332 17290
rect 11394 17238 11406 17290
rect 11468 17238 11470 17290
rect 11308 17236 11332 17238
rect 11388 17236 11412 17238
rect 11468 17236 11492 17238
rect 11252 17216 11548 17236
rect 11624 16990 11652 18134
rect 11716 17398 11744 18762
rect 11888 18616 11940 18622
rect 11888 18558 11940 18564
rect 11704 17392 11756 17398
rect 11704 17334 11756 17340
rect 11704 17052 11756 17058
rect 11704 16994 11756 17000
rect 11612 16984 11664 16990
rect 11612 16926 11664 16932
rect 11716 16650 11744 16994
rect 11704 16644 11756 16650
rect 11704 16586 11756 16592
rect 11252 16204 11548 16224
rect 11308 16202 11332 16204
rect 11388 16202 11412 16204
rect 11468 16202 11492 16204
rect 11330 16150 11332 16202
rect 11394 16150 11406 16202
rect 11468 16150 11470 16202
rect 11308 16148 11332 16150
rect 11388 16148 11412 16150
rect 11468 16148 11492 16150
rect 11252 16128 11548 16148
rect 11716 15834 11744 16586
rect 11704 15828 11756 15834
rect 11704 15770 11756 15776
rect 11252 15116 11548 15136
rect 11308 15114 11332 15116
rect 11388 15114 11412 15116
rect 11468 15114 11492 15116
rect 11330 15062 11332 15114
rect 11394 15062 11406 15114
rect 11468 15062 11470 15114
rect 11308 15060 11332 15062
rect 11388 15060 11412 15062
rect 11468 15060 11492 15062
rect 11252 15040 11548 15060
rect 11252 14028 11548 14048
rect 11308 14026 11332 14028
rect 11388 14026 11412 14028
rect 11468 14026 11492 14028
rect 11330 13974 11332 14026
rect 11394 13974 11406 14026
rect 11468 13974 11470 14026
rect 11308 13972 11332 13974
rect 11388 13972 11412 13974
rect 11468 13972 11492 13974
rect 11252 13952 11548 13972
rect 11252 12940 11548 12960
rect 11308 12938 11332 12940
rect 11388 12938 11412 12940
rect 11468 12938 11492 12940
rect 11330 12886 11332 12938
rect 11394 12886 11406 12938
rect 11468 12886 11470 12938
rect 11308 12884 11332 12886
rect 11388 12884 11412 12886
rect 11468 12884 11492 12886
rect 11252 12864 11548 12884
rect 11252 11852 11548 11872
rect 11308 11850 11332 11852
rect 11388 11850 11412 11852
rect 11468 11850 11492 11852
rect 11330 11798 11332 11850
rect 11394 11798 11406 11850
rect 11468 11798 11470 11850
rect 11308 11796 11332 11798
rect 11388 11796 11412 11798
rect 11468 11796 11492 11798
rect 11252 11776 11548 11796
rect 11252 10764 11548 10784
rect 11308 10762 11332 10764
rect 11388 10762 11412 10764
rect 11468 10762 11492 10764
rect 11330 10710 11332 10762
rect 11394 10710 11406 10762
rect 11468 10710 11470 10762
rect 11308 10708 11332 10710
rect 11388 10708 11412 10710
rect 11468 10708 11492 10710
rect 11252 10688 11548 10708
rect 11072 10382 11192 10410
rect 11244 10456 11296 10462
rect 11244 10398 11296 10404
rect 11072 8490 11100 10382
rect 11152 10320 11204 10326
rect 11152 10262 11204 10268
rect 11164 9850 11192 10262
rect 11256 10122 11284 10398
rect 11336 10320 11388 10326
rect 11336 10262 11388 10268
rect 11348 10122 11376 10262
rect 11244 10116 11296 10122
rect 11244 10058 11296 10064
rect 11336 10116 11388 10122
rect 11336 10058 11388 10064
rect 11796 10048 11848 10054
rect 11796 9990 11848 9996
rect 11612 9912 11664 9918
rect 11612 9854 11664 9860
rect 11704 9912 11756 9918
rect 11704 9854 11756 9860
rect 11152 9844 11204 9850
rect 11152 9786 11204 9792
rect 11252 9676 11548 9696
rect 11308 9674 11332 9676
rect 11388 9674 11412 9676
rect 11468 9674 11492 9676
rect 11330 9622 11332 9674
rect 11394 9622 11406 9674
rect 11468 9622 11470 9674
rect 11308 9620 11332 9622
rect 11388 9620 11412 9622
rect 11468 9620 11492 9622
rect 11252 9600 11548 9620
rect 11624 9034 11652 9854
rect 11612 9028 11664 9034
rect 11612 8970 11664 8976
rect 11716 8830 11744 9854
rect 11808 9442 11836 9990
rect 11796 9436 11848 9442
rect 11796 9378 11848 9384
rect 11900 9306 11928 18558
rect 11992 17942 12020 22176
rect 12164 19024 12216 19030
rect 12164 18966 12216 18972
rect 12440 19024 12492 19030
rect 12440 18966 12492 18972
rect 12072 18208 12124 18214
rect 12072 18150 12124 18156
rect 12084 17942 12112 18150
rect 12176 18146 12204 18966
rect 12452 18826 12480 18966
rect 12544 18826 12572 22176
rect 12624 19160 12676 19166
rect 12624 19102 12676 19108
rect 12440 18820 12492 18826
rect 12440 18762 12492 18768
rect 12532 18820 12584 18826
rect 12532 18762 12584 18768
rect 12636 18486 12664 19102
rect 12992 18820 13044 18826
rect 12992 18762 13044 18768
rect 12624 18480 12676 18486
rect 12624 18422 12676 18428
rect 12716 18480 12768 18486
rect 12716 18422 12768 18428
rect 12164 18140 12216 18146
rect 12164 18082 12216 18088
rect 11980 17936 12032 17942
rect 11980 17878 12032 17884
rect 12072 17936 12124 17942
rect 12072 17878 12124 17884
rect 12164 17732 12216 17738
rect 12164 17674 12216 17680
rect 12176 17126 12204 17674
rect 12348 17392 12400 17398
rect 12348 17334 12400 17340
rect 12360 17126 12388 17334
rect 12164 17120 12216 17126
rect 12164 17062 12216 17068
rect 12348 17120 12400 17126
rect 12348 17062 12400 17068
rect 12532 16848 12584 16854
rect 12532 16790 12584 16796
rect 12544 16650 12572 16790
rect 12532 16644 12584 16650
rect 12532 16586 12584 16592
rect 12532 16508 12584 16514
rect 12532 16450 12584 16456
rect 12544 16106 12572 16450
rect 12636 16446 12664 18422
rect 12728 18282 12756 18422
rect 12716 18276 12768 18282
rect 12716 18218 12768 18224
rect 12714 18040 12770 18049
rect 12714 17975 12716 17984
rect 12768 17975 12770 17984
rect 12716 17946 12768 17952
rect 12716 17052 12768 17058
rect 12716 16994 12768 17000
rect 12728 16514 12756 16994
rect 12716 16508 12768 16514
rect 12716 16450 12768 16456
rect 12624 16440 12676 16446
rect 12624 16382 12676 16388
rect 12636 16106 12664 16382
rect 12532 16100 12584 16106
rect 12532 16042 12584 16048
rect 12624 16100 12676 16106
rect 12624 16042 12676 16048
rect 12162 15320 12218 15329
rect 12162 15255 12218 15264
rect 12176 14950 12204 15255
rect 12164 14944 12216 14950
rect 12164 14886 12216 14892
rect 12808 14876 12860 14882
rect 12808 14818 12860 14824
rect 12256 14808 12308 14814
rect 12256 14750 12308 14756
rect 12268 14406 12296 14750
rect 12624 14672 12676 14678
rect 12624 14614 12676 14620
rect 12716 14672 12768 14678
rect 12716 14614 12768 14620
rect 12256 14400 12308 14406
rect 12256 14342 12308 14348
rect 12532 14196 12584 14202
rect 12532 14138 12584 14144
rect 12072 14128 12124 14134
rect 12072 14070 12124 14076
rect 11980 10524 12032 10530
rect 11980 10466 12032 10472
rect 11992 10054 12020 10466
rect 11980 10048 12032 10054
rect 11980 9990 12032 9996
rect 12084 9374 12112 14070
rect 12544 13930 12572 14138
rect 12636 13930 12664 14614
rect 12728 14474 12756 14614
rect 12716 14468 12768 14474
rect 12716 14410 12768 14416
rect 12820 14134 12848 14818
rect 12808 14128 12860 14134
rect 12808 14070 12860 14076
rect 12532 13924 12584 13930
rect 12532 13866 12584 13872
rect 12624 13924 12676 13930
rect 12624 13866 12676 13872
rect 12544 13794 12572 13866
rect 12532 13788 12584 13794
rect 12532 13730 12584 13736
rect 12440 12088 12492 12094
rect 12440 12030 12492 12036
rect 12452 11754 12480 12030
rect 12440 11748 12492 11754
rect 12440 11690 12492 11696
rect 12808 9980 12860 9986
rect 12808 9922 12860 9928
rect 12820 9510 12848 9922
rect 12808 9504 12860 9510
rect 12808 9446 12860 9452
rect 12072 9368 12124 9374
rect 12072 9310 12124 9316
rect 11888 9300 11940 9306
rect 11888 9242 11940 9248
rect 12084 9034 12112 9310
rect 12532 9232 12584 9238
rect 12532 9174 12584 9180
rect 12072 9028 12124 9034
rect 12072 8970 12124 8976
rect 12544 8966 12572 9174
rect 12532 8960 12584 8966
rect 12532 8902 12584 8908
rect 11704 8824 11756 8830
rect 11704 8766 11756 8772
rect 11252 8588 11548 8608
rect 11308 8586 11332 8588
rect 11388 8586 11412 8588
rect 11468 8586 11492 8588
rect 11330 8534 11332 8586
rect 11394 8534 11406 8586
rect 11468 8534 11470 8586
rect 11308 8532 11332 8534
rect 11388 8532 11412 8534
rect 11468 8532 11492 8534
rect 11252 8512 11548 8532
rect 11060 8484 11112 8490
rect 11060 8426 11112 8432
rect 11244 8280 11296 8286
rect 11244 8222 11296 8228
rect 11256 7878 11284 8222
rect 11244 7872 11296 7878
rect 11244 7814 11296 7820
rect 11252 7500 11548 7520
rect 11308 7498 11332 7500
rect 11388 7498 11412 7500
rect 11468 7498 11492 7500
rect 11330 7446 11332 7498
rect 11394 7446 11406 7498
rect 11468 7446 11470 7498
rect 11308 7444 11332 7446
rect 11388 7444 11412 7446
rect 11468 7444 11492 7446
rect 11252 7424 11548 7444
rect 10784 6716 10836 6722
rect 10784 6658 10836 6664
rect 9312 6580 9364 6586
rect 9312 6522 9364 6528
rect 4388 6412 4684 6432
rect 4444 6410 4468 6412
rect 4524 6410 4548 6412
rect 4604 6410 4628 6412
rect 4466 6358 4468 6410
rect 4530 6358 4542 6410
rect 4604 6358 4606 6410
rect 4444 6356 4468 6358
rect 4524 6356 4548 6358
rect 4604 6356 4628 6358
rect 4388 6336 4684 6356
rect 11252 6412 11548 6432
rect 11308 6410 11332 6412
rect 11388 6410 11412 6412
rect 11468 6410 11492 6412
rect 11330 6358 11332 6410
rect 11394 6358 11406 6410
rect 11468 6358 11470 6410
rect 11308 6356 11332 6358
rect 11388 6356 11412 6358
rect 11468 6356 11492 6358
rect 11252 6336 11548 6356
rect 7820 5868 8116 5888
rect 7876 5866 7900 5868
rect 7956 5866 7980 5868
rect 8036 5866 8060 5868
rect 7898 5814 7900 5866
rect 7962 5814 7974 5866
rect 8036 5814 8038 5866
rect 7876 5812 7900 5814
rect 7956 5812 7980 5814
rect 8036 5812 8060 5814
rect 7820 5792 8116 5812
rect 13004 5770 13032 18762
rect 13096 17942 13124 22176
rect 13648 18214 13676 22176
rect 14200 20338 14228 22176
rect 14108 20310 14228 20338
rect 13820 19092 13872 19098
rect 13820 19034 13872 19040
rect 13832 18826 13860 19034
rect 14108 18826 14136 20310
rect 14752 20202 14780 22176
rect 14200 20174 14780 20202
rect 13820 18820 13872 18826
rect 13820 18762 13872 18768
rect 14096 18820 14148 18826
rect 14096 18762 14148 18768
rect 13636 18208 13688 18214
rect 13636 18150 13688 18156
rect 13832 18146 13860 18762
rect 14096 18616 14148 18622
rect 14096 18558 14148 18564
rect 13820 18140 13872 18146
rect 13820 18082 13872 18088
rect 14108 18078 14136 18558
rect 14096 18072 14148 18078
rect 13358 18040 13414 18049
rect 14096 18014 14148 18020
rect 13358 17975 13360 17984
rect 13412 17975 13414 17984
rect 13360 17946 13412 17952
rect 13084 17936 13136 17942
rect 13084 17878 13136 17884
rect 13636 17936 13688 17942
rect 13636 17878 13688 17884
rect 13452 15964 13504 15970
rect 13452 15906 13504 15912
rect 13464 14678 13492 15906
rect 13452 14672 13504 14678
rect 13452 14614 13504 14620
rect 13464 14406 13492 14614
rect 13452 14400 13504 14406
rect 13452 14342 13504 14348
rect 13452 14264 13504 14270
rect 13452 14206 13504 14212
rect 13464 13726 13492 14206
rect 13452 13720 13504 13726
rect 13452 13662 13504 13668
rect 13176 13176 13228 13182
rect 13176 13118 13228 13124
rect 13188 12842 13216 13118
rect 13176 12836 13228 12842
rect 13176 12778 13228 12784
rect 13544 12836 13596 12842
rect 13544 12778 13596 12784
rect 13556 12706 13584 12778
rect 13544 12700 13596 12706
rect 13544 12642 13596 12648
rect 13084 11748 13136 11754
rect 13084 11690 13136 11696
rect 13096 10530 13124 11690
rect 13084 10524 13136 10530
rect 13084 10466 13136 10472
rect 13096 9986 13124 10466
rect 13084 9980 13136 9986
rect 13084 9922 13136 9928
rect 13648 9510 13676 17878
rect 14096 17052 14148 17058
rect 14096 16994 14148 17000
rect 14004 16848 14056 16854
rect 14004 16790 14056 16796
rect 14016 16650 14044 16790
rect 14004 16644 14056 16650
rect 14004 16586 14056 16592
rect 14108 16378 14136 16994
rect 14096 16372 14148 16378
rect 14096 16314 14148 16320
rect 14108 15902 14136 16314
rect 14096 15896 14148 15902
rect 14096 15838 14148 15844
rect 13912 14808 13964 14814
rect 13912 14750 13964 14756
rect 13820 13108 13872 13114
rect 13820 13050 13872 13056
rect 13728 12700 13780 12706
rect 13728 12642 13780 12648
rect 13740 12230 13768 12642
rect 13728 12224 13780 12230
rect 13728 12166 13780 12172
rect 13832 11958 13860 13050
rect 13924 12570 13952 14750
rect 14096 13244 14148 13250
rect 14096 13186 14148 13192
rect 13912 12564 13964 12570
rect 13912 12506 13964 12512
rect 13820 11952 13872 11958
rect 13820 11894 13872 11900
rect 13832 11618 13860 11894
rect 13820 11612 13872 11618
rect 13820 11554 13872 11560
rect 13832 10462 13860 11554
rect 13924 11550 13952 12506
rect 14108 12298 14136 13186
rect 14096 12292 14148 12298
rect 14096 12234 14148 12240
rect 13912 11544 13964 11550
rect 13912 11486 13964 11492
rect 13820 10456 13872 10462
rect 13820 10398 13872 10404
rect 14096 9776 14148 9782
rect 14096 9718 14148 9724
rect 13636 9504 13688 9510
rect 13636 9446 13688 9452
rect 13452 9368 13504 9374
rect 13452 9310 13504 9316
rect 13464 8354 13492 9310
rect 13452 8348 13504 8354
rect 13452 8290 13504 8296
rect 13176 8280 13228 8286
rect 13176 8222 13228 8228
rect 13188 7946 13216 8222
rect 13912 8144 13964 8150
rect 13912 8086 13964 8092
rect 13924 7946 13952 8086
rect 13176 7940 13228 7946
rect 13176 7882 13228 7888
rect 13912 7940 13964 7946
rect 13912 7882 13964 7888
rect 14004 7804 14056 7810
rect 14004 7746 14056 7752
rect 13636 7736 13688 7742
rect 13636 7678 13688 7684
rect 13648 6858 13676 7678
rect 14016 7402 14044 7746
rect 14108 7742 14136 9718
rect 14200 7946 14228 20174
rect 14684 20012 14980 20032
rect 14740 20010 14764 20012
rect 14820 20010 14844 20012
rect 14900 20010 14924 20012
rect 14762 19958 14764 20010
rect 14826 19958 14838 20010
rect 14900 19958 14902 20010
rect 14740 19956 14764 19958
rect 14820 19956 14844 19958
rect 14900 19956 14924 19958
rect 14684 19936 14980 19956
rect 14372 19160 14424 19166
rect 14372 19102 14424 19108
rect 14384 18690 14412 19102
rect 14464 19024 14516 19030
rect 14464 18966 14516 18972
rect 14476 18758 14504 18966
rect 14684 18924 14980 18944
rect 14740 18922 14764 18924
rect 14820 18922 14844 18924
rect 14900 18922 14924 18924
rect 14762 18870 14764 18922
rect 14826 18870 14838 18922
rect 14900 18870 14902 18922
rect 14740 18868 14764 18870
rect 14820 18868 14844 18870
rect 14900 18868 14924 18870
rect 14684 18848 14980 18868
rect 14556 18820 14608 18826
rect 14556 18762 14608 18768
rect 14464 18752 14516 18758
rect 14464 18694 14516 18700
rect 14372 18684 14424 18690
rect 14372 18626 14424 18632
rect 14280 18208 14332 18214
rect 14280 18150 14332 18156
rect 14188 7940 14240 7946
rect 14188 7882 14240 7888
rect 14096 7736 14148 7742
rect 14096 7678 14148 7684
rect 14004 7396 14056 7402
rect 14004 7338 14056 7344
rect 14108 7198 14136 7678
rect 14096 7192 14148 7198
rect 14096 7134 14148 7140
rect 14188 7192 14240 7198
rect 14188 7134 14240 7140
rect 13636 6852 13688 6858
rect 13636 6794 13688 6800
rect 14096 6648 14148 6654
rect 14200 6636 14228 7134
rect 14148 6608 14228 6636
rect 14096 6590 14148 6596
rect 14292 6314 14320 18150
rect 14476 18146 14504 18694
rect 14464 18140 14516 18146
rect 14464 18082 14516 18088
rect 14372 16848 14424 16854
rect 14372 16790 14424 16796
rect 14384 15834 14412 16790
rect 14568 16394 14596 18762
rect 15304 17942 15332 22176
rect 15384 19092 15436 19098
rect 15384 19034 15436 19040
rect 15200 17936 15252 17942
rect 15200 17878 15252 17884
rect 15292 17936 15344 17942
rect 15292 17878 15344 17884
rect 14684 17836 14980 17856
rect 14740 17834 14764 17836
rect 14820 17834 14844 17836
rect 14900 17834 14924 17836
rect 14762 17782 14764 17834
rect 14826 17782 14838 17834
rect 14900 17782 14902 17834
rect 14740 17780 14764 17782
rect 14820 17780 14844 17782
rect 14900 17780 14924 17782
rect 14684 17760 14980 17780
rect 14684 16748 14980 16768
rect 14740 16746 14764 16748
rect 14820 16746 14844 16748
rect 14900 16746 14924 16748
rect 14762 16694 14764 16746
rect 14826 16694 14838 16746
rect 14900 16694 14902 16746
rect 14740 16692 14764 16694
rect 14820 16692 14844 16694
rect 14900 16692 14924 16694
rect 14684 16672 14980 16692
rect 15108 16440 15160 16446
rect 14568 16366 15056 16394
rect 15108 16382 15160 16388
rect 14372 15828 14424 15834
rect 14372 15770 14424 15776
rect 14556 15760 14608 15766
rect 14556 15702 14608 15708
rect 14568 14406 14596 15702
rect 14684 15660 14980 15680
rect 14740 15658 14764 15660
rect 14820 15658 14844 15660
rect 14900 15658 14924 15660
rect 14762 15606 14764 15658
rect 14826 15606 14838 15658
rect 14900 15606 14902 15658
rect 14740 15604 14764 15606
rect 14820 15604 14844 15606
rect 14900 15604 14924 15606
rect 14684 15584 14980 15604
rect 14684 14572 14980 14592
rect 14740 14570 14764 14572
rect 14820 14570 14844 14572
rect 14900 14570 14924 14572
rect 14762 14518 14764 14570
rect 14826 14518 14838 14570
rect 14900 14518 14902 14570
rect 14740 14516 14764 14518
rect 14820 14516 14844 14518
rect 14900 14516 14924 14518
rect 14684 14496 14980 14516
rect 14556 14400 14608 14406
rect 14556 14342 14608 14348
rect 14372 13584 14424 13590
rect 14372 13526 14424 13532
rect 14384 12774 14412 13526
rect 14684 13484 14980 13504
rect 14740 13482 14764 13484
rect 14820 13482 14844 13484
rect 14900 13482 14924 13484
rect 14762 13430 14764 13482
rect 14826 13430 14838 13482
rect 14900 13430 14902 13482
rect 14740 13428 14764 13430
rect 14820 13428 14844 13430
rect 14900 13428 14924 13430
rect 14684 13408 14980 13428
rect 14832 13040 14884 13046
rect 14832 12982 14884 12988
rect 14372 12768 14424 12774
rect 14372 12710 14424 12716
rect 14384 12502 14412 12710
rect 14844 12706 14872 12982
rect 14740 12700 14792 12706
rect 14740 12642 14792 12648
rect 14832 12700 14884 12706
rect 14832 12642 14884 12648
rect 14752 12586 14780 12642
rect 14476 12558 14780 12586
rect 14372 12496 14424 12502
rect 14372 12438 14424 12444
rect 14476 10666 14504 12558
rect 14556 12496 14608 12502
rect 14556 12438 14608 12444
rect 14568 11754 14596 12438
rect 14684 12396 14980 12416
rect 14740 12394 14764 12396
rect 14820 12394 14844 12396
rect 14900 12394 14924 12396
rect 14762 12342 14764 12394
rect 14826 12342 14838 12394
rect 14900 12342 14902 12394
rect 14740 12340 14764 12342
rect 14820 12340 14844 12342
rect 14900 12340 14924 12342
rect 14684 12320 14980 12340
rect 14556 11748 14608 11754
rect 14556 11690 14608 11696
rect 14556 11408 14608 11414
rect 14556 11350 14608 11356
rect 14464 10660 14516 10666
rect 14464 10602 14516 10608
rect 14476 9986 14504 10602
rect 14464 9980 14516 9986
rect 14464 9922 14516 9928
rect 14372 7124 14424 7130
rect 14372 7066 14424 7072
rect 14384 6654 14412 7066
rect 14372 6648 14424 6654
rect 14372 6590 14424 6596
rect 14280 6308 14332 6314
rect 14280 6250 14332 6256
rect 12992 5764 13044 5770
rect 12992 5706 13044 5712
rect 3606 5664 3662 5673
rect 3606 5599 3662 5608
rect 13820 5628 13872 5634
rect 13820 5570 13872 5576
rect 4388 5324 4684 5344
rect 4444 5322 4468 5324
rect 4524 5322 4548 5324
rect 4604 5322 4628 5324
rect 4466 5270 4468 5322
rect 4530 5270 4542 5322
rect 4604 5270 4606 5322
rect 4444 5268 4468 5270
rect 4524 5268 4548 5270
rect 4604 5268 4628 5270
rect 4388 5248 4684 5268
rect 11252 5324 11548 5344
rect 11308 5322 11332 5324
rect 11388 5322 11412 5324
rect 11468 5322 11492 5324
rect 11330 5270 11332 5322
rect 11394 5270 11406 5322
rect 11468 5270 11470 5322
rect 11308 5268 11332 5270
rect 11388 5268 11412 5270
rect 11468 5268 11492 5270
rect 11252 5248 11548 5268
rect 13832 5226 13860 5570
rect 13820 5220 13872 5226
rect 13820 5162 13872 5168
rect 7820 4780 8116 4800
rect 7876 4778 7900 4780
rect 7956 4778 7980 4780
rect 8036 4778 8060 4780
rect 7898 4726 7900 4778
rect 7962 4726 7974 4778
rect 8036 4726 8038 4778
rect 7876 4724 7900 4726
rect 7956 4724 7980 4726
rect 8036 4724 8060 4726
rect 7820 4704 8116 4724
rect 4388 4236 4684 4256
rect 4444 4234 4468 4236
rect 4524 4234 4548 4236
rect 4604 4234 4628 4236
rect 4466 4182 4468 4234
rect 4530 4182 4542 4234
rect 4604 4182 4606 4234
rect 4444 4180 4468 4182
rect 4524 4180 4548 4182
rect 4604 4180 4628 4182
rect 4388 4160 4684 4180
rect 11252 4236 11548 4256
rect 11308 4234 11332 4236
rect 11388 4234 11412 4236
rect 11468 4234 11492 4236
rect 11330 4182 11332 4234
rect 11394 4182 11406 4234
rect 11468 4182 11470 4234
rect 11308 4180 11332 4182
rect 11388 4180 11412 4182
rect 11468 4180 11492 4182
rect 11252 4160 11548 4180
rect 14568 4002 14596 11350
rect 14684 11308 14980 11328
rect 14740 11306 14764 11308
rect 14820 11306 14844 11308
rect 14900 11306 14924 11308
rect 14762 11254 14764 11306
rect 14826 11254 14838 11306
rect 14900 11254 14902 11306
rect 14740 11252 14764 11254
rect 14820 11252 14844 11254
rect 14900 11252 14924 11254
rect 14684 11232 14980 11252
rect 14684 10220 14980 10240
rect 14740 10218 14764 10220
rect 14820 10218 14844 10220
rect 14900 10218 14924 10220
rect 14762 10166 14764 10218
rect 14826 10166 14838 10218
rect 14900 10166 14902 10218
rect 14740 10164 14764 10166
rect 14820 10164 14844 10166
rect 14900 10164 14924 10166
rect 14684 10144 14980 10164
rect 15028 9510 15056 16366
rect 15120 15766 15148 16382
rect 15212 15902 15240 17878
rect 15200 15896 15252 15902
rect 15200 15838 15252 15844
rect 15108 15760 15160 15766
rect 15108 15702 15160 15708
rect 15200 15760 15252 15766
rect 15200 15702 15252 15708
rect 15108 15284 15160 15290
rect 15108 15226 15160 15232
rect 15120 15018 15148 15226
rect 15108 15012 15160 15018
rect 15108 14954 15160 14960
rect 15108 12496 15160 12502
rect 15108 12438 15160 12444
rect 15120 12094 15148 12438
rect 15212 12162 15240 15702
rect 15396 14882 15424 19034
rect 15856 18010 15884 22176
rect 16304 19024 16356 19030
rect 16304 18966 16356 18972
rect 15936 18684 15988 18690
rect 15936 18626 15988 18632
rect 15844 18004 15896 18010
rect 15844 17946 15896 17952
rect 15948 17058 15976 18626
rect 16120 17664 16172 17670
rect 16120 17606 16172 17612
rect 16132 17398 16160 17606
rect 16316 17602 16344 18966
rect 16304 17596 16356 17602
rect 16304 17538 16356 17544
rect 16120 17392 16172 17398
rect 16120 17334 16172 17340
rect 16408 17210 16436 22176
rect 16488 19228 16540 19234
rect 16488 19170 16540 19176
rect 16500 18758 16528 19170
rect 16488 18752 16540 18758
rect 16488 18694 16540 18700
rect 16960 17942 16988 22176
rect 17224 19704 17276 19710
rect 17224 19646 17276 19652
rect 17236 19166 17264 19646
rect 17512 19386 17540 22176
rect 17972 20594 18000 22327
rect 18050 22176 18106 22656
rect 18602 22176 18658 22656
rect 19154 22176 19210 22656
rect 19706 22176 19762 22656
rect 20258 22176 20314 22656
rect 20810 22176 20866 22656
rect 21362 22176 21418 22656
rect 21914 22176 21970 22656
rect 22466 22176 22522 22656
rect 17960 20588 18012 20594
rect 17960 20530 18012 20536
rect 18064 19658 18092 22176
rect 18616 19930 18644 22176
rect 18786 21440 18842 21449
rect 18786 21375 18842 21384
rect 18616 19902 18736 19930
rect 18800 19914 18828 21375
rect 18970 21032 19026 21041
rect 18970 20967 19026 20976
rect 18604 19772 18656 19778
rect 18604 19714 18656 19720
rect 17972 19630 18092 19658
rect 17512 19358 17724 19386
rect 17500 19228 17552 19234
rect 17552 19188 17632 19216
rect 17500 19170 17552 19176
rect 17224 19160 17276 19166
rect 17224 19102 17276 19108
rect 17604 18486 17632 19188
rect 17696 18622 17724 19358
rect 17972 18826 18000 19630
rect 18116 19468 18412 19488
rect 18172 19466 18196 19468
rect 18252 19466 18276 19468
rect 18332 19466 18356 19468
rect 18194 19414 18196 19466
rect 18258 19414 18270 19466
rect 18332 19414 18334 19466
rect 18172 19412 18196 19414
rect 18252 19412 18276 19414
rect 18332 19412 18356 19414
rect 18116 19392 18412 19412
rect 18616 19234 18644 19714
rect 18604 19228 18656 19234
rect 18604 19170 18656 19176
rect 17960 18820 18012 18826
rect 17960 18762 18012 18768
rect 17960 18684 18012 18690
rect 17960 18626 18012 18632
rect 17684 18616 17736 18622
rect 17684 18558 17736 18564
rect 17592 18480 17644 18486
rect 17592 18422 17644 18428
rect 16488 17936 16540 17942
rect 16488 17878 16540 17884
rect 16948 17936 17000 17942
rect 16948 17878 17000 17884
rect 16224 17182 16436 17210
rect 15936 17052 15988 17058
rect 15936 16994 15988 17000
rect 15948 16514 15976 16994
rect 15936 16508 15988 16514
rect 15936 16450 15988 16456
rect 15948 16106 15976 16450
rect 15936 16100 15988 16106
rect 15936 16042 15988 16048
rect 15384 14876 15436 14882
rect 15384 14818 15436 14824
rect 15476 14672 15528 14678
rect 15476 14614 15528 14620
rect 15488 14474 15516 14614
rect 15476 14468 15528 14474
rect 15476 14410 15528 14416
rect 15568 13176 15620 13182
rect 15568 13118 15620 13124
rect 15580 12706 15608 13118
rect 15568 12700 15620 12706
rect 15568 12642 15620 12648
rect 16028 12632 16080 12638
rect 16028 12574 16080 12580
rect 16040 12178 16068 12574
rect 15200 12156 15252 12162
rect 15200 12098 15252 12104
rect 15856 12150 16068 12178
rect 15108 12088 15160 12094
rect 15108 12030 15160 12036
rect 15212 11414 15240 12098
rect 15856 12094 15884 12150
rect 15844 12088 15896 12094
rect 15844 12030 15896 12036
rect 15200 11408 15252 11414
rect 15200 11350 15252 11356
rect 15856 9918 15884 12030
rect 16028 11476 16080 11482
rect 16028 11418 16080 11424
rect 16040 10394 16068 11418
rect 16120 11408 16172 11414
rect 16120 11350 16172 11356
rect 16132 11210 16160 11350
rect 16120 11204 16172 11210
rect 16120 11146 16172 11152
rect 16028 10388 16080 10394
rect 16028 10330 16080 10336
rect 15844 9912 15896 9918
rect 15844 9854 15896 9860
rect 15016 9504 15068 9510
rect 15016 9446 15068 9452
rect 15568 9368 15620 9374
rect 15568 9310 15620 9316
rect 14684 9132 14980 9152
rect 14740 9130 14764 9132
rect 14820 9130 14844 9132
rect 14900 9130 14924 9132
rect 14762 9078 14764 9130
rect 14826 9078 14838 9130
rect 14900 9078 14902 9130
rect 14740 9076 14764 9078
rect 14820 9076 14844 9078
rect 14900 9076 14924 9078
rect 14684 9056 14980 9076
rect 15580 8966 15608 9310
rect 15568 8960 15620 8966
rect 15568 8902 15620 8908
rect 14684 8044 14980 8064
rect 14740 8042 14764 8044
rect 14820 8042 14844 8044
rect 14900 8042 14924 8044
rect 14762 7990 14764 8042
rect 14826 7990 14838 8042
rect 14900 7990 14902 8042
rect 14740 7988 14764 7990
rect 14820 7988 14844 7990
rect 14900 7988 14924 7990
rect 14684 7968 14980 7988
rect 14684 6956 14980 6976
rect 14740 6954 14764 6956
rect 14820 6954 14844 6956
rect 14900 6954 14924 6956
rect 14762 6902 14764 6954
rect 14826 6902 14838 6954
rect 14900 6902 14902 6954
rect 14740 6900 14764 6902
rect 14820 6900 14844 6902
rect 14900 6900 14924 6902
rect 14684 6880 14980 6900
rect 14684 5868 14980 5888
rect 14740 5866 14764 5868
rect 14820 5866 14844 5868
rect 14900 5866 14924 5868
rect 14762 5814 14764 5866
rect 14826 5814 14838 5866
rect 14900 5814 14902 5866
rect 14740 5812 14764 5814
rect 14820 5812 14844 5814
rect 14900 5812 14924 5814
rect 14684 5792 14980 5812
rect 14684 4780 14980 4800
rect 14740 4778 14764 4780
rect 14820 4778 14844 4780
rect 14900 4778 14924 4780
rect 14762 4726 14764 4778
rect 14826 4726 14838 4778
rect 14900 4726 14902 4778
rect 14740 4724 14764 4726
rect 14820 4724 14844 4726
rect 14900 4724 14924 4726
rect 14684 4704 14980 4724
rect 14556 3996 14608 4002
rect 14556 3938 14608 3944
rect 7820 3692 8116 3712
rect 7876 3690 7900 3692
rect 7956 3690 7980 3692
rect 8036 3690 8060 3692
rect 7898 3638 7900 3690
rect 7962 3638 7974 3690
rect 8036 3638 8038 3690
rect 7876 3636 7900 3638
rect 7956 3636 7980 3638
rect 8036 3636 8060 3638
rect 7820 3616 8116 3636
rect 14684 3692 14980 3712
rect 14740 3690 14764 3692
rect 14820 3690 14844 3692
rect 14900 3690 14924 3692
rect 14762 3638 14764 3690
rect 14826 3638 14838 3690
rect 14900 3638 14902 3690
rect 14740 3636 14764 3638
rect 14820 3636 14844 3638
rect 14900 3636 14924 3638
rect 14684 3616 14980 3636
rect 4388 3148 4684 3168
rect 4444 3146 4468 3148
rect 4524 3146 4548 3148
rect 4604 3146 4628 3148
rect 4466 3094 4468 3146
rect 4530 3094 4542 3146
rect 4604 3094 4606 3146
rect 4444 3092 4468 3094
rect 4524 3092 4548 3094
rect 4604 3092 4628 3094
rect 4388 3072 4684 3092
rect 11252 3148 11548 3168
rect 11308 3146 11332 3148
rect 11388 3146 11412 3148
rect 11468 3146 11492 3148
rect 11330 3094 11332 3146
rect 11394 3094 11406 3146
rect 11468 3094 11470 3146
rect 11308 3092 11332 3094
rect 11388 3092 11412 3094
rect 11468 3092 11492 3094
rect 11252 3072 11548 3092
rect 7820 2604 8116 2624
rect 7876 2602 7900 2604
rect 7956 2602 7980 2604
rect 8036 2602 8060 2604
rect 7898 2550 7900 2602
rect 7962 2550 7974 2602
rect 8036 2550 8038 2602
rect 7876 2548 7900 2550
rect 7956 2548 7980 2550
rect 8036 2548 8060 2550
rect 7820 2528 8116 2548
rect 14684 2604 14980 2624
rect 14740 2602 14764 2604
rect 14820 2602 14844 2604
rect 14900 2602 14924 2604
rect 14762 2550 14764 2602
rect 14826 2550 14838 2602
rect 14900 2550 14902 2602
rect 14740 2548 14764 2550
rect 14820 2548 14844 2550
rect 14900 2548 14924 2550
rect 14684 2528 14980 2548
rect 4388 2060 4684 2080
rect 4444 2058 4468 2060
rect 4524 2058 4548 2060
rect 4604 2058 4628 2060
rect 4466 2006 4468 2058
rect 4530 2006 4542 2058
rect 4604 2006 4606 2058
rect 4444 2004 4468 2006
rect 4524 2004 4548 2006
rect 4604 2004 4628 2006
rect 4388 1984 4684 2004
rect 11252 2060 11548 2080
rect 11308 2058 11332 2060
rect 11388 2058 11412 2060
rect 11468 2058 11492 2060
rect 11330 2006 11332 2058
rect 11394 2006 11406 2058
rect 11468 2006 11470 2058
rect 11308 2004 11332 2006
rect 11388 2004 11412 2006
rect 11468 2004 11492 2006
rect 11252 1984 11548 2004
rect 16040 1214 16068 10330
rect 16224 9034 16252 17182
rect 16500 17074 16528 17878
rect 17224 17596 17276 17602
rect 17224 17538 17276 17544
rect 17236 17194 17264 17538
rect 17408 17460 17460 17466
rect 17408 17402 17460 17408
rect 17224 17188 17276 17194
rect 17224 17130 17276 17136
rect 16408 17046 16528 17074
rect 16304 14672 16356 14678
rect 16304 14614 16356 14620
rect 16316 11770 16344 14614
rect 16408 11906 16436 17046
rect 16580 15420 16632 15426
rect 16580 15362 16632 15368
rect 16592 13930 16620 15362
rect 16672 15352 16724 15358
rect 16764 15352 16816 15358
rect 16672 15294 16724 15300
rect 16762 15320 16764 15329
rect 16816 15320 16818 15329
rect 16684 15018 16712 15294
rect 16818 15278 16896 15306
rect 16762 15255 16818 15264
rect 16672 15012 16724 15018
rect 16672 14954 16724 14960
rect 16764 14876 16816 14882
rect 16764 14818 16816 14824
rect 16776 14406 16804 14818
rect 16868 14474 16896 15278
rect 16856 14468 16908 14474
rect 16856 14410 16908 14416
rect 16764 14400 16816 14406
rect 16764 14342 16816 14348
rect 16580 13924 16632 13930
rect 16580 13866 16632 13872
rect 16672 13924 16724 13930
rect 16672 13866 16724 13872
rect 16684 13810 16712 13866
rect 16500 13782 16712 13810
rect 16776 13794 16804 14342
rect 16764 13788 16816 13794
rect 16500 12842 16528 13782
rect 16764 13730 16816 13736
rect 16488 12836 16540 12842
rect 16488 12778 16540 12784
rect 17040 12156 17092 12162
rect 17040 12098 17092 12104
rect 16408 11878 16528 11906
rect 16316 11742 16436 11770
rect 16304 11680 16356 11686
rect 16304 11622 16356 11628
rect 16316 10462 16344 11622
rect 16408 11482 16436 11742
rect 16396 11476 16448 11482
rect 16396 11418 16448 11424
rect 16304 10456 16356 10462
rect 16304 10398 16356 10404
rect 16316 10054 16344 10398
rect 16304 10048 16356 10054
rect 16304 9990 16356 9996
rect 16212 9028 16264 9034
rect 16212 8970 16264 8976
rect 16120 8892 16172 8898
rect 16120 8834 16172 8840
rect 16132 8490 16160 8834
rect 16120 8484 16172 8490
rect 16120 8426 16172 8432
rect 16120 7804 16172 7810
rect 16120 7746 16172 7752
rect 16132 7266 16160 7746
rect 16500 7606 16528 11878
rect 17052 11618 17080 12098
rect 17040 11612 17092 11618
rect 17040 11554 17092 11560
rect 16764 11068 16816 11074
rect 16764 11010 16816 11016
rect 16776 10666 16804 11010
rect 17052 11006 17080 11554
rect 17236 11006 17264 17130
rect 17316 16848 17368 16854
rect 17316 16790 17368 16796
rect 17328 16514 17356 16790
rect 17420 16514 17448 17402
rect 17604 16990 17632 18422
rect 17972 17194 18000 18626
rect 18116 18380 18412 18400
rect 18172 18378 18196 18380
rect 18252 18378 18276 18380
rect 18332 18378 18356 18380
rect 18194 18326 18196 18378
rect 18258 18326 18270 18378
rect 18332 18326 18334 18378
rect 18172 18324 18196 18326
rect 18252 18324 18276 18326
rect 18332 18324 18356 18326
rect 18116 18304 18412 18324
rect 18512 17392 18564 17398
rect 18512 17334 18564 17340
rect 18116 17292 18412 17312
rect 18172 17290 18196 17292
rect 18252 17290 18276 17292
rect 18332 17290 18356 17292
rect 18194 17238 18196 17290
rect 18258 17238 18270 17290
rect 18332 17238 18334 17290
rect 18172 17236 18196 17238
rect 18252 17236 18276 17238
rect 18332 17236 18356 17238
rect 18116 17216 18412 17236
rect 17960 17188 18012 17194
rect 17960 17130 18012 17136
rect 17684 17052 17736 17058
rect 17684 16994 17736 17000
rect 17592 16984 17644 16990
rect 17592 16926 17644 16932
rect 17316 16508 17368 16514
rect 17316 16450 17368 16456
rect 17408 16508 17460 16514
rect 17408 16450 17460 16456
rect 17328 15970 17356 16450
rect 17696 16310 17724 16994
rect 17960 16848 18012 16854
rect 17960 16790 18012 16796
rect 17684 16304 17736 16310
rect 17684 16246 17736 16252
rect 17972 16106 18000 16790
rect 18524 16650 18552 17334
rect 18512 16644 18564 16650
rect 18512 16586 18564 16592
rect 18116 16204 18412 16224
rect 18172 16202 18196 16204
rect 18252 16202 18276 16204
rect 18332 16202 18356 16204
rect 18194 16150 18196 16202
rect 18258 16150 18270 16202
rect 18332 16150 18334 16202
rect 18172 16148 18196 16150
rect 18252 16148 18276 16150
rect 18332 16148 18356 16150
rect 18116 16128 18412 16148
rect 17960 16100 18012 16106
rect 17960 16042 18012 16048
rect 17316 15964 17368 15970
rect 17316 15906 17368 15912
rect 17868 15216 17920 15222
rect 17868 15158 17920 15164
rect 17880 14814 17908 15158
rect 18116 15116 18412 15136
rect 18172 15114 18196 15116
rect 18252 15114 18276 15116
rect 18332 15114 18356 15116
rect 18194 15062 18196 15114
rect 18258 15062 18270 15114
rect 18332 15062 18334 15114
rect 18172 15060 18196 15062
rect 18252 15060 18276 15062
rect 18332 15060 18356 15062
rect 18116 15040 18412 15060
rect 17776 14808 17828 14814
rect 17776 14750 17828 14756
rect 17868 14808 17920 14814
rect 17868 14750 17920 14756
rect 17788 14406 17816 14750
rect 18708 14474 18736 19902
rect 18788 19908 18840 19914
rect 18788 19850 18840 19856
rect 18878 19264 18934 19273
rect 18878 19199 18934 19208
rect 18788 19160 18840 19166
rect 18788 19102 18840 19108
rect 18800 18758 18828 19102
rect 18788 18752 18840 18758
rect 18788 18694 18840 18700
rect 18892 16106 18920 19199
rect 18984 19030 19012 20967
rect 19168 19930 19196 22176
rect 19338 21984 19394 21993
rect 19338 21919 19394 21928
rect 19076 19902 19196 19930
rect 19352 19914 19380 21919
rect 19340 19908 19392 19914
rect 18972 19024 19024 19030
rect 18972 18966 19024 18972
rect 19076 18486 19104 19902
rect 19340 19850 19392 19856
rect 19156 19772 19208 19778
rect 19156 19714 19208 19720
rect 19168 18690 19196 19714
rect 19432 18820 19484 18826
rect 19432 18762 19484 18768
rect 19156 18684 19208 18690
rect 19156 18626 19208 18632
rect 19340 18684 19392 18690
rect 19340 18626 19392 18632
rect 19064 18480 19116 18486
rect 19064 18422 19116 18428
rect 19352 18282 19380 18626
rect 19340 18276 19392 18282
rect 19340 18218 19392 18224
rect 19340 18004 19392 18010
rect 19340 17946 19392 17952
rect 19352 17890 19380 17946
rect 19260 17862 19380 17890
rect 19260 16802 19288 17862
rect 19340 17732 19392 17738
rect 19340 17674 19392 17680
rect 19352 16990 19380 17674
rect 19444 17210 19472 18762
rect 19524 18684 19576 18690
rect 19524 18626 19576 18632
rect 19536 17534 19564 18626
rect 19614 18312 19670 18321
rect 19614 18247 19670 18256
rect 19628 17738 19656 18247
rect 19720 18010 19748 22176
rect 20272 20746 20300 22176
rect 19996 20718 20300 20746
rect 19892 18208 19944 18214
rect 19892 18150 19944 18156
rect 19800 18140 19852 18146
rect 19800 18082 19852 18088
rect 19708 18004 19760 18010
rect 19708 17946 19760 17952
rect 19616 17732 19668 17738
rect 19616 17674 19668 17680
rect 19708 17732 19760 17738
rect 19708 17674 19760 17680
rect 19524 17528 19576 17534
rect 19524 17470 19576 17476
rect 19444 17182 19656 17210
rect 19340 16984 19392 16990
rect 19340 16926 19392 16932
rect 19432 16984 19484 16990
rect 19432 16926 19484 16932
rect 19260 16774 19380 16802
rect 18880 16100 18932 16106
rect 18880 16042 18932 16048
rect 19156 15896 19208 15902
rect 19156 15838 19208 15844
rect 19168 15494 19196 15838
rect 19156 15488 19208 15494
rect 19156 15430 19208 15436
rect 19352 14898 19380 16774
rect 19444 16582 19472 16926
rect 19432 16576 19484 16582
rect 19432 16518 19484 16524
rect 19628 16394 19656 17182
rect 19720 16650 19748 17674
rect 19708 16644 19760 16650
rect 19708 16586 19760 16592
rect 19536 16366 19656 16394
rect 19352 14870 19472 14898
rect 19340 14808 19392 14814
rect 19340 14750 19392 14756
rect 18696 14468 18748 14474
rect 18696 14410 18748 14416
rect 19352 14406 19380 14750
rect 17776 14400 17828 14406
rect 17776 14342 17828 14348
rect 19340 14400 19392 14406
rect 19340 14342 19392 14348
rect 18512 14332 18564 14338
rect 18512 14274 18564 14280
rect 17500 14264 17552 14270
rect 17500 14206 17552 14212
rect 17512 13726 17540 14206
rect 18116 14028 18412 14048
rect 18172 14026 18196 14028
rect 18252 14026 18276 14028
rect 18332 14026 18356 14028
rect 18194 13974 18196 14026
rect 18258 13974 18270 14026
rect 18332 13974 18334 14026
rect 18172 13972 18196 13974
rect 18252 13972 18276 13974
rect 18332 13972 18356 13974
rect 18116 13952 18412 13972
rect 18524 13794 18552 14274
rect 18512 13788 18564 13794
rect 18512 13730 18564 13736
rect 17500 13720 17552 13726
rect 17500 13662 17552 13668
rect 17408 13652 17460 13658
rect 17408 13594 17460 13600
rect 18512 13652 18564 13658
rect 18512 13594 18564 13600
rect 17316 12632 17368 12638
rect 17316 12574 17368 12580
rect 17040 11000 17092 11006
rect 17040 10942 17092 10948
rect 17224 11000 17276 11006
rect 17224 10942 17276 10948
rect 16764 10660 16816 10666
rect 16764 10602 16816 10608
rect 16856 10388 16908 10394
rect 16856 10330 16908 10336
rect 16868 9306 16896 10330
rect 16948 10320 17000 10326
rect 16948 10262 17000 10268
rect 16960 9306 16988 10262
rect 17052 10122 17080 10942
rect 17040 10116 17092 10122
rect 17040 10058 17092 10064
rect 16856 9300 16908 9306
rect 16856 9242 16908 9248
rect 16948 9300 17000 9306
rect 16948 9242 17000 9248
rect 16868 8966 16896 9242
rect 16856 8960 16908 8966
rect 16856 8902 16908 8908
rect 16960 8898 16988 9242
rect 16948 8892 17000 8898
rect 16948 8834 17000 8840
rect 17224 8348 17276 8354
rect 17224 8290 17276 8296
rect 16580 8144 16632 8150
rect 16580 8086 16632 8092
rect 16488 7600 16540 7606
rect 16488 7542 16540 7548
rect 16592 7402 16620 8086
rect 17236 7878 17264 8290
rect 17224 7872 17276 7878
rect 17224 7814 17276 7820
rect 17236 7674 17264 7814
rect 17224 7668 17276 7674
rect 17224 7610 17276 7616
rect 16580 7396 16632 7402
rect 16580 7338 16632 7344
rect 16120 7260 16172 7266
rect 16120 7202 16172 7208
rect 16488 6852 16540 6858
rect 16488 6794 16540 6800
rect 16500 5158 16528 6794
rect 16488 5152 16540 5158
rect 16488 5094 16540 5100
rect 16028 1208 16080 1214
rect 16028 1150 16080 1156
rect 17328 505 17356 12574
rect 17420 12298 17448 13594
rect 18116 12940 18412 12960
rect 18172 12938 18196 12940
rect 18252 12938 18276 12940
rect 18332 12938 18356 12940
rect 18194 12886 18196 12938
rect 18258 12886 18270 12938
rect 18332 12886 18334 12938
rect 18172 12884 18196 12886
rect 18252 12884 18276 12886
rect 18332 12884 18356 12886
rect 18116 12864 18412 12884
rect 17684 12564 17736 12570
rect 17684 12506 17736 12512
rect 17408 12292 17460 12298
rect 17408 12234 17460 12240
rect 17408 12088 17460 12094
rect 17408 12030 17460 12036
rect 17420 10938 17448 12030
rect 17696 12026 17724 12506
rect 17776 12292 17828 12298
rect 17776 12234 17828 12240
rect 17684 12020 17736 12026
rect 17684 11962 17736 11968
rect 17788 11074 17816 12234
rect 17960 12224 18012 12230
rect 17960 12166 18012 12172
rect 17776 11068 17828 11074
rect 17776 11010 17828 11016
rect 17408 10932 17460 10938
rect 17408 10874 17460 10880
rect 17788 9442 17816 11010
rect 17868 11000 17920 11006
rect 17868 10942 17920 10948
rect 17776 9436 17828 9442
rect 17776 9378 17828 9384
rect 17788 3633 17816 9378
rect 17880 9238 17908 10942
rect 17868 9232 17920 9238
rect 17868 9174 17920 9180
rect 17774 3624 17830 3633
rect 17774 3559 17830 3568
rect 17880 2817 17908 9174
rect 17972 7062 18000 12166
rect 18116 11852 18412 11872
rect 18172 11850 18196 11852
rect 18252 11850 18276 11852
rect 18332 11850 18356 11852
rect 18194 11798 18196 11850
rect 18258 11798 18270 11850
rect 18332 11798 18334 11850
rect 18172 11796 18196 11798
rect 18252 11796 18276 11798
rect 18332 11796 18356 11798
rect 18116 11776 18412 11796
rect 18116 10764 18412 10784
rect 18172 10762 18196 10764
rect 18252 10762 18276 10764
rect 18332 10762 18356 10764
rect 18194 10710 18196 10762
rect 18258 10710 18270 10762
rect 18332 10710 18334 10762
rect 18172 10708 18196 10710
rect 18252 10708 18276 10710
rect 18332 10708 18356 10710
rect 18116 10688 18412 10708
rect 18524 10666 18552 13594
rect 18972 13244 19024 13250
rect 18972 13186 19024 13192
rect 18984 12706 19012 13186
rect 18972 12700 19024 12706
rect 18972 12642 19024 12648
rect 18696 12632 18748 12638
rect 18696 12574 18748 12580
rect 19444 12586 19472 14870
rect 19536 12722 19564 16366
rect 19616 16304 19668 16310
rect 19616 16246 19668 16252
rect 19628 12842 19656 16246
rect 19812 15306 19840 18082
rect 19904 16310 19932 18150
rect 19892 16304 19944 16310
rect 19892 16246 19944 16252
rect 19892 15896 19944 15902
rect 19892 15838 19944 15844
rect 19904 15494 19932 15838
rect 19892 15488 19944 15494
rect 19892 15430 19944 15436
rect 19812 15278 19932 15306
rect 19800 14332 19852 14338
rect 19800 14274 19852 14280
rect 19812 13833 19840 14274
rect 19904 13862 19932 15278
rect 19892 13856 19944 13862
rect 19798 13824 19854 13833
rect 19892 13798 19944 13804
rect 19798 13759 19854 13768
rect 19800 13720 19852 13726
rect 19800 13662 19852 13668
rect 19708 13380 19760 13386
rect 19708 13322 19760 13328
rect 19720 13289 19748 13322
rect 19706 13280 19762 13289
rect 19706 13215 19762 13224
rect 19812 12881 19840 13662
rect 19798 12872 19854 12881
rect 19616 12836 19668 12842
rect 19798 12807 19854 12816
rect 19616 12778 19668 12784
rect 19536 12694 19656 12722
rect 18708 12298 18736 12574
rect 19444 12558 19564 12586
rect 18696 12292 18748 12298
rect 18696 12234 18748 12240
rect 18604 12224 18656 12230
rect 18604 12166 18656 12172
rect 18616 11754 18644 12166
rect 18696 11952 18748 11958
rect 18696 11894 18748 11900
rect 18604 11748 18656 11754
rect 18604 11690 18656 11696
rect 18512 10660 18564 10666
rect 18512 10602 18564 10608
rect 18236 10320 18288 10326
rect 18236 10262 18288 10268
rect 18248 10122 18276 10262
rect 18236 10116 18288 10122
rect 18236 10058 18288 10064
rect 18116 9676 18412 9696
rect 18172 9674 18196 9676
rect 18252 9674 18276 9676
rect 18332 9674 18356 9676
rect 18194 9622 18196 9674
rect 18258 9622 18270 9674
rect 18332 9622 18334 9674
rect 18172 9620 18196 9622
rect 18252 9620 18276 9622
rect 18332 9620 18356 9622
rect 18116 9600 18412 9620
rect 18116 8588 18412 8608
rect 18172 8586 18196 8588
rect 18252 8586 18276 8588
rect 18332 8586 18356 8588
rect 18194 8534 18196 8586
rect 18258 8534 18270 8586
rect 18332 8534 18334 8586
rect 18172 8532 18196 8534
rect 18252 8532 18276 8534
rect 18332 8532 18356 8534
rect 18116 8512 18412 8532
rect 18052 8280 18104 8286
rect 18052 8222 18104 8228
rect 18064 7810 18092 8222
rect 18052 7804 18104 7810
rect 18052 7746 18104 7752
rect 18116 7500 18412 7520
rect 18172 7498 18196 7500
rect 18252 7498 18276 7500
rect 18332 7498 18356 7500
rect 18194 7446 18196 7498
rect 18258 7446 18270 7498
rect 18332 7446 18334 7498
rect 18172 7444 18196 7446
rect 18252 7444 18276 7446
rect 18332 7444 18356 7446
rect 18116 7424 18412 7444
rect 18604 7124 18656 7130
rect 18604 7066 18656 7072
rect 17960 7056 18012 7062
rect 17960 6998 18012 7004
rect 18512 6716 18564 6722
rect 18512 6658 18564 6664
rect 18116 6412 18412 6432
rect 18172 6410 18196 6412
rect 18252 6410 18276 6412
rect 18332 6410 18356 6412
rect 18194 6358 18196 6410
rect 18258 6358 18270 6410
rect 18332 6358 18334 6410
rect 18172 6356 18196 6358
rect 18252 6356 18276 6358
rect 18332 6356 18356 6358
rect 18116 6336 18412 6356
rect 17960 6104 18012 6110
rect 17960 6046 18012 6052
rect 17972 5945 18000 6046
rect 17958 5936 18014 5945
rect 17958 5871 18014 5880
rect 18524 5537 18552 6658
rect 18616 6489 18644 7066
rect 18602 6480 18658 6489
rect 18602 6415 18658 6424
rect 18510 5528 18566 5537
rect 18510 5463 18566 5472
rect 18116 5324 18412 5344
rect 18172 5322 18196 5324
rect 18252 5322 18276 5324
rect 18332 5322 18356 5324
rect 18194 5270 18196 5322
rect 18258 5270 18270 5322
rect 18332 5270 18334 5322
rect 18172 5268 18196 5270
rect 18252 5268 18276 5270
rect 18332 5268 18356 5270
rect 18116 5248 18412 5268
rect 17960 5220 18012 5226
rect 17960 5162 18012 5168
rect 17972 4993 18000 5162
rect 18052 5152 18104 5158
rect 18052 5094 18104 5100
rect 17958 4984 18014 4993
rect 17958 4919 18014 4928
rect 18064 4585 18092 5094
rect 18050 4576 18106 4585
rect 18050 4511 18106 4520
rect 18116 4236 18412 4256
rect 18172 4234 18196 4236
rect 18252 4234 18276 4236
rect 18332 4234 18356 4236
rect 18194 4182 18196 4234
rect 18258 4182 18270 4234
rect 18332 4182 18334 4234
rect 18172 4180 18196 4182
rect 18252 4180 18276 4182
rect 18332 4180 18356 4182
rect 18116 4160 18412 4180
rect 18512 3996 18564 4002
rect 18512 3938 18564 3944
rect 18524 3225 18552 3938
rect 18510 3216 18566 3225
rect 18116 3148 18412 3168
rect 18510 3151 18566 3160
rect 18172 3146 18196 3148
rect 18252 3146 18276 3148
rect 18332 3146 18356 3148
rect 18194 3094 18196 3146
rect 18258 3094 18270 3146
rect 18332 3094 18334 3146
rect 18172 3092 18196 3094
rect 18252 3092 18276 3094
rect 18332 3092 18356 3094
rect 18116 3072 18412 3092
rect 17866 2808 17922 2817
rect 17866 2743 17922 2752
rect 18116 2060 18412 2080
rect 18172 2058 18196 2060
rect 18252 2058 18276 2060
rect 18332 2058 18356 2060
rect 18194 2006 18196 2058
rect 18258 2006 18270 2058
rect 18332 2006 18334 2058
rect 18172 2004 18196 2006
rect 18252 2004 18276 2006
rect 18332 2004 18356 2006
rect 18116 1984 18412 2004
rect 18708 1457 18736 11894
rect 19156 11408 19208 11414
rect 19156 11350 19208 11356
rect 19168 11210 19196 11350
rect 19156 11204 19208 11210
rect 19156 11146 19208 11152
rect 19340 10524 19392 10530
rect 19340 10466 19392 10472
rect 18972 10320 19024 10326
rect 18972 10262 19024 10268
rect 18786 10016 18842 10025
rect 18786 9951 18842 9960
rect 18800 9374 18828 9951
rect 18984 9578 19012 10262
rect 19352 9986 19380 10466
rect 19340 9980 19392 9986
rect 19340 9922 19392 9928
rect 18972 9572 19024 9578
rect 18972 9514 19024 9520
rect 18788 9368 18840 9374
rect 18788 9310 18840 9316
rect 19064 9300 19116 9306
rect 19064 9242 19116 9248
rect 18880 9232 18932 9238
rect 18880 9174 18932 9180
rect 18788 8960 18840 8966
rect 18788 8902 18840 8908
rect 18800 1865 18828 8902
rect 18892 7198 18920 9174
rect 18880 7192 18932 7198
rect 18880 7134 18932 7140
rect 18880 7056 18932 7062
rect 18880 6998 18932 7004
rect 18892 2273 18920 6998
rect 18878 2264 18934 2273
rect 18878 2199 18934 2208
rect 18786 1856 18842 1865
rect 18786 1791 18842 1800
rect 18694 1448 18750 1457
rect 18694 1383 18750 1392
rect 18144 1208 18196 1214
rect 18144 1150 18196 1156
rect 17314 496 17370 505
rect 17314 431 17370 440
rect 18156 97 18184 1150
rect 19076 913 19104 9242
rect 19352 8490 19380 9922
rect 19432 9436 19484 9442
rect 19432 9378 19484 9384
rect 19340 8484 19392 8490
rect 19340 8426 19392 8432
rect 19444 8218 19472 9378
rect 19536 8422 19564 12558
rect 19628 10666 19656 12694
rect 19708 12632 19760 12638
rect 19708 12574 19760 12580
rect 19720 12337 19748 12574
rect 19706 12328 19762 12337
rect 19996 12298 20024 20718
rect 20074 20624 20130 20633
rect 20074 20559 20130 20568
rect 20088 19914 20116 20559
rect 20626 20080 20682 20089
rect 20626 20015 20682 20024
rect 20640 19914 20668 20015
rect 20076 19908 20128 19914
rect 20076 19850 20128 19856
rect 20628 19908 20680 19914
rect 20628 19850 20680 19856
rect 20260 19772 20312 19778
rect 20260 19714 20312 19720
rect 20444 19772 20496 19778
rect 20444 19714 20496 19720
rect 20272 19234 20300 19714
rect 20260 19228 20312 19234
rect 20260 19170 20312 19176
rect 20076 19160 20128 19166
rect 20076 19102 20128 19108
rect 20088 18554 20116 19102
rect 20456 19098 20484 19714
rect 20718 19672 20774 19681
rect 20718 19607 20774 19616
rect 20444 19092 20496 19098
rect 20444 19034 20496 19040
rect 20732 18826 20760 19607
rect 20720 18820 20772 18826
rect 20720 18762 20772 18768
rect 20534 18720 20590 18729
rect 20534 18655 20590 18664
rect 20076 18548 20128 18554
rect 20076 18490 20128 18496
rect 20260 18072 20312 18078
rect 20260 18014 20312 18020
rect 20076 17936 20128 17942
rect 20076 17878 20128 17884
rect 20088 17738 20116 17878
rect 20076 17732 20128 17738
rect 20076 17674 20128 17680
rect 20076 17596 20128 17602
rect 20076 17538 20128 17544
rect 20088 16582 20116 17538
rect 20168 17392 20220 17398
rect 20168 17334 20220 17340
rect 20180 16961 20208 17334
rect 20272 17058 20300 18014
rect 20352 18004 20404 18010
rect 20352 17946 20404 17952
rect 20260 17052 20312 17058
rect 20260 16994 20312 17000
rect 20166 16952 20222 16961
rect 20166 16887 20222 16896
rect 20364 16802 20392 17946
rect 20444 17936 20496 17942
rect 20442 17904 20444 17913
rect 20496 17904 20498 17913
rect 20442 17839 20498 17848
rect 20444 17732 20496 17738
rect 20444 17674 20496 17680
rect 20180 16774 20392 16802
rect 20076 16576 20128 16582
rect 20076 16518 20128 16524
rect 20076 15420 20128 15426
rect 20076 15362 20128 15368
rect 20088 14406 20116 15362
rect 20076 14400 20128 14406
rect 20076 14342 20128 14348
rect 19706 12263 19762 12272
rect 19984 12292 20036 12298
rect 19984 12234 20036 12240
rect 19984 12156 20036 12162
rect 19984 12098 20036 12104
rect 20076 12156 20128 12162
rect 20076 12098 20128 12104
rect 19996 11521 20024 12098
rect 20088 11550 20116 12098
rect 20180 11754 20208 16774
rect 20260 16644 20312 16650
rect 20260 16586 20312 16592
rect 20272 12722 20300 16586
rect 20456 16122 20484 17674
rect 20364 16094 20484 16122
rect 20364 12842 20392 16094
rect 20444 16032 20496 16038
rect 20442 16000 20444 16009
rect 20496 16000 20498 16009
rect 20442 15935 20498 15944
rect 20442 15048 20498 15057
rect 20442 14983 20444 14992
rect 20496 14983 20498 14992
rect 20444 14954 20496 14960
rect 20548 14898 20576 18655
rect 20628 18480 20680 18486
rect 20628 18422 20680 18428
rect 20640 16802 20668 18422
rect 20824 17738 20852 22176
rect 21180 18616 21232 18622
rect 21180 18558 21232 18564
rect 20996 17936 21048 17942
rect 20996 17878 21048 17884
rect 20812 17732 20864 17738
rect 20812 17674 20864 17680
rect 20812 17528 20864 17534
rect 20812 17470 20864 17476
rect 20720 17392 20772 17398
rect 20718 17360 20720 17369
rect 20772 17360 20774 17369
rect 20718 17295 20774 17304
rect 20824 17058 20852 17470
rect 20812 17052 20864 17058
rect 20812 16994 20864 17000
rect 20640 16774 20760 16802
rect 20628 16644 20680 16650
rect 20628 16586 20680 16592
rect 20640 16417 20668 16586
rect 20626 16408 20682 16417
rect 20626 16343 20682 16352
rect 20732 16258 20760 16774
rect 20640 16230 20760 16258
rect 20640 15034 20668 16230
rect 20718 15592 20774 15601
rect 20718 15527 20720 15536
rect 20772 15527 20774 15536
rect 20720 15498 20772 15504
rect 20640 15006 20760 15034
rect 20548 14870 20668 14898
rect 20536 14740 20588 14746
rect 20536 14682 20588 14688
rect 20442 14640 20498 14649
rect 20442 14575 20498 14584
rect 20456 13930 20484 14575
rect 20548 14338 20576 14682
rect 20640 14474 20668 14870
rect 20628 14468 20680 14474
rect 20628 14410 20680 14416
rect 20732 14354 20760 15006
rect 20536 14332 20588 14338
rect 20536 14274 20588 14280
rect 20640 14326 20760 14354
rect 20444 13924 20496 13930
rect 20444 13866 20496 13872
rect 20352 12836 20404 12842
rect 20352 12778 20404 12784
rect 20272 12694 20392 12722
rect 20260 12632 20312 12638
rect 20260 12574 20312 12580
rect 20272 11929 20300 12574
rect 20258 11920 20314 11929
rect 20258 11855 20314 11864
rect 20168 11748 20220 11754
rect 20168 11690 20220 11696
rect 20076 11544 20128 11550
rect 19982 11512 20038 11521
rect 20076 11486 20128 11492
rect 20260 11544 20312 11550
rect 20260 11486 20312 11492
rect 19982 11447 20038 11456
rect 19800 11000 19852 11006
rect 20272 10977 20300 11486
rect 19800 10942 19852 10948
rect 20258 10968 20314 10977
rect 19616 10660 19668 10666
rect 19616 10602 19668 10608
rect 19812 10462 19840 10942
rect 20258 10903 20314 10912
rect 19800 10456 19852 10462
rect 19800 10398 19852 10404
rect 20260 10456 20312 10462
rect 20260 10398 20312 10404
rect 19812 10122 19840 10398
rect 19800 10116 19852 10122
rect 19800 10058 19852 10064
rect 20272 9617 20300 10398
rect 20258 9608 20314 9617
rect 20258 9543 20314 9552
rect 20364 9510 20392 12694
rect 20640 11210 20668 14326
rect 20718 13688 20774 13697
rect 20718 13623 20774 13632
rect 20732 13386 20760 13623
rect 20720 13380 20772 13386
rect 20720 13322 20772 13328
rect 20628 11204 20680 11210
rect 20628 11146 20680 11152
rect 20536 11068 20588 11074
rect 20536 11010 20588 11016
rect 20548 10569 20576 11010
rect 20534 10560 20590 10569
rect 20534 10495 20590 10504
rect 20536 9980 20588 9986
rect 20536 9922 20588 9928
rect 20352 9504 20404 9510
rect 20352 9446 20404 9452
rect 20260 9368 20312 9374
rect 20260 9310 20312 9316
rect 20272 8665 20300 9310
rect 20548 9209 20576 9922
rect 20534 9200 20590 9209
rect 20534 9135 20590 9144
rect 20536 8892 20588 8898
rect 20536 8834 20588 8840
rect 20258 8656 20314 8665
rect 20258 8591 20314 8600
rect 19524 8416 19576 8422
rect 19524 8358 19576 8364
rect 20260 8280 20312 8286
rect 20548 8257 20576 8834
rect 20260 8222 20312 8228
rect 20534 8248 20590 8257
rect 19432 8212 19484 8218
rect 19432 8154 19484 8160
rect 19444 7946 19472 8154
rect 19432 7940 19484 7946
rect 19432 7882 19484 7888
rect 20272 7849 20300 8222
rect 20534 8183 20590 8192
rect 20258 7840 20314 7849
rect 19984 7804 20036 7810
rect 20258 7775 20314 7784
rect 20536 7804 20588 7810
rect 19984 7746 20036 7752
rect 20536 7746 20588 7752
rect 19996 7305 20024 7746
rect 19982 7296 20038 7305
rect 19982 7231 20038 7240
rect 20548 6897 20576 7746
rect 20534 6888 20590 6897
rect 20534 6823 20590 6832
rect 21008 4682 21036 17878
rect 21086 14232 21142 14241
rect 21086 14167 21142 14176
rect 21100 12298 21128 14167
rect 21088 12292 21140 12298
rect 21088 12234 21140 12240
rect 21192 10122 21220 18558
rect 21376 18214 21404 22176
rect 21364 18208 21416 18214
rect 21364 18150 21416 18156
rect 21928 18146 21956 22176
rect 21916 18140 21968 18146
rect 21916 18082 21968 18088
rect 22480 17942 22508 22176
rect 22468 17936 22520 17942
rect 22468 17878 22520 17884
rect 21180 10116 21232 10122
rect 21180 10058 21232 10064
rect 20996 4676 21048 4682
rect 20996 4618 21048 4624
rect 20536 4540 20588 4546
rect 20536 4482 20588 4488
rect 20548 4177 20576 4482
rect 20534 4168 20590 4177
rect 20534 4103 20590 4112
rect 19062 904 19118 913
rect 19062 839 19118 848
rect 18142 88 18198 97
rect 18142 23 18198 32
<< via2 >>
rect 17958 22336 18014 22392
rect 4388 19466 4444 19468
rect 4468 19466 4524 19468
rect 4548 19466 4604 19468
rect 4628 19466 4684 19468
rect 4388 19414 4414 19466
rect 4414 19414 4444 19466
rect 4468 19414 4478 19466
rect 4478 19414 4524 19466
rect 4548 19414 4594 19466
rect 4594 19414 4604 19466
rect 4628 19414 4658 19466
rect 4658 19414 4684 19466
rect 4388 19412 4444 19414
rect 4468 19412 4524 19414
rect 4548 19412 4604 19414
rect 4628 19412 4684 19414
rect 4388 18378 4444 18380
rect 4468 18378 4524 18380
rect 4548 18378 4604 18380
rect 4628 18378 4684 18380
rect 4388 18326 4414 18378
rect 4414 18326 4444 18378
rect 4468 18326 4478 18378
rect 4478 18326 4524 18378
rect 4548 18326 4594 18378
rect 4594 18326 4604 18378
rect 4628 18326 4658 18378
rect 4658 18326 4684 18378
rect 4388 18324 4444 18326
rect 4468 18324 4524 18326
rect 4548 18324 4604 18326
rect 4628 18324 4684 18326
rect 4388 17290 4444 17292
rect 4468 17290 4524 17292
rect 4548 17290 4604 17292
rect 4628 17290 4684 17292
rect 4388 17238 4414 17290
rect 4414 17238 4444 17290
rect 4468 17238 4478 17290
rect 4478 17238 4524 17290
rect 4548 17238 4594 17290
rect 4594 17238 4604 17290
rect 4628 17238 4658 17290
rect 4658 17238 4684 17290
rect 4388 17236 4444 17238
rect 4468 17236 4524 17238
rect 4548 17236 4604 17238
rect 4628 17236 4684 17238
rect 4388 16202 4444 16204
rect 4468 16202 4524 16204
rect 4548 16202 4604 16204
rect 4628 16202 4684 16204
rect 4388 16150 4414 16202
rect 4414 16150 4444 16202
rect 4468 16150 4478 16202
rect 4478 16150 4524 16202
rect 4548 16150 4594 16202
rect 4594 16150 4604 16202
rect 4628 16150 4658 16202
rect 4658 16150 4684 16202
rect 4388 16148 4444 16150
rect 4468 16148 4524 16150
rect 4548 16148 4604 16150
rect 4628 16148 4684 16150
rect 4388 15114 4444 15116
rect 4468 15114 4524 15116
rect 4548 15114 4604 15116
rect 4628 15114 4684 15116
rect 4388 15062 4414 15114
rect 4414 15062 4444 15114
rect 4468 15062 4478 15114
rect 4478 15062 4524 15114
rect 4548 15062 4594 15114
rect 4594 15062 4604 15114
rect 4628 15062 4658 15114
rect 4658 15062 4684 15114
rect 4388 15060 4444 15062
rect 4468 15060 4524 15062
rect 4548 15060 4604 15062
rect 4628 15060 4684 15062
rect 4388 14026 4444 14028
rect 4468 14026 4524 14028
rect 4548 14026 4604 14028
rect 4628 14026 4684 14028
rect 4388 13974 4414 14026
rect 4414 13974 4444 14026
rect 4468 13974 4478 14026
rect 4478 13974 4524 14026
rect 4548 13974 4594 14026
rect 4594 13974 4604 14026
rect 4628 13974 4658 14026
rect 4658 13974 4684 14026
rect 4388 13972 4444 13974
rect 4468 13972 4524 13974
rect 4548 13972 4604 13974
rect 4628 13972 4684 13974
rect 4388 12938 4444 12940
rect 4468 12938 4524 12940
rect 4548 12938 4604 12940
rect 4628 12938 4684 12940
rect 4388 12886 4414 12938
rect 4414 12886 4444 12938
rect 4468 12886 4478 12938
rect 4478 12886 4524 12938
rect 4548 12886 4594 12938
rect 4594 12886 4604 12938
rect 4628 12886 4658 12938
rect 4658 12886 4684 12938
rect 4388 12884 4444 12886
rect 4468 12884 4524 12886
rect 4548 12884 4604 12886
rect 4628 12884 4684 12886
rect 7820 20010 7876 20012
rect 7900 20010 7956 20012
rect 7980 20010 8036 20012
rect 8060 20010 8116 20012
rect 7820 19958 7846 20010
rect 7846 19958 7876 20010
rect 7900 19958 7910 20010
rect 7910 19958 7956 20010
rect 7980 19958 8026 20010
rect 8026 19958 8036 20010
rect 8060 19958 8090 20010
rect 8090 19958 8116 20010
rect 7820 19956 7876 19958
rect 7900 19956 7956 19958
rect 7980 19956 8036 19958
rect 8060 19956 8116 19958
rect 7820 18922 7876 18924
rect 7900 18922 7956 18924
rect 7980 18922 8036 18924
rect 8060 18922 8116 18924
rect 7820 18870 7846 18922
rect 7846 18870 7876 18922
rect 7900 18870 7910 18922
rect 7910 18870 7956 18922
rect 7980 18870 8026 18922
rect 8026 18870 8036 18922
rect 8060 18870 8090 18922
rect 8090 18870 8116 18922
rect 7820 18868 7876 18870
rect 7900 18868 7956 18870
rect 7980 18868 8036 18870
rect 8060 18868 8116 18870
rect 7820 17834 7876 17836
rect 7900 17834 7956 17836
rect 7980 17834 8036 17836
rect 8060 17834 8116 17836
rect 7820 17782 7846 17834
rect 7846 17782 7876 17834
rect 7900 17782 7910 17834
rect 7910 17782 7956 17834
rect 7980 17782 8026 17834
rect 8026 17782 8036 17834
rect 8060 17782 8090 17834
rect 8090 17782 8116 17834
rect 7820 17780 7876 17782
rect 7900 17780 7956 17782
rect 7980 17780 8036 17782
rect 8060 17780 8116 17782
rect 7820 16746 7876 16748
rect 7900 16746 7956 16748
rect 7980 16746 8036 16748
rect 8060 16746 8116 16748
rect 7820 16694 7846 16746
rect 7846 16694 7876 16746
rect 7900 16694 7910 16746
rect 7910 16694 7956 16746
rect 7980 16694 8026 16746
rect 8026 16694 8036 16746
rect 8060 16694 8090 16746
rect 8090 16694 8116 16746
rect 7820 16692 7876 16694
rect 7900 16692 7956 16694
rect 7980 16692 8036 16694
rect 8060 16692 8116 16694
rect 7820 15658 7876 15660
rect 7900 15658 7956 15660
rect 7980 15658 8036 15660
rect 8060 15658 8116 15660
rect 7820 15606 7846 15658
rect 7846 15606 7876 15658
rect 7900 15606 7910 15658
rect 7910 15606 7956 15658
rect 7980 15606 8026 15658
rect 8026 15606 8036 15658
rect 8060 15606 8090 15658
rect 8090 15606 8116 15658
rect 7820 15604 7876 15606
rect 7900 15604 7956 15606
rect 7980 15604 8036 15606
rect 8060 15604 8116 15606
rect 7820 14570 7876 14572
rect 7900 14570 7956 14572
rect 7980 14570 8036 14572
rect 8060 14570 8116 14572
rect 7820 14518 7846 14570
rect 7846 14518 7876 14570
rect 7900 14518 7910 14570
rect 7910 14518 7956 14570
rect 7980 14518 8026 14570
rect 8026 14518 8036 14570
rect 8060 14518 8090 14570
rect 8090 14518 8116 14570
rect 7820 14516 7876 14518
rect 7900 14516 7956 14518
rect 7980 14516 8036 14518
rect 8060 14516 8116 14518
rect 7820 13482 7876 13484
rect 7900 13482 7956 13484
rect 7980 13482 8036 13484
rect 8060 13482 8116 13484
rect 7820 13430 7846 13482
rect 7846 13430 7876 13482
rect 7900 13430 7910 13482
rect 7910 13430 7956 13482
rect 7980 13430 8026 13482
rect 8026 13430 8036 13482
rect 8060 13430 8090 13482
rect 8090 13430 8116 13482
rect 7820 13428 7876 13430
rect 7900 13428 7956 13430
rect 7980 13428 8036 13430
rect 8060 13428 8116 13430
rect 4388 11850 4444 11852
rect 4468 11850 4524 11852
rect 4548 11850 4604 11852
rect 4628 11850 4684 11852
rect 4388 11798 4414 11850
rect 4414 11798 4444 11850
rect 4468 11798 4478 11850
rect 4478 11798 4524 11850
rect 4548 11798 4594 11850
rect 4594 11798 4604 11850
rect 4628 11798 4658 11850
rect 4658 11798 4684 11850
rect 4388 11796 4444 11798
rect 4468 11796 4524 11798
rect 4548 11796 4604 11798
rect 4628 11796 4684 11798
rect 4388 10762 4444 10764
rect 4468 10762 4524 10764
rect 4548 10762 4604 10764
rect 4628 10762 4684 10764
rect 4388 10710 4414 10762
rect 4414 10710 4444 10762
rect 4468 10710 4478 10762
rect 4478 10710 4524 10762
rect 4548 10710 4594 10762
rect 4594 10710 4604 10762
rect 4628 10710 4658 10762
rect 4658 10710 4684 10762
rect 4388 10708 4444 10710
rect 4468 10708 4524 10710
rect 4548 10708 4604 10710
rect 4628 10708 4684 10710
rect 7820 12394 7876 12396
rect 7900 12394 7956 12396
rect 7980 12394 8036 12396
rect 8060 12394 8116 12396
rect 7820 12342 7846 12394
rect 7846 12342 7876 12394
rect 7900 12342 7910 12394
rect 7910 12342 7956 12394
rect 7980 12342 8026 12394
rect 8026 12342 8036 12394
rect 8060 12342 8090 12394
rect 8090 12342 8116 12394
rect 7820 12340 7876 12342
rect 7900 12340 7956 12342
rect 7980 12340 8036 12342
rect 8060 12340 8116 12342
rect 9586 17032 9642 17088
rect 7820 11306 7876 11308
rect 7900 11306 7956 11308
rect 7980 11306 8036 11308
rect 8060 11306 8116 11308
rect 7820 11254 7846 11306
rect 7846 11254 7876 11306
rect 7900 11254 7910 11306
rect 7910 11254 7956 11306
rect 7980 11254 8026 11306
rect 8026 11254 8036 11306
rect 8060 11254 8090 11306
rect 8090 11254 8116 11306
rect 7820 11252 7876 11254
rect 7900 11252 7956 11254
rect 7980 11252 8036 11254
rect 8060 11252 8116 11254
rect 9862 13804 9864 13824
rect 9864 13804 9916 13824
rect 9916 13804 9918 13824
rect 9862 13768 9918 13804
rect 7820 10218 7876 10220
rect 7900 10218 7956 10220
rect 7980 10218 8036 10220
rect 8060 10218 8116 10220
rect 7820 10166 7846 10218
rect 7846 10166 7876 10218
rect 7900 10166 7910 10218
rect 7910 10166 7956 10218
rect 7980 10166 8026 10218
rect 8026 10166 8036 10218
rect 8060 10166 8090 10218
rect 8090 10166 8116 10218
rect 7820 10164 7876 10166
rect 7900 10164 7956 10166
rect 7980 10164 8036 10166
rect 8060 10164 8116 10166
rect 4388 9674 4444 9676
rect 4468 9674 4524 9676
rect 4548 9674 4604 9676
rect 4628 9674 4684 9676
rect 4388 9622 4414 9674
rect 4414 9622 4444 9674
rect 4468 9622 4478 9674
rect 4478 9622 4524 9674
rect 4548 9622 4594 9674
rect 4594 9622 4604 9674
rect 4628 9622 4658 9674
rect 4658 9622 4684 9674
rect 4388 9620 4444 9622
rect 4468 9620 4524 9622
rect 4548 9620 4604 9622
rect 4628 9620 4684 9622
rect 7820 9130 7876 9132
rect 7900 9130 7956 9132
rect 7980 9130 8036 9132
rect 8060 9130 8116 9132
rect 7820 9078 7846 9130
rect 7846 9078 7876 9130
rect 7900 9078 7910 9130
rect 7910 9078 7956 9130
rect 7980 9078 8026 9130
rect 8026 9078 8036 9130
rect 8060 9078 8090 9130
rect 8090 9078 8116 9130
rect 7820 9076 7876 9078
rect 7900 9076 7956 9078
rect 7980 9076 8036 9078
rect 8060 9076 8116 9078
rect 4388 8586 4444 8588
rect 4468 8586 4524 8588
rect 4548 8586 4604 8588
rect 4628 8586 4684 8588
rect 4388 8534 4414 8586
rect 4414 8534 4444 8586
rect 4468 8534 4478 8586
rect 4478 8534 4524 8586
rect 4548 8534 4594 8586
rect 4594 8534 4604 8586
rect 4628 8534 4658 8586
rect 4658 8534 4684 8586
rect 4388 8532 4444 8534
rect 4468 8532 4524 8534
rect 4548 8532 4604 8534
rect 4628 8532 4684 8534
rect 7820 8042 7876 8044
rect 7900 8042 7956 8044
rect 7980 8042 8036 8044
rect 8060 8042 8116 8044
rect 7820 7990 7846 8042
rect 7846 7990 7876 8042
rect 7900 7990 7910 8042
rect 7910 7990 7956 8042
rect 7980 7990 8026 8042
rect 8026 7990 8036 8042
rect 8060 7990 8090 8042
rect 8090 7990 8116 8042
rect 7820 7988 7876 7990
rect 7900 7988 7956 7990
rect 7980 7988 8036 7990
rect 8060 7988 8116 7990
rect 4388 7498 4444 7500
rect 4468 7498 4524 7500
rect 4548 7498 4604 7500
rect 4628 7498 4684 7500
rect 4388 7446 4414 7498
rect 4414 7446 4444 7498
rect 4468 7446 4478 7498
rect 4478 7446 4524 7498
rect 4548 7446 4594 7498
rect 4594 7446 4604 7498
rect 4628 7446 4658 7498
rect 4658 7446 4684 7498
rect 4388 7444 4444 7446
rect 4468 7444 4524 7446
rect 4548 7444 4604 7446
rect 4628 7444 4684 7446
rect 7820 6954 7876 6956
rect 7900 6954 7956 6956
rect 7980 6954 8036 6956
rect 8060 6954 8116 6956
rect 7820 6902 7846 6954
rect 7846 6902 7876 6954
rect 7900 6902 7910 6954
rect 7910 6902 7956 6954
rect 7980 6902 8026 6954
rect 8026 6902 8036 6954
rect 8060 6902 8090 6954
rect 8090 6902 8116 6954
rect 7820 6900 7876 6902
rect 7900 6900 7956 6902
rect 7980 6900 8036 6902
rect 8060 6900 8116 6902
rect 11252 19466 11308 19468
rect 11332 19466 11388 19468
rect 11412 19466 11468 19468
rect 11492 19466 11548 19468
rect 11252 19414 11278 19466
rect 11278 19414 11308 19466
rect 11332 19414 11342 19466
rect 11342 19414 11388 19466
rect 11412 19414 11458 19466
rect 11458 19414 11468 19466
rect 11492 19414 11522 19466
rect 11522 19414 11548 19466
rect 11252 19412 11308 19414
rect 11332 19412 11388 19414
rect 11412 19412 11468 19414
rect 11492 19412 11548 19414
rect 11252 18378 11308 18380
rect 11332 18378 11388 18380
rect 11412 18378 11468 18380
rect 11492 18378 11548 18380
rect 11252 18326 11278 18378
rect 11278 18326 11308 18378
rect 11332 18326 11342 18378
rect 11342 18326 11388 18378
rect 11412 18326 11458 18378
rect 11458 18326 11468 18378
rect 11492 18326 11522 18378
rect 11522 18326 11548 18378
rect 11252 18324 11308 18326
rect 11332 18324 11388 18326
rect 11412 18324 11468 18326
rect 11492 18324 11548 18326
rect 11252 17290 11308 17292
rect 11332 17290 11388 17292
rect 11412 17290 11468 17292
rect 11492 17290 11548 17292
rect 11252 17238 11278 17290
rect 11278 17238 11308 17290
rect 11332 17238 11342 17290
rect 11342 17238 11388 17290
rect 11412 17238 11458 17290
rect 11458 17238 11468 17290
rect 11492 17238 11522 17290
rect 11522 17238 11548 17290
rect 11252 17236 11308 17238
rect 11332 17236 11388 17238
rect 11412 17236 11468 17238
rect 11492 17236 11548 17238
rect 11252 16202 11308 16204
rect 11332 16202 11388 16204
rect 11412 16202 11468 16204
rect 11492 16202 11548 16204
rect 11252 16150 11278 16202
rect 11278 16150 11308 16202
rect 11332 16150 11342 16202
rect 11342 16150 11388 16202
rect 11412 16150 11458 16202
rect 11458 16150 11468 16202
rect 11492 16150 11522 16202
rect 11522 16150 11548 16202
rect 11252 16148 11308 16150
rect 11332 16148 11388 16150
rect 11412 16148 11468 16150
rect 11492 16148 11548 16150
rect 11252 15114 11308 15116
rect 11332 15114 11388 15116
rect 11412 15114 11468 15116
rect 11492 15114 11548 15116
rect 11252 15062 11278 15114
rect 11278 15062 11308 15114
rect 11332 15062 11342 15114
rect 11342 15062 11388 15114
rect 11412 15062 11458 15114
rect 11458 15062 11468 15114
rect 11492 15062 11522 15114
rect 11522 15062 11548 15114
rect 11252 15060 11308 15062
rect 11332 15060 11388 15062
rect 11412 15060 11468 15062
rect 11492 15060 11548 15062
rect 11252 14026 11308 14028
rect 11332 14026 11388 14028
rect 11412 14026 11468 14028
rect 11492 14026 11548 14028
rect 11252 13974 11278 14026
rect 11278 13974 11308 14026
rect 11332 13974 11342 14026
rect 11342 13974 11388 14026
rect 11412 13974 11458 14026
rect 11458 13974 11468 14026
rect 11492 13974 11522 14026
rect 11522 13974 11548 14026
rect 11252 13972 11308 13974
rect 11332 13972 11388 13974
rect 11412 13972 11468 13974
rect 11492 13972 11548 13974
rect 11252 12938 11308 12940
rect 11332 12938 11388 12940
rect 11412 12938 11468 12940
rect 11492 12938 11548 12940
rect 11252 12886 11278 12938
rect 11278 12886 11308 12938
rect 11332 12886 11342 12938
rect 11342 12886 11388 12938
rect 11412 12886 11458 12938
rect 11458 12886 11468 12938
rect 11492 12886 11522 12938
rect 11522 12886 11548 12938
rect 11252 12884 11308 12886
rect 11332 12884 11388 12886
rect 11412 12884 11468 12886
rect 11492 12884 11548 12886
rect 11252 11850 11308 11852
rect 11332 11850 11388 11852
rect 11412 11850 11468 11852
rect 11492 11850 11548 11852
rect 11252 11798 11278 11850
rect 11278 11798 11308 11850
rect 11332 11798 11342 11850
rect 11342 11798 11388 11850
rect 11412 11798 11458 11850
rect 11458 11798 11468 11850
rect 11492 11798 11522 11850
rect 11522 11798 11548 11850
rect 11252 11796 11308 11798
rect 11332 11796 11388 11798
rect 11412 11796 11468 11798
rect 11492 11796 11548 11798
rect 11252 10762 11308 10764
rect 11332 10762 11388 10764
rect 11412 10762 11468 10764
rect 11492 10762 11548 10764
rect 11252 10710 11278 10762
rect 11278 10710 11308 10762
rect 11332 10710 11342 10762
rect 11342 10710 11388 10762
rect 11412 10710 11458 10762
rect 11458 10710 11468 10762
rect 11492 10710 11522 10762
rect 11522 10710 11548 10762
rect 11252 10708 11308 10710
rect 11332 10708 11388 10710
rect 11412 10708 11468 10710
rect 11492 10708 11548 10710
rect 11252 9674 11308 9676
rect 11332 9674 11388 9676
rect 11412 9674 11468 9676
rect 11492 9674 11548 9676
rect 11252 9622 11278 9674
rect 11278 9622 11308 9674
rect 11332 9622 11342 9674
rect 11342 9622 11388 9674
rect 11412 9622 11458 9674
rect 11458 9622 11468 9674
rect 11492 9622 11522 9674
rect 11522 9622 11548 9674
rect 11252 9620 11308 9622
rect 11332 9620 11388 9622
rect 11412 9620 11468 9622
rect 11492 9620 11548 9622
rect 12714 18004 12770 18040
rect 12714 17984 12716 18004
rect 12716 17984 12768 18004
rect 12768 17984 12770 18004
rect 12162 15264 12218 15320
rect 11252 8586 11308 8588
rect 11332 8586 11388 8588
rect 11412 8586 11468 8588
rect 11492 8586 11548 8588
rect 11252 8534 11278 8586
rect 11278 8534 11308 8586
rect 11332 8534 11342 8586
rect 11342 8534 11388 8586
rect 11412 8534 11458 8586
rect 11458 8534 11468 8586
rect 11492 8534 11522 8586
rect 11522 8534 11548 8586
rect 11252 8532 11308 8534
rect 11332 8532 11388 8534
rect 11412 8532 11468 8534
rect 11492 8532 11548 8534
rect 11252 7498 11308 7500
rect 11332 7498 11388 7500
rect 11412 7498 11468 7500
rect 11492 7498 11548 7500
rect 11252 7446 11278 7498
rect 11278 7446 11308 7498
rect 11332 7446 11342 7498
rect 11342 7446 11388 7498
rect 11412 7446 11458 7498
rect 11458 7446 11468 7498
rect 11492 7446 11522 7498
rect 11522 7446 11548 7498
rect 11252 7444 11308 7446
rect 11332 7444 11388 7446
rect 11412 7444 11468 7446
rect 11492 7444 11548 7446
rect 4388 6410 4444 6412
rect 4468 6410 4524 6412
rect 4548 6410 4604 6412
rect 4628 6410 4684 6412
rect 4388 6358 4414 6410
rect 4414 6358 4444 6410
rect 4468 6358 4478 6410
rect 4478 6358 4524 6410
rect 4548 6358 4594 6410
rect 4594 6358 4604 6410
rect 4628 6358 4658 6410
rect 4658 6358 4684 6410
rect 4388 6356 4444 6358
rect 4468 6356 4524 6358
rect 4548 6356 4604 6358
rect 4628 6356 4684 6358
rect 11252 6410 11308 6412
rect 11332 6410 11388 6412
rect 11412 6410 11468 6412
rect 11492 6410 11548 6412
rect 11252 6358 11278 6410
rect 11278 6358 11308 6410
rect 11332 6358 11342 6410
rect 11342 6358 11388 6410
rect 11412 6358 11458 6410
rect 11458 6358 11468 6410
rect 11492 6358 11522 6410
rect 11522 6358 11548 6410
rect 11252 6356 11308 6358
rect 11332 6356 11388 6358
rect 11412 6356 11468 6358
rect 11492 6356 11548 6358
rect 7820 5866 7876 5868
rect 7900 5866 7956 5868
rect 7980 5866 8036 5868
rect 8060 5866 8116 5868
rect 7820 5814 7846 5866
rect 7846 5814 7876 5866
rect 7900 5814 7910 5866
rect 7910 5814 7956 5866
rect 7980 5814 8026 5866
rect 8026 5814 8036 5866
rect 8060 5814 8090 5866
rect 8090 5814 8116 5866
rect 7820 5812 7876 5814
rect 7900 5812 7956 5814
rect 7980 5812 8036 5814
rect 8060 5812 8116 5814
rect 13358 18004 13414 18040
rect 13358 17984 13360 18004
rect 13360 17984 13412 18004
rect 13412 17984 13414 18004
rect 14684 20010 14740 20012
rect 14764 20010 14820 20012
rect 14844 20010 14900 20012
rect 14924 20010 14980 20012
rect 14684 19958 14710 20010
rect 14710 19958 14740 20010
rect 14764 19958 14774 20010
rect 14774 19958 14820 20010
rect 14844 19958 14890 20010
rect 14890 19958 14900 20010
rect 14924 19958 14954 20010
rect 14954 19958 14980 20010
rect 14684 19956 14740 19958
rect 14764 19956 14820 19958
rect 14844 19956 14900 19958
rect 14924 19956 14980 19958
rect 14684 18922 14740 18924
rect 14764 18922 14820 18924
rect 14844 18922 14900 18924
rect 14924 18922 14980 18924
rect 14684 18870 14710 18922
rect 14710 18870 14740 18922
rect 14764 18870 14774 18922
rect 14774 18870 14820 18922
rect 14844 18870 14890 18922
rect 14890 18870 14900 18922
rect 14924 18870 14954 18922
rect 14954 18870 14980 18922
rect 14684 18868 14740 18870
rect 14764 18868 14820 18870
rect 14844 18868 14900 18870
rect 14924 18868 14980 18870
rect 14684 17834 14740 17836
rect 14764 17834 14820 17836
rect 14844 17834 14900 17836
rect 14924 17834 14980 17836
rect 14684 17782 14710 17834
rect 14710 17782 14740 17834
rect 14764 17782 14774 17834
rect 14774 17782 14820 17834
rect 14844 17782 14890 17834
rect 14890 17782 14900 17834
rect 14924 17782 14954 17834
rect 14954 17782 14980 17834
rect 14684 17780 14740 17782
rect 14764 17780 14820 17782
rect 14844 17780 14900 17782
rect 14924 17780 14980 17782
rect 14684 16746 14740 16748
rect 14764 16746 14820 16748
rect 14844 16746 14900 16748
rect 14924 16746 14980 16748
rect 14684 16694 14710 16746
rect 14710 16694 14740 16746
rect 14764 16694 14774 16746
rect 14774 16694 14820 16746
rect 14844 16694 14890 16746
rect 14890 16694 14900 16746
rect 14924 16694 14954 16746
rect 14954 16694 14980 16746
rect 14684 16692 14740 16694
rect 14764 16692 14820 16694
rect 14844 16692 14900 16694
rect 14924 16692 14980 16694
rect 14684 15658 14740 15660
rect 14764 15658 14820 15660
rect 14844 15658 14900 15660
rect 14924 15658 14980 15660
rect 14684 15606 14710 15658
rect 14710 15606 14740 15658
rect 14764 15606 14774 15658
rect 14774 15606 14820 15658
rect 14844 15606 14890 15658
rect 14890 15606 14900 15658
rect 14924 15606 14954 15658
rect 14954 15606 14980 15658
rect 14684 15604 14740 15606
rect 14764 15604 14820 15606
rect 14844 15604 14900 15606
rect 14924 15604 14980 15606
rect 14684 14570 14740 14572
rect 14764 14570 14820 14572
rect 14844 14570 14900 14572
rect 14924 14570 14980 14572
rect 14684 14518 14710 14570
rect 14710 14518 14740 14570
rect 14764 14518 14774 14570
rect 14774 14518 14820 14570
rect 14844 14518 14890 14570
rect 14890 14518 14900 14570
rect 14924 14518 14954 14570
rect 14954 14518 14980 14570
rect 14684 14516 14740 14518
rect 14764 14516 14820 14518
rect 14844 14516 14900 14518
rect 14924 14516 14980 14518
rect 14684 13482 14740 13484
rect 14764 13482 14820 13484
rect 14844 13482 14900 13484
rect 14924 13482 14980 13484
rect 14684 13430 14710 13482
rect 14710 13430 14740 13482
rect 14764 13430 14774 13482
rect 14774 13430 14820 13482
rect 14844 13430 14890 13482
rect 14890 13430 14900 13482
rect 14924 13430 14954 13482
rect 14954 13430 14980 13482
rect 14684 13428 14740 13430
rect 14764 13428 14820 13430
rect 14844 13428 14900 13430
rect 14924 13428 14980 13430
rect 14684 12394 14740 12396
rect 14764 12394 14820 12396
rect 14844 12394 14900 12396
rect 14924 12394 14980 12396
rect 14684 12342 14710 12394
rect 14710 12342 14740 12394
rect 14764 12342 14774 12394
rect 14774 12342 14820 12394
rect 14844 12342 14890 12394
rect 14890 12342 14900 12394
rect 14924 12342 14954 12394
rect 14954 12342 14980 12394
rect 14684 12340 14740 12342
rect 14764 12340 14820 12342
rect 14844 12340 14900 12342
rect 14924 12340 14980 12342
rect 3606 5608 3662 5664
rect 4388 5322 4444 5324
rect 4468 5322 4524 5324
rect 4548 5322 4604 5324
rect 4628 5322 4684 5324
rect 4388 5270 4414 5322
rect 4414 5270 4444 5322
rect 4468 5270 4478 5322
rect 4478 5270 4524 5322
rect 4548 5270 4594 5322
rect 4594 5270 4604 5322
rect 4628 5270 4658 5322
rect 4658 5270 4684 5322
rect 4388 5268 4444 5270
rect 4468 5268 4524 5270
rect 4548 5268 4604 5270
rect 4628 5268 4684 5270
rect 11252 5322 11308 5324
rect 11332 5322 11388 5324
rect 11412 5322 11468 5324
rect 11492 5322 11548 5324
rect 11252 5270 11278 5322
rect 11278 5270 11308 5322
rect 11332 5270 11342 5322
rect 11342 5270 11388 5322
rect 11412 5270 11458 5322
rect 11458 5270 11468 5322
rect 11492 5270 11522 5322
rect 11522 5270 11548 5322
rect 11252 5268 11308 5270
rect 11332 5268 11388 5270
rect 11412 5268 11468 5270
rect 11492 5268 11548 5270
rect 7820 4778 7876 4780
rect 7900 4778 7956 4780
rect 7980 4778 8036 4780
rect 8060 4778 8116 4780
rect 7820 4726 7846 4778
rect 7846 4726 7876 4778
rect 7900 4726 7910 4778
rect 7910 4726 7956 4778
rect 7980 4726 8026 4778
rect 8026 4726 8036 4778
rect 8060 4726 8090 4778
rect 8090 4726 8116 4778
rect 7820 4724 7876 4726
rect 7900 4724 7956 4726
rect 7980 4724 8036 4726
rect 8060 4724 8116 4726
rect 4388 4234 4444 4236
rect 4468 4234 4524 4236
rect 4548 4234 4604 4236
rect 4628 4234 4684 4236
rect 4388 4182 4414 4234
rect 4414 4182 4444 4234
rect 4468 4182 4478 4234
rect 4478 4182 4524 4234
rect 4548 4182 4594 4234
rect 4594 4182 4604 4234
rect 4628 4182 4658 4234
rect 4658 4182 4684 4234
rect 4388 4180 4444 4182
rect 4468 4180 4524 4182
rect 4548 4180 4604 4182
rect 4628 4180 4684 4182
rect 11252 4234 11308 4236
rect 11332 4234 11388 4236
rect 11412 4234 11468 4236
rect 11492 4234 11548 4236
rect 11252 4182 11278 4234
rect 11278 4182 11308 4234
rect 11332 4182 11342 4234
rect 11342 4182 11388 4234
rect 11412 4182 11458 4234
rect 11458 4182 11468 4234
rect 11492 4182 11522 4234
rect 11522 4182 11548 4234
rect 11252 4180 11308 4182
rect 11332 4180 11388 4182
rect 11412 4180 11468 4182
rect 11492 4180 11548 4182
rect 14684 11306 14740 11308
rect 14764 11306 14820 11308
rect 14844 11306 14900 11308
rect 14924 11306 14980 11308
rect 14684 11254 14710 11306
rect 14710 11254 14740 11306
rect 14764 11254 14774 11306
rect 14774 11254 14820 11306
rect 14844 11254 14890 11306
rect 14890 11254 14900 11306
rect 14924 11254 14954 11306
rect 14954 11254 14980 11306
rect 14684 11252 14740 11254
rect 14764 11252 14820 11254
rect 14844 11252 14900 11254
rect 14924 11252 14980 11254
rect 14684 10218 14740 10220
rect 14764 10218 14820 10220
rect 14844 10218 14900 10220
rect 14924 10218 14980 10220
rect 14684 10166 14710 10218
rect 14710 10166 14740 10218
rect 14764 10166 14774 10218
rect 14774 10166 14820 10218
rect 14844 10166 14890 10218
rect 14890 10166 14900 10218
rect 14924 10166 14954 10218
rect 14954 10166 14980 10218
rect 14684 10164 14740 10166
rect 14764 10164 14820 10166
rect 14844 10164 14900 10166
rect 14924 10164 14980 10166
rect 18786 21384 18842 21440
rect 18970 20976 19026 21032
rect 18116 19466 18172 19468
rect 18196 19466 18252 19468
rect 18276 19466 18332 19468
rect 18356 19466 18412 19468
rect 18116 19414 18142 19466
rect 18142 19414 18172 19466
rect 18196 19414 18206 19466
rect 18206 19414 18252 19466
rect 18276 19414 18322 19466
rect 18322 19414 18332 19466
rect 18356 19414 18386 19466
rect 18386 19414 18412 19466
rect 18116 19412 18172 19414
rect 18196 19412 18252 19414
rect 18276 19412 18332 19414
rect 18356 19412 18412 19414
rect 14684 9130 14740 9132
rect 14764 9130 14820 9132
rect 14844 9130 14900 9132
rect 14924 9130 14980 9132
rect 14684 9078 14710 9130
rect 14710 9078 14740 9130
rect 14764 9078 14774 9130
rect 14774 9078 14820 9130
rect 14844 9078 14890 9130
rect 14890 9078 14900 9130
rect 14924 9078 14954 9130
rect 14954 9078 14980 9130
rect 14684 9076 14740 9078
rect 14764 9076 14820 9078
rect 14844 9076 14900 9078
rect 14924 9076 14980 9078
rect 14684 8042 14740 8044
rect 14764 8042 14820 8044
rect 14844 8042 14900 8044
rect 14924 8042 14980 8044
rect 14684 7990 14710 8042
rect 14710 7990 14740 8042
rect 14764 7990 14774 8042
rect 14774 7990 14820 8042
rect 14844 7990 14890 8042
rect 14890 7990 14900 8042
rect 14924 7990 14954 8042
rect 14954 7990 14980 8042
rect 14684 7988 14740 7990
rect 14764 7988 14820 7990
rect 14844 7988 14900 7990
rect 14924 7988 14980 7990
rect 14684 6954 14740 6956
rect 14764 6954 14820 6956
rect 14844 6954 14900 6956
rect 14924 6954 14980 6956
rect 14684 6902 14710 6954
rect 14710 6902 14740 6954
rect 14764 6902 14774 6954
rect 14774 6902 14820 6954
rect 14844 6902 14890 6954
rect 14890 6902 14900 6954
rect 14924 6902 14954 6954
rect 14954 6902 14980 6954
rect 14684 6900 14740 6902
rect 14764 6900 14820 6902
rect 14844 6900 14900 6902
rect 14924 6900 14980 6902
rect 14684 5866 14740 5868
rect 14764 5866 14820 5868
rect 14844 5866 14900 5868
rect 14924 5866 14980 5868
rect 14684 5814 14710 5866
rect 14710 5814 14740 5866
rect 14764 5814 14774 5866
rect 14774 5814 14820 5866
rect 14844 5814 14890 5866
rect 14890 5814 14900 5866
rect 14924 5814 14954 5866
rect 14954 5814 14980 5866
rect 14684 5812 14740 5814
rect 14764 5812 14820 5814
rect 14844 5812 14900 5814
rect 14924 5812 14980 5814
rect 14684 4778 14740 4780
rect 14764 4778 14820 4780
rect 14844 4778 14900 4780
rect 14924 4778 14980 4780
rect 14684 4726 14710 4778
rect 14710 4726 14740 4778
rect 14764 4726 14774 4778
rect 14774 4726 14820 4778
rect 14844 4726 14890 4778
rect 14890 4726 14900 4778
rect 14924 4726 14954 4778
rect 14954 4726 14980 4778
rect 14684 4724 14740 4726
rect 14764 4724 14820 4726
rect 14844 4724 14900 4726
rect 14924 4724 14980 4726
rect 7820 3690 7876 3692
rect 7900 3690 7956 3692
rect 7980 3690 8036 3692
rect 8060 3690 8116 3692
rect 7820 3638 7846 3690
rect 7846 3638 7876 3690
rect 7900 3638 7910 3690
rect 7910 3638 7956 3690
rect 7980 3638 8026 3690
rect 8026 3638 8036 3690
rect 8060 3638 8090 3690
rect 8090 3638 8116 3690
rect 7820 3636 7876 3638
rect 7900 3636 7956 3638
rect 7980 3636 8036 3638
rect 8060 3636 8116 3638
rect 14684 3690 14740 3692
rect 14764 3690 14820 3692
rect 14844 3690 14900 3692
rect 14924 3690 14980 3692
rect 14684 3638 14710 3690
rect 14710 3638 14740 3690
rect 14764 3638 14774 3690
rect 14774 3638 14820 3690
rect 14844 3638 14890 3690
rect 14890 3638 14900 3690
rect 14924 3638 14954 3690
rect 14954 3638 14980 3690
rect 14684 3636 14740 3638
rect 14764 3636 14820 3638
rect 14844 3636 14900 3638
rect 14924 3636 14980 3638
rect 4388 3146 4444 3148
rect 4468 3146 4524 3148
rect 4548 3146 4604 3148
rect 4628 3146 4684 3148
rect 4388 3094 4414 3146
rect 4414 3094 4444 3146
rect 4468 3094 4478 3146
rect 4478 3094 4524 3146
rect 4548 3094 4594 3146
rect 4594 3094 4604 3146
rect 4628 3094 4658 3146
rect 4658 3094 4684 3146
rect 4388 3092 4444 3094
rect 4468 3092 4524 3094
rect 4548 3092 4604 3094
rect 4628 3092 4684 3094
rect 11252 3146 11308 3148
rect 11332 3146 11388 3148
rect 11412 3146 11468 3148
rect 11492 3146 11548 3148
rect 11252 3094 11278 3146
rect 11278 3094 11308 3146
rect 11332 3094 11342 3146
rect 11342 3094 11388 3146
rect 11412 3094 11458 3146
rect 11458 3094 11468 3146
rect 11492 3094 11522 3146
rect 11522 3094 11548 3146
rect 11252 3092 11308 3094
rect 11332 3092 11388 3094
rect 11412 3092 11468 3094
rect 11492 3092 11548 3094
rect 7820 2602 7876 2604
rect 7900 2602 7956 2604
rect 7980 2602 8036 2604
rect 8060 2602 8116 2604
rect 7820 2550 7846 2602
rect 7846 2550 7876 2602
rect 7900 2550 7910 2602
rect 7910 2550 7956 2602
rect 7980 2550 8026 2602
rect 8026 2550 8036 2602
rect 8060 2550 8090 2602
rect 8090 2550 8116 2602
rect 7820 2548 7876 2550
rect 7900 2548 7956 2550
rect 7980 2548 8036 2550
rect 8060 2548 8116 2550
rect 14684 2602 14740 2604
rect 14764 2602 14820 2604
rect 14844 2602 14900 2604
rect 14924 2602 14980 2604
rect 14684 2550 14710 2602
rect 14710 2550 14740 2602
rect 14764 2550 14774 2602
rect 14774 2550 14820 2602
rect 14844 2550 14890 2602
rect 14890 2550 14900 2602
rect 14924 2550 14954 2602
rect 14954 2550 14980 2602
rect 14684 2548 14740 2550
rect 14764 2548 14820 2550
rect 14844 2548 14900 2550
rect 14924 2548 14980 2550
rect 4388 2058 4444 2060
rect 4468 2058 4524 2060
rect 4548 2058 4604 2060
rect 4628 2058 4684 2060
rect 4388 2006 4414 2058
rect 4414 2006 4444 2058
rect 4468 2006 4478 2058
rect 4478 2006 4524 2058
rect 4548 2006 4594 2058
rect 4594 2006 4604 2058
rect 4628 2006 4658 2058
rect 4658 2006 4684 2058
rect 4388 2004 4444 2006
rect 4468 2004 4524 2006
rect 4548 2004 4604 2006
rect 4628 2004 4684 2006
rect 11252 2058 11308 2060
rect 11332 2058 11388 2060
rect 11412 2058 11468 2060
rect 11492 2058 11548 2060
rect 11252 2006 11278 2058
rect 11278 2006 11308 2058
rect 11332 2006 11342 2058
rect 11342 2006 11388 2058
rect 11412 2006 11458 2058
rect 11458 2006 11468 2058
rect 11492 2006 11522 2058
rect 11522 2006 11548 2058
rect 11252 2004 11308 2006
rect 11332 2004 11388 2006
rect 11412 2004 11468 2006
rect 11492 2004 11548 2006
rect 16762 15300 16764 15320
rect 16764 15300 16816 15320
rect 16816 15300 16818 15320
rect 16762 15264 16818 15300
rect 18116 18378 18172 18380
rect 18196 18378 18252 18380
rect 18276 18378 18332 18380
rect 18356 18378 18412 18380
rect 18116 18326 18142 18378
rect 18142 18326 18172 18378
rect 18196 18326 18206 18378
rect 18206 18326 18252 18378
rect 18276 18326 18322 18378
rect 18322 18326 18332 18378
rect 18356 18326 18386 18378
rect 18386 18326 18412 18378
rect 18116 18324 18172 18326
rect 18196 18324 18252 18326
rect 18276 18324 18332 18326
rect 18356 18324 18412 18326
rect 18116 17290 18172 17292
rect 18196 17290 18252 17292
rect 18276 17290 18332 17292
rect 18356 17290 18412 17292
rect 18116 17238 18142 17290
rect 18142 17238 18172 17290
rect 18196 17238 18206 17290
rect 18206 17238 18252 17290
rect 18276 17238 18322 17290
rect 18322 17238 18332 17290
rect 18356 17238 18386 17290
rect 18386 17238 18412 17290
rect 18116 17236 18172 17238
rect 18196 17236 18252 17238
rect 18276 17236 18332 17238
rect 18356 17236 18412 17238
rect 18116 16202 18172 16204
rect 18196 16202 18252 16204
rect 18276 16202 18332 16204
rect 18356 16202 18412 16204
rect 18116 16150 18142 16202
rect 18142 16150 18172 16202
rect 18196 16150 18206 16202
rect 18206 16150 18252 16202
rect 18276 16150 18322 16202
rect 18322 16150 18332 16202
rect 18356 16150 18386 16202
rect 18386 16150 18412 16202
rect 18116 16148 18172 16150
rect 18196 16148 18252 16150
rect 18276 16148 18332 16150
rect 18356 16148 18412 16150
rect 18116 15114 18172 15116
rect 18196 15114 18252 15116
rect 18276 15114 18332 15116
rect 18356 15114 18412 15116
rect 18116 15062 18142 15114
rect 18142 15062 18172 15114
rect 18196 15062 18206 15114
rect 18206 15062 18252 15114
rect 18276 15062 18322 15114
rect 18322 15062 18332 15114
rect 18356 15062 18386 15114
rect 18386 15062 18412 15114
rect 18116 15060 18172 15062
rect 18196 15060 18252 15062
rect 18276 15060 18332 15062
rect 18356 15060 18412 15062
rect 18878 19208 18934 19264
rect 19338 21928 19394 21984
rect 19614 18256 19670 18312
rect 18116 14026 18172 14028
rect 18196 14026 18252 14028
rect 18276 14026 18332 14028
rect 18356 14026 18412 14028
rect 18116 13974 18142 14026
rect 18142 13974 18172 14026
rect 18196 13974 18206 14026
rect 18206 13974 18252 14026
rect 18276 13974 18322 14026
rect 18322 13974 18332 14026
rect 18356 13974 18386 14026
rect 18386 13974 18412 14026
rect 18116 13972 18172 13974
rect 18196 13972 18252 13974
rect 18276 13972 18332 13974
rect 18356 13972 18412 13974
rect 18116 12938 18172 12940
rect 18196 12938 18252 12940
rect 18276 12938 18332 12940
rect 18356 12938 18412 12940
rect 18116 12886 18142 12938
rect 18142 12886 18172 12938
rect 18196 12886 18206 12938
rect 18206 12886 18252 12938
rect 18276 12886 18322 12938
rect 18322 12886 18332 12938
rect 18356 12886 18386 12938
rect 18386 12886 18412 12938
rect 18116 12884 18172 12886
rect 18196 12884 18252 12886
rect 18276 12884 18332 12886
rect 18356 12884 18412 12886
rect 17774 3568 17830 3624
rect 18116 11850 18172 11852
rect 18196 11850 18252 11852
rect 18276 11850 18332 11852
rect 18356 11850 18412 11852
rect 18116 11798 18142 11850
rect 18142 11798 18172 11850
rect 18196 11798 18206 11850
rect 18206 11798 18252 11850
rect 18276 11798 18322 11850
rect 18322 11798 18332 11850
rect 18356 11798 18386 11850
rect 18386 11798 18412 11850
rect 18116 11796 18172 11798
rect 18196 11796 18252 11798
rect 18276 11796 18332 11798
rect 18356 11796 18412 11798
rect 18116 10762 18172 10764
rect 18196 10762 18252 10764
rect 18276 10762 18332 10764
rect 18356 10762 18412 10764
rect 18116 10710 18142 10762
rect 18142 10710 18172 10762
rect 18196 10710 18206 10762
rect 18206 10710 18252 10762
rect 18276 10710 18322 10762
rect 18322 10710 18332 10762
rect 18356 10710 18386 10762
rect 18386 10710 18412 10762
rect 18116 10708 18172 10710
rect 18196 10708 18252 10710
rect 18276 10708 18332 10710
rect 18356 10708 18412 10710
rect 19798 13768 19854 13824
rect 19706 13224 19762 13280
rect 19798 12816 19854 12872
rect 18116 9674 18172 9676
rect 18196 9674 18252 9676
rect 18276 9674 18332 9676
rect 18356 9674 18412 9676
rect 18116 9622 18142 9674
rect 18142 9622 18172 9674
rect 18196 9622 18206 9674
rect 18206 9622 18252 9674
rect 18276 9622 18322 9674
rect 18322 9622 18332 9674
rect 18356 9622 18386 9674
rect 18386 9622 18412 9674
rect 18116 9620 18172 9622
rect 18196 9620 18252 9622
rect 18276 9620 18332 9622
rect 18356 9620 18412 9622
rect 18116 8586 18172 8588
rect 18196 8586 18252 8588
rect 18276 8586 18332 8588
rect 18356 8586 18412 8588
rect 18116 8534 18142 8586
rect 18142 8534 18172 8586
rect 18196 8534 18206 8586
rect 18206 8534 18252 8586
rect 18276 8534 18322 8586
rect 18322 8534 18332 8586
rect 18356 8534 18386 8586
rect 18386 8534 18412 8586
rect 18116 8532 18172 8534
rect 18196 8532 18252 8534
rect 18276 8532 18332 8534
rect 18356 8532 18412 8534
rect 18116 7498 18172 7500
rect 18196 7498 18252 7500
rect 18276 7498 18332 7500
rect 18356 7498 18412 7500
rect 18116 7446 18142 7498
rect 18142 7446 18172 7498
rect 18196 7446 18206 7498
rect 18206 7446 18252 7498
rect 18276 7446 18322 7498
rect 18322 7446 18332 7498
rect 18356 7446 18386 7498
rect 18386 7446 18412 7498
rect 18116 7444 18172 7446
rect 18196 7444 18252 7446
rect 18276 7444 18332 7446
rect 18356 7444 18412 7446
rect 18116 6410 18172 6412
rect 18196 6410 18252 6412
rect 18276 6410 18332 6412
rect 18356 6410 18412 6412
rect 18116 6358 18142 6410
rect 18142 6358 18172 6410
rect 18196 6358 18206 6410
rect 18206 6358 18252 6410
rect 18276 6358 18322 6410
rect 18322 6358 18332 6410
rect 18356 6358 18386 6410
rect 18386 6358 18412 6410
rect 18116 6356 18172 6358
rect 18196 6356 18252 6358
rect 18276 6356 18332 6358
rect 18356 6356 18412 6358
rect 17958 5880 18014 5936
rect 18602 6424 18658 6480
rect 18510 5472 18566 5528
rect 18116 5322 18172 5324
rect 18196 5322 18252 5324
rect 18276 5322 18332 5324
rect 18356 5322 18412 5324
rect 18116 5270 18142 5322
rect 18142 5270 18172 5322
rect 18196 5270 18206 5322
rect 18206 5270 18252 5322
rect 18276 5270 18322 5322
rect 18322 5270 18332 5322
rect 18356 5270 18386 5322
rect 18386 5270 18412 5322
rect 18116 5268 18172 5270
rect 18196 5268 18252 5270
rect 18276 5268 18332 5270
rect 18356 5268 18412 5270
rect 17958 4928 18014 4984
rect 18050 4520 18106 4576
rect 18116 4234 18172 4236
rect 18196 4234 18252 4236
rect 18276 4234 18332 4236
rect 18356 4234 18412 4236
rect 18116 4182 18142 4234
rect 18142 4182 18172 4234
rect 18196 4182 18206 4234
rect 18206 4182 18252 4234
rect 18276 4182 18322 4234
rect 18322 4182 18332 4234
rect 18356 4182 18386 4234
rect 18386 4182 18412 4234
rect 18116 4180 18172 4182
rect 18196 4180 18252 4182
rect 18276 4180 18332 4182
rect 18356 4180 18412 4182
rect 18510 3160 18566 3216
rect 18116 3146 18172 3148
rect 18196 3146 18252 3148
rect 18276 3146 18332 3148
rect 18356 3146 18412 3148
rect 18116 3094 18142 3146
rect 18142 3094 18172 3146
rect 18196 3094 18206 3146
rect 18206 3094 18252 3146
rect 18276 3094 18322 3146
rect 18322 3094 18332 3146
rect 18356 3094 18386 3146
rect 18386 3094 18412 3146
rect 18116 3092 18172 3094
rect 18196 3092 18252 3094
rect 18276 3092 18332 3094
rect 18356 3092 18412 3094
rect 17866 2752 17922 2808
rect 18116 2058 18172 2060
rect 18196 2058 18252 2060
rect 18276 2058 18332 2060
rect 18356 2058 18412 2060
rect 18116 2006 18142 2058
rect 18142 2006 18172 2058
rect 18196 2006 18206 2058
rect 18206 2006 18252 2058
rect 18276 2006 18322 2058
rect 18322 2006 18332 2058
rect 18356 2006 18386 2058
rect 18386 2006 18412 2058
rect 18116 2004 18172 2006
rect 18196 2004 18252 2006
rect 18276 2004 18332 2006
rect 18356 2004 18412 2006
rect 18786 9960 18842 10016
rect 18878 2208 18934 2264
rect 18786 1800 18842 1856
rect 18694 1392 18750 1448
rect 17314 440 17370 496
rect 19706 12272 19762 12328
rect 20074 20568 20130 20624
rect 20626 20024 20682 20080
rect 20718 19616 20774 19672
rect 20534 18664 20590 18720
rect 20166 16896 20222 16952
rect 20442 17884 20444 17904
rect 20444 17884 20496 17904
rect 20496 17884 20498 17904
rect 20442 17848 20498 17884
rect 20442 15980 20444 16000
rect 20444 15980 20496 16000
rect 20496 15980 20498 16000
rect 20442 15944 20498 15980
rect 20442 15012 20498 15048
rect 20442 14992 20444 15012
rect 20444 14992 20496 15012
rect 20496 14992 20498 15012
rect 20718 17340 20720 17360
rect 20720 17340 20772 17360
rect 20772 17340 20774 17360
rect 20718 17304 20774 17340
rect 20626 16352 20682 16408
rect 20718 15556 20774 15592
rect 20718 15536 20720 15556
rect 20720 15536 20772 15556
rect 20772 15536 20774 15556
rect 20442 14584 20498 14640
rect 20258 11864 20314 11920
rect 19982 11456 20038 11512
rect 20258 10912 20314 10968
rect 20258 9552 20314 9608
rect 20718 13632 20774 13688
rect 20534 10504 20590 10560
rect 20534 9144 20590 9200
rect 20258 8600 20314 8656
rect 20534 8192 20590 8248
rect 20258 7784 20314 7840
rect 19982 7240 20038 7296
rect 20534 6832 20590 6888
rect 21086 14176 21142 14232
rect 20534 4112 20590 4168
rect 19062 848 19118 904
rect 18142 32 18198 88
<< metal3 >>
rect 17953 22394 18019 22397
rect 22320 22394 22800 22424
rect 17953 22392 22800 22394
rect 17953 22336 17958 22392
rect 18014 22336 22800 22392
rect 17953 22334 22800 22336
rect 17953 22331 18019 22334
rect 22320 22304 22800 22334
rect 19333 21986 19399 21989
rect 22320 21986 22800 22016
rect 19333 21984 22800 21986
rect 19333 21928 19338 21984
rect 19394 21928 22800 21984
rect 19333 21926 22800 21928
rect 19333 21923 19399 21926
rect 22320 21896 22800 21926
rect 18781 21442 18847 21445
rect 22320 21442 22800 21472
rect 18781 21440 22800 21442
rect 18781 21384 18786 21440
rect 18842 21384 22800 21440
rect 18781 21382 22800 21384
rect 18781 21379 18847 21382
rect 22320 21352 22800 21382
rect 18965 21034 19031 21037
rect 22320 21034 22800 21064
rect 18965 21032 22800 21034
rect 18965 20976 18970 21032
rect 19026 20976 22800 21032
rect 18965 20974 22800 20976
rect 18965 20971 19031 20974
rect 22320 20944 22800 20974
rect 20069 20626 20135 20629
rect 22320 20626 22800 20656
rect 20069 20624 22800 20626
rect 20069 20568 20074 20624
rect 20130 20568 22800 20624
rect 20069 20566 22800 20568
rect 20069 20563 20135 20566
rect 22320 20536 22800 20566
rect 20621 20082 20687 20085
rect 22320 20082 22800 20112
rect 20621 20080 22800 20082
rect 20621 20024 20626 20080
rect 20682 20024 22800 20080
rect 20621 20022 22800 20024
rect 20621 20019 20687 20022
rect 7808 20016 8128 20017
rect 7808 19952 7816 20016
rect 7880 19952 7896 20016
rect 7960 19952 7976 20016
rect 8040 19952 8056 20016
rect 8120 19952 8128 20016
rect 7808 19951 8128 19952
rect 14672 20016 14992 20017
rect 14672 19952 14680 20016
rect 14744 19952 14760 20016
rect 14824 19952 14840 20016
rect 14904 19952 14920 20016
rect 14984 19952 14992 20016
rect 22320 19992 22800 20022
rect 14672 19951 14992 19952
rect 20713 19674 20779 19677
rect 22320 19674 22800 19704
rect 20713 19672 22800 19674
rect 20713 19616 20718 19672
rect 20774 19616 22800 19672
rect 20713 19614 22800 19616
rect 20713 19611 20779 19614
rect 22320 19584 22800 19614
rect 4376 19472 4696 19473
rect 4376 19408 4384 19472
rect 4448 19408 4464 19472
rect 4528 19408 4544 19472
rect 4608 19408 4624 19472
rect 4688 19408 4696 19472
rect 4376 19407 4696 19408
rect 11240 19472 11560 19473
rect 11240 19408 11248 19472
rect 11312 19408 11328 19472
rect 11392 19408 11408 19472
rect 11472 19408 11488 19472
rect 11552 19408 11560 19472
rect 11240 19407 11560 19408
rect 18104 19472 18424 19473
rect 18104 19408 18112 19472
rect 18176 19408 18192 19472
rect 18256 19408 18272 19472
rect 18336 19408 18352 19472
rect 18416 19408 18424 19472
rect 18104 19407 18424 19408
rect 18873 19266 18939 19269
rect 22320 19266 22800 19296
rect 18873 19264 22800 19266
rect 18873 19208 18878 19264
rect 18934 19208 22800 19264
rect 18873 19206 22800 19208
rect 18873 19203 18939 19206
rect 22320 19176 22800 19206
rect 7808 18928 8128 18929
rect 7808 18864 7816 18928
rect 7880 18864 7896 18928
rect 7960 18864 7976 18928
rect 8040 18864 8056 18928
rect 8120 18864 8128 18928
rect 7808 18863 8128 18864
rect 14672 18928 14992 18929
rect 14672 18864 14680 18928
rect 14744 18864 14760 18928
rect 14824 18864 14840 18928
rect 14904 18864 14920 18928
rect 14984 18864 14992 18928
rect 14672 18863 14992 18864
rect 20529 18722 20595 18725
rect 22320 18722 22800 18752
rect 20529 18720 22800 18722
rect 20529 18664 20534 18720
rect 20590 18664 22800 18720
rect 20529 18662 22800 18664
rect 20529 18659 20595 18662
rect 22320 18632 22800 18662
rect 4376 18384 4696 18385
rect 4376 18320 4384 18384
rect 4448 18320 4464 18384
rect 4528 18320 4544 18384
rect 4608 18320 4624 18384
rect 4688 18320 4696 18384
rect 4376 18319 4696 18320
rect 11240 18384 11560 18385
rect 11240 18320 11248 18384
rect 11312 18320 11328 18384
rect 11392 18320 11408 18384
rect 11472 18320 11488 18384
rect 11552 18320 11560 18384
rect 11240 18319 11560 18320
rect 18104 18384 18424 18385
rect 18104 18320 18112 18384
rect 18176 18320 18192 18384
rect 18256 18320 18272 18384
rect 18336 18320 18352 18384
rect 18416 18320 18424 18384
rect 18104 18319 18424 18320
rect 19609 18314 19675 18317
rect 22320 18314 22800 18344
rect 19609 18312 22800 18314
rect 19609 18256 19614 18312
rect 19670 18256 22800 18312
rect 19609 18254 22800 18256
rect 19609 18251 19675 18254
rect 22320 18224 22800 18254
rect 12709 18042 12775 18045
rect 13353 18042 13419 18045
rect 12709 18040 13419 18042
rect 12709 17984 12714 18040
rect 12770 17984 13358 18040
rect 13414 17984 13419 18040
rect 12709 17982 13419 17984
rect 12709 17979 12775 17982
rect 13353 17979 13419 17982
rect 20437 17906 20503 17909
rect 22320 17906 22800 17936
rect 20437 17904 22800 17906
rect 20437 17848 20442 17904
rect 20498 17848 22800 17904
rect 20437 17846 22800 17848
rect 20437 17843 20503 17846
rect 7808 17840 8128 17841
rect 7808 17776 7816 17840
rect 7880 17776 7896 17840
rect 7960 17776 7976 17840
rect 8040 17776 8056 17840
rect 8120 17776 8128 17840
rect 7808 17775 8128 17776
rect 14672 17840 14992 17841
rect 14672 17776 14680 17840
rect 14744 17776 14760 17840
rect 14824 17776 14840 17840
rect 14904 17776 14920 17840
rect 14984 17776 14992 17840
rect 22320 17816 22800 17846
rect 14672 17775 14992 17776
rect 20713 17362 20779 17365
rect 22320 17362 22800 17392
rect 20713 17360 22800 17362
rect 20713 17304 20718 17360
rect 20774 17304 22800 17360
rect 20713 17302 22800 17304
rect 20713 17299 20779 17302
rect 4376 17296 4696 17297
rect 4376 17232 4384 17296
rect 4448 17232 4464 17296
rect 4528 17232 4544 17296
rect 4608 17232 4624 17296
rect 4688 17232 4696 17296
rect 4376 17231 4696 17232
rect 11240 17296 11560 17297
rect 11240 17232 11248 17296
rect 11312 17232 11328 17296
rect 11392 17232 11408 17296
rect 11472 17232 11488 17296
rect 11552 17232 11560 17296
rect 11240 17231 11560 17232
rect 18104 17296 18424 17297
rect 18104 17232 18112 17296
rect 18176 17232 18192 17296
rect 18256 17232 18272 17296
rect 18336 17232 18352 17296
rect 18416 17232 18424 17296
rect 22320 17272 22800 17302
rect 18104 17231 18424 17232
rect 0 17090 480 17120
rect 9581 17090 9647 17093
rect 0 17088 9647 17090
rect 0 17032 9586 17088
rect 9642 17032 9647 17088
rect 0 17030 9647 17032
rect 0 17000 480 17030
rect 9581 17027 9647 17030
rect 20161 16954 20227 16957
rect 22320 16954 22800 16984
rect 20161 16952 22800 16954
rect 20161 16896 20166 16952
rect 20222 16896 22800 16952
rect 20161 16894 22800 16896
rect 20161 16891 20227 16894
rect 22320 16864 22800 16894
rect 7808 16752 8128 16753
rect 7808 16688 7816 16752
rect 7880 16688 7896 16752
rect 7960 16688 7976 16752
rect 8040 16688 8056 16752
rect 8120 16688 8128 16752
rect 7808 16687 8128 16688
rect 14672 16752 14992 16753
rect 14672 16688 14680 16752
rect 14744 16688 14760 16752
rect 14824 16688 14840 16752
rect 14904 16688 14920 16752
rect 14984 16688 14992 16752
rect 14672 16687 14992 16688
rect 20621 16410 20687 16413
rect 22320 16410 22800 16440
rect 20621 16408 22800 16410
rect 20621 16352 20626 16408
rect 20682 16352 22800 16408
rect 20621 16350 22800 16352
rect 20621 16347 20687 16350
rect 22320 16320 22800 16350
rect 4376 16208 4696 16209
rect 4376 16144 4384 16208
rect 4448 16144 4464 16208
rect 4528 16144 4544 16208
rect 4608 16144 4624 16208
rect 4688 16144 4696 16208
rect 4376 16143 4696 16144
rect 11240 16208 11560 16209
rect 11240 16144 11248 16208
rect 11312 16144 11328 16208
rect 11392 16144 11408 16208
rect 11472 16144 11488 16208
rect 11552 16144 11560 16208
rect 11240 16143 11560 16144
rect 18104 16208 18424 16209
rect 18104 16144 18112 16208
rect 18176 16144 18192 16208
rect 18256 16144 18272 16208
rect 18336 16144 18352 16208
rect 18416 16144 18424 16208
rect 18104 16143 18424 16144
rect 20437 16002 20503 16005
rect 22320 16002 22800 16032
rect 20437 16000 22800 16002
rect 20437 15944 20442 16000
rect 20498 15944 22800 16000
rect 20437 15942 22800 15944
rect 20437 15939 20503 15942
rect 22320 15912 22800 15942
rect 7808 15664 8128 15665
rect 7808 15600 7816 15664
rect 7880 15600 7896 15664
rect 7960 15600 7976 15664
rect 8040 15600 8056 15664
rect 8120 15600 8128 15664
rect 7808 15599 8128 15600
rect 14672 15664 14992 15665
rect 14672 15600 14680 15664
rect 14744 15600 14760 15664
rect 14824 15600 14840 15664
rect 14904 15600 14920 15664
rect 14984 15600 14992 15664
rect 14672 15599 14992 15600
rect 20713 15594 20779 15597
rect 22320 15594 22800 15624
rect 20713 15592 22800 15594
rect 20713 15536 20718 15592
rect 20774 15536 22800 15592
rect 20713 15534 22800 15536
rect 20713 15531 20779 15534
rect 22320 15504 22800 15534
rect 12157 15322 12223 15325
rect 16757 15322 16823 15325
rect 12157 15320 16823 15322
rect 12157 15264 12162 15320
rect 12218 15264 16762 15320
rect 16818 15264 16823 15320
rect 12157 15262 16823 15264
rect 12157 15259 12223 15262
rect 16757 15259 16823 15262
rect 4376 15120 4696 15121
rect 4376 15056 4384 15120
rect 4448 15056 4464 15120
rect 4528 15056 4544 15120
rect 4608 15056 4624 15120
rect 4688 15056 4696 15120
rect 4376 15055 4696 15056
rect 11240 15120 11560 15121
rect 11240 15056 11248 15120
rect 11312 15056 11328 15120
rect 11392 15056 11408 15120
rect 11472 15056 11488 15120
rect 11552 15056 11560 15120
rect 11240 15055 11560 15056
rect 18104 15120 18424 15121
rect 18104 15056 18112 15120
rect 18176 15056 18192 15120
rect 18256 15056 18272 15120
rect 18336 15056 18352 15120
rect 18416 15056 18424 15120
rect 18104 15055 18424 15056
rect 20437 15050 20503 15053
rect 22320 15050 22800 15080
rect 20437 15048 22800 15050
rect 20437 14992 20442 15048
rect 20498 14992 22800 15048
rect 20437 14990 22800 14992
rect 20437 14987 20503 14990
rect 22320 14960 22800 14990
rect 20437 14642 20503 14645
rect 22320 14642 22800 14672
rect 20437 14640 22800 14642
rect 20437 14584 20442 14640
rect 20498 14584 22800 14640
rect 20437 14582 22800 14584
rect 20437 14579 20503 14582
rect 7808 14576 8128 14577
rect 7808 14512 7816 14576
rect 7880 14512 7896 14576
rect 7960 14512 7976 14576
rect 8040 14512 8056 14576
rect 8120 14512 8128 14576
rect 7808 14511 8128 14512
rect 14672 14576 14992 14577
rect 14672 14512 14680 14576
rect 14744 14512 14760 14576
rect 14824 14512 14840 14576
rect 14904 14512 14920 14576
rect 14984 14512 14992 14576
rect 22320 14552 22800 14582
rect 14672 14511 14992 14512
rect 21081 14234 21147 14237
rect 22320 14234 22800 14264
rect 21081 14232 22800 14234
rect 21081 14176 21086 14232
rect 21142 14176 22800 14232
rect 21081 14174 22800 14176
rect 21081 14171 21147 14174
rect 22320 14144 22800 14174
rect 4376 14032 4696 14033
rect 4376 13968 4384 14032
rect 4448 13968 4464 14032
rect 4528 13968 4544 14032
rect 4608 13968 4624 14032
rect 4688 13968 4696 14032
rect 4376 13967 4696 13968
rect 11240 14032 11560 14033
rect 11240 13968 11248 14032
rect 11312 13968 11328 14032
rect 11392 13968 11408 14032
rect 11472 13968 11488 14032
rect 11552 13968 11560 14032
rect 11240 13967 11560 13968
rect 18104 14032 18424 14033
rect 18104 13968 18112 14032
rect 18176 13968 18192 14032
rect 18256 13968 18272 14032
rect 18336 13968 18352 14032
rect 18416 13968 18424 14032
rect 18104 13967 18424 13968
rect 9857 13826 9923 13829
rect 19793 13826 19859 13829
rect 9857 13824 19859 13826
rect 9857 13768 9862 13824
rect 9918 13768 19798 13824
rect 19854 13768 19859 13824
rect 9857 13766 19859 13768
rect 9857 13763 9923 13766
rect 19793 13763 19859 13766
rect 20713 13690 20779 13693
rect 22320 13690 22800 13720
rect 20713 13688 22800 13690
rect 20713 13632 20718 13688
rect 20774 13632 22800 13688
rect 20713 13630 22800 13632
rect 20713 13627 20779 13630
rect 22320 13600 22800 13630
rect 7808 13488 8128 13489
rect 7808 13424 7816 13488
rect 7880 13424 7896 13488
rect 7960 13424 7976 13488
rect 8040 13424 8056 13488
rect 8120 13424 8128 13488
rect 7808 13423 8128 13424
rect 14672 13488 14992 13489
rect 14672 13424 14680 13488
rect 14744 13424 14760 13488
rect 14824 13424 14840 13488
rect 14904 13424 14920 13488
rect 14984 13424 14992 13488
rect 14672 13423 14992 13424
rect 19701 13282 19767 13285
rect 22320 13282 22800 13312
rect 19701 13280 22800 13282
rect 19701 13224 19706 13280
rect 19762 13224 22800 13280
rect 19701 13222 22800 13224
rect 19701 13219 19767 13222
rect 22320 13192 22800 13222
rect 4376 12944 4696 12945
rect 4376 12880 4384 12944
rect 4448 12880 4464 12944
rect 4528 12880 4544 12944
rect 4608 12880 4624 12944
rect 4688 12880 4696 12944
rect 4376 12879 4696 12880
rect 11240 12944 11560 12945
rect 11240 12880 11248 12944
rect 11312 12880 11328 12944
rect 11392 12880 11408 12944
rect 11472 12880 11488 12944
rect 11552 12880 11560 12944
rect 11240 12879 11560 12880
rect 18104 12944 18424 12945
rect 18104 12880 18112 12944
rect 18176 12880 18192 12944
rect 18256 12880 18272 12944
rect 18336 12880 18352 12944
rect 18416 12880 18424 12944
rect 18104 12879 18424 12880
rect 19793 12874 19859 12877
rect 22320 12874 22800 12904
rect 19793 12872 22800 12874
rect 19793 12816 19798 12872
rect 19854 12816 22800 12872
rect 19793 12814 22800 12816
rect 19793 12811 19859 12814
rect 22320 12784 22800 12814
rect 7808 12400 8128 12401
rect 7808 12336 7816 12400
rect 7880 12336 7896 12400
rect 7960 12336 7976 12400
rect 8040 12336 8056 12400
rect 8120 12336 8128 12400
rect 7808 12335 8128 12336
rect 14672 12400 14992 12401
rect 14672 12336 14680 12400
rect 14744 12336 14760 12400
rect 14824 12336 14840 12400
rect 14904 12336 14920 12400
rect 14984 12336 14992 12400
rect 14672 12335 14992 12336
rect 19701 12330 19767 12333
rect 22320 12330 22800 12360
rect 19701 12328 22800 12330
rect 19701 12272 19706 12328
rect 19762 12272 22800 12328
rect 19701 12270 22800 12272
rect 19701 12267 19767 12270
rect 22320 12240 22800 12270
rect 20253 11922 20319 11925
rect 22320 11922 22800 11952
rect 20253 11920 22800 11922
rect 20253 11864 20258 11920
rect 20314 11864 22800 11920
rect 20253 11862 22800 11864
rect 20253 11859 20319 11862
rect 4376 11856 4696 11857
rect 4376 11792 4384 11856
rect 4448 11792 4464 11856
rect 4528 11792 4544 11856
rect 4608 11792 4624 11856
rect 4688 11792 4696 11856
rect 4376 11791 4696 11792
rect 11240 11856 11560 11857
rect 11240 11792 11248 11856
rect 11312 11792 11328 11856
rect 11392 11792 11408 11856
rect 11472 11792 11488 11856
rect 11552 11792 11560 11856
rect 11240 11791 11560 11792
rect 18104 11856 18424 11857
rect 18104 11792 18112 11856
rect 18176 11792 18192 11856
rect 18256 11792 18272 11856
rect 18336 11792 18352 11856
rect 18416 11792 18424 11856
rect 22320 11832 22800 11862
rect 18104 11791 18424 11792
rect 19977 11514 20043 11517
rect 22320 11514 22800 11544
rect 19977 11512 22800 11514
rect 19977 11456 19982 11512
rect 20038 11456 22800 11512
rect 19977 11454 22800 11456
rect 19977 11451 20043 11454
rect 22320 11424 22800 11454
rect 7808 11312 8128 11313
rect 7808 11248 7816 11312
rect 7880 11248 7896 11312
rect 7960 11248 7976 11312
rect 8040 11248 8056 11312
rect 8120 11248 8128 11312
rect 7808 11247 8128 11248
rect 14672 11312 14992 11313
rect 14672 11248 14680 11312
rect 14744 11248 14760 11312
rect 14824 11248 14840 11312
rect 14904 11248 14920 11312
rect 14984 11248 14992 11312
rect 14672 11247 14992 11248
rect 20253 10970 20319 10973
rect 22320 10970 22800 11000
rect 20253 10968 22800 10970
rect 20253 10912 20258 10968
rect 20314 10912 22800 10968
rect 20253 10910 22800 10912
rect 20253 10907 20319 10910
rect 22320 10880 22800 10910
rect 4376 10768 4696 10769
rect 4376 10704 4384 10768
rect 4448 10704 4464 10768
rect 4528 10704 4544 10768
rect 4608 10704 4624 10768
rect 4688 10704 4696 10768
rect 4376 10703 4696 10704
rect 11240 10768 11560 10769
rect 11240 10704 11248 10768
rect 11312 10704 11328 10768
rect 11392 10704 11408 10768
rect 11472 10704 11488 10768
rect 11552 10704 11560 10768
rect 11240 10703 11560 10704
rect 18104 10768 18424 10769
rect 18104 10704 18112 10768
rect 18176 10704 18192 10768
rect 18256 10704 18272 10768
rect 18336 10704 18352 10768
rect 18416 10704 18424 10768
rect 18104 10703 18424 10704
rect 20529 10562 20595 10565
rect 22320 10562 22800 10592
rect 20529 10560 22800 10562
rect 20529 10504 20534 10560
rect 20590 10504 22800 10560
rect 20529 10502 22800 10504
rect 20529 10499 20595 10502
rect 22320 10472 22800 10502
rect 7808 10224 8128 10225
rect 7808 10160 7816 10224
rect 7880 10160 7896 10224
rect 7960 10160 7976 10224
rect 8040 10160 8056 10224
rect 8120 10160 8128 10224
rect 7808 10159 8128 10160
rect 14672 10224 14992 10225
rect 14672 10160 14680 10224
rect 14744 10160 14760 10224
rect 14824 10160 14840 10224
rect 14904 10160 14920 10224
rect 14984 10160 14992 10224
rect 14672 10159 14992 10160
rect 18781 10018 18847 10021
rect 22320 10018 22800 10048
rect 18781 10016 22800 10018
rect 18781 9960 18786 10016
rect 18842 9960 22800 10016
rect 18781 9958 22800 9960
rect 18781 9955 18847 9958
rect 22320 9928 22800 9958
rect 4376 9680 4696 9681
rect 4376 9616 4384 9680
rect 4448 9616 4464 9680
rect 4528 9616 4544 9680
rect 4608 9616 4624 9680
rect 4688 9616 4696 9680
rect 4376 9615 4696 9616
rect 11240 9680 11560 9681
rect 11240 9616 11248 9680
rect 11312 9616 11328 9680
rect 11392 9616 11408 9680
rect 11472 9616 11488 9680
rect 11552 9616 11560 9680
rect 11240 9615 11560 9616
rect 18104 9680 18424 9681
rect 18104 9616 18112 9680
rect 18176 9616 18192 9680
rect 18256 9616 18272 9680
rect 18336 9616 18352 9680
rect 18416 9616 18424 9680
rect 18104 9615 18424 9616
rect 20253 9610 20319 9613
rect 22320 9610 22800 9640
rect 20253 9608 22800 9610
rect 20253 9552 20258 9608
rect 20314 9552 22800 9608
rect 20253 9550 22800 9552
rect 20253 9547 20319 9550
rect 22320 9520 22800 9550
rect 20529 9202 20595 9205
rect 22320 9202 22800 9232
rect 20529 9200 22800 9202
rect 20529 9144 20534 9200
rect 20590 9144 22800 9200
rect 20529 9142 22800 9144
rect 20529 9139 20595 9142
rect 7808 9136 8128 9137
rect 7808 9072 7816 9136
rect 7880 9072 7896 9136
rect 7960 9072 7976 9136
rect 8040 9072 8056 9136
rect 8120 9072 8128 9136
rect 7808 9071 8128 9072
rect 14672 9136 14992 9137
rect 14672 9072 14680 9136
rect 14744 9072 14760 9136
rect 14824 9072 14840 9136
rect 14904 9072 14920 9136
rect 14984 9072 14992 9136
rect 22320 9112 22800 9142
rect 14672 9071 14992 9072
rect 20253 8658 20319 8661
rect 22320 8658 22800 8688
rect 20253 8656 22800 8658
rect 20253 8600 20258 8656
rect 20314 8600 22800 8656
rect 20253 8598 22800 8600
rect 20253 8595 20319 8598
rect 4376 8592 4696 8593
rect 4376 8528 4384 8592
rect 4448 8528 4464 8592
rect 4528 8528 4544 8592
rect 4608 8528 4624 8592
rect 4688 8528 4696 8592
rect 4376 8527 4696 8528
rect 11240 8592 11560 8593
rect 11240 8528 11248 8592
rect 11312 8528 11328 8592
rect 11392 8528 11408 8592
rect 11472 8528 11488 8592
rect 11552 8528 11560 8592
rect 11240 8527 11560 8528
rect 18104 8592 18424 8593
rect 18104 8528 18112 8592
rect 18176 8528 18192 8592
rect 18256 8528 18272 8592
rect 18336 8528 18352 8592
rect 18416 8528 18424 8592
rect 22320 8568 22800 8598
rect 18104 8527 18424 8528
rect 20529 8250 20595 8253
rect 22320 8250 22800 8280
rect 20529 8248 22800 8250
rect 20529 8192 20534 8248
rect 20590 8192 22800 8248
rect 20529 8190 22800 8192
rect 20529 8187 20595 8190
rect 22320 8160 22800 8190
rect 7808 8048 8128 8049
rect 7808 7984 7816 8048
rect 7880 7984 7896 8048
rect 7960 7984 7976 8048
rect 8040 7984 8056 8048
rect 8120 7984 8128 8048
rect 7808 7983 8128 7984
rect 14672 8048 14992 8049
rect 14672 7984 14680 8048
rect 14744 7984 14760 8048
rect 14824 7984 14840 8048
rect 14904 7984 14920 8048
rect 14984 7984 14992 8048
rect 14672 7983 14992 7984
rect 20253 7842 20319 7845
rect 22320 7842 22800 7872
rect 20253 7840 22800 7842
rect 20253 7784 20258 7840
rect 20314 7784 22800 7840
rect 20253 7782 22800 7784
rect 20253 7779 20319 7782
rect 22320 7752 22800 7782
rect 4376 7504 4696 7505
rect 4376 7440 4384 7504
rect 4448 7440 4464 7504
rect 4528 7440 4544 7504
rect 4608 7440 4624 7504
rect 4688 7440 4696 7504
rect 4376 7439 4696 7440
rect 11240 7504 11560 7505
rect 11240 7440 11248 7504
rect 11312 7440 11328 7504
rect 11392 7440 11408 7504
rect 11472 7440 11488 7504
rect 11552 7440 11560 7504
rect 11240 7439 11560 7440
rect 18104 7504 18424 7505
rect 18104 7440 18112 7504
rect 18176 7440 18192 7504
rect 18256 7440 18272 7504
rect 18336 7440 18352 7504
rect 18416 7440 18424 7504
rect 18104 7439 18424 7440
rect 19977 7298 20043 7301
rect 22320 7298 22800 7328
rect 19977 7296 22800 7298
rect 19977 7240 19982 7296
rect 20038 7240 22800 7296
rect 19977 7238 22800 7240
rect 19977 7235 20043 7238
rect 22320 7208 22800 7238
rect 7808 6960 8128 6961
rect 7808 6896 7816 6960
rect 7880 6896 7896 6960
rect 7960 6896 7976 6960
rect 8040 6896 8056 6960
rect 8120 6896 8128 6960
rect 7808 6895 8128 6896
rect 14672 6960 14992 6961
rect 14672 6896 14680 6960
rect 14744 6896 14760 6960
rect 14824 6896 14840 6960
rect 14904 6896 14920 6960
rect 14984 6896 14992 6960
rect 14672 6895 14992 6896
rect 20529 6890 20595 6893
rect 22320 6890 22800 6920
rect 20529 6888 22800 6890
rect 20529 6832 20534 6888
rect 20590 6832 22800 6888
rect 20529 6830 22800 6832
rect 20529 6827 20595 6830
rect 22320 6800 22800 6830
rect 18597 6482 18663 6485
rect 22320 6482 22800 6512
rect 18597 6480 22800 6482
rect 18597 6424 18602 6480
rect 18658 6424 22800 6480
rect 18597 6422 22800 6424
rect 18597 6419 18663 6422
rect 4376 6416 4696 6417
rect 4376 6352 4384 6416
rect 4448 6352 4464 6416
rect 4528 6352 4544 6416
rect 4608 6352 4624 6416
rect 4688 6352 4696 6416
rect 4376 6351 4696 6352
rect 11240 6416 11560 6417
rect 11240 6352 11248 6416
rect 11312 6352 11328 6416
rect 11392 6352 11408 6416
rect 11472 6352 11488 6416
rect 11552 6352 11560 6416
rect 11240 6351 11560 6352
rect 18104 6416 18424 6417
rect 18104 6352 18112 6416
rect 18176 6352 18192 6416
rect 18256 6352 18272 6416
rect 18336 6352 18352 6416
rect 18416 6352 18424 6416
rect 22320 6392 22800 6422
rect 18104 6351 18424 6352
rect 17953 5938 18019 5941
rect 22320 5938 22800 5968
rect 17953 5936 22800 5938
rect 17953 5880 17958 5936
rect 18014 5880 22800 5936
rect 17953 5878 22800 5880
rect 17953 5875 18019 5878
rect 7808 5872 8128 5873
rect 7808 5808 7816 5872
rect 7880 5808 7896 5872
rect 7960 5808 7976 5872
rect 8040 5808 8056 5872
rect 8120 5808 8128 5872
rect 7808 5807 8128 5808
rect 14672 5872 14992 5873
rect 14672 5808 14680 5872
rect 14744 5808 14760 5872
rect 14824 5808 14840 5872
rect 14904 5808 14920 5872
rect 14984 5808 14992 5872
rect 22320 5848 22800 5878
rect 14672 5807 14992 5808
rect 0 5666 480 5696
rect 3601 5666 3667 5669
rect 0 5664 3667 5666
rect 0 5608 3606 5664
rect 3662 5608 3667 5664
rect 0 5606 3667 5608
rect 0 5576 480 5606
rect 3601 5603 3667 5606
rect 18505 5530 18571 5533
rect 22320 5530 22800 5560
rect 18505 5528 22800 5530
rect 18505 5472 18510 5528
rect 18566 5472 22800 5528
rect 18505 5470 22800 5472
rect 18505 5467 18571 5470
rect 22320 5440 22800 5470
rect 4376 5328 4696 5329
rect 4376 5264 4384 5328
rect 4448 5264 4464 5328
rect 4528 5264 4544 5328
rect 4608 5264 4624 5328
rect 4688 5264 4696 5328
rect 4376 5263 4696 5264
rect 11240 5328 11560 5329
rect 11240 5264 11248 5328
rect 11312 5264 11328 5328
rect 11392 5264 11408 5328
rect 11472 5264 11488 5328
rect 11552 5264 11560 5328
rect 11240 5263 11560 5264
rect 18104 5328 18424 5329
rect 18104 5264 18112 5328
rect 18176 5264 18192 5328
rect 18256 5264 18272 5328
rect 18336 5264 18352 5328
rect 18416 5264 18424 5328
rect 18104 5263 18424 5264
rect 17953 4986 18019 4989
rect 22320 4986 22800 5016
rect 17953 4984 22800 4986
rect 17953 4928 17958 4984
rect 18014 4928 22800 4984
rect 17953 4926 22800 4928
rect 17953 4923 18019 4926
rect 22320 4896 22800 4926
rect 7808 4784 8128 4785
rect 7808 4720 7816 4784
rect 7880 4720 7896 4784
rect 7960 4720 7976 4784
rect 8040 4720 8056 4784
rect 8120 4720 8128 4784
rect 7808 4719 8128 4720
rect 14672 4784 14992 4785
rect 14672 4720 14680 4784
rect 14744 4720 14760 4784
rect 14824 4720 14840 4784
rect 14904 4720 14920 4784
rect 14984 4720 14992 4784
rect 14672 4719 14992 4720
rect 18045 4578 18111 4581
rect 22320 4578 22800 4608
rect 18045 4576 22800 4578
rect 18045 4520 18050 4576
rect 18106 4520 22800 4576
rect 18045 4518 22800 4520
rect 18045 4515 18111 4518
rect 22320 4488 22800 4518
rect 4376 4240 4696 4241
rect 4376 4176 4384 4240
rect 4448 4176 4464 4240
rect 4528 4176 4544 4240
rect 4608 4176 4624 4240
rect 4688 4176 4696 4240
rect 4376 4175 4696 4176
rect 11240 4240 11560 4241
rect 11240 4176 11248 4240
rect 11312 4176 11328 4240
rect 11392 4176 11408 4240
rect 11472 4176 11488 4240
rect 11552 4176 11560 4240
rect 11240 4175 11560 4176
rect 18104 4240 18424 4241
rect 18104 4176 18112 4240
rect 18176 4176 18192 4240
rect 18256 4176 18272 4240
rect 18336 4176 18352 4240
rect 18416 4176 18424 4240
rect 18104 4175 18424 4176
rect 20529 4170 20595 4173
rect 22320 4170 22800 4200
rect 20529 4168 22800 4170
rect 20529 4112 20534 4168
rect 20590 4112 22800 4168
rect 20529 4110 22800 4112
rect 20529 4107 20595 4110
rect 22320 4080 22800 4110
rect 7808 3696 8128 3697
rect 7808 3632 7816 3696
rect 7880 3632 7896 3696
rect 7960 3632 7976 3696
rect 8040 3632 8056 3696
rect 8120 3632 8128 3696
rect 7808 3631 8128 3632
rect 14672 3696 14992 3697
rect 14672 3632 14680 3696
rect 14744 3632 14760 3696
rect 14824 3632 14840 3696
rect 14904 3632 14920 3696
rect 14984 3632 14992 3696
rect 14672 3631 14992 3632
rect 17769 3626 17835 3629
rect 22320 3626 22800 3656
rect 17769 3624 22800 3626
rect 17769 3568 17774 3624
rect 17830 3568 22800 3624
rect 17769 3566 22800 3568
rect 17769 3563 17835 3566
rect 22320 3536 22800 3566
rect 18505 3218 18571 3221
rect 22320 3218 22800 3248
rect 18505 3216 22800 3218
rect 18505 3160 18510 3216
rect 18566 3160 22800 3216
rect 18505 3158 22800 3160
rect 18505 3155 18571 3158
rect 4376 3152 4696 3153
rect 4376 3088 4384 3152
rect 4448 3088 4464 3152
rect 4528 3088 4544 3152
rect 4608 3088 4624 3152
rect 4688 3088 4696 3152
rect 4376 3087 4696 3088
rect 11240 3152 11560 3153
rect 11240 3088 11248 3152
rect 11312 3088 11328 3152
rect 11392 3088 11408 3152
rect 11472 3088 11488 3152
rect 11552 3088 11560 3152
rect 11240 3087 11560 3088
rect 18104 3152 18424 3153
rect 18104 3088 18112 3152
rect 18176 3088 18192 3152
rect 18256 3088 18272 3152
rect 18336 3088 18352 3152
rect 18416 3088 18424 3152
rect 22320 3128 22800 3158
rect 18104 3087 18424 3088
rect 17861 2810 17927 2813
rect 22320 2810 22800 2840
rect 17861 2808 22800 2810
rect 17861 2752 17866 2808
rect 17922 2752 22800 2808
rect 17861 2750 22800 2752
rect 17861 2747 17927 2750
rect 22320 2720 22800 2750
rect 7808 2608 8128 2609
rect 7808 2544 7816 2608
rect 7880 2544 7896 2608
rect 7960 2544 7976 2608
rect 8040 2544 8056 2608
rect 8120 2544 8128 2608
rect 7808 2543 8128 2544
rect 14672 2608 14992 2609
rect 14672 2544 14680 2608
rect 14744 2544 14760 2608
rect 14824 2544 14840 2608
rect 14904 2544 14920 2608
rect 14984 2544 14992 2608
rect 14672 2543 14992 2544
rect 18873 2266 18939 2269
rect 22320 2266 22800 2296
rect 18873 2264 22800 2266
rect 18873 2208 18878 2264
rect 18934 2208 22800 2264
rect 18873 2206 22800 2208
rect 18873 2203 18939 2206
rect 22320 2176 22800 2206
rect 4376 2064 4696 2065
rect 4376 2000 4384 2064
rect 4448 2000 4464 2064
rect 4528 2000 4544 2064
rect 4608 2000 4624 2064
rect 4688 2000 4696 2064
rect 4376 1999 4696 2000
rect 11240 2064 11560 2065
rect 11240 2000 11248 2064
rect 11312 2000 11328 2064
rect 11392 2000 11408 2064
rect 11472 2000 11488 2064
rect 11552 2000 11560 2064
rect 11240 1999 11560 2000
rect 18104 2064 18424 2065
rect 18104 2000 18112 2064
rect 18176 2000 18192 2064
rect 18256 2000 18272 2064
rect 18336 2000 18352 2064
rect 18416 2000 18424 2064
rect 18104 1999 18424 2000
rect 18781 1858 18847 1861
rect 22320 1858 22800 1888
rect 18781 1856 22800 1858
rect 18781 1800 18786 1856
rect 18842 1800 22800 1856
rect 18781 1798 22800 1800
rect 18781 1795 18847 1798
rect 22320 1768 22800 1798
rect 18689 1450 18755 1453
rect 22320 1450 22800 1480
rect 18689 1448 22800 1450
rect 18689 1392 18694 1448
rect 18750 1392 22800 1448
rect 18689 1390 22800 1392
rect 18689 1387 18755 1390
rect 22320 1360 22800 1390
rect 19057 906 19123 909
rect 22320 906 22800 936
rect 19057 904 22800 906
rect 19057 848 19062 904
rect 19118 848 22800 904
rect 19057 846 22800 848
rect 19057 843 19123 846
rect 22320 816 22800 846
rect 17309 498 17375 501
rect 22320 498 22800 528
rect 17309 496 22800 498
rect 17309 440 17314 496
rect 17370 440 22800 496
rect 17309 438 22800 440
rect 17309 435 17375 438
rect 22320 408 22800 438
rect 18137 90 18203 93
rect 22320 90 22800 120
rect 18137 88 22800 90
rect 18137 32 18142 88
rect 18198 32 22800 88
rect 18137 30 22800 32
rect 18137 27 18203 30
rect 22320 0 22800 30
<< via3 >>
rect 7816 20012 7880 20016
rect 7816 19956 7820 20012
rect 7820 19956 7876 20012
rect 7876 19956 7880 20012
rect 7816 19952 7880 19956
rect 7896 20012 7960 20016
rect 7896 19956 7900 20012
rect 7900 19956 7956 20012
rect 7956 19956 7960 20012
rect 7896 19952 7960 19956
rect 7976 20012 8040 20016
rect 7976 19956 7980 20012
rect 7980 19956 8036 20012
rect 8036 19956 8040 20012
rect 7976 19952 8040 19956
rect 8056 20012 8120 20016
rect 8056 19956 8060 20012
rect 8060 19956 8116 20012
rect 8116 19956 8120 20012
rect 8056 19952 8120 19956
rect 14680 20012 14744 20016
rect 14680 19956 14684 20012
rect 14684 19956 14740 20012
rect 14740 19956 14744 20012
rect 14680 19952 14744 19956
rect 14760 20012 14824 20016
rect 14760 19956 14764 20012
rect 14764 19956 14820 20012
rect 14820 19956 14824 20012
rect 14760 19952 14824 19956
rect 14840 20012 14904 20016
rect 14840 19956 14844 20012
rect 14844 19956 14900 20012
rect 14900 19956 14904 20012
rect 14840 19952 14904 19956
rect 14920 20012 14984 20016
rect 14920 19956 14924 20012
rect 14924 19956 14980 20012
rect 14980 19956 14984 20012
rect 14920 19952 14984 19956
rect 4384 19468 4448 19472
rect 4384 19412 4388 19468
rect 4388 19412 4444 19468
rect 4444 19412 4448 19468
rect 4384 19408 4448 19412
rect 4464 19468 4528 19472
rect 4464 19412 4468 19468
rect 4468 19412 4524 19468
rect 4524 19412 4528 19468
rect 4464 19408 4528 19412
rect 4544 19468 4608 19472
rect 4544 19412 4548 19468
rect 4548 19412 4604 19468
rect 4604 19412 4608 19468
rect 4544 19408 4608 19412
rect 4624 19468 4688 19472
rect 4624 19412 4628 19468
rect 4628 19412 4684 19468
rect 4684 19412 4688 19468
rect 4624 19408 4688 19412
rect 11248 19468 11312 19472
rect 11248 19412 11252 19468
rect 11252 19412 11308 19468
rect 11308 19412 11312 19468
rect 11248 19408 11312 19412
rect 11328 19468 11392 19472
rect 11328 19412 11332 19468
rect 11332 19412 11388 19468
rect 11388 19412 11392 19468
rect 11328 19408 11392 19412
rect 11408 19468 11472 19472
rect 11408 19412 11412 19468
rect 11412 19412 11468 19468
rect 11468 19412 11472 19468
rect 11408 19408 11472 19412
rect 11488 19468 11552 19472
rect 11488 19412 11492 19468
rect 11492 19412 11548 19468
rect 11548 19412 11552 19468
rect 11488 19408 11552 19412
rect 18112 19468 18176 19472
rect 18112 19412 18116 19468
rect 18116 19412 18172 19468
rect 18172 19412 18176 19468
rect 18112 19408 18176 19412
rect 18192 19468 18256 19472
rect 18192 19412 18196 19468
rect 18196 19412 18252 19468
rect 18252 19412 18256 19468
rect 18192 19408 18256 19412
rect 18272 19468 18336 19472
rect 18272 19412 18276 19468
rect 18276 19412 18332 19468
rect 18332 19412 18336 19468
rect 18272 19408 18336 19412
rect 18352 19468 18416 19472
rect 18352 19412 18356 19468
rect 18356 19412 18412 19468
rect 18412 19412 18416 19468
rect 18352 19408 18416 19412
rect 7816 18924 7880 18928
rect 7816 18868 7820 18924
rect 7820 18868 7876 18924
rect 7876 18868 7880 18924
rect 7816 18864 7880 18868
rect 7896 18924 7960 18928
rect 7896 18868 7900 18924
rect 7900 18868 7956 18924
rect 7956 18868 7960 18924
rect 7896 18864 7960 18868
rect 7976 18924 8040 18928
rect 7976 18868 7980 18924
rect 7980 18868 8036 18924
rect 8036 18868 8040 18924
rect 7976 18864 8040 18868
rect 8056 18924 8120 18928
rect 8056 18868 8060 18924
rect 8060 18868 8116 18924
rect 8116 18868 8120 18924
rect 8056 18864 8120 18868
rect 14680 18924 14744 18928
rect 14680 18868 14684 18924
rect 14684 18868 14740 18924
rect 14740 18868 14744 18924
rect 14680 18864 14744 18868
rect 14760 18924 14824 18928
rect 14760 18868 14764 18924
rect 14764 18868 14820 18924
rect 14820 18868 14824 18924
rect 14760 18864 14824 18868
rect 14840 18924 14904 18928
rect 14840 18868 14844 18924
rect 14844 18868 14900 18924
rect 14900 18868 14904 18924
rect 14840 18864 14904 18868
rect 14920 18924 14984 18928
rect 14920 18868 14924 18924
rect 14924 18868 14980 18924
rect 14980 18868 14984 18924
rect 14920 18864 14984 18868
rect 4384 18380 4448 18384
rect 4384 18324 4388 18380
rect 4388 18324 4444 18380
rect 4444 18324 4448 18380
rect 4384 18320 4448 18324
rect 4464 18380 4528 18384
rect 4464 18324 4468 18380
rect 4468 18324 4524 18380
rect 4524 18324 4528 18380
rect 4464 18320 4528 18324
rect 4544 18380 4608 18384
rect 4544 18324 4548 18380
rect 4548 18324 4604 18380
rect 4604 18324 4608 18380
rect 4544 18320 4608 18324
rect 4624 18380 4688 18384
rect 4624 18324 4628 18380
rect 4628 18324 4684 18380
rect 4684 18324 4688 18380
rect 4624 18320 4688 18324
rect 11248 18380 11312 18384
rect 11248 18324 11252 18380
rect 11252 18324 11308 18380
rect 11308 18324 11312 18380
rect 11248 18320 11312 18324
rect 11328 18380 11392 18384
rect 11328 18324 11332 18380
rect 11332 18324 11388 18380
rect 11388 18324 11392 18380
rect 11328 18320 11392 18324
rect 11408 18380 11472 18384
rect 11408 18324 11412 18380
rect 11412 18324 11468 18380
rect 11468 18324 11472 18380
rect 11408 18320 11472 18324
rect 11488 18380 11552 18384
rect 11488 18324 11492 18380
rect 11492 18324 11548 18380
rect 11548 18324 11552 18380
rect 11488 18320 11552 18324
rect 18112 18380 18176 18384
rect 18112 18324 18116 18380
rect 18116 18324 18172 18380
rect 18172 18324 18176 18380
rect 18112 18320 18176 18324
rect 18192 18380 18256 18384
rect 18192 18324 18196 18380
rect 18196 18324 18252 18380
rect 18252 18324 18256 18380
rect 18192 18320 18256 18324
rect 18272 18380 18336 18384
rect 18272 18324 18276 18380
rect 18276 18324 18332 18380
rect 18332 18324 18336 18380
rect 18272 18320 18336 18324
rect 18352 18380 18416 18384
rect 18352 18324 18356 18380
rect 18356 18324 18412 18380
rect 18412 18324 18416 18380
rect 18352 18320 18416 18324
rect 7816 17836 7880 17840
rect 7816 17780 7820 17836
rect 7820 17780 7876 17836
rect 7876 17780 7880 17836
rect 7816 17776 7880 17780
rect 7896 17836 7960 17840
rect 7896 17780 7900 17836
rect 7900 17780 7956 17836
rect 7956 17780 7960 17836
rect 7896 17776 7960 17780
rect 7976 17836 8040 17840
rect 7976 17780 7980 17836
rect 7980 17780 8036 17836
rect 8036 17780 8040 17836
rect 7976 17776 8040 17780
rect 8056 17836 8120 17840
rect 8056 17780 8060 17836
rect 8060 17780 8116 17836
rect 8116 17780 8120 17836
rect 8056 17776 8120 17780
rect 14680 17836 14744 17840
rect 14680 17780 14684 17836
rect 14684 17780 14740 17836
rect 14740 17780 14744 17836
rect 14680 17776 14744 17780
rect 14760 17836 14824 17840
rect 14760 17780 14764 17836
rect 14764 17780 14820 17836
rect 14820 17780 14824 17836
rect 14760 17776 14824 17780
rect 14840 17836 14904 17840
rect 14840 17780 14844 17836
rect 14844 17780 14900 17836
rect 14900 17780 14904 17836
rect 14840 17776 14904 17780
rect 14920 17836 14984 17840
rect 14920 17780 14924 17836
rect 14924 17780 14980 17836
rect 14980 17780 14984 17836
rect 14920 17776 14984 17780
rect 4384 17292 4448 17296
rect 4384 17236 4388 17292
rect 4388 17236 4444 17292
rect 4444 17236 4448 17292
rect 4384 17232 4448 17236
rect 4464 17292 4528 17296
rect 4464 17236 4468 17292
rect 4468 17236 4524 17292
rect 4524 17236 4528 17292
rect 4464 17232 4528 17236
rect 4544 17292 4608 17296
rect 4544 17236 4548 17292
rect 4548 17236 4604 17292
rect 4604 17236 4608 17292
rect 4544 17232 4608 17236
rect 4624 17292 4688 17296
rect 4624 17236 4628 17292
rect 4628 17236 4684 17292
rect 4684 17236 4688 17292
rect 4624 17232 4688 17236
rect 11248 17292 11312 17296
rect 11248 17236 11252 17292
rect 11252 17236 11308 17292
rect 11308 17236 11312 17292
rect 11248 17232 11312 17236
rect 11328 17292 11392 17296
rect 11328 17236 11332 17292
rect 11332 17236 11388 17292
rect 11388 17236 11392 17292
rect 11328 17232 11392 17236
rect 11408 17292 11472 17296
rect 11408 17236 11412 17292
rect 11412 17236 11468 17292
rect 11468 17236 11472 17292
rect 11408 17232 11472 17236
rect 11488 17292 11552 17296
rect 11488 17236 11492 17292
rect 11492 17236 11548 17292
rect 11548 17236 11552 17292
rect 11488 17232 11552 17236
rect 18112 17292 18176 17296
rect 18112 17236 18116 17292
rect 18116 17236 18172 17292
rect 18172 17236 18176 17292
rect 18112 17232 18176 17236
rect 18192 17292 18256 17296
rect 18192 17236 18196 17292
rect 18196 17236 18252 17292
rect 18252 17236 18256 17292
rect 18192 17232 18256 17236
rect 18272 17292 18336 17296
rect 18272 17236 18276 17292
rect 18276 17236 18332 17292
rect 18332 17236 18336 17292
rect 18272 17232 18336 17236
rect 18352 17292 18416 17296
rect 18352 17236 18356 17292
rect 18356 17236 18412 17292
rect 18412 17236 18416 17292
rect 18352 17232 18416 17236
rect 7816 16748 7880 16752
rect 7816 16692 7820 16748
rect 7820 16692 7876 16748
rect 7876 16692 7880 16748
rect 7816 16688 7880 16692
rect 7896 16748 7960 16752
rect 7896 16692 7900 16748
rect 7900 16692 7956 16748
rect 7956 16692 7960 16748
rect 7896 16688 7960 16692
rect 7976 16748 8040 16752
rect 7976 16692 7980 16748
rect 7980 16692 8036 16748
rect 8036 16692 8040 16748
rect 7976 16688 8040 16692
rect 8056 16748 8120 16752
rect 8056 16692 8060 16748
rect 8060 16692 8116 16748
rect 8116 16692 8120 16748
rect 8056 16688 8120 16692
rect 14680 16748 14744 16752
rect 14680 16692 14684 16748
rect 14684 16692 14740 16748
rect 14740 16692 14744 16748
rect 14680 16688 14744 16692
rect 14760 16748 14824 16752
rect 14760 16692 14764 16748
rect 14764 16692 14820 16748
rect 14820 16692 14824 16748
rect 14760 16688 14824 16692
rect 14840 16748 14904 16752
rect 14840 16692 14844 16748
rect 14844 16692 14900 16748
rect 14900 16692 14904 16748
rect 14840 16688 14904 16692
rect 14920 16748 14984 16752
rect 14920 16692 14924 16748
rect 14924 16692 14980 16748
rect 14980 16692 14984 16748
rect 14920 16688 14984 16692
rect 4384 16204 4448 16208
rect 4384 16148 4388 16204
rect 4388 16148 4444 16204
rect 4444 16148 4448 16204
rect 4384 16144 4448 16148
rect 4464 16204 4528 16208
rect 4464 16148 4468 16204
rect 4468 16148 4524 16204
rect 4524 16148 4528 16204
rect 4464 16144 4528 16148
rect 4544 16204 4608 16208
rect 4544 16148 4548 16204
rect 4548 16148 4604 16204
rect 4604 16148 4608 16204
rect 4544 16144 4608 16148
rect 4624 16204 4688 16208
rect 4624 16148 4628 16204
rect 4628 16148 4684 16204
rect 4684 16148 4688 16204
rect 4624 16144 4688 16148
rect 11248 16204 11312 16208
rect 11248 16148 11252 16204
rect 11252 16148 11308 16204
rect 11308 16148 11312 16204
rect 11248 16144 11312 16148
rect 11328 16204 11392 16208
rect 11328 16148 11332 16204
rect 11332 16148 11388 16204
rect 11388 16148 11392 16204
rect 11328 16144 11392 16148
rect 11408 16204 11472 16208
rect 11408 16148 11412 16204
rect 11412 16148 11468 16204
rect 11468 16148 11472 16204
rect 11408 16144 11472 16148
rect 11488 16204 11552 16208
rect 11488 16148 11492 16204
rect 11492 16148 11548 16204
rect 11548 16148 11552 16204
rect 11488 16144 11552 16148
rect 18112 16204 18176 16208
rect 18112 16148 18116 16204
rect 18116 16148 18172 16204
rect 18172 16148 18176 16204
rect 18112 16144 18176 16148
rect 18192 16204 18256 16208
rect 18192 16148 18196 16204
rect 18196 16148 18252 16204
rect 18252 16148 18256 16204
rect 18192 16144 18256 16148
rect 18272 16204 18336 16208
rect 18272 16148 18276 16204
rect 18276 16148 18332 16204
rect 18332 16148 18336 16204
rect 18272 16144 18336 16148
rect 18352 16204 18416 16208
rect 18352 16148 18356 16204
rect 18356 16148 18412 16204
rect 18412 16148 18416 16204
rect 18352 16144 18416 16148
rect 7816 15660 7880 15664
rect 7816 15604 7820 15660
rect 7820 15604 7876 15660
rect 7876 15604 7880 15660
rect 7816 15600 7880 15604
rect 7896 15660 7960 15664
rect 7896 15604 7900 15660
rect 7900 15604 7956 15660
rect 7956 15604 7960 15660
rect 7896 15600 7960 15604
rect 7976 15660 8040 15664
rect 7976 15604 7980 15660
rect 7980 15604 8036 15660
rect 8036 15604 8040 15660
rect 7976 15600 8040 15604
rect 8056 15660 8120 15664
rect 8056 15604 8060 15660
rect 8060 15604 8116 15660
rect 8116 15604 8120 15660
rect 8056 15600 8120 15604
rect 14680 15660 14744 15664
rect 14680 15604 14684 15660
rect 14684 15604 14740 15660
rect 14740 15604 14744 15660
rect 14680 15600 14744 15604
rect 14760 15660 14824 15664
rect 14760 15604 14764 15660
rect 14764 15604 14820 15660
rect 14820 15604 14824 15660
rect 14760 15600 14824 15604
rect 14840 15660 14904 15664
rect 14840 15604 14844 15660
rect 14844 15604 14900 15660
rect 14900 15604 14904 15660
rect 14840 15600 14904 15604
rect 14920 15660 14984 15664
rect 14920 15604 14924 15660
rect 14924 15604 14980 15660
rect 14980 15604 14984 15660
rect 14920 15600 14984 15604
rect 4384 15116 4448 15120
rect 4384 15060 4388 15116
rect 4388 15060 4444 15116
rect 4444 15060 4448 15116
rect 4384 15056 4448 15060
rect 4464 15116 4528 15120
rect 4464 15060 4468 15116
rect 4468 15060 4524 15116
rect 4524 15060 4528 15116
rect 4464 15056 4528 15060
rect 4544 15116 4608 15120
rect 4544 15060 4548 15116
rect 4548 15060 4604 15116
rect 4604 15060 4608 15116
rect 4544 15056 4608 15060
rect 4624 15116 4688 15120
rect 4624 15060 4628 15116
rect 4628 15060 4684 15116
rect 4684 15060 4688 15116
rect 4624 15056 4688 15060
rect 11248 15116 11312 15120
rect 11248 15060 11252 15116
rect 11252 15060 11308 15116
rect 11308 15060 11312 15116
rect 11248 15056 11312 15060
rect 11328 15116 11392 15120
rect 11328 15060 11332 15116
rect 11332 15060 11388 15116
rect 11388 15060 11392 15116
rect 11328 15056 11392 15060
rect 11408 15116 11472 15120
rect 11408 15060 11412 15116
rect 11412 15060 11468 15116
rect 11468 15060 11472 15116
rect 11408 15056 11472 15060
rect 11488 15116 11552 15120
rect 11488 15060 11492 15116
rect 11492 15060 11548 15116
rect 11548 15060 11552 15116
rect 11488 15056 11552 15060
rect 18112 15116 18176 15120
rect 18112 15060 18116 15116
rect 18116 15060 18172 15116
rect 18172 15060 18176 15116
rect 18112 15056 18176 15060
rect 18192 15116 18256 15120
rect 18192 15060 18196 15116
rect 18196 15060 18252 15116
rect 18252 15060 18256 15116
rect 18192 15056 18256 15060
rect 18272 15116 18336 15120
rect 18272 15060 18276 15116
rect 18276 15060 18332 15116
rect 18332 15060 18336 15116
rect 18272 15056 18336 15060
rect 18352 15116 18416 15120
rect 18352 15060 18356 15116
rect 18356 15060 18412 15116
rect 18412 15060 18416 15116
rect 18352 15056 18416 15060
rect 7816 14572 7880 14576
rect 7816 14516 7820 14572
rect 7820 14516 7876 14572
rect 7876 14516 7880 14572
rect 7816 14512 7880 14516
rect 7896 14572 7960 14576
rect 7896 14516 7900 14572
rect 7900 14516 7956 14572
rect 7956 14516 7960 14572
rect 7896 14512 7960 14516
rect 7976 14572 8040 14576
rect 7976 14516 7980 14572
rect 7980 14516 8036 14572
rect 8036 14516 8040 14572
rect 7976 14512 8040 14516
rect 8056 14572 8120 14576
rect 8056 14516 8060 14572
rect 8060 14516 8116 14572
rect 8116 14516 8120 14572
rect 8056 14512 8120 14516
rect 14680 14572 14744 14576
rect 14680 14516 14684 14572
rect 14684 14516 14740 14572
rect 14740 14516 14744 14572
rect 14680 14512 14744 14516
rect 14760 14572 14824 14576
rect 14760 14516 14764 14572
rect 14764 14516 14820 14572
rect 14820 14516 14824 14572
rect 14760 14512 14824 14516
rect 14840 14572 14904 14576
rect 14840 14516 14844 14572
rect 14844 14516 14900 14572
rect 14900 14516 14904 14572
rect 14840 14512 14904 14516
rect 14920 14572 14984 14576
rect 14920 14516 14924 14572
rect 14924 14516 14980 14572
rect 14980 14516 14984 14572
rect 14920 14512 14984 14516
rect 4384 14028 4448 14032
rect 4384 13972 4388 14028
rect 4388 13972 4444 14028
rect 4444 13972 4448 14028
rect 4384 13968 4448 13972
rect 4464 14028 4528 14032
rect 4464 13972 4468 14028
rect 4468 13972 4524 14028
rect 4524 13972 4528 14028
rect 4464 13968 4528 13972
rect 4544 14028 4608 14032
rect 4544 13972 4548 14028
rect 4548 13972 4604 14028
rect 4604 13972 4608 14028
rect 4544 13968 4608 13972
rect 4624 14028 4688 14032
rect 4624 13972 4628 14028
rect 4628 13972 4684 14028
rect 4684 13972 4688 14028
rect 4624 13968 4688 13972
rect 11248 14028 11312 14032
rect 11248 13972 11252 14028
rect 11252 13972 11308 14028
rect 11308 13972 11312 14028
rect 11248 13968 11312 13972
rect 11328 14028 11392 14032
rect 11328 13972 11332 14028
rect 11332 13972 11388 14028
rect 11388 13972 11392 14028
rect 11328 13968 11392 13972
rect 11408 14028 11472 14032
rect 11408 13972 11412 14028
rect 11412 13972 11468 14028
rect 11468 13972 11472 14028
rect 11408 13968 11472 13972
rect 11488 14028 11552 14032
rect 11488 13972 11492 14028
rect 11492 13972 11548 14028
rect 11548 13972 11552 14028
rect 11488 13968 11552 13972
rect 18112 14028 18176 14032
rect 18112 13972 18116 14028
rect 18116 13972 18172 14028
rect 18172 13972 18176 14028
rect 18112 13968 18176 13972
rect 18192 14028 18256 14032
rect 18192 13972 18196 14028
rect 18196 13972 18252 14028
rect 18252 13972 18256 14028
rect 18192 13968 18256 13972
rect 18272 14028 18336 14032
rect 18272 13972 18276 14028
rect 18276 13972 18332 14028
rect 18332 13972 18336 14028
rect 18272 13968 18336 13972
rect 18352 14028 18416 14032
rect 18352 13972 18356 14028
rect 18356 13972 18412 14028
rect 18412 13972 18416 14028
rect 18352 13968 18416 13972
rect 7816 13484 7880 13488
rect 7816 13428 7820 13484
rect 7820 13428 7876 13484
rect 7876 13428 7880 13484
rect 7816 13424 7880 13428
rect 7896 13484 7960 13488
rect 7896 13428 7900 13484
rect 7900 13428 7956 13484
rect 7956 13428 7960 13484
rect 7896 13424 7960 13428
rect 7976 13484 8040 13488
rect 7976 13428 7980 13484
rect 7980 13428 8036 13484
rect 8036 13428 8040 13484
rect 7976 13424 8040 13428
rect 8056 13484 8120 13488
rect 8056 13428 8060 13484
rect 8060 13428 8116 13484
rect 8116 13428 8120 13484
rect 8056 13424 8120 13428
rect 14680 13484 14744 13488
rect 14680 13428 14684 13484
rect 14684 13428 14740 13484
rect 14740 13428 14744 13484
rect 14680 13424 14744 13428
rect 14760 13484 14824 13488
rect 14760 13428 14764 13484
rect 14764 13428 14820 13484
rect 14820 13428 14824 13484
rect 14760 13424 14824 13428
rect 14840 13484 14904 13488
rect 14840 13428 14844 13484
rect 14844 13428 14900 13484
rect 14900 13428 14904 13484
rect 14840 13424 14904 13428
rect 14920 13484 14984 13488
rect 14920 13428 14924 13484
rect 14924 13428 14980 13484
rect 14980 13428 14984 13484
rect 14920 13424 14984 13428
rect 4384 12940 4448 12944
rect 4384 12884 4388 12940
rect 4388 12884 4444 12940
rect 4444 12884 4448 12940
rect 4384 12880 4448 12884
rect 4464 12940 4528 12944
rect 4464 12884 4468 12940
rect 4468 12884 4524 12940
rect 4524 12884 4528 12940
rect 4464 12880 4528 12884
rect 4544 12940 4608 12944
rect 4544 12884 4548 12940
rect 4548 12884 4604 12940
rect 4604 12884 4608 12940
rect 4544 12880 4608 12884
rect 4624 12940 4688 12944
rect 4624 12884 4628 12940
rect 4628 12884 4684 12940
rect 4684 12884 4688 12940
rect 4624 12880 4688 12884
rect 11248 12940 11312 12944
rect 11248 12884 11252 12940
rect 11252 12884 11308 12940
rect 11308 12884 11312 12940
rect 11248 12880 11312 12884
rect 11328 12940 11392 12944
rect 11328 12884 11332 12940
rect 11332 12884 11388 12940
rect 11388 12884 11392 12940
rect 11328 12880 11392 12884
rect 11408 12940 11472 12944
rect 11408 12884 11412 12940
rect 11412 12884 11468 12940
rect 11468 12884 11472 12940
rect 11408 12880 11472 12884
rect 11488 12940 11552 12944
rect 11488 12884 11492 12940
rect 11492 12884 11548 12940
rect 11548 12884 11552 12940
rect 11488 12880 11552 12884
rect 18112 12940 18176 12944
rect 18112 12884 18116 12940
rect 18116 12884 18172 12940
rect 18172 12884 18176 12940
rect 18112 12880 18176 12884
rect 18192 12940 18256 12944
rect 18192 12884 18196 12940
rect 18196 12884 18252 12940
rect 18252 12884 18256 12940
rect 18192 12880 18256 12884
rect 18272 12940 18336 12944
rect 18272 12884 18276 12940
rect 18276 12884 18332 12940
rect 18332 12884 18336 12940
rect 18272 12880 18336 12884
rect 18352 12940 18416 12944
rect 18352 12884 18356 12940
rect 18356 12884 18412 12940
rect 18412 12884 18416 12940
rect 18352 12880 18416 12884
rect 7816 12396 7880 12400
rect 7816 12340 7820 12396
rect 7820 12340 7876 12396
rect 7876 12340 7880 12396
rect 7816 12336 7880 12340
rect 7896 12396 7960 12400
rect 7896 12340 7900 12396
rect 7900 12340 7956 12396
rect 7956 12340 7960 12396
rect 7896 12336 7960 12340
rect 7976 12396 8040 12400
rect 7976 12340 7980 12396
rect 7980 12340 8036 12396
rect 8036 12340 8040 12396
rect 7976 12336 8040 12340
rect 8056 12396 8120 12400
rect 8056 12340 8060 12396
rect 8060 12340 8116 12396
rect 8116 12340 8120 12396
rect 8056 12336 8120 12340
rect 14680 12396 14744 12400
rect 14680 12340 14684 12396
rect 14684 12340 14740 12396
rect 14740 12340 14744 12396
rect 14680 12336 14744 12340
rect 14760 12396 14824 12400
rect 14760 12340 14764 12396
rect 14764 12340 14820 12396
rect 14820 12340 14824 12396
rect 14760 12336 14824 12340
rect 14840 12396 14904 12400
rect 14840 12340 14844 12396
rect 14844 12340 14900 12396
rect 14900 12340 14904 12396
rect 14840 12336 14904 12340
rect 14920 12396 14984 12400
rect 14920 12340 14924 12396
rect 14924 12340 14980 12396
rect 14980 12340 14984 12396
rect 14920 12336 14984 12340
rect 4384 11852 4448 11856
rect 4384 11796 4388 11852
rect 4388 11796 4444 11852
rect 4444 11796 4448 11852
rect 4384 11792 4448 11796
rect 4464 11852 4528 11856
rect 4464 11796 4468 11852
rect 4468 11796 4524 11852
rect 4524 11796 4528 11852
rect 4464 11792 4528 11796
rect 4544 11852 4608 11856
rect 4544 11796 4548 11852
rect 4548 11796 4604 11852
rect 4604 11796 4608 11852
rect 4544 11792 4608 11796
rect 4624 11852 4688 11856
rect 4624 11796 4628 11852
rect 4628 11796 4684 11852
rect 4684 11796 4688 11852
rect 4624 11792 4688 11796
rect 11248 11852 11312 11856
rect 11248 11796 11252 11852
rect 11252 11796 11308 11852
rect 11308 11796 11312 11852
rect 11248 11792 11312 11796
rect 11328 11852 11392 11856
rect 11328 11796 11332 11852
rect 11332 11796 11388 11852
rect 11388 11796 11392 11852
rect 11328 11792 11392 11796
rect 11408 11852 11472 11856
rect 11408 11796 11412 11852
rect 11412 11796 11468 11852
rect 11468 11796 11472 11852
rect 11408 11792 11472 11796
rect 11488 11852 11552 11856
rect 11488 11796 11492 11852
rect 11492 11796 11548 11852
rect 11548 11796 11552 11852
rect 11488 11792 11552 11796
rect 18112 11852 18176 11856
rect 18112 11796 18116 11852
rect 18116 11796 18172 11852
rect 18172 11796 18176 11852
rect 18112 11792 18176 11796
rect 18192 11852 18256 11856
rect 18192 11796 18196 11852
rect 18196 11796 18252 11852
rect 18252 11796 18256 11852
rect 18192 11792 18256 11796
rect 18272 11852 18336 11856
rect 18272 11796 18276 11852
rect 18276 11796 18332 11852
rect 18332 11796 18336 11852
rect 18272 11792 18336 11796
rect 18352 11852 18416 11856
rect 18352 11796 18356 11852
rect 18356 11796 18412 11852
rect 18412 11796 18416 11852
rect 18352 11792 18416 11796
rect 7816 11308 7880 11312
rect 7816 11252 7820 11308
rect 7820 11252 7876 11308
rect 7876 11252 7880 11308
rect 7816 11248 7880 11252
rect 7896 11308 7960 11312
rect 7896 11252 7900 11308
rect 7900 11252 7956 11308
rect 7956 11252 7960 11308
rect 7896 11248 7960 11252
rect 7976 11308 8040 11312
rect 7976 11252 7980 11308
rect 7980 11252 8036 11308
rect 8036 11252 8040 11308
rect 7976 11248 8040 11252
rect 8056 11308 8120 11312
rect 8056 11252 8060 11308
rect 8060 11252 8116 11308
rect 8116 11252 8120 11308
rect 8056 11248 8120 11252
rect 14680 11308 14744 11312
rect 14680 11252 14684 11308
rect 14684 11252 14740 11308
rect 14740 11252 14744 11308
rect 14680 11248 14744 11252
rect 14760 11308 14824 11312
rect 14760 11252 14764 11308
rect 14764 11252 14820 11308
rect 14820 11252 14824 11308
rect 14760 11248 14824 11252
rect 14840 11308 14904 11312
rect 14840 11252 14844 11308
rect 14844 11252 14900 11308
rect 14900 11252 14904 11308
rect 14840 11248 14904 11252
rect 14920 11308 14984 11312
rect 14920 11252 14924 11308
rect 14924 11252 14980 11308
rect 14980 11252 14984 11308
rect 14920 11248 14984 11252
rect 4384 10764 4448 10768
rect 4384 10708 4388 10764
rect 4388 10708 4444 10764
rect 4444 10708 4448 10764
rect 4384 10704 4448 10708
rect 4464 10764 4528 10768
rect 4464 10708 4468 10764
rect 4468 10708 4524 10764
rect 4524 10708 4528 10764
rect 4464 10704 4528 10708
rect 4544 10764 4608 10768
rect 4544 10708 4548 10764
rect 4548 10708 4604 10764
rect 4604 10708 4608 10764
rect 4544 10704 4608 10708
rect 4624 10764 4688 10768
rect 4624 10708 4628 10764
rect 4628 10708 4684 10764
rect 4684 10708 4688 10764
rect 4624 10704 4688 10708
rect 11248 10764 11312 10768
rect 11248 10708 11252 10764
rect 11252 10708 11308 10764
rect 11308 10708 11312 10764
rect 11248 10704 11312 10708
rect 11328 10764 11392 10768
rect 11328 10708 11332 10764
rect 11332 10708 11388 10764
rect 11388 10708 11392 10764
rect 11328 10704 11392 10708
rect 11408 10764 11472 10768
rect 11408 10708 11412 10764
rect 11412 10708 11468 10764
rect 11468 10708 11472 10764
rect 11408 10704 11472 10708
rect 11488 10764 11552 10768
rect 11488 10708 11492 10764
rect 11492 10708 11548 10764
rect 11548 10708 11552 10764
rect 11488 10704 11552 10708
rect 18112 10764 18176 10768
rect 18112 10708 18116 10764
rect 18116 10708 18172 10764
rect 18172 10708 18176 10764
rect 18112 10704 18176 10708
rect 18192 10764 18256 10768
rect 18192 10708 18196 10764
rect 18196 10708 18252 10764
rect 18252 10708 18256 10764
rect 18192 10704 18256 10708
rect 18272 10764 18336 10768
rect 18272 10708 18276 10764
rect 18276 10708 18332 10764
rect 18332 10708 18336 10764
rect 18272 10704 18336 10708
rect 18352 10764 18416 10768
rect 18352 10708 18356 10764
rect 18356 10708 18412 10764
rect 18412 10708 18416 10764
rect 18352 10704 18416 10708
rect 7816 10220 7880 10224
rect 7816 10164 7820 10220
rect 7820 10164 7876 10220
rect 7876 10164 7880 10220
rect 7816 10160 7880 10164
rect 7896 10220 7960 10224
rect 7896 10164 7900 10220
rect 7900 10164 7956 10220
rect 7956 10164 7960 10220
rect 7896 10160 7960 10164
rect 7976 10220 8040 10224
rect 7976 10164 7980 10220
rect 7980 10164 8036 10220
rect 8036 10164 8040 10220
rect 7976 10160 8040 10164
rect 8056 10220 8120 10224
rect 8056 10164 8060 10220
rect 8060 10164 8116 10220
rect 8116 10164 8120 10220
rect 8056 10160 8120 10164
rect 14680 10220 14744 10224
rect 14680 10164 14684 10220
rect 14684 10164 14740 10220
rect 14740 10164 14744 10220
rect 14680 10160 14744 10164
rect 14760 10220 14824 10224
rect 14760 10164 14764 10220
rect 14764 10164 14820 10220
rect 14820 10164 14824 10220
rect 14760 10160 14824 10164
rect 14840 10220 14904 10224
rect 14840 10164 14844 10220
rect 14844 10164 14900 10220
rect 14900 10164 14904 10220
rect 14840 10160 14904 10164
rect 14920 10220 14984 10224
rect 14920 10164 14924 10220
rect 14924 10164 14980 10220
rect 14980 10164 14984 10220
rect 14920 10160 14984 10164
rect 4384 9676 4448 9680
rect 4384 9620 4388 9676
rect 4388 9620 4444 9676
rect 4444 9620 4448 9676
rect 4384 9616 4448 9620
rect 4464 9676 4528 9680
rect 4464 9620 4468 9676
rect 4468 9620 4524 9676
rect 4524 9620 4528 9676
rect 4464 9616 4528 9620
rect 4544 9676 4608 9680
rect 4544 9620 4548 9676
rect 4548 9620 4604 9676
rect 4604 9620 4608 9676
rect 4544 9616 4608 9620
rect 4624 9676 4688 9680
rect 4624 9620 4628 9676
rect 4628 9620 4684 9676
rect 4684 9620 4688 9676
rect 4624 9616 4688 9620
rect 11248 9676 11312 9680
rect 11248 9620 11252 9676
rect 11252 9620 11308 9676
rect 11308 9620 11312 9676
rect 11248 9616 11312 9620
rect 11328 9676 11392 9680
rect 11328 9620 11332 9676
rect 11332 9620 11388 9676
rect 11388 9620 11392 9676
rect 11328 9616 11392 9620
rect 11408 9676 11472 9680
rect 11408 9620 11412 9676
rect 11412 9620 11468 9676
rect 11468 9620 11472 9676
rect 11408 9616 11472 9620
rect 11488 9676 11552 9680
rect 11488 9620 11492 9676
rect 11492 9620 11548 9676
rect 11548 9620 11552 9676
rect 11488 9616 11552 9620
rect 18112 9676 18176 9680
rect 18112 9620 18116 9676
rect 18116 9620 18172 9676
rect 18172 9620 18176 9676
rect 18112 9616 18176 9620
rect 18192 9676 18256 9680
rect 18192 9620 18196 9676
rect 18196 9620 18252 9676
rect 18252 9620 18256 9676
rect 18192 9616 18256 9620
rect 18272 9676 18336 9680
rect 18272 9620 18276 9676
rect 18276 9620 18332 9676
rect 18332 9620 18336 9676
rect 18272 9616 18336 9620
rect 18352 9676 18416 9680
rect 18352 9620 18356 9676
rect 18356 9620 18412 9676
rect 18412 9620 18416 9676
rect 18352 9616 18416 9620
rect 7816 9132 7880 9136
rect 7816 9076 7820 9132
rect 7820 9076 7876 9132
rect 7876 9076 7880 9132
rect 7816 9072 7880 9076
rect 7896 9132 7960 9136
rect 7896 9076 7900 9132
rect 7900 9076 7956 9132
rect 7956 9076 7960 9132
rect 7896 9072 7960 9076
rect 7976 9132 8040 9136
rect 7976 9076 7980 9132
rect 7980 9076 8036 9132
rect 8036 9076 8040 9132
rect 7976 9072 8040 9076
rect 8056 9132 8120 9136
rect 8056 9076 8060 9132
rect 8060 9076 8116 9132
rect 8116 9076 8120 9132
rect 8056 9072 8120 9076
rect 14680 9132 14744 9136
rect 14680 9076 14684 9132
rect 14684 9076 14740 9132
rect 14740 9076 14744 9132
rect 14680 9072 14744 9076
rect 14760 9132 14824 9136
rect 14760 9076 14764 9132
rect 14764 9076 14820 9132
rect 14820 9076 14824 9132
rect 14760 9072 14824 9076
rect 14840 9132 14904 9136
rect 14840 9076 14844 9132
rect 14844 9076 14900 9132
rect 14900 9076 14904 9132
rect 14840 9072 14904 9076
rect 14920 9132 14984 9136
rect 14920 9076 14924 9132
rect 14924 9076 14980 9132
rect 14980 9076 14984 9132
rect 14920 9072 14984 9076
rect 4384 8588 4448 8592
rect 4384 8532 4388 8588
rect 4388 8532 4444 8588
rect 4444 8532 4448 8588
rect 4384 8528 4448 8532
rect 4464 8588 4528 8592
rect 4464 8532 4468 8588
rect 4468 8532 4524 8588
rect 4524 8532 4528 8588
rect 4464 8528 4528 8532
rect 4544 8588 4608 8592
rect 4544 8532 4548 8588
rect 4548 8532 4604 8588
rect 4604 8532 4608 8588
rect 4544 8528 4608 8532
rect 4624 8588 4688 8592
rect 4624 8532 4628 8588
rect 4628 8532 4684 8588
rect 4684 8532 4688 8588
rect 4624 8528 4688 8532
rect 11248 8588 11312 8592
rect 11248 8532 11252 8588
rect 11252 8532 11308 8588
rect 11308 8532 11312 8588
rect 11248 8528 11312 8532
rect 11328 8588 11392 8592
rect 11328 8532 11332 8588
rect 11332 8532 11388 8588
rect 11388 8532 11392 8588
rect 11328 8528 11392 8532
rect 11408 8588 11472 8592
rect 11408 8532 11412 8588
rect 11412 8532 11468 8588
rect 11468 8532 11472 8588
rect 11408 8528 11472 8532
rect 11488 8588 11552 8592
rect 11488 8532 11492 8588
rect 11492 8532 11548 8588
rect 11548 8532 11552 8588
rect 11488 8528 11552 8532
rect 18112 8588 18176 8592
rect 18112 8532 18116 8588
rect 18116 8532 18172 8588
rect 18172 8532 18176 8588
rect 18112 8528 18176 8532
rect 18192 8588 18256 8592
rect 18192 8532 18196 8588
rect 18196 8532 18252 8588
rect 18252 8532 18256 8588
rect 18192 8528 18256 8532
rect 18272 8588 18336 8592
rect 18272 8532 18276 8588
rect 18276 8532 18332 8588
rect 18332 8532 18336 8588
rect 18272 8528 18336 8532
rect 18352 8588 18416 8592
rect 18352 8532 18356 8588
rect 18356 8532 18412 8588
rect 18412 8532 18416 8588
rect 18352 8528 18416 8532
rect 7816 8044 7880 8048
rect 7816 7988 7820 8044
rect 7820 7988 7876 8044
rect 7876 7988 7880 8044
rect 7816 7984 7880 7988
rect 7896 8044 7960 8048
rect 7896 7988 7900 8044
rect 7900 7988 7956 8044
rect 7956 7988 7960 8044
rect 7896 7984 7960 7988
rect 7976 8044 8040 8048
rect 7976 7988 7980 8044
rect 7980 7988 8036 8044
rect 8036 7988 8040 8044
rect 7976 7984 8040 7988
rect 8056 8044 8120 8048
rect 8056 7988 8060 8044
rect 8060 7988 8116 8044
rect 8116 7988 8120 8044
rect 8056 7984 8120 7988
rect 14680 8044 14744 8048
rect 14680 7988 14684 8044
rect 14684 7988 14740 8044
rect 14740 7988 14744 8044
rect 14680 7984 14744 7988
rect 14760 8044 14824 8048
rect 14760 7988 14764 8044
rect 14764 7988 14820 8044
rect 14820 7988 14824 8044
rect 14760 7984 14824 7988
rect 14840 8044 14904 8048
rect 14840 7988 14844 8044
rect 14844 7988 14900 8044
rect 14900 7988 14904 8044
rect 14840 7984 14904 7988
rect 14920 8044 14984 8048
rect 14920 7988 14924 8044
rect 14924 7988 14980 8044
rect 14980 7988 14984 8044
rect 14920 7984 14984 7988
rect 4384 7500 4448 7504
rect 4384 7444 4388 7500
rect 4388 7444 4444 7500
rect 4444 7444 4448 7500
rect 4384 7440 4448 7444
rect 4464 7500 4528 7504
rect 4464 7444 4468 7500
rect 4468 7444 4524 7500
rect 4524 7444 4528 7500
rect 4464 7440 4528 7444
rect 4544 7500 4608 7504
rect 4544 7444 4548 7500
rect 4548 7444 4604 7500
rect 4604 7444 4608 7500
rect 4544 7440 4608 7444
rect 4624 7500 4688 7504
rect 4624 7444 4628 7500
rect 4628 7444 4684 7500
rect 4684 7444 4688 7500
rect 4624 7440 4688 7444
rect 11248 7500 11312 7504
rect 11248 7444 11252 7500
rect 11252 7444 11308 7500
rect 11308 7444 11312 7500
rect 11248 7440 11312 7444
rect 11328 7500 11392 7504
rect 11328 7444 11332 7500
rect 11332 7444 11388 7500
rect 11388 7444 11392 7500
rect 11328 7440 11392 7444
rect 11408 7500 11472 7504
rect 11408 7444 11412 7500
rect 11412 7444 11468 7500
rect 11468 7444 11472 7500
rect 11408 7440 11472 7444
rect 11488 7500 11552 7504
rect 11488 7444 11492 7500
rect 11492 7444 11548 7500
rect 11548 7444 11552 7500
rect 11488 7440 11552 7444
rect 18112 7500 18176 7504
rect 18112 7444 18116 7500
rect 18116 7444 18172 7500
rect 18172 7444 18176 7500
rect 18112 7440 18176 7444
rect 18192 7500 18256 7504
rect 18192 7444 18196 7500
rect 18196 7444 18252 7500
rect 18252 7444 18256 7500
rect 18192 7440 18256 7444
rect 18272 7500 18336 7504
rect 18272 7444 18276 7500
rect 18276 7444 18332 7500
rect 18332 7444 18336 7500
rect 18272 7440 18336 7444
rect 18352 7500 18416 7504
rect 18352 7444 18356 7500
rect 18356 7444 18412 7500
rect 18412 7444 18416 7500
rect 18352 7440 18416 7444
rect 7816 6956 7880 6960
rect 7816 6900 7820 6956
rect 7820 6900 7876 6956
rect 7876 6900 7880 6956
rect 7816 6896 7880 6900
rect 7896 6956 7960 6960
rect 7896 6900 7900 6956
rect 7900 6900 7956 6956
rect 7956 6900 7960 6956
rect 7896 6896 7960 6900
rect 7976 6956 8040 6960
rect 7976 6900 7980 6956
rect 7980 6900 8036 6956
rect 8036 6900 8040 6956
rect 7976 6896 8040 6900
rect 8056 6956 8120 6960
rect 8056 6900 8060 6956
rect 8060 6900 8116 6956
rect 8116 6900 8120 6956
rect 8056 6896 8120 6900
rect 14680 6956 14744 6960
rect 14680 6900 14684 6956
rect 14684 6900 14740 6956
rect 14740 6900 14744 6956
rect 14680 6896 14744 6900
rect 14760 6956 14824 6960
rect 14760 6900 14764 6956
rect 14764 6900 14820 6956
rect 14820 6900 14824 6956
rect 14760 6896 14824 6900
rect 14840 6956 14904 6960
rect 14840 6900 14844 6956
rect 14844 6900 14900 6956
rect 14900 6900 14904 6956
rect 14840 6896 14904 6900
rect 14920 6956 14984 6960
rect 14920 6900 14924 6956
rect 14924 6900 14980 6956
rect 14980 6900 14984 6956
rect 14920 6896 14984 6900
rect 4384 6412 4448 6416
rect 4384 6356 4388 6412
rect 4388 6356 4444 6412
rect 4444 6356 4448 6412
rect 4384 6352 4448 6356
rect 4464 6412 4528 6416
rect 4464 6356 4468 6412
rect 4468 6356 4524 6412
rect 4524 6356 4528 6412
rect 4464 6352 4528 6356
rect 4544 6412 4608 6416
rect 4544 6356 4548 6412
rect 4548 6356 4604 6412
rect 4604 6356 4608 6412
rect 4544 6352 4608 6356
rect 4624 6412 4688 6416
rect 4624 6356 4628 6412
rect 4628 6356 4684 6412
rect 4684 6356 4688 6412
rect 4624 6352 4688 6356
rect 11248 6412 11312 6416
rect 11248 6356 11252 6412
rect 11252 6356 11308 6412
rect 11308 6356 11312 6412
rect 11248 6352 11312 6356
rect 11328 6412 11392 6416
rect 11328 6356 11332 6412
rect 11332 6356 11388 6412
rect 11388 6356 11392 6412
rect 11328 6352 11392 6356
rect 11408 6412 11472 6416
rect 11408 6356 11412 6412
rect 11412 6356 11468 6412
rect 11468 6356 11472 6412
rect 11408 6352 11472 6356
rect 11488 6412 11552 6416
rect 11488 6356 11492 6412
rect 11492 6356 11548 6412
rect 11548 6356 11552 6412
rect 11488 6352 11552 6356
rect 18112 6412 18176 6416
rect 18112 6356 18116 6412
rect 18116 6356 18172 6412
rect 18172 6356 18176 6412
rect 18112 6352 18176 6356
rect 18192 6412 18256 6416
rect 18192 6356 18196 6412
rect 18196 6356 18252 6412
rect 18252 6356 18256 6412
rect 18192 6352 18256 6356
rect 18272 6412 18336 6416
rect 18272 6356 18276 6412
rect 18276 6356 18332 6412
rect 18332 6356 18336 6412
rect 18272 6352 18336 6356
rect 18352 6412 18416 6416
rect 18352 6356 18356 6412
rect 18356 6356 18412 6412
rect 18412 6356 18416 6412
rect 18352 6352 18416 6356
rect 7816 5868 7880 5872
rect 7816 5812 7820 5868
rect 7820 5812 7876 5868
rect 7876 5812 7880 5868
rect 7816 5808 7880 5812
rect 7896 5868 7960 5872
rect 7896 5812 7900 5868
rect 7900 5812 7956 5868
rect 7956 5812 7960 5868
rect 7896 5808 7960 5812
rect 7976 5868 8040 5872
rect 7976 5812 7980 5868
rect 7980 5812 8036 5868
rect 8036 5812 8040 5868
rect 7976 5808 8040 5812
rect 8056 5868 8120 5872
rect 8056 5812 8060 5868
rect 8060 5812 8116 5868
rect 8116 5812 8120 5868
rect 8056 5808 8120 5812
rect 14680 5868 14744 5872
rect 14680 5812 14684 5868
rect 14684 5812 14740 5868
rect 14740 5812 14744 5868
rect 14680 5808 14744 5812
rect 14760 5868 14824 5872
rect 14760 5812 14764 5868
rect 14764 5812 14820 5868
rect 14820 5812 14824 5868
rect 14760 5808 14824 5812
rect 14840 5868 14904 5872
rect 14840 5812 14844 5868
rect 14844 5812 14900 5868
rect 14900 5812 14904 5868
rect 14840 5808 14904 5812
rect 14920 5868 14984 5872
rect 14920 5812 14924 5868
rect 14924 5812 14980 5868
rect 14980 5812 14984 5868
rect 14920 5808 14984 5812
rect 4384 5324 4448 5328
rect 4384 5268 4388 5324
rect 4388 5268 4444 5324
rect 4444 5268 4448 5324
rect 4384 5264 4448 5268
rect 4464 5324 4528 5328
rect 4464 5268 4468 5324
rect 4468 5268 4524 5324
rect 4524 5268 4528 5324
rect 4464 5264 4528 5268
rect 4544 5324 4608 5328
rect 4544 5268 4548 5324
rect 4548 5268 4604 5324
rect 4604 5268 4608 5324
rect 4544 5264 4608 5268
rect 4624 5324 4688 5328
rect 4624 5268 4628 5324
rect 4628 5268 4684 5324
rect 4684 5268 4688 5324
rect 4624 5264 4688 5268
rect 11248 5324 11312 5328
rect 11248 5268 11252 5324
rect 11252 5268 11308 5324
rect 11308 5268 11312 5324
rect 11248 5264 11312 5268
rect 11328 5324 11392 5328
rect 11328 5268 11332 5324
rect 11332 5268 11388 5324
rect 11388 5268 11392 5324
rect 11328 5264 11392 5268
rect 11408 5324 11472 5328
rect 11408 5268 11412 5324
rect 11412 5268 11468 5324
rect 11468 5268 11472 5324
rect 11408 5264 11472 5268
rect 11488 5324 11552 5328
rect 11488 5268 11492 5324
rect 11492 5268 11548 5324
rect 11548 5268 11552 5324
rect 11488 5264 11552 5268
rect 18112 5324 18176 5328
rect 18112 5268 18116 5324
rect 18116 5268 18172 5324
rect 18172 5268 18176 5324
rect 18112 5264 18176 5268
rect 18192 5324 18256 5328
rect 18192 5268 18196 5324
rect 18196 5268 18252 5324
rect 18252 5268 18256 5324
rect 18192 5264 18256 5268
rect 18272 5324 18336 5328
rect 18272 5268 18276 5324
rect 18276 5268 18332 5324
rect 18332 5268 18336 5324
rect 18272 5264 18336 5268
rect 18352 5324 18416 5328
rect 18352 5268 18356 5324
rect 18356 5268 18412 5324
rect 18412 5268 18416 5324
rect 18352 5264 18416 5268
rect 7816 4780 7880 4784
rect 7816 4724 7820 4780
rect 7820 4724 7876 4780
rect 7876 4724 7880 4780
rect 7816 4720 7880 4724
rect 7896 4780 7960 4784
rect 7896 4724 7900 4780
rect 7900 4724 7956 4780
rect 7956 4724 7960 4780
rect 7896 4720 7960 4724
rect 7976 4780 8040 4784
rect 7976 4724 7980 4780
rect 7980 4724 8036 4780
rect 8036 4724 8040 4780
rect 7976 4720 8040 4724
rect 8056 4780 8120 4784
rect 8056 4724 8060 4780
rect 8060 4724 8116 4780
rect 8116 4724 8120 4780
rect 8056 4720 8120 4724
rect 14680 4780 14744 4784
rect 14680 4724 14684 4780
rect 14684 4724 14740 4780
rect 14740 4724 14744 4780
rect 14680 4720 14744 4724
rect 14760 4780 14824 4784
rect 14760 4724 14764 4780
rect 14764 4724 14820 4780
rect 14820 4724 14824 4780
rect 14760 4720 14824 4724
rect 14840 4780 14904 4784
rect 14840 4724 14844 4780
rect 14844 4724 14900 4780
rect 14900 4724 14904 4780
rect 14840 4720 14904 4724
rect 14920 4780 14984 4784
rect 14920 4724 14924 4780
rect 14924 4724 14980 4780
rect 14980 4724 14984 4780
rect 14920 4720 14984 4724
rect 4384 4236 4448 4240
rect 4384 4180 4388 4236
rect 4388 4180 4444 4236
rect 4444 4180 4448 4236
rect 4384 4176 4448 4180
rect 4464 4236 4528 4240
rect 4464 4180 4468 4236
rect 4468 4180 4524 4236
rect 4524 4180 4528 4236
rect 4464 4176 4528 4180
rect 4544 4236 4608 4240
rect 4544 4180 4548 4236
rect 4548 4180 4604 4236
rect 4604 4180 4608 4236
rect 4544 4176 4608 4180
rect 4624 4236 4688 4240
rect 4624 4180 4628 4236
rect 4628 4180 4684 4236
rect 4684 4180 4688 4236
rect 4624 4176 4688 4180
rect 11248 4236 11312 4240
rect 11248 4180 11252 4236
rect 11252 4180 11308 4236
rect 11308 4180 11312 4236
rect 11248 4176 11312 4180
rect 11328 4236 11392 4240
rect 11328 4180 11332 4236
rect 11332 4180 11388 4236
rect 11388 4180 11392 4236
rect 11328 4176 11392 4180
rect 11408 4236 11472 4240
rect 11408 4180 11412 4236
rect 11412 4180 11468 4236
rect 11468 4180 11472 4236
rect 11408 4176 11472 4180
rect 11488 4236 11552 4240
rect 11488 4180 11492 4236
rect 11492 4180 11548 4236
rect 11548 4180 11552 4236
rect 11488 4176 11552 4180
rect 18112 4236 18176 4240
rect 18112 4180 18116 4236
rect 18116 4180 18172 4236
rect 18172 4180 18176 4236
rect 18112 4176 18176 4180
rect 18192 4236 18256 4240
rect 18192 4180 18196 4236
rect 18196 4180 18252 4236
rect 18252 4180 18256 4236
rect 18192 4176 18256 4180
rect 18272 4236 18336 4240
rect 18272 4180 18276 4236
rect 18276 4180 18332 4236
rect 18332 4180 18336 4236
rect 18272 4176 18336 4180
rect 18352 4236 18416 4240
rect 18352 4180 18356 4236
rect 18356 4180 18412 4236
rect 18412 4180 18416 4236
rect 18352 4176 18416 4180
rect 7816 3692 7880 3696
rect 7816 3636 7820 3692
rect 7820 3636 7876 3692
rect 7876 3636 7880 3692
rect 7816 3632 7880 3636
rect 7896 3692 7960 3696
rect 7896 3636 7900 3692
rect 7900 3636 7956 3692
rect 7956 3636 7960 3692
rect 7896 3632 7960 3636
rect 7976 3692 8040 3696
rect 7976 3636 7980 3692
rect 7980 3636 8036 3692
rect 8036 3636 8040 3692
rect 7976 3632 8040 3636
rect 8056 3692 8120 3696
rect 8056 3636 8060 3692
rect 8060 3636 8116 3692
rect 8116 3636 8120 3692
rect 8056 3632 8120 3636
rect 14680 3692 14744 3696
rect 14680 3636 14684 3692
rect 14684 3636 14740 3692
rect 14740 3636 14744 3692
rect 14680 3632 14744 3636
rect 14760 3692 14824 3696
rect 14760 3636 14764 3692
rect 14764 3636 14820 3692
rect 14820 3636 14824 3692
rect 14760 3632 14824 3636
rect 14840 3692 14904 3696
rect 14840 3636 14844 3692
rect 14844 3636 14900 3692
rect 14900 3636 14904 3692
rect 14840 3632 14904 3636
rect 14920 3692 14984 3696
rect 14920 3636 14924 3692
rect 14924 3636 14980 3692
rect 14980 3636 14984 3692
rect 14920 3632 14984 3636
rect 4384 3148 4448 3152
rect 4384 3092 4388 3148
rect 4388 3092 4444 3148
rect 4444 3092 4448 3148
rect 4384 3088 4448 3092
rect 4464 3148 4528 3152
rect 4464 3092 4468 3148
rect 4468 3092 4524 3148
rect 4524 3092 4528 3148
rect 4464 3088 4528 3092
rect 4544 3148 4608 3152
rect 4544 3092 4548 3148
rect 4548 3092 4604 3148
rect 4604 3092 4608 3148
rect 4544 3088 4608 3092
rect 4624 3148 4688 3152
rect 4624 3092 4628 3148
rect 4628 3092 4684 3148
rect 4684 3092 4688 3148
rect 4624 3088 4688 3092
rect 11248 3148 11312 3152
rect 11248 3092 11252 3148
rect 11252 3092 11308 3148
rect 11308 3092 11312 3148
rect 11248 3088 11312 3092
rect 11328 3148 11392 3152
rect 11328 3092 11332 3148
rect 11332 3092 11388 3148
rect 11388 3092 11392 3148
rect 11328 3088 11392 3092
rect 11408 3148 11472 3152
rect 11408 3092 11412 3148
rect 11412 3092 11468 3148
rect 11468 3092 11472 3148
rect 11408 3088 11472 3092
rect 11488 3148 11552 3152
rect 11488 3092 11492 3148
rect 11492 3092 11548 3148
rect 11548 3092 11552 3148
rect 11488 3088 11552 3092
rect 18112 3148 18176 3152
rect 18112 3092 18116 3148
rect 18116 3092 18172 3148
rect 18172 3092 18176 3148
rect 18112 3088 18176 3092
rect 18192 3148 18256 3152
rect 18192 3092 18196 3148
rect 18196 3092 18252 3148
rect 18252 3092 18256 3148
rect 18192 3088 18256 3092
rect 18272 3148 18336 3152
rect 18272 3092 18276 3148
rect 18276 3092 18332 3148
rect 18332 3092 18336 3148
rect 18272 3088 18336 3092
rect 18352 3148 18416 3152
rect 18352 3092 18356 3148
rect 18356 3092 18412 3148
rect 18412 3092 18416 3148
rect 18352 3088 18416 3092
rect 7816 2604 7880 2608
rect 7816 2548 7820 2604
rect 7820 2548 7876 2604
rect 7876 2548 7880 2604
rect 7816 2544 7880 2548
rect 7896 2604 7960 2608
rect 7896 2548 7900 2604
rect 7900 2548 7956 2604
rect 7956 2548 7960 2604
rect 7896 2544 7960 2548
rect 7976 2604 8040 2608
rect 7976 2548 7980 2604
rect 7980 2548 8036 2604
rect 8036 2548 8040 2604
rect 7976 2544 8040 2548
rect 8056 2604 8120 2608
rect 8056 2548 8060 2604
rect 8060 2548 8116 2604
rect 8116 2548 8120 2604
rect 8056 2544 8120 2548
rect 14680 2604 14744 2608
rect 14680 2548 14684 2604
rect 14684 2548 14740 2604
rect 14740 2548 14744 2604
rect 14680 2544 14744 2548
rect 14760 2604 14824 2608
rect 14760 2548 14764 2604
rect 14764 2548 14820 2604
rect 14820 2548 14824 2604
rect 14760 2544 14824 2548
rect 14840 2604 14904 2608
rect 14840 2548 14844 2604
rect 14844 2548 14900 2604
rect 14900 2548 14904 2604
rect 14840 2544 14904 2548
rect 14920 2604 14984 2608
rect 14920 2548 14924 2604
rect 14924 2548 14980 2604
rect 14980 2548 14984 2604
rect 14920 2544 14984 2548
rect 4384 2060 4448 2064
rect 4384 2004 4388 2060
rect 4388 2004 4444 2060
rect 4444 2004 4448 2060
rect 4384 2000 4448 2004
rect 4464 2060 4528 2064
rect 4464 2004 4468 2060
rect 4468 2004 4524 2060
rect 4524 2004 4528 2060
rect 4464 2000 4528 2004
rect 4544 2060 4608 2064
rect 4544 2004 4548 2060
rect 4548 2004 4604 2060
rect 4604 2004 4608 2060
rect 4544 2000 4608 2004
rect 4624 2060 4688 2064
rect 4624 2004 4628 2060
rect 4628 2004 4684 2060
rect 4684 2004 4688 2060
rect 4624 2000 4688 2004
rect 11248 2060 11312 2064
rect 11248 2004 11252 2060
rect 11252 2004 11308 2060
rect 11308 2004 11312 2060
rect 11248 2000 11312 2004
rect 11328 2060 11392 2064
rect 11328 2004 11332 2060
rect 11332 2004 11388 2060
rect 11388 2004 11392 2060
rect 11328 2000 11392 2004
rect 11408 2060 11472 2064
rect 11408 2004 11412 2060
rect 11412 2004 11468 2060
rect 11468 2004 11472 2060
rect 11408 2000 11472 2004
rect 11488 2060 11552 2064
rect 11488 2004 11492 2060
rect 11492 2004 11548 2060
rect 11548 2004 11552 2060
rect 11488 2000 11552 2004
rect 18112 2060 18176 2064
rect 18112 2004 18116 2060
rect 18116 2004 18172 2060
rect 18172 2004 18176 2060
rect 18112 2000 18176 2004
rect 18192 2060 18256 2064
rect 18192 2004 18196 2060
rect 18196 2004 18252 2060
rect 18252 2004 18256 2060
rect 18192 2000 18256 2004
rect 18272 2060 18336 2064
rect 18272 2004 18276 2060
rect 18276 2004 18332 2060
rect 18332 2004 18336 2060
rect 18272 2000 18336 2004
rect 18352 2060 18416 2064
rect 18352 2004 18356 2060
rect 18356 2004 18412 2060
rect 18412 2004 18416 2060
rect 18352 2000 18416 2004
<< metal4 >>
rect 4376 19472 4696 20032
rect 4376 19408 4384 19472
rect 4448 19408 4464 19472
rect 4528 19408 4544 19472
rect 4608 19408 4624 19472
rect 4688 19408 4696 19472
rect 4376 18384 4696 19408
rect 4376 18320 4384 18384
rect 4448 18320 4464 18384
rect 4528 18320 4544 18384
rect 4608 18320 4624 18384
rect 4688 18320 4696 18384
rect 4376 17296 4696 18320
rect 4376 17232 4384 17296
rect 4448 17232 4464 17296
rect 4528 17232 4544 17296
rect 4608 17232 4624 17296
rect 4688 17232 4696 17296
rect 4376 16208 4696 17232
rect 4376 16144 4384 16208
rect 4448 16144 4464 16208
rect 4528 16144 4544 16208
rect 4608 16144 4624 16208
rect 4688 16144 4696 16208
rect 4376 15120 4696 16144
rect 4376 15056 4384 15120
rect 4448 15056 4464 15120
rect 4528 15056 4544 15120
rect 4608 15056 4624 15120
rect 4688 15056 4696 15120
rect 4376 14032 4696 15056
rect 4376 13968 4384 14032
rect 4448 13968 4464 14032
rect 4528 13968 4544 14032
rect 4608 13968 4624 14032
rect 4688 13968 4696 14032
rect 4376 12944 4696 13968
rect 4376 12880 4384 12944
rect 4448 12880 4464 12944
rect 4528 12880 4544 12944
rect 4608 12880 4624 12944
rect 4688 12880 4696 12944
rect 4376 11856 4696 12880
rect 4376 11792 4384 11856
rect 4448 11792 4464 11856
rect 4528 11792 4544 11856
rect 4608 11792 4624 11856
rect 4688 11792 4696 11856
rect 4376 10768 4696 11792
rect 4376 10704 4384 10768
rect 4448 10704 4464 10768
rect 4528 10704 4544 10768
rect 4608 10704 4624 10768
rect 4688 10704 4696 10768
rect 4376 9680 4696 10704
rect 4376 9616 4384 9680
rect 4448 9616 4464 9680
rect 4528 9616 4544 9680
rect 4608 9616 4624 9680
rect 4688 9616 4696 9680
rect 4376 8592 4696 9616
rect 4376 8528 4384 8592
rect 4448 8528 4464 8592
rect 4528 8528 4544 8592
rect 4608 8528 4624 8592
rect 4688 8528 4696 8592
rect 4376 7504 4696 8528
rect 4376 7440 4384 7504
rect 4448 7440 4464 7504
rect 4528 7440 4544 7504
rect 4608 7440 4624 7504
rect 4688 7440 4696 7504
rect 4376 6416 4696 7440
rect 4376 6352 4384 6416
rect 4448 6352 4464 6416
rect 4528 6352 4544 6416
rect 4608 6352 4624 6416
rect 4688 6352 4696 6416
rect 4376 5328 4696 6352
rect 4376 5264 4384 5328
rect 4448 5264 4464 5328
rect 4528 5264 4544 5328
rect 4608 5264 4624 5328
rect 4688 5264 4696 5328
rect 4376 4240 4696 5264
rect 4376 4176 4384 4240
rect 4448 4176 4464 4240
rect 4528 4176 4544 4240
rect 4608 4176 4624 4240
rect 4688 4176 4696 4240
rect 4376 3152 4696 4176
rect 4376 3088 4384 3152
rect 4448 3088 4464 3152
rect 4528 3088 4544 3152
rect 4608 3088 4624 3152
rect 4688 3088 4696 3152
rect 4376 2064 4696 3088
rect 4376 2000 4384 2064
rect 4448 2000 4464 2064
rect 4528 2000 4544 2064
rect 4608 2000 4624 2064
rect 4688 2000 4696 2064
rect 4376 1984 4696 2000
rect 7808 20016 8128 20032
rect 7808 19952 7816 20016
rect 7880 19952 7896 20016
rect 7960 19952 7976 20016
rect 8040 19952 8056 20016
rect 8120 19952 8128 20016
rect 7808 18928 8128 19952
rect 7808 18864 7816 18928
rect 7880 18864 7896 18928
rect 7960 18864 7976 18928
rect 8040 18864 8056 18928
rect 8120 18864 8128 18928
rect 7808 17840 8128 18864
rect 7808 17776 7816 17840
rect 7880 17776 7896 17840
rect 7960 17776 7976 17840
rect 8040 17776 8056 17840
rect 8120 17776 8128 17840
rect 7808 16752 8128 17776
rect 7808 16688 7816 16752
rect 7880 16688 7896 16752
rect 7960 16688 7976 16752
rect 8040 16688 8056 16752
rect 8120 16688 8128 16752
rect 7808 15664 8128 16688
rect 7808 15600 7816 15664
rect 7880 15600 7896 15664
rect 7960 15600 7976 15664
rect 8040 15600 8056 15664
rect 8120 15600 8128 15664
rect 7808 14576 8128 15600
rect 7808 14512 7816 14576
rect 7880 14512 7896 14576
rect 7960 14512 7976 14576
rect 8040 14512 8056 14576
rect 8120 14512 8128 14576
rect 7808 13488 8128 14512
rect 7808 13424 7816 13488
rect 7880 13424 7896 13488
rect 7960 13424 7976 13488
rect 8040 13424 8056 13488
rect 8120 13424 8128 13488
rect 7808 12400 8128 13424
rect 7808 12336 7816 12400
rect 7880 12336 7896 12400
rect 7960 12336 7976 12400
rect 8040 12336 8056 12400
rect 8120 12336 8128 12400
rect 7808 11312 8128 12336
rect 7808 11248 7816 11312
rect 7880 11248 7896 11312
rect 7960 11248 7976 11312
rect 8040 11248 8056 11312
rect 8120 11248 8128 11312
rect 7808 10224 8128 11248
rect 7808 10160 7816 10224
rect 7880 10160 7896 10224
rect 7960 10160 7976 10224
rect 8040 10160 8056 10224
rect 8120 10160 8128 10224
rect 7808 9136 8128 10160
rect 7808 9072 7816 9136
rect 7880 9072 7896 9136
rect 7960 9072 7976 9136
rect 8040 9072 8056 9136
rect 8120 9072 8128 9136
rect 7808 8048 8128 9072
rect 7808 7984 7816 8048
rect 7880 7984 7896 8048
rect 7960 7984 7976 8048
rect 8040 7984 8056 8048
rect 8120 7984 8128 8048
rect 7808 6960 8128 7984
rect 7808 6896 7816 6960
rect 7880 6896 7896 6960
rect 7960 6896 7976 6960
rect 8040 6896 8056 6960
rect 8120 6896 8128 6960
rect 7808 5872 8128 6896
rect 7808 5808 7816 5872
rect 7880 5808 7896 5872
rect 7960 5808 7976 5872
rect 8040 5808 8056 5872
rect 8120 5808 8128 5872
rect 7808 4784 8128 5808
rect 7808 4720 7816 4784
rect 7880 4720 7896 4784
rect 7960 4720 7976 4784
rect 8040 4720 8056 4784
rect 8120 4720 8128 4784
rect 7808 3696 8128 4720
rect 7808 3632 7816 3696
rect 7880 3632 7896 3696
rect 7960 3632 7976 3696
rect 8040 3632 8056 3696
rect 8120 3632 8128 3696
rect 7808 2608 8128 3632
rect 7808 2544 7816 2608
rect 7880 2544 7896 2608
rect 7960 2544 7976 2608
rect 8040 2544 8056 2608
rect 8120 2544 8128 2608
rect 7808 1984 8128 2544
rect 11240 19472 11560 20032
rect 11240 19408 11248 19472
rect 11312 19408 11328 19472
rect 11392 19408 11408 19472
rect 11472 19408 11488 19472
rect 11552 19408 11560 19472
rect 11240 18384 11560 19408
rect 11240 18320 11248 18384
rect 11312 18320 11328 18384
rect 11392 18320 11408 18384
rect 11472 18320 11488 18384
rect 11552 18320 11560 18384
rect 11240 17296 11560 18320
rect 11240 17232 11248 17296
rect 11312 17232 11328 17296
rect 11392 17232 11408 17296
rect 11472 17232 11488 17296
rect 11552 17232 11560 17296
rect 11240 16208 11560 17232
rect 11240 16144 11248 16208
rect 11312 16144 11328 16208
rect 11392 16144 11408 16208
rect 11472 16144 11488 16208
rect 11552 16144 11560 16208
rect 11240 15120 11560 16144
rect 11240 15056 11248 15120
rect 11312 15056 11328 15120
rect 11392 15056 11408 15120
rect 11472 15056 11488 15120
rect 11552 15056 11560 15120
rect 11240 14032 11560 15056
rect 11240 13968 11248 14032
rect 11312 13968 11328 14032
rect 11392 13968 11408 14032
rect 11472 13968 11488 14032
rect 11552 13968 11560 14032
rect 11240 12944 11560 13968
rect 11240 12880 11248 12944
rect 11312 12880 11328 12944
rect 11392 12880 11408 12944
rect 11472 12880 11488 12944
rect 11552 12880 11560 12944
rect 11240 11856 11560 12880
rect 11240 11792 11248 11856
rect 11312 11792 11328 11856
rect 11392 11792 11408 11856
rect 11472 11792 11488 11856
rect 11552 11792 11560 11856
rect 11240 10768 11560 11792
rect 11240 10704 11248 10768
rect 11312 10704 11328 10768
rect 11392 10704 11408 10768
rect 11472 10704 11488 10768
rect 11552 10704 11560 10768
rect 11240 9680 11560 10704
rect 11240 9616 11248 9680
rect 11312 9616 11328 9680
rect 11392 9616 11408 9680
rect 11472 9616 11488 9680
rect 11552 9616 11560 9680
rect 11240 8592 11560 9616
rect 11240 8528 11248 8592
rect 11312 8528 11328 8592
rect 11392 8528 11408 8592
rect 11472 8528 11488 8592
rect 11552 8528 11560 8592
rect 11240 7504 11560 8528
rect 11240 7440 11248 7504
rect 11312 7440 11328 7504
rect 11392 7440 11408 7504
rect 11472 7440 11488 7504
rect 11552 7440 11560 7504
rect 11240 6416 11560 7440
rect 11240 6352 11248 6416
rect 11312 6352 11328 6416
rect 11392 6352 11408 6416
rect 11472 6352 11488 6416
rect 11552 6352 11560 6416
rect 11240 5328 11560 6352
rect 11240 5264 11248 5328
rect 11312 5264 11328 5328
rect 11392 5264 11408 5328
rect 11472 5264 11488 5328
rect 11552 5264 11560 5328
rect 11240 4240 11560 5264
rect 11240 4176 11248 4240
rect 11312 4176 11328 4240
rect 11392 4176 11408 4240
rect 11472 4176 11488 4240
rect 11552 4176 11560 4240
rect 11240 3152 11560 4176
rect 11240 3088 11248 3152
rect 11312 3088 11328 3152
rect 11392 3088 11408 3152
rect 11472 3088 11488 3152
rect 11552 3088 11560 3152
rect 11240 2064 11560 3088
rect 11240 2000 11248 2064
rect 11312 2000 11328 2064
rect 11392 2000 11408 2064
rect 11472 2000 11488 2064
rect 11552 2000 11560 2064
rect 11240 1984 11560 2000
rect 14672 20016 14992 20032
rect 14672 19952 14680 20016
rect 14744 19952 14760 20016
rect 14824 19952 14840 20016
rect 14904 19952 14920 20016
rect 14984 19952 14992 20016
rect 14672 18928 14992 19952
rect 14672 18864 14680 18928
rect 14744 18864 14760 18928
rect 14824 18864 14840 18928
rect 14904 18864 14920 18928
rect 14984 18864 14992 18928
rect 14672 17840 14992 18864
rect 14672 17776 14680 17840
rect 14744 17776 14760 17840
rect 14824 17776 14840 17840
rect 14904 17776 14920 17840
rect 14984 17776 14992 17840
rect 14672 16752 14992 17776
rect 14672 16688 14680 16752
rect 14744 16688 14760 16752
rect 14824 16688 14840 16752
rect 14904 16688 14920 16752
rect 14984 16688 14992 16752
rect 14672 15664 14992 16688
rect 14672 15600 14680 15664
rect 14744 15600 14760 15664
rect 14824 15600 14840 15664
rect 14904 15600 14920 15664
rect 14984 15600 14992 15664
rect 14672 14576 14992 15600
rect 14672 14512 14680 14576
rect 14744 14512 14760 14576
rect 14824 14512 14840 14576
rect 14904 14512 14920 14576
rect 14984 14512 14992 14576
rect 14672 13488 14992 14512
rect 14672 13424 14680 13488
rect 14744 13424 14760 13488
rect 14824 13424 14840 13488
rect 14904 13424 14920 13488
rect 14984 13424 14992 13488
rect 14672 12400 14992 13424
rect 14672 12336 14680 12400
rect 14744 12336 14760 12400
rect 14824 12336 14840 12400
rect 14904 12336 14920 12400
rect 14984 12336 14992 12400
rect 14672 11312 14992 12336
rect 14672 11248 14680 11312
rect 14744 11248 14760 11312
rect 14824 11248 14840 11312
rect 14904 11248 14920 11312
rect 14984 11248 14992 11312
rect 14672 10224 14992 11248
rect 14672 10160 14680 10224
rect 14744 10160 14760 10224
rect 14824 10160 14840 10224
rect 14904 10160 14920 10224
rect 14984 10160 14992 10224
rect 14672 9136 14992 10160
rect 14672 9072 14680 9136
rect 14744 9072 14760 9136
rect 14824 9072 14840 9136
rect 14904 9072 14920 9136
rect 14984 9072 14992 9136
rect 14672 8048 14992 9072
rect 14672 7984 14680 8048
rect 14744 7984 14760 8048
rect 14824 7984 14840 8048
rect 14904 7984 14920 8048
rect 14984 7984 14992 8048
rect 14672 6960 14992 7984
rect 14672 6896 14680 6960
rect 14744 6896 14760 6960
rect 14824 6896 14840 6960
rect 14904 6896 14920 6960
rect 14984 6896 14992 6960
rect 14672 5872 14992 6896
rect 14672 5808 14680 5872
rect 14744 5808 14760 5872
rect 14824 5808 14840 5872
rect 14904 5808 14920 5872
rect 14984 5808 14992 5872
rect 14672 4784 14992 5808
rect 14672 4720 14680 4784
rect 14744 4720 14760 4784
rect 14824 4720 14840 4784
rect 14904 4720 14920 4784
rect 14984 4720 14992 4784
rect 14672 3696 14992 4720
rect 14672 3632 14680 3696
rect 14744 3632 14760 3696
rect 14824 3632 14840 3696
rect 14904 3632 14920 3696
rect 14984 3632 14992 3696
rect 14672 2608 14992 3632
rect 14672 2544 14680 2608
rect 14744 2544 14760 2608
rect 14824 2544 14840 2608
rect 14904 2544 14920 2608
rect 14984 2544 14992 2608
rect 14672 1984 14992 2544
rect 18104 19472 18424 20032
rect 18104 19408 18112 19472
rect 18176 19408 18192 19472
rect 18256 19408 18272 19472
rect 18336 19408 18352 19472
rect 18416 19408 18424 19472
rect 18104 18384 18424 19408
rect 18104 18320 18112 18384
rect 18176 18320 18192 18384
rect 18256 18320 18272 18384
rect 18336 18320 18352 18384
rect 18416 18320 18424 18384
rect 18104 17296 18424 18320
rect 18104 17232 18112 17296
rect 18176 17232 18192 17296
rect 18256 17232 18272 17296
rect 18336 17232 18352 17296
rect 18416 17232 18424 17296
rect 18104 16208 18424 17232
rect 18104 16144 18112 16208
rect 18176 16144 18192 16208
rect 18256 16144 18272 16208
rect 18336 16144 18352 16208
rect 18416 16144 18424 16208
rect 18104 15120 18424 16144
rect 18104 15056 18112 15120
rect 18176 15056 18192 15120
rect 18256 15056 18272 15120
rect 18336 15056 18352 15120
rect 18416 15056 18424 15120
rect 18104 14032 18424 15056
rect 18104 13968 18112 14032
rect 18176 13968 18192 14032
rect 18256 13968 18272 14032
rect 18336 13968 18352 14032
rect 18416 13968 18424 14032
rect 18104 12944 18424 13968
rect 18104 12880 18112 12944
rect 18176 12880 18192 12944
rect 18256 12880 18272 12944
rect 18336 12880 18352 12944
rect 18416 12880 18424 12944
rect 18104 11856 18424 12880
rect 18104 11792 18112 11856
rect 18176 11792 18192 11856
rect 18256 11792 18272 11856
rect 18336 11792 18352 11856
rect 18416 11792 18424 11856
rect 18104 10768 18424 11792
rect 18104 10704 18112 10768
rect 18176 10704 18192 10768
rect 18256 10704 18272 10768
rect 18336 10704 18352 10768
rect 18416 10704 18424 10768
rect 18104 9680 18424 10704
rect 18104 9616 18112 9680
rect 18176 9616 18192 9680
rect 18256 9616 18272 9680
rect 18336 9616 18352 9680
rect 18416 9616 18424 9680
rect 18104 8592 18424 9616
rect 18104 8528 18112 8592
rect 18176 8528 18192 8592
rect 18256 8528 18272 8592
rect 18336 8528 18352 8592
rect 18416 8528 18424 8592
rect 18104 7504 18424 8528
rect 18104 7440 18112 7504
rect 18176 7440 18192 7504
rect 18256 7440 18272 7504
rect 18336 7440 18352 7504
rect 18416 7440 18424 7504
rect 18104 6416 18424 7440
rect 18104 6352 18112 6416
rect 18176 6352 18192 6416
rect 18256 6352 18272 6416
rect 18336 6352 18352 6416
rect 18416 6352 18424 6416
rect 18104 5328 18424 6352
rect 18104 5264 18112 5328
rect 18176 5264 18192 5328
rect 18256 5264 18272 5328
rect 18336 5264 18352 5328
rect 18416 5264 18424 5328
rect 18104 4240 18424 5264
rect 18104 4176 18112 4240
rect 18176 4176 18192 4240
rect 18256 4176 18272 4240
rect 18336 4176 18352 4240
rect 18416 4176 18424 4240
rect 18104 3152 18424 4176
rect 18104 3088 18112 3152
rect 18176 3088 18192 3152
rect 18256 3088 18272 3152
rect 18336 3088 18352 3152
rect 18416 3088 18424 3152
rect 18104 2064 18424 3088
rect 18104 2000 18112 2064
rect 18176 2000 18192 2064
rect 18256 2000 18272 2064
rect 18336 2000 18352 2064
rect 18416 2000 18424 2064
rect 18104 1984 18424 2000
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1605641404
transform 1 0 2484 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1605641404
transform 1 0 1380 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1605641404
transform 1 0 2484 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 3956 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3588 0 -1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1605641404
transform 1 0 4048 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1605641404
transform 1 0 3588 0 1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1605641404
transform 1 0 4048 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 6808 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 5152 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6256 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1605641404
transform 1 0 5152 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1605641404
transform 1 0 6256 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1605641404
transform 1 0 8004 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1605641404
transform 1 0 7360 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1605641404
transform 1 0 8464 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9660 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 9568 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1605641404
transform 1 0 9108 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1605641404
transform 1 0 9752 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1605641404
transform 1 0 9660 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 12512 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1605641404
transform 1 0 10856 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1605641404
transform 1 0 11960 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1605641404
transform 1 0 12604 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_105
timestamp 1605641404
transform 1 0 10764 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1605641404
transform 1 0 11868 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1605641404
transform 1 0 13708 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1605641404
transform 1 0 12972 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_141
timestamp 1605641404
transform 1 0 14076 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15364 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 15180 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1605641404
transform 1 0 14812 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1605641404
transform 1 0 15456 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1605641404
transform 1 0 15272 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_166
timestamp 1605641404
transform 1 0 16376 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 18216 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1605641404
transform 1 0 16560 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1605641404
transform 1 0 17664 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1605641404
transform 1 0 18308 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_178
timestamp 1605641404
transform 1 0 17480 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1605641404
transform 1 0 19412 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1605641404
transform 1 0 18584 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_202
timestamp 1605641404
transform 1 0 19688 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 21620 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 21620 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 21068 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 20792 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1605641404
transform 1 0 20516 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 21160 0 -1 2576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1605641404
transform 1 0 20884 0 1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 21252 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1605641404
transform 1 0 2484 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_27
timestamp 1605641404
transform 1 0 3588 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1605641404
transform 1 0 4692 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 6716 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5796 0 -1 3664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59
timestamp 1605641404
transform 1 0 6532 0 -1 3664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1605641404
transform 1 0 6808 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_74
timestamp 1605641404
transform 1 0 7912 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_86
timestamp 1605641404
transform 1 0 9016 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_98
timestamp 1605641404
transform 1 0 10120 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 12328 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_110
timestamp 1605641404
transform 1 0 11224 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1605641404
transform 1 0 12420 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_135
timestamp 1605641404
transform 1 0 13524 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_147
timestamp 1605641404
transform 1 0 14628 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_159
timestamp 1605641404
transform 1 0 15732 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 17940 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1605641404
transform 1 0 16836 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1605641404
transform 1 0 18032 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_196
timestamp 1605641404
transform 1 0 19136 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_208
timestamp 1605641404
transform 1 0 20240 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 21620 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1605641404
transform 1 0 2484 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 3956 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1605641404
transform 1 0 3588 0 1 3664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1605641404
transform 1 0 4048 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1605641404
transform 1 0 5152 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_56
timestamp 1605641404
transform 1 0 6256 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1605641404
transform 1 0 7360 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1605641404
transform 1 0 8464 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 9568 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1605641404
transform 1 0 9660 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_105
timestamp 1605641404
transform 1 0 10764 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_117
timestamp 1605641404
transform 1 0 11868 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_129
timestamp 1605641404
transform 1 0 12972 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_141
timestamp 1605641404
transform 1 0 14076 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 15180 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_154
timestamp 1605641404
transform 1 0 15272 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_166
timestamp 1605641404
transform 1 0 16376 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_178
timestamp 1605641404
transform 1 0 17480 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_190
timestamp 1605641404
transform 1 0 18584 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_202
timestamp 1605641404
transform 1 0 19688 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 21620 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 20792 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_215
timestamp 1605641404
transform 1 0 20884 0 1 3664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_219
timestamp 1605641404
transform 1 0 21252 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1605641404
transform 1 0 2484 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_27
timestamp 1605641404
transform 1 0 3588 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_39
timestamp 1605641404
transform 1 0 4692 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 6716 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_51
timestamp 1605641404
transform 1 0 5796 0 -1 4752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1605641404
transform 1 0 6532 0 -1 4752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1605641404
transform 1 0 6808 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_74
timestamp 1605641404
transform 1 0 7912 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_86
timestamp 1605641404
transform 1 0 9016 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1605641404
transform 1 0 10120 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 12328 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1605641404
transform 1 0 11224 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1605641404
transform 1 0 12420 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_135
timestamp 1605641404
transform 1 0 13524 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_147
timestamp 1605641404
transform 1 0 14628 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_159
timestamp 1605641404
transform 1 0 15732 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 17940 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_171
timestamp 1605641404
transform 1 0 16836 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1605641404
transform 1 0 18032 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1605641404
transform 1 0 19136 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_208
timestamp 1605641404
transform 1 0 20240 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 20516 0 -1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 21620 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1605641404
transform 1 0 20884 0 -1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1605641404
transform 1 0 21252 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1605641404
transform 1 0 2484 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 3956 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1605641404
transform 1 0 3588 0 1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1605641404
transform 1 0 4048 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1605641404
transform 1 0 5152 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_56
timestamp 1605641404
transform 1 0 6256 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_68
timestamp 1605641404
transform 1 0 7360 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_80
timestamp 1605641404
transform 1 0 8464 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 9568 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1605641404
transform 1 0 9660 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_105
timestamp 1605641404
transform 1 0 10764 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_117
timestamp 1605641404
transform 1 0 11868 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_129
timestamp 1605641404
transform 1 0 12972 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_141
timestamp 1605641404
transform 1 0 14076 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 15180 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_154
timestamp 1605641404
transform 1 0 15272 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_166
timestamp 1605641404
transform 1 0 16376 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_178
timestamp 1605641404
transform 1 0 17480 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_190
timestamp 1605641404
transform 1 0 18584 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_202
timestamp 1605641404
transform 1 0 19688 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 21620 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 20792 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1605641404
transform 1 0 20884 0 1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1605641404
transform 1 0 21252 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1605641404
transform 1 0 2484 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1605641404
transform 1 0 2484 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 3956 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_27
timestamp 1605641404
transform 1 0 3588 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1605641404
transform 1 0 4692 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1605641404
transform 1 0 3588 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1605641404
transform 1 0 4048 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 6716 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1605641404
transform 1 0 5796 0 -1 5840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1605641404
transform 1 0 6532 0 -1 5840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_62
timestamp 1605641404
transform 1 0 6808 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1605641404
transform 1 0 5152 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_56
timestamp 1605641404
transform 1 0 6256 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1605641404
transform 1 0 7912 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1605641404
transform 1 0 7360 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1605641404
transform 1 0 8464 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 9568 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_86
timestamp 1605641404
transform 1 0 9016 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_98
timestamp 1605641404
transform 1 0 10120 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1605641404
transform 1 0 9660 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 12328 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_110
timestamp 1605641404
transform 1 0 11224 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_123
timestamp 1605641404
transform 1 0 12420 0 -1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_105
timestamp 1605641404
transform 1 0 10764 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_117
timestamp 1605641404
transform 1 0 11868 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1605641404
transform 1 0 13984 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1605641404
transform 1 0 12880 0 -1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_127
timestamp 1605641404
transform 1 0 12788 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_132
timestamp 1605641404
transform 1 0 13248 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1605641404
transform 1 0 14352 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_129
timestamp 1605641404
transform 1 0 12972 0 1 5840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_137
timestamp 1605641404
transform 1 0 13708 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_144
timestamp 1605641404
transform 1 0 14352 0 1 5840
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 15180 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_156
timestamp 1605641404
transform 1 0 15456 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_152
timestamp 1605641404
transform 1 0 15088 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_154
timestamp 1605641404
transform 1 0 15272 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_166
timestamp 1605641404
transform 1 0 16376 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 17940 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_168
timestamp 1605641404
transform 1 0 16560 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_180
timestamp 1605641404
transform 1 0 17664 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1605641404
transform 1 0 18032 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_178
timestamp 1605641404
transform 1 0 17480 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1605641404
transform 1 0 19136 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_208
timestamp 1605641404
transform 1 0 20240 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_190
timestamp 1605641404
transform 1 0 18584 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_202
timestamp 1605641404
transform 1 0 19688 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 21620 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 21620 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 20792 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1605641404
transform 1 0 20884 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1605641404
transform 1 0 21252 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1605641404
transform 1 0 2484 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_27
timestamp 1605641404
transform 1 0 3588 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_39
timestamp 1605641404
transform 1 0 4692 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 6716 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1605641404
transform 1 0 5796 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1605641404
transform 1 0 6532 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_62
timestamp 1605641404
transform 1 0 6808 0 -1 6928
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7452 0 -1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_68
timestamp 1605641404
transform 1 0 7360 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10488 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1605641404
transform 1 0 8924 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_97
timestamp 1605641404
transform 1 0 10028 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp 1605641404
transform 1 0 10396 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 12328 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_111
timestamp 1605641404
transform 1 0 11316 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_119
timestamp 1605641404
transform 1 0 12052 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1605641404
transform 1 0 12420 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13616 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_135
timestamp 1605641404
transform 1 0 13524 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_145
timestamp 1605641404
transform 1 0 14444 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_157
timestamp 1605641404
transform 1 0 15548 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 17940 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_169
timestamp 1605641404
transform 1 0 16652 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_181
timestamp 1605641404
transform 1 0 17756 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1605641404
transform 1 0 18032 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_196
timestamp 1605641404
transform 1 0 19136 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_208
timestamp 1605641404
transform 1 0 20240 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 21620 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1605641404
transform 1 0 2484 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 3956 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1605641404
transform 1 0 3588 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1605641404
transform 1 0 4048 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1605641404
transform 1 0 5152 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_56
timestamp 1605641404
transform 1 0 6256 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_68
timestamp 1605641404
transform 1 0 7360 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_80
timestamp 1605641404
transform 1 0 8464 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9936 0 1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 9568 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_93
timestamp 1605641404
transform 1 0 9660 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10948 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12604 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_105
timestamp 1605641404
transform 1 0 10764 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1605641404
transform 1 0 12420 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_141
timestamp 1605641404
transform 1 0 14076 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 15180 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_154
timestamp 1605641404
transform 1 0 15272 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1605641404
transform 1 0 16376 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16560 0 1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_177
timestamp 1605641404
transform 1 0 17388 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_189
timestamp 1605641404
transform 1 0 18492 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_201
timestamp 1605641404
transform 1 0 19596 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 21620 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 20792 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_213
timestamp 1605641404
transform 1 0 20700 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1605641404
transform 1 0 20884 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1605641404
transform 1 0 21252 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1605641404
transform 1 0 2484 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1605641404
transform 1 0 3588 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1605641404
transform 1 0 4692 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 6716 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1605641404
transform 1 0 5796 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1605641404
transform 1 0 6532 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_62
timestamp 1605641404
transform 1 0 6808 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1605641404
transform 1 0 7912 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9016 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10672 0 -1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1605641404
transform 1 0 10488 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11408 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 12328 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_110
timestamp 1605641404
transform 1 0 11224 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_115
timestamp 1605641404
transform 1 0 11684 0 -1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1605641404
transform 1 0 12236 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_123
timestamp 1605641404
transform 1 0 12420 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14168 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13156 0 -1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_140
timestamp 1605641404
transform 1 0 13984 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15824 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_158
timestamp 1605641404
transform 1 0 15640 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18032 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 17940 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_176
timestamp 1605641404
transform 1 0 17296 0 -1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_182
timestamp 1605641404
transform 1 0 17848 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1605641404
transform 1 0 19964 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_200
timestamp 1605641404
transform 1 0 19504 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_204
timestamp 1605641404
transform 1 0 19872 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1605641404
transform 1 0 20516 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 21620 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_209
timestamp 1605641404
transform 1 0 20332 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1605641404
transform 1 0 20884 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1605641404
transform 1 0 21252 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1605641404
transform 1 0 2484 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 3956 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1605641404
transform 1 0 3588 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1605641404
transform 1 0 4048 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1605641404
transform 1 0 5152 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_56
timestamp 1605641404
transform 1 0 6256 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1605641404
transform 1 0 7360 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1605641404
transform 1 0 8464 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 9568 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1605641404
transform 1 0 9660 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1605641404
transform 1 0 11224 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_105
timestamp 1605641404
transform 1 0 10764 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_109
timestamp 1605641404
transform 1 0 11132 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_114
timestamp 1605641404
transform 1 0 11592 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1605641404
transform 1 0 13892 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13156 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_126
timestamp 1605641404
transform 1 0 12696 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_130
timestamp 1605641404
transform 1 0 13064 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_137
timestamp 1605641404
transform 1 0 13708 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_142
timestamp 1605641404
transform 1 0 14168 0 1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16100 0 1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 15180 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_150
timestamp 1605641404
transform 1 0 14904 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_154
timestamp 1605641404
transform 1 0 15272 0 1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_162
timestamp 1605641404
transform 1 0 16008 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1605641404
transform 1 0 17112 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18216 0 1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1605641404
transform 1 0 16928 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_177
timestamp 1605641404
transform 1 0 17388 0 1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_185
timestamp 1605641404
transform 1 0 18124 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1605641404
transform 1 0 20240 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_202
timestamp 1605641404
transform 1 0 19688 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 21620 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 20792 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1605641404
transform 1 0 20608 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1605641404
transform 1 0 20884 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_219
timestamp 1605641404
transform 1 0 21252 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1605641404
transform 1 0 2484 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1605641404
transform 1 0 3588 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1605641404
transform 1 0 4692 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 6716 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_51
timestamp 1605641404
transform 1 0 5796 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1605641404
transform 1 0 6532 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1605641404
transform 1 0 6808 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_74
timestamp 1605641404
transform 1 0 7912 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_86
timestamp 1605641404
transform 1 0 9016 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_98
timestamp 1605641404
transform 1 0 10120 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10948 0 -1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 12328 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_106
timestamp 1605641404
transform 1 0 10856 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_116
timestamp 1605641404
transform 1 0 11776 0 -1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1605641404
transform 1 0 12420 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_135
timestamp 1605641404
transform 1 0 13524 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15272 0 -1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_147
timestamp 1605641404
transform 1 0 14628 0 -1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_153
timestamp 1605641404
transform 1 0 15180 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_160
timestamp 1605641404
transform 1 0 15824 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 17940 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_172
timestamp 1605641404
transform 1 0 16928 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_180
timestamp 1605641404
transform 1 0 17664 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_184
timestamp 1605641404
transform 1 0 18032 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_196
timestamp 1605641404
transform 1 0 19136 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_208
timestamp 1605641404
transform 1 0 20240 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1605641404
transform 1 0 20516 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 21620 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1605641404
transform 1 0 20884 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1605641404
transform 1 0 21252 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1605641404
transform 1 0 2484 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1605641404
transform 1 0 2484 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 3956 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1605641404
transform 1 0 3588 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1605641404
transform 1 0 4048 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_27
timestamp 1605641404
transform 1 0 3588 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_39
timestamp 1605641404
transform 1 0 4692 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1605641404
transform 1 0 6716 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1605641404
transform 1 0 5152 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_56
timestamp 1605641404
transform 1 0 6256 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51
timestamp 1605641404
transform 1 0 5796 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1605641404
transform 1 0 6532 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_62
timestamp 1605641404
transform 1 0 6808 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8188 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_13_68
timestamp 1605641404
transform 1 0 7360 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_80
timestamp 1605641404
transform 1 0 8464 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_74
timestamp 1605641404
transform 1 0 7912 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9844 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 9568 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1605641404
transform 1 0 9660 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1605641404
transform 1 0 9660 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1605641404
transform 1 0 11500 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 11132 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12512 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12420 0 -1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1605641404
transform 1 0 12328 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_105
timestamp 1605641404
transform 1 0 10764 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_118
timestamp 1605641404
transform 1 0 11960 0 1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_111
timestamp 1605641404
transform 1 0 11316 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_116
timestamp 1605641404
transform 1 0 11776 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1605641404
transform 1 0 13524 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13708 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_13_133
timestamp 1605641404
transform 1 0 13340 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1605641404
transform 1 0 13892 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_132
timestamp 1605641404
transform 1 0 13248 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_136
timestamp 1605641404
transform 1 0 13616 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1605641404
transform 1 0 15272 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16008 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1605641404
transform 1 0 15180 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1605641404
transform 1 0 14996 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_158
timestamp 1605641404
transform 1 0 15640 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_153
timestamp 1605641404
transform 1 0 15180 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_161
timestamp 1605641404
transform 1 0 15916 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1605641404
transform 1 0 18216 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1605641404
transform 1 0 17940 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_170
timestamp 1605641404
transform 1 0 16744 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_182
timestamp 1605641404
transform 1 0 17848 0 1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_178
timestamp 1605641404
transform 1 0 17480 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_182
timestamp 1605641404
transform 1 0 17848 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_184
timestamp 1605641404
transform 1 0 18032 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1605641404
transform 1 0 20240 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18676 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18400 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_197
timestamp 1605641404
transform 1 0 19228 0 1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_205
timestamp 1605641404
transform 1 0 19964 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1605641404
transform 1 0 18492 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_207
timestamp 1605641404
transform 1 0 20148 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1605641404
transform 1 0 20516 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 21620 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 21620 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1605641404
transform 1 0 20792 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1605641404
transform 1 0 20608 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1605641404
transform 1 0 20884 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1605641404
transform 1 0 21252 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1605641404
transform 1 0 20884 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1605641404
transform 1 0 21252 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1605641404
transform 1 0 2484 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1605641404
transform 1 0 3956 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1605641404
transform 1 0 3588 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1605641404
transform 1 0 4048 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6624 0 1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1605641404
transform 1 0 5152 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_56
timestamp 1605641404
transform 1 0 6256 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_76
timestamp 1605641404
transform 1 0 8096 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 10304 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1605641404
transform 1 0 9568 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1605641404
transform 1 0 9200 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_93
timestamp 1605641404
transform 1 0 9660 0 1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_99
timestamp 1605641404
transform 1 0 10212 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_109
timestamp 1605641404
transform 1 0 11132 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_120
timestamp 1605641404
transform 1 0 12144 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 13064 0 1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_128
timestamp 1605641404
transform 1 0 12880 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1605641404
transform 1 0 15180 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_146
timestamp 1605641404
transform 1 0 14536 0 1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_152
timestamp 1605641404
transform 1 0 15088 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_154
timestamp 1605641404
transform 1 0 15272 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_166
timestamp 1605641404
transform 1 0 16376 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16468 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_176
timestamp 1605641404
transform 1 0 17296 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1605641404
transform 1 0 20240 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18492 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_188
timestamp 1605641404
transform 1 0 18400 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_198
timestamp 1605641404
transform 1 0 19320 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_206
timestamp 1605641404
transform 1 0 20056 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 21620 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1605641404
transform 1 0 20792 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1605641404
transform 1 0 20608 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_215
timestamp 1605641404
transform 1 0 20884 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_219
timestamp 1605641404
transform 1 0 21252 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1605641404
transform 1 0 2484 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_27
timestamp 1605641404
transform 1 0 3588 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_39
timestamp 1605641404
transform 1 0 4692 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1605641404
transform 1 0 6716 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1605641404
transform 1 0 5796 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1605641404
transform 1 0 6532 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_62
timestamp 1605641404
transform 1 0 6808 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 8372 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_74
timestamp 1605641404
transform 1 0 7912 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_78
timestamp 1605641404
transform 1 0 8280 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_82
timestamp 1605641404
transform 1 0 8648 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_94
timestamp 1605641404
transform 1 0 9752 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1605641404
transform 1 0 12328 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_106
timestamp 1605641404
transform 1 0 10856 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp 1605641404
transform 1 0 11960 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1605641404
transform 1 0 12420 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_135
timestamp 1605641404
transform 1 0 13524 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16376 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_147
timestamp 1605641404
transform 1 0 14628 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_159
timestamp 1605641404
transform 1 0 15732 0 -1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_165
timestamp 1605641404
transform 1 0 16284 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1605641404
transform 1 0 17940 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_175
timestamp 1605641404
transform 1 0 17204 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_184
timestamp 1605641404
transform 1 0 18032 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 19136 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_205
timestamp 1605641404
transform 1 0 19964 0 -1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1605641404
transform 1 0 20516 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 21620 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1605641404
transform 1 0 20884 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1605641404
transform 1 0 21252 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1605641404
transform 1 0 2484 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1605641404
transform 1 0 3956 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1605641404
transform 1 0 3588 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1605641404
transform 1 0 4048 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1605641404
transform 1 0 5152 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_56
timestamp 1605641404
transform 1 0 6256 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1605641404
transform 1 0 7912 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_68
timestamp 1605641404
transform 1 0 7360 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_83
timestamp 1605641404
transform 1 0 8740 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1605641404
transform 1 0 9568 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_91
timestamp 1605641404
transform 1 0 9476 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1605641404
transform 1 0 9660 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11040 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_105
timestamp 1605641404
transform 1 0 10764 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_114
timestamp 1605641404
transform 1 0 11592 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 14076 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 13800 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_126
timestamp 1605641404
transform 1 0 12696 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1605641404
transform 1 0 15272 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16100 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1605641404
transform 1 0 15180 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_150
timestamp 1605641404
transform 1 0 14904 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_157
timestamp 1605641404
transform 1 0 15548 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1605641404
transform 1 0 16928 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_184
timestamp 1605641404
transform 1 0 18032 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1605641404
transform 1 0 19596 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1605641404
transform 1 0 20240 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 18584 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1605641404
transform 1 0 19412 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_204
timestamp 1605641404
transform 1 0 19872 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 21620 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1605641404
transform 1 0 20792 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1605641404
transform 1 0 20608 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_215
timestamp 1605641404
transform 1 0 20884 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_219
timestamp 1605641404
transform 1 0 21252 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1605641404
transform 1 0 2484 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_27
timestamp 1605641404
transform 1 0 3588 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_39
timestamp 1605641404
transform 1 0 4692 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1605641404
transform 1 0 6716 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_51
timestamp 1605641404
transform 1 0 5796 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1605641404
transform 1 0 6532 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8648 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_78
timestamp 1605641404
transform 1 0 8280 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10396 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_98
timestamp 1605641404
transform 1 0 10120 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1605641404
transform 1 0 11408 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12420 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1605641404
transform 1 0 12328 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_110
timestamp 1605641404
transform 1 0 11224 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_115
timestamp 1605641404
transform 1 0 11684 0 -1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1605641404
transform 1 0 12236 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14444 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_139
timestamp 1605641404
transform 1 0 13892 0 -1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 16284 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_154
timestamp 1605641404
transform 1 0 15272 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_162
timestamp 1605641404
transform 1 0 16008 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 18032 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1605641404
transform 1 0 17940 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_181
timestamp 1605641404
transform 1 0 17756 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1605641404
transform 1 0 19964 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_193
timestamp 1605641404
transform 1 0 18860 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1605641404
transform 1 0 20516 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 21620 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_209
timestamp 1605641404
transform 1 0 20332 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1605641404
transform 1 0 20884 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1605641404
transform 1 0 21252 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1605641404
transform 1 0 2484 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1605641404
transform 1 0 2484 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1605641404
transform 1 0 3956 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1605641404
transform 1 0 3588 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1605641404
transform 1 0 4048 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_27
timestamp 1605641404
transform 1 0 3588 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_39
timestamp 1605641404
transform 1 0 4692 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1605641404
transform 1 0 6072 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6624 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1605641404
transform 1 0 6716 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1605641404
transform 1 0 5152 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_56
timestamp 1605641404
transform 1 0 6256 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_51
timestamp 1605641404
transform 1 0 5796 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_57
timestamp 1605641404
transform 1 0 6348 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_62
timestamp 1605641404
transform 1 0 6808 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7636 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1605641404
transform 1 0 7452 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_80
timestamp 1605641404
transform 1 0 8464 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_74
timestamp 1605641404
transform 1 0 7912 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9844 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1605641404
transform 1 0 9568 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10120 0 -1 13456
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1605641404
transform 1 0 9660 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_104
timestamp 1605641404
transform 1 0 10672 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_86
timestamp 1605641404
transform 1 0 9016 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 10856 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1605641404
transform 1 0 12328 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_112
timestamp 1605641404
transform 1 0 11408 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_124
timestamp 1605641404
transform 1 0 12512 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_118
timestamp 1605641404
transform 1 0 11960 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1605641404
transform 1 0 12420 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13156 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13708 0 -1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 14168 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 12696 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_129
timestamp 1605641404
transform 1 0 12972 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_140
timestamp 1605641404
transform 1 0 13984 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_135
timestamp 1605641404
transform 1 0 13524 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16100 0 1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15272 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1605641404
transform 1 0 15180 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_151
timestamp 1605641404
transform 1 0 14996 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_160
timestamp 1605641404
transform 1 0 15824 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_146
timestamp 1605641404
transform 1 0 14536 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_158
timestamp 1605641404
transform 1 0 15640 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1605641404
transform 1 0 17940 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_179
timestamp 1605641404
transform 1 0 17572 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_170
timestamp 1605641404
transform 1 0 16744 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_182
timestamp 1605641404
transform 1 0 17848 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_184
timestamp 1605641404
transform 1 0 18032 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1605641404
transform 1 0 19504 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1605641404
transform 1 0 19688 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1605641404
transform 1 0 20240 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18676 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_197
timestamp 1605641404
transform 1 0 19228 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_201
timestamp 1605641404
transform 1 0 19596 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_206
timestamp 1605641404
transform 1 0 20056 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_196
timestamp 1605641404
transform 1 0 19136 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_204
timestamp 1605641404
transform 1 0 19872 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_210
timestamp 1605641404
transform 1 0 20424 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_212
timestamp 1605641404
transform 1 0 20608 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1605641404
transform 1 0 20516 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1605641404
transform 1 0 20884 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_215
timestamp 1605641404
transform 1 0 20884 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1605641404
transform 1 0 20792 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1605641404
transform 1 0 21252 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_219
timestamp 1605641404
transform 1 0 21252 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 21620 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 21620 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2300 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1605641404
transform 1 0 2116 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4784 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1605641404
transform 1 0 3956 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1605641404
transform 1 0 3772 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_32
timestamp 1605641404
transform 1 0 4048 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6440 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_56
timestamp 1605641404
transform 1 0 6256 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8004 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_67
timestamp 1605641404
transform 1 0 7268 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9844 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1605641404
transform 1 0 9568 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 9016 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_84
timestamp 1605641404
transform 1 0 8832 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_89
timestamp 1605641404
transform 1 0 9292 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1605641404
transform 1 0 9660 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_111
timestamp 1605641404
transform 1 0 11316 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_123
timestamp 1605641404
transform 1 0 12420 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1605641404
transform 1 0 12696 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1605641404
transform 1 0 13524 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1605641404
transform 1 0 15180 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_147
timestamp 1605641404
transform 1 0 14628 0 1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_154
timestamp 1605641404
transform 1 0 15272 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1605641404
transform 1 0 16376 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16560 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18124 0 1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_177
timestamp 1605641404
transform 1 0 17388 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1605641404
transform 1 0 20240 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1605641404
transform 1 0 19688 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_191
timestamp 1605641404
transform 1 0 18676 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_199
timestamp 1605641404
transform 1 0 19412 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1605641404
transform 1 0 20056 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 21620 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1605641404
transform 1 0 20792 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1605641404
transform 1 0 20608 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_215
timestamp 1605641404
transform 1 0 20884 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_219
timestamp 1605641404
transform 1 0 21252 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1605641404
transform 1 0 2484 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3864 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_22_27
timestamp 1605641404
transform 1 0 3588 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5612 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1605641404
transform 1 0 6716 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_46
timestamp 1605641404
transform 1 0 5336 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_58
timestamp 1605641404
transform 1 0 6440 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_62
timestamp 1605641404
transform 1 0 6808 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7268 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_66
timestamp 1605641404
transform 1 0 7176 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_83
timestamp 1605641404
transform 1 0 8740 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1605641404
transform 1 0 9752 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10672 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_22_91
timestamp 1605641404
transform 1 0 9476 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_97
timestamp 1605641404
transform 1 0 10028 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_103
timestamp 1605641404
transform 1 0 10580 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12420 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1605641404
transform 1 0 12328 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_120
timestamp 1605641404
transform 1 0 12144 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1605641404
transform 1 0 13432 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14168 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1605641404
transform 1 0 13248 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_137
timestamp 1605641404
transform 1 0 13708 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1605641404
transform 1 0 14076 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15824 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_158
timestamp 1605641404
transform 1 0 15640 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1605641404
transform 1 0 17480 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1605641404
transform 1 0 17940 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_176
timestamp 1605641404
transform 1 0 17296 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_181
timestamp 1605641404
transform 1 0 17756 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_184
timestamp 1605641404
transform 1 0 18032 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1605641404
transform 1 0 18492 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19780 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19044 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_188
timestamp 1605641404
transform 1 0 18400 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_193
timestamp 1605641404
transform 1 0 18860 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_201
timestamp 1605641404
transform 1 0 19596 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1605641404
transform 1 0 20516 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 21620 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_209
timestamp 1605641404
transform 1 0 20332 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1605641404
transform 1 0 20884 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1605641404
transform 1 0 21252 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1564 0 1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4048 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1605641404
transform 1 0 3956 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_21
timestamp 1605641404
transform 1 0 3036 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_29
timestamp 1605641404
transform 1 0 3772 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_41
timestamp 1605641404
transform 1 0 4876 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_53
timestamp 1605641404
transform 1 0 5980 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_61
timestamp 1605641404
transform 1 0 6716 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7912 0 1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 6992 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_67
timestamp 1605641404
transform 1 0 7268 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_73
timestamp 1605641404
transform 1 0 7820 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9660 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1605641404
transform 1 0 9568 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_90
timestamp 1605641404
transform 1 0 9384 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_102
timestamp 1605641404
transform 1 0 10488 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12236 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_23_114
timestamp 1605641404
transform 1 0 11592 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_120
timestamp 1605641404
transform 1 0 12144 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 13432 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_130
timestamp 1605641404
transform 1 0 13064 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1605641404
transform 1 0 13708 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16100 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1605641404
transform 1 0 15180 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_149
timestamp 1605641404
transform 1 0 14812 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_154
timestamp 1605641404
transform 1 0 15272 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_162
timestamp 1605641404
transform 1 0 16008 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1605641404
transform 1 0 16928 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_184
timestamp 1605641404
transform 1 0 18032 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1605641404
transform 1 0 20240 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18860 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_192
timestamp 1605641404
transform 1 0 18768 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_199
timestamp 1605641404
transform 1 0 19412 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_207
timestamp 1605641404
transform 1 0 20148 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 21620 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1605641404
transform 1 0 20792 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_212
timestamp 1605641404
transform 1 0 20608 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1605641404
transform 1 0 20884 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1605641404
transform 1 0 21252 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1605641404
transform 1 0 1380 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_15
timestamp 1605641404
transform 1 0 2484 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_19
timestamp 1605641404
transform 1 0 2852 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1605641404
transform 1 0 3956 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4876 0 -1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1605641404
transform 1 0 3772 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_34
timestamp 1605641404
transform 1 0 4232 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_40
timestamp 1605641404
transform 1 0 4784 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1605641404
transform 1 0 6716 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1605641404
transform 1 0 6348 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_62
timestamp 1605641404
transform 1 0 6808 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_74
timestamp 1605641404
transform 1 0 7912 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_86
timestamp 1605641404
transform 1 0 9016 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_98
timestamp 1605641404
transform 1 0 10120 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1605641404
transform 1 0 12328 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_110
timestamp 1605641404
transform 1 0 11224 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1605641404
transform 1 0 12420 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_135
timestamp 1605641404
transform 1 0 13524 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16192 0 -1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_147
timestamp 1605641404
transform 1 0 14628 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1605641404
transform 1 0 15732 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_163
timestamp 1605641404
transform 1 0 16100 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1605641404
transform 1 0 17940 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_173
timestamp 1605641404
transform 1 0 17020 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_181
timestamp 1605641404
transform 1 0 17756 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_184
timestamp 1605641404
transform 1 0 18032 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19596 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18860 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_192
timestamp 1605641404
transform 1 0 18768 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_199
timestamp 1605641404
transform 1 0 19412 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1605641404
transform 1 0 20148 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1605641404
transform 1 0 20516 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 21620 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1605641404
transform 1 0 20884 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1605641404
transform 1 0 21252 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 1748 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1605641404
transform 1 0 1104 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1605641404
transform 1 0 1380 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1605641404
transform 1 0 3956 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_23
timestamp 1605641404
transform 1 0 3220 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_32
timestamp 1605641404
transform 1 0 4048 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5428 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_44
timestamp 1605641404
transform 1 0 5152 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7084 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_63
timestamp 1605641404
transform 1 0 6900 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1605641404
transform 1 0 7912 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1605641404
transform 1 0 9844 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1605641404
transform 1 0 9568 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_86
timestamp 1605641404
transform 1 0 9016 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_93
timestamp 1605641404
transform 1 0 9660 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_98
timestamp 1605641404
transform 1 0 10120 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 11132 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_106
timestamp 1605641404
transform 1 0 10856 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_125
timestamp 1605641404
transform 1 0 12604 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13524 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_133
timestamp 1605641404
transform 1 0 13340 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1605641404
transform 1 0 15180 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_151
timestamp 1605641404
transform 1 0 14996 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_154
timestamp 1605641404
transform 1 0 15272 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_166
timestamp 1605641404
transform 1 0 16376 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16744 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_179
timestamp 1605641404
transform 1 0 17572 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1605641404
transform 1 0 19688 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1605641404
transform 1 0 20240 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_191
timestamp 1605641404
transform 1 0 18676 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_199
timestamp 1605641404
transform 1 0 19412 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_206
timestamp 1605641404
transform 1 0 20056 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1605641404
transform -1 0 21620 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1605641404
transform 1 0 20792 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_212
timestamp 1605641404
transform 1 0 20608 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1605641404
transform 1 0 20884 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1605641404
transform 1 0 21252 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1605641404
transform 1 0 1104 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1605641404
transform 1 0 1104 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1605641404
transform 1 0 1380 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1605641404
transform 1 0 2484 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1605641404
transform 1 0 1380 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_15
timestamp 1605641404
transform 1 0 2484 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_19
timestamp 1605641404
transform 1 0 2852 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4048 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3864 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1605641404
transform 1 0 3956 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_27
timestamp 1605641404
transform 1 0 3588 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_36
timestamp 1605641404
transform 1 0 4416 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1605641404
transform 1 0 3772 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_41
timestamp 1605641404
transform 1 0 4876 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1605641404
transform 1 0 6256 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6808 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1605641404
transform 1 0 6716 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_48
timestamp 1605641404
transform 1 0 5520 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_59
timestamp 1605641404
transform 1 0 6532 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_53
timestamp 1605641404
transform 1 0 5980 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8188 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8096 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 7176 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_71
timestamp 1605641404
transform 1 0 7636 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_65
timestamp 1605641404
transform 1 0 7084 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_72
timestamp 1605641404
transform 1 0 7728 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9844 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9660 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1605641404
transform 1 0 9568 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1605641404
transform 1 0 9660 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_85
timestamp 1605641404
transform 1 0 8924 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_91
timestamp 1605641404
transform 1 0 9476 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_102
timestamp 1605641404
transform 1 0 10488 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_108
timestamp 1605641404
transform 1 0 11040 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_111
timestamp 1605641404
transform 1 0 11316 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11132 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1605641404
transform 1 0 11960 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_123
timestamp 1605641404
transform 1 0 12420 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1605641404
transform 1 0 12144 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1605641404
transform 1 0 12328 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12144 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1605641404
transform 1 0 11868 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12604 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13984 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1605641404
transform 1 0 14076 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1605641404
transform 1 0 14444 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_129
timestamp 1605641404
transform 1 0 12972 0 1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_137
timestamp 1605641404
transform 1 0 13708 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_154
timestamp 1605641404
transform 1 0 15272 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_149
timestamp 1605641404
transform 1 0 14812 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_155
timestamp 1605641404
transform 1 0 15364 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1605641404
transform 1 0 15180 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14536 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_160
timestamp 1605641404
transform 1 0 15824 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_164
timestamp 1605641404
transform 1 0 16192 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_160
timestamp 1605641404
transform 1 0 15824 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1605641404
transform 1 0 15548 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16284 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15916 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1605641404
transform 1 0 17664 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1605641404
transform 1 0 17940 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_181
timestamp 1605641404
transform 1 0 17756 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_184
timestamp 1605641404
transform 1 0 18032 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_177
timestamp 1605641404
transform 1 0 17388 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1605641404
transform 1 0 18676 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19320 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19320 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20056 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_196
timestamp 1605641404
transform 1 0 19136 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_204
timestamp 1605641404
transform 1 0 19872 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_189
timestamp 1605641404
transform 1 0 18492 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_194
timestamp 1605641404
transform 1 0 18952 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_204
timestamp 1605641404
transform 1 0 19872 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_212
timestamp 1605641404
transform 1 0 20608 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_210
timestamp 1605641404
transform 1 0 20424 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1605641404
transform 1 0 20516 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1605641404
transform 1 0 20884 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1605641404
transform 1 0 20884 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1605641404
transform 1 0 20792 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1605641404
transform 1 0 21252 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1605641404
transform 1 0 21252 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1605641404
transform -1 0 21620 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1605641404
transform -1 0 21620 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1564 0 -1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1605641404
transform 1 0 1104 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1605641404
transform 1 0 1380 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1605641404
transform 1 0 3312 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_21
timestamp 1605641404
transform 1 0 3036 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_27
timestamp 1605641404
transform 1 0 3588 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_39
timestamp 1605641404
transform 1 0 4692 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5060 0 -1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1605641404
transform 1 0 6716 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_59
timestamp 1605641404
transform 1 0 6532 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_62
timestamp 1605641404
transform 1 0 6808 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_74
timestamp 1605641404
transform 1 0 7912 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_86
timestamp 1605641404
transform 1 0 9016 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_98
timestamp 1605641404
transform 1 0 10120 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1605641404
transform 1 0 12328 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_110
timestamp 1605641404
transform 1 0 11224 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1605641404
transform 1 0 12420 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_135
timestamp 1605641404
transform 1 0 13524 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_147
timestamp 1605641404
transform 1 0 14628 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_159
timestamp 1605641404
transform 1 0 15732 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1605641404
transform 1 0 17940 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_171
timestamp 1605641404
transform 1 0 16836 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_184
timestamp 1605641404
transform 1 0 18032 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1605641404
transform 1 0 19412 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1605641404
transform 1 0 19964 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_196
timestamp 1605641404
transform 1 0 19136 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_203
timestamp 1605641404
transform 1 0 19780 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1605641404
transform 1 0 20516 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1605641404
transform -1 0 21620 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_209
timestamp 1605641404
transform 1 0 20332 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1605641404
transform 1 0 20884 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1605641404
transform 1 0 21252 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1605641404
transform 1 0 1104 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1605641404
transform 1 0 1380 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1605641404
transform 1 0 2484 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1605641404
transform 1 0 3956 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1605641404
transform 1 0 3588 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1605641404
transform 1 0 4048 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 5152 0 1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_50
timestamp 1605641404
transform 1 0 5704 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1605641404
transform 1 0 6808 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7912 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_83
timestamp 1605641404
transform 1 0 8740 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1605641404
transform 1 0 9568 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_91
timestamp 1605641404
transform 1 0 9476 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1605641404
transform 1 0 9660 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1605641404
transform 1 0 11684 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_105
timestamp 1605641404
transform 1 0 10764 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1605641404
transform 1 0 11500 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_118
timestamp 1605641404
transform 1 0 11960 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12880 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14168 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_126
timestamp 1605641404
transform 1 0 12696 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_137
timestamp 1605641404
transform 1 0 13708 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_141
timestamp 1605641404
transform 1 0 14076 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1605641404
transform 1 0 15180 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_151
timestamp 1605641404
transform 1 0 14996 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_154
timestamp 1605641404
transform 1 0 15272 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_166
timestamp 1605641404
transform 1 0 16376 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_178
timestamp 1605641404
transform 1 0 17480 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1605641404
transform 1 0 20240 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_190
timestamp 1605641404
transform 1 0 18584 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_202
timestamp 1605641404
transform 1 0 19688 0 1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1605641404
transform -1 0 21620 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1605641404
transform 1 0 20792 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_212
timestamp 1605641404
transform 1 0 20608 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1605641404
transform 1 0 20884 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1605641404
transform 1 0 21252 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2392 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1605641404
transform 1 0 1104 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1605641404
transform 1 0 1380 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_11
timestamp 1605641404
transform 1 0 2116 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4692 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_30
timestamp 1605641404
transform 1 0 3864 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1605641404
transform 1 0 4600 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1605641404
transform 1 0 5704 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1605641404
transform 1 0 6716 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_48
timestamp 1605641404
transform 1 0 5520 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_53
timestamp 1605641404
transform 1 0 5980 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8740 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_78
timestamp 1605641404
transform 1 0 8280 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_82
timestamp 1605641404
transform 1 0 8648 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10396 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_99
timestamp 1605641404
transform 1 0 10212 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1605641404
transform 1 0 12328 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_117
timestamp 1605641404
transform 1 0 11868 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_121
timestamp 1605641404
transform 1 0 12236 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1605641404
transform 1 0 14076 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_139
timestamp 1605641404
transform 1 0 13892 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_144
timestamp 1605641404
transform 1 0 14352 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14536 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16192 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_162
timestamp 1605641404
transform 1 0 16008 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18216 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1605641404
transform 1 0 17940 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_180
timestamp 1605641404
transform 1 0 17664 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_184
timestamp 1605641404
transform 1 0 18032 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19320 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_192
timestamp 1605641404
transform 1 0 18768 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_204
timestamp 1605641404
transform 1 0 19872 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1605641404
transform 1 0 20516 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1605641404
transform -1 0 21620 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_210
timestamp 1605641404
transform 1 0 20424 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1605641404
transform 1 0 20884 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1605641404
transform 1 0 21252 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1605641404
transform 1 0 1104 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1605641404
transform 1 0 1380 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1605641404
transform 1 0 2484 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4048 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1605641404
transform 1 0 3956 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_27
timestamp 1605641404
transform 1 0 3588 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_48
timestamp 1605641404
transform 1 0 5520 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_60
timestamp 1605641404
transform 1 0 6624 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1605641404
transform 1 0 8648 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6992 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_80
timestamp 1605641404
transform 1 0 8464 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9844 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1605641404
transform 1 0 9568 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_85
timestamp 1605641404
transform 1 0 8924 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_91
timestamp 1605641404
transform 1 0 9476 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_93
timestamp 1605641404
transform 1 0 9660 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_104
timestamp 1605641404
transform 1 0 10672 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_110
timestamp 1605641404
transform 1 0 11224 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_120
timestamp 1605641404
transform 1 0 12144 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13064 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_128
timestamp 1605641404
transform 1 0 12880 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15824 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1605641404
transform 1 0 15180 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_146
timestamp 1605641404
transform 1 0 14536 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_152
timestamp 1605641404
transform 1 0 15088 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_154
timestamp 1605641404
transform 1 0 15272 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16836 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17848 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1605641404
transform 1 0 16652 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_180
timestamp 1605641404
transform 1 0 17664 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1605641404
transform 1 0 18768 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19320 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20056 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_188
timestamp 1605641404
transform 1 0 18400 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_196
timestamp 1605641404
transform 1 0 19136 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_204
timestamp 1605641404
transform 1 0 19872 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1605641404
transform -1 0 21620 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1605641404
transform 1 0 20792 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1605641404
transform 1 0 20608 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1605641404
transform 1 0 20884 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1605641404
transform 1 0 21252 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1605641404
transform 1 0 1104 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1605641404
transform 1 0 1380 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1605641404
transform 1 0 2484 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4600 0 -1 19984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1605641404
transform 1 0 3956 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1605641404
transform 1 0 3588 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_32
timestamp 1605641404
transform 1 0 4048 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1605641404
transform 1 0 6808 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_47
timestamp 1605641404
transform 1 0 5428 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_59
timestamp 1605641404
transform 1 0 6532 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8096 0 -1 19984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1605641404
transform 1 0 6900 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_75
timestamp 1605641404
transform 1 0 8004 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1605641404
transform 1 0 9660 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1605641404
transform 1 0 8924 0 -1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1605641404
transform 1 0 9752 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1605641404
transform 1 0 12512 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1605641404
transform 1 0 10856 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1605641404
transform 1 0 11960 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1605641404
transform 1 0 12604 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1605641404
transform 1 0 13708 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1605641404
transform 1 0 15364 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1605641404
transform 1 0 14812 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1605641404
transform 1 0 15456 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1605641404
transform 1 0 17204 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1605641404
transform 1 0 18216 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_168
timestamp 1605641404
transform 1 0 16560 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_174
timestamp 1605641404
transform 1 0 17112 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_178
timestamp 1605641404
transform 1 0 17480 0 -1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_187
timestamp 1605641404
transform 1 0 18308 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1605641404
transform 1 0 19136 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1605641404
transform 1 0 18584 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1605641404
transform 1 0 19872 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1605641404
transform 1 0 18952 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_200
timestamp 1605641404
transform 1 0 19504 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_208
timestamp 1605641404
transform 1 0 20240 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1605641404
transform 1 0 20424 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1605641404
transform -1 0 21620 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1605641404
transform 1 0 21068 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_214
timestamp 1605641404
transform 1 0 20792 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1605641404
transform 1 0 21160 0 -1 19984
box -38 -48 222 592
<< labels >>
rlabel metal3 s 0 5576 480 5696 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 17000 480 17120 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 22320 4080 22800 4200 6 chanx_right_in[0]
port 2 nsew default input
rlabel metal3 s 22320 8568 22800 8688 6 chanx_right_in[10]
port 3 nsew default input
rlabel metal3 s 22320 9112 22800 9232 6 chanx_right_in[11]
port 4 nsew default input
rlabel metal3 s 22320 9520 22800 9640 6 chanx_right_in[12]
port 5 nsew default input
rlabel metal3 s 22320 9928 22800 10048 6 chanx_right_in[13]
port 6 nsew default input
rlabel metal3 s 22320 10472 22800 10592 6 chanx_right_in[14]
port 7 nsew default input
rlabel metal3 s 22320 10880 22800 11000 6 chanx_right_in[15]
port 8 nsew default input
rlabel metal3 s 22320 11424 22800 11544 6 chanx_right_in[16]
port 9 nsew default input
rlabel metal3 s 22320 11832 22800 11952 6 chanx_right_in[17]
port 10 nsew default input
rlabel metal3 s 22320 12240 22800 12360 6 chanx_right_in[18]
port 11 nsew default input
rlabel metal3 s 22320 12784 22800 12904 6 chanx_right_in[19]
port 12 nsew default input
rlabel metal3 s 22320 4488 22800 4608 6 chanx_right_in[1]
port 13 nsew default input
rlabel metal3 s 22320 4896 22800 5016 6 chanx_right_in[2]
port 14 nsew default input
rlabel metal3 s 22320 5440 22800 5560 6 chanx_right_in[3]
port 15 nsew default input
rlabel metal3 s 22320 5848 22800 5968 6 chanx_right_in[4]
port 16 nsew default input
rlabel metal3 s 22320 6392 22800 6512 6 chanx_right_in[5]
port 17 nsew default input
rlabel metal3 s 22320 6800 22800 6920 6 chanx_right_in[6]
port 18 nsew default input
rlabel metal3 s 22320 7208 22800 7328 6 chanx_right_in[7]
port 19 nsew default input
rlabel metal3 s 22320 7752 22800 7872 6 chanx_right_in[8]
port 20 nsew default input
rlabel metal3 s 22320 8160 22800 8280 6 chanx_right_in[9]
port 21 nsew default input
rlabel metal3 s 22320 13192 22800 13312 6 chanx_right_out[0]
port 22 nsew default tristate
rlabel metal3 s 22320 17816 22800 17936 6 chanx_right_out[10]
port 23 nsew default tristate
rlabel metal3 s 22320 18224 22800 18344 6 chanx_right_out[11]
port 24 nsew default tristate
rlabel metal3 s 22320 18632 22800 18752 6 chanx_right_out[12]
port 25 nsew default tristate
rlabel metal3 s 22320 19176 22800 19296 6 chanx_right_out[13]
port 26 nsew default tristate
rlabel metal3 s 22320 19584 22800 19704 6 chanx_right_out[14]
port 27 nsew default tristate
rlabel metal3 s 22320 19992 22800 20112 6 chanx_right_out[15]
port 28 nsew default tristate
rlabel metal3 s 22320 20536 22800 20656 6 chanx_right_out[16]
port 29 nsew default tristate
rlabel metal3 s 22320 20944 22800 21064 6 chanx_right_out[17]
port 30 nsew default tristate
rlabel metal3 s 22320 21352 22800 21472 6 chanx_right_out[18]
port 31 nsew default tristate
rlabel metal3 s 22320 21896 22800 22016 6 chanx_right_out[19]
port 32 nsew default tristate
rlabel metal3 s 22320 13600 22800 13720 6 chanx_right_out[1]
port 33 nsew default tristate
rlabel metal3 s 22320 14144 22800 14264 6 chanx_right_out[2]
port 34 nsew default tristate
rlabel metal3 s 22320 14552 22800 14672 6 chanx_right_out[3]
port 35 nsew default tristate
rlabel metal3 s 22320 14960 22800 15080 6 chanx_right_out[4]
port 36 nsew default tristate
rlabel metal3 s 22320 15504 22800 15624 6 chanx_right_out[5]
port 37 nsew default tristate
rlabel metal3 s 22320 15912 22800 16032 6 chanx_right_out[6]
port 38 nsew default tristate
rlabel metal3 s 22320 16320 22800 16440 6 chanx_right_out[7]
port 39 nsew default tristate
rlabel metal3 s 22320 16864 22800 16984 6 chanx_right_out[8]
port 40 nsew default tristate
rlabel metal3 s 22320 17272 22800 17392 6 chanx_right_out[9]
port 41 nsew default tristate
rlabel metal2 s 846 22176 902 22656 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 6366 22176 6422 22656 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 6918 22176 6974 22656 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 7470 22176 7526 22656 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 8022 22176 8078 22656 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 8574 22176 8630 22656 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 9126 22176 9182 22656 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 9678 22176 9734 22656 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 10230 22176 10286 22656 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 10782 22176 10838 22656 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 11334 22176 11390 22656 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 1398 22176 1454 22656 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 1950 22176 2006 22656 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 2502 22176 2558 22656 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 3054 22176 3110 22656 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 3606 22176 3662 22656 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 4158 22176 4214 22656 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 4710 22176 4766 22656 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 5262 22176 5318 22656 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 5814 22176 5870 22656 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 11978 22176 12034 22656 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 17498 22176 17554 22656 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 18050 22176 18106 22656 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 18602 22176 18658 22656 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 19154 22176 19210 22656 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 19706 22176 19762 22656 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 20258 22176 20314 22656 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 20810 22176 20866 22656 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 21362 22176 21418 22656 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 21914 22176 21970 22656 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 22466 22176 22522 22656 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 12530 22176 12586 22656 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 13082 22176 13138 22656 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 13634 22176 13690 22656 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 14186 22176 14242 22656 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 14738 22176 14794 22656 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 15290 22176 15346 22656 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 15842 22176 15898 22656 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 16394 22176 16450 22656 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 16946 22176 17002 22656 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 22320 22304 22800 22424 6 prog_clk
port 82 nsew default input
rlabel metal3 s 22320 2176 22800 2296 6 right_bottom_grid_pin_11_
port 83 nsew default input
rlabel metal3 s 22320 2720 22800 2840 6 right_bottom_grid_pin_13_
port 84 nsew default input
rlabel metal3 s 22320 3128 22800 3248 6 right_bottom_grid_pin_15_
port 85 nsew default input
rlabel metal3 s 22320 3536 22800 3656 6 right_bottom_grid_pin_17_
port 86 nsew default input
rlabel metal3 s 22320 0 22800 120 6 right_bottom_grid_pin_1_
port 87 nsew default input
rlabel metal3 s 22320 408 22800 528 6 right_bottom_grid_pin_3_
port 88 nsew default input
rlabel metal3 s 22320 816 22800 936 6 right_bottom_grid_pin_5_
port 89 nsew default input
rlabel metal3 s 22320 1360 22800 1480 6 right_bottom_grid_pin_7_
port 90 nsew default input
rlabel metal3 s 22320 1768 22800 1888 6 right_bottom_grid_pin_9_
port 91 nsew default input
rlabel metal2 s 294 22176 350 22656 6 top_left_grid_pin_1_
port 92 nsew default input
rlabel metal4 s 4376 1984 4696 20032 6 VPWR
port 93 nsew default input
rlabel metal4 s 7808 1984 8128 20032 6 VGND
port 94 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22656
<< end >>
