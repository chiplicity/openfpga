VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_top
  CLASS BLOCK ;
  FOREIGN fpga_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 1568.660 BY 1557.040 ;
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.110 44.120 141.390 46.520 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 324.650 44.120 324.930 46.520 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1517.080 105.360 1519.480 105.960 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 125.760 51.880 126.360 ;
    END
  END clk
  PIN gfpga_pad_GPIO_A[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 508.650 44.120 508.930 46.520 ;
    END
  END gfpga_pad_GPIO_A[0]
  PIN gfpga_pad_GPIO_A[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 288.960 51.880 289.560 ;
    END
  END gfpga_pad_GPIO_A[1]
  PIN gfpga_pad_GPIO_A[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1517.080 227.760 1519.480 228.360 ;
    END
  END gfpga_pad_GPIO_A[2]
  PIN gfpga_pad_GPIO_A[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1517.080 350.160 1519.480 350.760 ;
    END
  END gfpga_pad_GPIO_A[3]
  PIN gfpga_pad_GPIO_A[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1517.080 472.560 1519.480 473.160 ;
    END
  END gfpga_pad_GPIO_A[4]
  PIN gfpga_pad_GPIO_A[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1517.080 594.960 1519.480 595.560 ;
    END
  END gfpga_pad_GPIO_A[5]
  PIN gfpga_pad_GPIO_A[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 452.160 51.880 452.760 ;
    END
  END gfpga_pad_GPIO_A[6]
  PIN gfpga_pad_GPIO_A[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 141.110 1511.720 141.390 1514.120 ;
    END
  END gfpga_pad_GPIO_A[7]
  PIN gfpga_pad_GPIO_IE[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 324.650 1511.720 324.930 1514.120 ;
    END
  END gfpga_pad_GPIO_IE[0]
  PIN gfpga_pad_GPIO_IE[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 615.360 51.880 615.960 ;
    END
  END gfpga_pad_GPIO_IE[1]
  PIN gfpga_pad_GPIO_IE[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 508.650 1511.720 508.930 1514.120 ;
    END
  END gfpga_pad_GPIO_IE[2]
  PIN gfpga_pad_GPIO_IE[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1517.080 717.360 1519.480 717.960 ;
    END
  END gfpga_pad_GPIO_IE[3]
  PIN gfpga_pad_GPIO_IE[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 778.560 51.880 779.160 ;
    END
  END gfpga_pad_GPIO_IE[4]
  PIN gfpga_pad_GPIO_IE[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1517.080 840.440 1519.480 841.040 ;
    END
  END gfpga_pad_GPIO_IE[5]
  PIN gfpga_pad_GPIO_IE[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.190 44.120 692.470 46.520 ;
    END
  END gfpga_pad_GPIO_IE[6]
  PIN gfpga_pad_GPIO_IE[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1517.080 962.840 1519.480 963.440 ;
    END
  END gfpga_pad_GPIO_IE[7]
  PIN gfpga_pad_GPIO_OE[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1517.080 1085.240 1519.480 1085.840 ;
    END
  END gfpga_pad_GPIO_OE[0]
  PIN gfpga_pad_GPIO_OE[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.190 1511.720 692.470 1514.120 ;
    END
  END gfpga_pad_GPIO_OE[1]
  PIN gfpga_pad_GPIO_OE[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 876.190 44.120 876.470 46.520 ;
    END
  END gfpga_pad_GPIO_OE[2]
  PIN gfpga_pad_GPIO_OE[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 876.190 1511.720 876.470 1514.120 ;
    END
  END gfpga_pad_GPIO_OE[3]
  PIN gfpga_pad_GPIO_OE[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 942.440 51.880 943.040 ;
    END
  END gfpga_pad_GPIO_OE[4]
  PIN gfpga_pad_GPIO_OE[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1059.730 44.120 1060.010 46.520 ;
    END
  END gfpga_pad_GPIO_OE[5]
  PIN gfpga_pad_GPIO_OE[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1059.730 1511.720 1060.010 1514.120 ;
    END
  END gfpga_pad_GPIO_OE[6]
  PIN gfpga_pad_GPIO_OE[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1105.640 51.880 1106.240 ;
    END
  END gfpga_pad_GPIO_OE[7]
  PIN gfpga_pad_GPIO_Y[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1517.080 1207.640 1519.480 1208.240 ;
    END
  END gfpga_pad_GPIO_Y[0]
  PIN gfpga_pad_GPIO_Y[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1517.080 1330.040 1519.480 1330.640 ;
    END
  END gfpga_pad_GPIO_Y[1]
  PIN gfpga_pad_GPIO_Y[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1268.840 51.880 1269.440 ;
    END
  END gfpga_pad_GPIO_Y[2]
  PIN gfpga_pad_GPIO_Y[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1243.730 1511.720 1244.010 1514.120 ;
    END
  END gfpga_pad_GPIO_Y[3]
  PIN gfpga_pad_GPIO_Y[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1243.730 44.120 1244.010 46.520 ;
    END
  END gfpga_pad_GPIO_Y[4]
  PIN gfpga_pad_GPIO_Y[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1517.080 1452.440 1519.480 1453.040 ;
    END
  END gfpga_pad_GPIO_Y[5]
  PIN gfpga_pad_GPIO_Y[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1427.270 1511.720 1427.550 1514.120 ;
    END
  END gfpga_pad_GPIO_Y[6]
  PIN gfpga_pad_GPIO_Y[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1432.040 51.880 1432.640 ;
    END
  END gfpga_pad_GPIO_Y[7]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1427.270 44.120 1427.550 46.520 ;
    END
  END prog_clk
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 1543.660 45.000 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 1568.660 20.000 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 105.000 104.915 1464.295 1452.205 ;
      LAYER met1 ;
        RECT 64.730 46.880 1502.090 1497.240 ;
      LAYER met2 ;
        RECT 64.750 1511.440 140.830 1511.720 ;
        RECT 141.670 1511.440 324.370 1511.720 ;
        RECT 325.210 1511.440 508.370 1511.720 ;
        RECT 509.210 1511.440 691.910 1511.720 ;
        RECT 692.750 1511.440 875.910 1511.720 ;
        RECT 876.750 1511.440 1059.450 1511.720 ;
        RECT 1060.290 1511.440 1243.450 1511.720 ;
        RECT 1244.290 1511.440 1426.990 1511.720 ;
        RECT 1427.830 1511.440 1502.530 1511.720 ;
        RECT 64.750 46.800 1502.530 1511.440 ;
        RECT 64.750 46.520 140.830 46.800 ;
        RECT 141.670 46.520 324.370 46.800 ;
        RECT 325.210 46.520 508.370 46.800 ;
        RECT 509.210 46.520 691.910 46.800 ;
        RECT 692.750 46.520 875.910 46.800 ;
        RECT 876.750 46.520 1059.450 46.800 ;
        RECT 1060.290 46.520 1243.450 46.800 ;
        RECT 1244.290 46.520 1426.990 46.800 ;
        RECT 1427.830 46.520 1502.530 46.800 ;
      LAYER met3 ;
        RECT 51.880 1452.040 1516.680 1452.905 ;
        RECT 51.880 1433.040 1517.080 1452.040 ;
        RECT 52.280 1431.640 1517.080 1433.040 ;
        RECT 51.880 1331.040 1517.080 1431.640 ;
        RECT 51.880 1329.640 1516.680 1331.040 ;
        RECT 51.880 1269.840 1517.080 1329.640 ;
        RECT 52.280 1268.440 1517.080 1269.840 ;
        RECT 51.880 1208.640 1517.080 1268.440 ;
        RECT 51.880 1207.240 1516.680 1208.640 ;
        RECT 51.880 1106.640 1517.080 1207.240 ;
        RECT 52.280 1105.240 1517.080 1106.640 ;
        RECT 51.880 1086.240 1517.080 1105.240 ;
        RECT 51.880 1084.840 1516.680 1086.240 ;
        RECT 51.880 963.840 1517.080 1084.840 ;
        RECT 51.880 962.440 1516.680 963.840 ;
        RECT 51.880 943.440 1517.080 962.440 ;
        RECT 52.280 942.040 1517.080 943.440 ;
        RECT 51.880 841.440 1517.080 942.040 ;
        RECT 51.880 840.040 1516.680 841.440 ;
        RECT 51.880 779.560 1517.080 840.040 ;
        RECT 52.280 778.160 1517.080 779.560 ;
        RECT 51.880 718.360 1517.080 778.160 ;
        RECT 51.880 716.960 1516.680 718.360 ;
        RECT 51.880 616.360 1517.080 716.960 ;
        RECT 52.280 614.960 1517.080 616.360 ;
        RECT 51.880 595.960 1517.080 614.960 ;
        RECT 51.880 594.560 1516.680 595.960 ;
        RECT 51.880 473.560 1517.080 594.560 ;
        RECT 51.880 472.160 1516.680 473.560 ;
        RECT 51.880 453.160 1517.080 472.160 ;
        RECT 52.280 451.760 1517.080 453.160 ;
        RECT 51.880 351.160 1517.080 451.760 ;
        RECT 51.880 349.760 1516.680 351.160 ;
        RECT 51.880 289.960 1517.080 349.760 ;
        RECT 52.280 288.560 1517.080 289.960 ;
        RECT 51.880 228.760 1517.080 288.560 ;
        RECT 51.880 227.360 1516.680 228.760 ;
        RECT 51.880 126.760 1517.080 227.360 ;
        RECT 52.280 125.360 1517.080 126.760 ;
        RECT 51.880 106.360 1517.080 125.360 ;
        RECT 51.880 104.960 1516.680 106.360 ;
        RECT 51.880 60.615 1517.080 104.960 ;
      LAYER met4 ;
        RECT 0.000 0.000 1568.660 1557.040 ;
      LAYER met5 ;
        RECT 0.000 119.200 1568.660 1557.040 ;
  END
END fpga_top
END LIBRARY

