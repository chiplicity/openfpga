magic
tech sky130A
magscale 1 2
timestamp 1606224231
<< locali >>
rect 9781 12155 9815 12257
rect 12633 12155 12667 12257
rect 5825 10999 5859 11237
rect 7573 11135 7607 11237
rect 12725 11135 12759 11237
rect 3065 9503 3099 9673
rect 9965 9367 9999 9537
rect 13001 8959 13035 9061
rect 4445 6171 4479 6341
rect 11897 5559 11931 5865
rect 10885 4471 10919 4709
rect 7573 3383 7607 3485
rect 7205 3043 7239 3145
rect 9137 3043 9171 3145
rect 6929 2431 6963 2601
<< viali >>
rect 4169 14569 4203 14603
rect 7389 14569 7423 14603
rect 10701 14569 10735 14603
rect 11713 14569 11747 14603
rect 13001 14569 13035 14603
rect 13645 14569 13679 14603
rect 15853 14569 15887 14603
rect 2513 14501 2547 14535
rect 14933 14501 14967 14535
rect 2421 14433 2455 14467
rect 4537 14433 4571 14467
rect 5549 14433 5583 14467
rect 5641 14433 5675 14467
rect 7297 14433 7331 14467
rect 9045 14433 9079 14467
rect 9137 14433 9171 14467
rect 10609 14433 10643 14467
rect 11621 14433 11655 14467
rect 14013 14433 14047 14467
rect 14105 14433 14139 14467
rect 14657 14433 14691 14467
rect 2605 14365 2639 14399
rect 4629 14365 4663 14399
rect 4721 14365 4755 14399
rect 5733 14365 5767 14399
rect 7481 14365 7515 14399
rect 9229 14365 9263 14399
rect 10793 14365 10827 14399
rect 11805 14365 11839 14399
rect 13093 14365 13127 14399
rect 13277 14365 13311 14399
rect 14197 14365 14231 14399
rect 15945 14365 15979 14399
rect 16129 14365 16163 14399
rect 2053 14229 2087 14263
rect 5181 14229 5215 14263
rect 6929 14229 6963 14263
rect 8677 14229 8711 14263
rect 10241 14229 10275 14263
rect 11253 14229 11287 14263
rect 12633 14229 12667 14263
rect 15485 14229 15519 14263
rect 4169 14025 4203 14059
rect 8217 14025 8251 14059
rect 8677 14025 8711 14059
rect 14105 14025 14139 14059
rect 15393 14025 15427 14059
rect 2053 13957 2087 13991
rect 3065 13957 3099 13991
rect 9689 13957 9723 13991
rect 11345 13957 11379 13991
rect 13829 13957 13863 13991
rect 2605 13889 2639 13923
rect 3525 13889 3559 13923
rect 3617 13889 3651 13923
rect 4813 13889 4847 13923
rect 5825 13889 5859 13923
rect 6837 13889 6871 13923
rect 9321 13889 9355 13923
rect 10333 13889 10367 13923
rect 11989 13889 12023 13923
rect 14657 13889 14691 13923
rect 15945 13889 15979 13923
rect 2513 13821 2547 13855
rect 5641 13821 5675 13855
rect 7104 13821 7138 13855
rect 9137 13821 9171 13855
rect 12449 13821 12483 13855
rect 14565 13821 14599 13855
rect 3433 13753 3467 13787
rect 4537 13753 4571 13787
rect 9045 13753 9079 13787
rect 10885 13753 10919 13787
rect 11713 13753 11747 13787
rect 12716 13753 12750 13787
rect 15853 13753 15887 13787
rect 2421 13685 2455 13719
rect 4629 13685 4663 13719
rect 5181 13685 5215 13719
rect 5549 13685 5583 13719
rect 6193 13685 6227 13719
rect 10057 13685 10091 13719
rect 10149 13685 10183 13719
rect 11805 13685 11839 13719
rect 14473 13685 14507 13719
rect 15761 13685 15795 13719
rect 4721 13481 4755 13515
rect 7113 13481 7147 13515
rect 7941 13481 7975 13515
rect 9689 13481 9723 13515
rect 10057 13481 10091 13515
rect 10149 13481 10183 13515
rect 13277 13481 13311 13515
rect 13921 13481 13955 13515
rect 16037 13481 16071 13515
rect 2596 13413 2630 13447
rect 5089 13413 5123 13447
rect 6000 13413 6034 13447
rect 9045 13413 9079 13447
rect 11520 13413 11554 13447
rect 13369 13413 13403 13447
rect 2329 13345 2363 13379
rect 8033 13345 8067 13379
rect 8953 13345 8987 13379
rect 10701 13345 10735 13379
rect 14289 13345 14323 13379
rect 15945 13345 15979 13379
rect 5181 13277 5215 13311
rect 5365 13277 5399 13311
rect 5733 13277 5767 13311
rect 8217 13277 8251 13311
rect 9229 13277 9263 13311
rect 10333 13277 10367 13311
rect 11253 13277 11287 13311
rect 13461 13277 13495 13311
rect 14381 13277 14415 13311
rect 14473 13277 14507 13311
rect 16129 13277 16163 13311
rect 12633 13209 12667 13243
rect 3709 13141 3743 13175
rect 7573 13141 7607 13175
rect 8585 13141 8619 13175
rect 10885 13141 10919 13175
rect 12909 13141 12943 13175
rect 15577 13141 15611 13175
rect 4353 12937 4387 12971
rect 4721 12937 4755 12971
rect 5733 12937 5767 12971
rect 9689 12937 9723 12971
rect 11345 12937 11379 12971
rect 8769 12869 8803 12903
rect 10977 12869 11011 12903
rect 2605 12801 2639 12835
rect 2973 12801 3007 12835
rect 5273 12801 5307 12835
rect 6193 12801 6227 12835
rect 6377 12801 6411 12835
rect 7389 12801 7423 12835
rect 9229 12801 9263 12835
rect 10149 12801 10183 12835
rect 10241 12801 10275 12835
rect 11989 12801 12023 12835
rect 13001 12801 13035 12835
rect 2329 12733 2363 12767
rect 3240 12733 3274 12767
rect 5181 12733 5215 12767
rect 10057 12733 10091 12767
rect 10793 12733 10827 12767
rect 12449 12733 12483 12767
rect 14933 12733 14967 12767
rect 7656 12665 7690 12699
rect 11713 12665 11747 12699
rect 13268 12665 13302 12699
rect 15200 12665 15234 12699
rect 1961 12597 1995 12631
rect 2421 12597 2455 12631
rect 5089 12597 5123 12631
rect 6101 12597 6135 12631
rect 11805 12597 11839 12631
rect 12633 12597 12667 12631
rect 14381 12597 14415 12631
rect 16313 12597 16347 12631
rect 1501 12393 1535 12427
rect 2973 12393 3007 12427
rect 8585 12393 8619 12427
rect 11805 12393 11839 12427
rect 12725 12393 12759 12427
rect 14565 12393 14599 12427
rect 15301 12393 15335 12427
rect 15669 12393 15703 12427
rect 4344 12325 4378 12359
rect 6653 12325 6687 12359
rect 7472 12325 7506 12359
rect 10670 12325 10704 12359
rect 2329 12257 2363 12291
rect 3341 12257 3375 12291
rect 6561 12257 6595 12291
rect 9045 12257 9079 12291
rect 9781 12257 9815 12291
rect 9873 12257 9907 12291
rect 10425 12257 10459 12291
rect 12173 12257 12207 12291
rect 12633 12257 12667 12291
rect 13093 12257 13127 12291
rect 2421 12189 2455 12223
rect 2513 12189 2547 12223
rect 3433 12189 3467 12223
rect 3525 12189 3559 12223
rect 4077 12189 4111 12223
rect 6745 12189 6779 12223
rect 7205 12189 7239 12223
rect 13185 12189 13219 12223
rect 13369 12189 13403 12223
rect 13737 12189 13771 12223
rect 14657 12189 14691 12223
rect 14841 12189 14875 12223
rect 15761 12189 15795 12223
rect 15853 12189 15887 12223
rect 9781 12121 9815 12155
rect 12357 12121 12391 12155
rect 12633 12121 12667 12155
rect 1961 12053 1995 12087
rect 5457 12053 5491 12087
rect 6193 12053 6227 12087
rect 9229 12053 9263 12087
rect 10057 12053 10091 12087
rect 14197 12053 14231 12087
rect 9229 11849 9263 11883
rect 10333 11849 10367 11883
rect 15761 11849 15795 11883
rect 8769 11781 8803 11815
rect 11345 11781 11379 11815
rect 6285 11713 6319 11747
rect 9689 11713 9723 11747
rect 9873 11713 9907 11747
rect 10977 11713 11011 11747
rect 11989 11713 12023 11747
rect 1777 11645 1811 11679
rect 3525 11645 3559 11679
rect 3792 11645 3826 11679
rect 7389 11645 7423 11679
rect 10793 11645 10827 11679
rect 11713 11645 11747 11679
rect 12725 11645 12759 11679
rect 14381 11645 14415 11679
rect 16037 11645 16071 11679
rect 2044 11577 2078 11611
rect 6101 11577 6135 11611
rect 6193 11577 6227 11611
rect 7634 11577 7668 11611
rect 10701 11577 10735 11611
rect 12992 11577 13026 11611
rect 14648 11577 14682 11611
rect 3157 11509 3191 11543
rect 4905 11509 4939 11543
rect 5733 11509 5767 11543
rect 6929 11509 6963 11543
rect 9597 11509 9631 11543
rect 11805 11509 11839 11543
rect 14105 11509 14139 11543
rect 16221 11509 16255 11543
rect 1961 11305 1995 11339
rect 2973 11305 3007 11339
rect 4997 11305 5031 11339
rect 7389 11305 7423 11339
rect 7665 11305 7699 11339
rect 10149 11305 10183 11339
rect 15669 11305 15703 11339
rect 3433 11237 3467 11271
rect 5825 11237 5859 11271
rect 1409 11169 1443 11203
rect 2329 11169 2363 11203
rect 3341 11169 3375 11203
rect 4077 11169 4111 11203
rect 4905 11169 4939 11203
rect 5365 11169 5399 11203
rect 2421 11101 2455 11135
rect 2605 11101 2639 11135
rect 3617 11101 3651 11135
rect 5457 11101 5491 11135
rect 5549 11101 5583 11135
rect 1593 11033 1627 11067
rect 7573 11237 7607 11271
rect 8208 11237 8242 11271
rect 9689 11237 9723 11271
rect 12725 11237 12759 11271
rect 15761 11237 15795 11271
rect 6276 11169 6310 11203
rect 7849 11169 7883 11203
rect 7941 11169 7975 11203
rect 10517 11169 10551 11203
rect 10609 11169 10643 11203
rect 11161 11169 11195 11203
rect 11428 11169 11462 11203
rect 13084 11169 13118 11203
rect 14657 11169 14691 11203
rect 16497 11169 16531 11203
rect 6009 11101 6043 11135
rect 7573 11101 7607 11135
rect 10793 11101 10827 11135
rect 12725 11101 12759 11135
rect 12817 11101 12851 11135
rect 15853 11101 15887 11135
rect 12541 11033 12575 11067
rect 15301 11033 15335 11067
rect 16313 11033 16347 11067
rect 4261 10965 4295 10999
rect 4721 10965 4755 10999
rect 5825 10965 5859 10999
rect 9321 10965 9355 10999
rect 14197 10965 14231 10999
rect 14841 10965 14875 10999
rect 2789 10761 2823 10795
rect 3065 10761 3099 10795
rect 4077 10761 4111 10795
rect 10057 10693 10091 10727
rect 11713 10693 11747 10727
rect 11989 10693 12023 10727
rect 12725 10693 12759 10727
rect 16313 10693 16347 10727
rect 3709 10625 3743 10659
rect 4629 10625 4663 10659
rect 5089 10625 5123 10659
rect 7481 10625 7515 10659
rect 8677 10625 8711 10659
rect 10333 10625 10367 10659
rect 13185 10625 13219 10659
rect 13277 10625 13311 10659
rect 14289 10625 14323 10659
rect 14933 10625 14967 10659
rect 1409 10557 1443 10591
rect 3525 10557 3559 10591
rect 4445 10557 4479 10591
rect 5356 10557 5390 10591
rect 8125 10557 8159 10591
rect 8944 10557 8978 10591
rect 10600 10557 10634 10591
rect 12173 10557 12207 10591
rect 15200 10557 15234 10591
rect 1676 10489 1710 10523
rect 7297 10489 7331 10523
rect 14105 10489 14139 10523
rect 3433 10421 3467 10455
rect 4537 10421 4571 10455
rect 6469 10421 6503 10455
rect 6837 10421 6871 10455
rect 7205 10421 7239 10455
rect 8309 10421 8343 10455
rect 13093 10421 13127 10455
rect 13737 10421 13771 10455
rect 14197 10421 14231 10455
rect 3617 10217 3651 10251
rect 4537 10217 4571 10251
rect 4997 10217 5031 10251
rect 5549 10217 5583 10251
rect 6009 10217 6043 10251
rect 6837 10217 6871 10251
rect 7205 10217 7239 10251
rect 7573 10217 7607 10251
rect 8217 10217 8251 10251
rect 8677 10217 8711 10251
rect 10149 10217 10183 10251
rect 15669 10217 15703 10251
rect 2228 10149 2262 10183
rect 5917 10149 5951 10183
rect 8585 10149 8619 10183
rect 9689 10149 9723 10183
rect 12725 10149 12759 10183
rect 12817 10149 12851 10183
rect 13820 10149 13854 10183
rect 1409 10081 1443 10115
rect 1961 10081 1995 10115
rect 3801 10081 3835 10115
rect 4905 10081 4939 10115
rect 6653 10081 6687 10115
rect 9505 10081 9539 10115
rect 10517 10081 10551 10115
rect 11529 10081 11563 10115
rect 13553 10081 13587 10115
rect 15761 10081 15795 10115
rect 5181 10013 5215 10047
rect 6193 10013 6227 10047
rect 7665 10013 7699 10047
rect 7757 10013 7791 10047
rect 8769 10013 8803 10047
rect 10609 10013 10643 10047
rect 10793 10013 10827 10047
rect 11621 10013 11655 10047
rect 11805 10013 11839 10047
rect 13001 10013 13035 10047
rect 15853 10013 15887 10047
rect 9321 9945 9355 9979
rect 1593 9877 1627 9911
rect 3341 9877 3375 9911
rect 11161 9877 11195 9911
rect 12357 9877 12391 9911
rect 14933 9877 14967 9911
rect 15301 9877 15335 9911
rect 3065 9673 3099 9707
rect 8217 9673 8251 9707
rect 10149 9673 10183 9707
rect 16221 9673 16255 9707
rect 2605 9537 2639 9571
rect 2789 9537 2823 9571
rect 5733 9605 5767 9639
rect 11161 9605 11195 9639
rect 13461 9605 13495 9639
rect 6377 9537 6411 9571
rect 9781 9537 9815 9571
rect 9965 9537 9999 9571
rect 10609 9537 10643 9571
rect 10793 9537 10827 9571
rect 11805 9537 11839 9571
rect 13001 9537 13035 9571
rect 14013 9537 14047 9571
rect 14841 9537 14875 9571
rect 1593 9469 1627 9503
rect 3065 9469 3099 9503
rect 3157 9469 3191 9503
rect 3424 9469 3458 9503
rect 4813 9469 4847 9503
rect 6193 9469 6227 9503
rect 6837 9469 6871 9503
rect 7104 9469 7138 9503
rect 8585 9469 8619 9503
rect 2513 9401 2547 9435
rect 9505 9401 9539 9435
rect 10517 9469 10551 9503
rect 12817 9469 12851 9503
rect 13921 9469 13955 9503
rect 12909 9401 12943 9435
rect 15086 9401 15120 9435
rect 1777 9333 1811 9367
rect 2145 9333 2179 9367
rect 4537 9333 4571 9367
rect 4997 9333 5031 9367
rect 6101 9333 6135 9367
rect 8769 9333 8803 9367
rect 9137 9333 9171 9367
rect 9597 9333 9631 9367
rect 9965 9333 9999 9367
rect 11529 9333 11563 9367
rect 11621 9333 11655 9367
rect 12449 9333 12483 9367
rect 13829 9333 13863 9367
rect 1961 9129 1995 9163
rect 3433 9129 3467 9163
rect 4077 9129 4111 9163
rect 4445 9129 4479 9163
rect 4537 9129 4571 9163
rect 14933 9129 14967 9163
rect 15761 9129 15795 9163
rect 9505 9061 9539 9095
rect 13001 9061 13035 9095
rect 1409 8993 1443 9027
rect 2329 8993 2363 9027
rect 2421 8993 2455 9027
rect 3341 8993 3375 9027
rect 5273 8993 5307 9027
rect 5632 8993 5666 9027
rect 7021 8993 7055 9027
rect 7757 8993 7791 9027
rect 9965 8993 9999 9027
rect 10885 8993 10919 9027
rect 11796 8993 11830 9027
rect 13369 8993 13403 9027
rect 13553 8993 13587 9027
rect 13820 8993 13854 9027
rect 15669 8993 15703 9027
rect 2605 8925 2639 8959
rect 3617 8925 3651 8959
rect 4629 8925 4663 8959
rect 5365 8925 5399 8959
rect 10977 8925 11011 8959
rect 11161 8925 11195 8959
rect 11529 8925 11563 8959
rect 13001 8925 13035 8959
rect 15853 8925 15887 8959
rect 6745 8857 6779 8891
rect 10149 8857 10183 8891
rect 13185 8857 13219 8891
rect 1593 8789 1627 8823
rect 2973 8789 3007 8823
rect 5089 8789 5123 8823
rect 7205 8789 7239 8823
rect 10517 8789 10551 8823
rect 12909 8789 12943 8823
rect 15301 8789 15335 8823
rect 9321 8585 9355 8619
rect 10333 8585 10367 8619
rect 14381 8585 14415 8619
rect 2789 8517 2823 8551
rect 5825 8517 5859 8551
rect 15393 8517 15427 8551
rect 3525 8449 3559 8483
rect 3709 8449 3743 8483
rect 7573 8449 7607 8483
rect 9781 8449 9815 8483
rect 9965 8449 9999 8483
rect 10977 8449 11011 8483
rect 11897 8449 11931 8483
rect 12725 8449 12759 8483
rect 14933 8449 14967 8483
rect 15945 8449 15979 8483
rect 1409 8381 1443 8415
rect 1676 8381 1710 8415
rect 3433 8381 3467 8415
rect 4077 8381 4111 8415
rect 4445 8381 4479 8415
rect 9689 8381 9723 8415
rect 10701 8381 10735 8415
rect 10793 8381 10827 8415
rect 11713 8381 11747 8415
rect 14749 8381 14783 8415
rect 14841 8381 14875 8415
rect 4712 8313 4746 8347
rect 6193 8313 6227 8347
rect 6285 8313 6319 8347
rect 7297 8313 7331 8347
rect 7840 8313 7874 8347
rect 11805 8313 11839 8347
rect 12992 8313 13026 8347
rect 15761 8313 15795 8347
rect 15853 8313 15887 8347
rect 3065 8245 3099 8279
rect 4261 8245 4295 8279
rect 8953 8245 8987 8279
rect 11345 8245 11379 8279
rect 14105 8245 14139 8279
rect 2329 8041 2363 8075
rect 2973 8041 3007 8075
rect 7021 8041 7055 8075
rect 7389 8041 7423 8075
rect 8309 8041 8343 8075
rect 8677 8041 8711 8075
rect 12817 8041 12851 8075
rect 13461 8041 13495 8075
rect 15301 8041 15335 8075
rect 2421 7973 2455 8007
rect 5150 7973 5184 8007
rect 7757 7973 7791 8007
rect 10057 7973 10091 8007
rect 1409 7905 1443 7939
rect 3341 7905 3375 7939
rect 4077 7905 4111 7939
rect 6929 7905 6963 7939
rect 7849 7905 7883 7939
rect 9505 7905 9539 7939
rect 10149 7905 10183 7939
rect 10784 7905 10818 7939
rect 13829 7905 13863 7939
rect 13921 7905 13955 7939
rect 14657 7905 14691 7939
rect 15669 7905 15703 7939
rect 2605 7837 2639 7871
rect 3433 7837 3467 7871
rect 3617 7837 3651 7871
rect 4905 7837 4939 7871
rect 7113 7837 7147 7871
rect 7941 7837 7975 7871
rect 8769 7837 8803 7871
rect 8953 7837 8987 7871
rect 10241 7837 10275 7871
rect 10517 7837 10551 7871
rect 12909 7837 12943 7871
rect 13093 7837 13127 7871
rect 14013 7837 14047 7871
rect 15761 7837 15795 7871
rect 15853 7837 15887 7871
rect 6561 7769 6595 7803
rect 9689 7769 9723 7803
rect 11897 7769 11931 7803
rect 1593 7701 1627 7735
rect 1961 7701 1995 7735
rect 4261 7701 4295 7735
rect 6285 7701 6319 7735
rect 9321 7701 9355 7735
rect 12449 7701 12483 7735
rect 14841 7701 14875 7735
rect 6837 7497 6871 7531
rect 11713 7497 11747 7531
rect 13001 7497 13035 7531
rect 15393 7497 15427 7531
rect 2973 7429 3007 7463
rect 13369 7429 13403 7463
rect 1593 7361 1627 7395
rect 3709 7361 3743 7395
rect 3801 7361 3835 7395
rect 4813 7361 4847 7395
rect 5733 7361 5767 7395
rect 5825 7361 5859 7395
rect 7389 7361 7423 7395
rect 7849 7361 7883 7395
rect 10333 7361 10367 7395
rect 13921 7361 13955 7395
rect 14841 7361 14875 7395
rect 15025 7361 15059 7395
rect 15853 7361 15887 7395
rect 15945 7361 15979 7395
rect 1860 7293 1894 7327
rect 7297 7293 7331 7327
rect 8309 7293 8343 7327
rect 9965 7293 9999 7327
rect 10600 7293 10634 7327
rect 12817 7293 12851 7327
rect 15761 7293 15795 7327
rect 3617 7225 3651 7259
rect 8576 7225 8610 7259
rect 13737 7225 13771 7259
rect 3249 7157 3283 7191
rect 4261 7157 4295 7191
rect 4629 7157 4663 7191
rect 4721 7157 4755 7191
rect 5273 7157 5307 7191
rect 5641 7157 5675 7191
rect 6285 7157 6319 7191
rect 7205 7157 7239 7191
rect 9689 7157 9723 7191
rect 10149 7157 10183 7191
rect 13829 7157 13863 7191
rect 14381 7157 14415 7191
rect 14749 7157 14783 7191
rect 4445 6953 4479 6987
rect 11345 6953 11379 6987
rect 13001 6953 13035 6987
rect 14197 6953 14231 6987
rect 14657 6953 14691 6987
rect 15669 6953 15703 6987
rect 8769 6885 8803 6919
rect 1501 6817 1535 6851
rect 2421 6817 2455 6851
rect 3065 6817 3099 6851
rect 3893 6817 3927 6851
rect 5540 6817 5574 6851
rect 6929 6817 6963 6851
rect 7196 6817 7230 6851
rect 9945 6817 9979 6851
rect 11529 6817 11563 6851
rect 11888 6817 11922 6851
rect 13461 6817 13495 6851
rect 13645 6817 13679 6851
rect 14565 6817 14599 6851
rect 2513 6749 2547 6783
rect 2605 6749 2639 6783
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 5273 6749 5307 6783
rect 8861 6749 8895 6783
rect 8953 6749 8987 6783
rect 9689 6749 9723 6783
rect 11621 6749 11655 6783
rect 14841 6749 14875 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 4077 6681 4111 6715
rect 8401 6681 8435 6715
rect 15301 6681 15335 6715
rect 1685 6613 1719 6647
rect 2053 6613 2087 6647
rect 3249 6613 3283 6647
rect 3709 6613 3743 6647
rect 6653 6613 6687 6647
rect 8309 6613 8343 6647
rect 11069 6613 11103 6647
rect 13277 6613 13311 6647
rect 13829 6613 13863 6647
rect 7113 6409 7147 6443
rect 9505 6409 9539 6443
rect 16221 6409 16255 6443
rect 4261 6341 4295 6375
rect 4445 6341 4479 6375
rect 11621 6341 11655 6375
rect 1409 6273 1443 6307
rect 2513 6273 2547 6307
rect 2881 6205 2915 6239
rect 3137 6205 3171 6239
rect 4537 6273 4571 6307
rect 7573 6273 7607 6307
rect 7757 6273 7791 6307
rect 13001 6273 13035 6307
rect 13093 6273 13127 6307
rect 14197 6273 14231 6307
rect 6193 6205 6227 6239
rect 7481 6205 7515 6239
rect 8125 6205 8159 6239
rect 10241 6205 10275 6239
rect 10508 6205 10542 6239
rect 14841 6205 14875 6239
rect 2237 6137 2271 6171
rect 4445 6137 4479 6171
rect 4782 6137 4816 6171
rect 8392 6137 8426 6171
rect 12909 6137 12943 6171
rect 14013 6137 14047 6171
rect 15108 6137 15142 6171
rect 1869 6069 1903 6103
rect 2329 6069 2363 6103
rect 5917 6069 5951 6103
rect 6377 6069 6411 6103
rect 9781 6069 9815 6103
rect 11897 6069 11931 6103
rect 12541 6069 12575 6103
rect 13645 6069 13679 6103
rect 14105 6069 14139 6103
rect 3709 5865 3743 5899
rect 4537 5865 4571 5899
rect 4629 5865 4663 5899
rect 5733 5865 5767 5899
rect 8125 5865 8159 5899
rect 8217 5865 8251 5899
rect 8585 5865 8619 5899
rect 8953 5865 8987 5899
rect 10425 5865 10459 5899
rect 10517 5865 10551 5899
rect 11069 5865 11103 5899
rect 11529 5865 11563 5899
rect 11897 5865 11931 5899
rect 12081 5865 12115 5899
rect 12449 5865 12483 5899
rect 15301 5865 15335 5899
rect 15761 5865 15795 5899
rect 2320 5797 2354 5831
rect 11437 5797 11471 5831
rect 1501 5729 1535 5763
rect 2053 5729 2087 5763
rect 3893 5729 3927 5763
rect 5181 5729 5215 5763
rect 5917 5729 5951 5763
rect 6009 5729 6043 5763
rect 6276 5729 6310 5763
rect 4721 5661 4755 5695
rect 8309 5661 8343 5695
rect 9045 5661 9079 5695
rect 9229 5661 9263 5695
rect 10701 5661 10735 5695
rect 11621 5661 11655 5695
rect 5365 5593 5399 5627
rect 7389 5593 7423 5627
rect 7757 5593 7791 5627
rect 12541 5797 12575 5831
rect 15669 5797 15703 5831
rect 13093 5729 13127 5763
rect 13360 5729 13394 5763
rect 12633 5661 12667 5695
rect 14749 5661 14783 5695
rect 15853 5661 15887 5695
rect 14473 5593 14507 5627
rect 1685 5525 1719 5559
rect 3433 5525 3467 5559
rect 4169 5525 4203 5559
rect 10057 5525 10091 5559
rect 11897 5525 11931 5559
rect 6837 5321 6871 5355
rect 8585 5321 8619 5355
rect 4169 5253 4203 5287
rect 10977 5253 11011 5287
rect 1685 5185 1719 5219
rect 2789 5185 2823 5219
rect 3801 5185 3835 5219
rect 4813 5185 4847 5219
rect 5733 5185 5767 5219
rect 7297 5185 7331 5219
rect 7481 5185 7515 5219
rect 9137 5185 9171 5219
rect 11805 5185 11839 5219
rect 14841 5185 14875 5219
rect 1409 5117 1443 5151
rect 2513 5117 2547 5151
rect 3617 5117 3651 5151
rect 4537 5117 4571 5151
rect 5549 5117 5583 5151
rect 6193 5117 6227 5151
rect 7665 5117 7699 5151
rect 8953 5117 8987 5151
rect 9597 5117 9631 5151
rect 9864 5117 9898 5151
rect 12449 5117 12483 5151
rect 14289 5117 14323 5151
rect 2605 5049 2639 5083
rect 7205 5049 7239 5083
rect 7941 5049 7975 5083
rect 11713 5049 11747 5083
rect 12716 5049 12750 5083
rect 15108 5049 15142 5083
rect 2145 4981 2179 5015
rect 3157 4981 3191 5015
rect 3525 4981 3559 5015
rect 4629 4981 4663 5015
rect 5181 4981 5215 5015
rect 5641 4981 5675 5015
rect 6377 4981 6411 5015
rect 9045 4981 9079 5015
rect 11253 4981 11287 5015
rect 11621 4981 11655 5015
rect 13829 4981 13863 5015
rect 14473 4981 14507 5015
rect 16221 4981 16255 5015
rect 10517 4777 10551 4811
rect 11437 4777 11471 4811
rect 12633 4777 12667 4811
rect 13185 4777 13219 4811
rect 13553 4777 13587 4811
rect 14197 4777 14231 4811
rect 14565 4777 14599 4811
rect 15301 4777 15335 4811
rect 15669 4777 15703 4811
rect 7656 4709 7690 4743
rect 10425 4709 10459 4743
rect 10885 4709 10919 4743
rect 14657 4709 14691 4743
rect 1501 4641 1535 4675
rect 1768 4641 1802 4675
rect 3249 4641 3283 4675
rect 4077 4641 4111 4675
rect 4344 4641 4378 4675
rect 5989 4641 6023 4675
rect 8861 4641 8895 4675
rect 9689 4641 9723 4675
rect 3525 4573 3559 4607
rect 5733 4573 5767 4607
rect 7389 4573 7423 4607
rect 9045 4573 9079 4607
rect 10701 4573 10735 4607
rect 9873 4505 9907 4539
rect 11529 4641 11563 4675
rect 12541 4641 12575 4675
rect 13645 4641 13679 4675
rect 11713 4573 11747 4607
rect 12817 4573 12851 4607
rect 13737 4573 13771 4607
rect 14841 4573 14875 4607
rect 15761 4573 15795 4607
rect 15853 4573 15887 4607
rect 2881 4437 2915 4471
rect 5457 4437 5491 4471
rect 7113 4437 7147 4471
rect 8769 4437 8803 4471
rect 10057 4437 10091 4471
rect 10885 4437 10919 4471
rect 11069 4437 11103 4471
rect 12173 4437 12207 4471
rect 8217 4233 8251 4267
rect 15485 4233 15519 4267
rect 5089 4165 5123 4199
rect 8493 4165 8527 4199
rect 1869 4097 1903 4131
rect 1961 4097 1995 4131
rect 2421 4097 2455 4131
rect 4537 4097 4571 4131
rect 4629 4097 4663 4131
rect 5641 4097 5675 4131
rect 6837 4097 6871 4131
rect 9045 4097 9079 4131
rect 10057 4097 10091 4131
rect 1777 4029 1811 4063
rect 6101 4029 6135 4063
rect 10609 4029 10643 4063
rect 10865 4029 10899 4063
rect 12449 4029 12483 4063
rect 14105 4029 14139 4063
rect 15761 4029 15795 4063
rect 2688 3961 2722 3995
rect 7082 3961 7116 3995
rect 12694 3961 12728 3995
rect 14350 3961 14384 3995
rect 16037 3961 16071 3995
rect 1409 3893 1443 3927
rect 3801 3893 3835 3927
rect 4077 3893 4111 3927
rect 4445 3893 4479 3927
rect 5457 3893 5491 3927
rect 5549 3893 5583 3927
rect 6285 3893 6319 3927
rect 8861 3893 8895 3927
rect 8953 3893 8987 3927
rect 9505 3893 9539 3927
rect 9873 3893 9907 3927
rect 9965 3893 9999 3927
rect 11989 3893 12023 3927
rect 13829 3893 13863 3927
rect 2697 3689 2731 3723
rect 2789 3689 2823 3723
rect 5457 3689 5491 3723
rect 6745 3689 6779 3723
rect 8401 3689 8435 3723
rect 8861 3689 8895 3723
rect 12725 3689 12759 3723
rect 12817 3689 12851 3723
rect 13829 3689 13863 3723
rect 4322 3621 4356 3655
rect 12173 3621 12207 3655
rect 1501 3553 1535 3587
rect 3341 3553 3375 3587
rect 6101 3553 6135 3587
rect 7113 3553 7147 3587
rect 7757 3553 7791 3587
rect 8769 3553 8803 3587
rect 10057 3553 10091 3587
rect 10149 3553 10183 3587
rect 10793 3553 10827 3587
rect 11529 3553 11563 3587
rect 14197 3553 14231 3587
rect 15301 3553 15335 3587
rect 16037 3553 16071 3587
rect 1685 3485 1719 3519
rect 2881 3485 2915 3519
rect 4077 3485 4111 3519
rect 6193 3485 6227 3519
rect 6285 3485 6319 3519
rect 7205 3485 7239 3519
rect 7389 3485 7423 3519
rect 7573 3485 7607 3519
rect 8953 3485 8987 3519
rect 10241 3485 10275 3519
rect 11621 3485 11655 3519
rect 11805 3485 11839 3519
rect 12909 3485 12943 3519
rect 14289 3485 14323 3519
rect 14473 3485 14507 3519
rect 15485 3485 15519 3519
rect 2329 3417 2363 3451
rect 7941 3417 7975 3451
rect 3525 3349 3559 3383
rect 5733 3349 5767 3383
rect 7573 3349 7607 3383
rect 9689 3349 9723 3383
rect 10977 3349 11011 3383
rect 11161 3349 11195 3383
rect 12357 3349 12391 3383
rect 16221 3349 16255 3383
rect 2237 3145 2271 3179
rect 3249 3145 3283 3179
rect 4261 3145 4295 3179
rect 7205 3145 7239 3179
rect 5457 3077 5491 3111
rect 9137 3145 9171 3179
rect 9321 3145 9355 3179
rect 11345 3145 11379 3179
rect 12449 3145 12483 3179
rect 13737 3145 13771 3179
rect 2789 3009 2823 3043
rect 3893 3009 3927 3043
rect 4905 3009 4939 3043
rect 6009 3009 6043 3043
rect 7205 3009 7239 3043
rect 7941 3009 7975 3043
rect 8769 3009 8803 3043
rect 8953 3009 8987 3043
rect 9137 3009 9171 3043
rect 9873 3009 9907 3043
rect 10885 3009 10919 3043
rect 11805 3009 11839 3043
rect 11989 3009 12023 3043
rect 13001 3009 13035 3043
rect 14197 3009 14231 3043
rect 14381 3009 14415 3043
rect 1501 2941 1535 2975
rect 3617 2941 3651 2975
rect 3709 2941 3743 2975
rect 6837 2941 6871 2975
rect 7665 2941 7699 2975
rect 7757 2941 7791 2975
rect 10701 2941 10735 2975
rect 12817 2941 12851 2975
rect 14749 2941 14783 2975
rect 15485 2941 15519 2975
rect 1777 2873 1811 2907
rect 2605 2873 2639 2907
rect 4721 2873 4755 2907
rect 5917 2873 5951 2907
rect 9781 2873 9815 2907
rect 11713 2873 11747 2907
rect 12909 2873 12943 2907
rect 15025 2873 15059 2907
rect 15761 2873 15795 2907
rect 2697 2805 2731 2839
rect 4629 2805 4663 2839
rect 5825 2805 5859 2839
rect 7297 2805 7331 2839
rect 8309 2805 8343 2839
rect 8677 2805 8711 2839
rect 9689 2805 9723 2839
rect 10333 2805 10367 2839
rect 10793 2805 10827 2839
rect 14105 2805 14139 2839
rect 2973 2601 3007 2635
rect 4445 2601 4479 2635
rect 4813 2601 4847 2635
rect 5917 2601 5951 2635
rect 6929 2601 6963 2635
rect 7113 2601 7147 2635
rect 7481 2601 7515 2635
rect 9781 2601 9815 2635
rect 10241 2601 10275 2635
rect 10793 2601 10827 2635
rect 11161 2601 11195 2635
rect 12633 2601 12667 2635
rect 13093 2601 13127 2635
rect 4905 2533 4939 2567
rect 5825 2533 5859 2567
rect 1501 2465 1535 2499
rect 2237 2465 2271 2499
rect 3341 2465 3375 2499
rect 3433 2465 3467 2499
rect 7573 2533 7607 2567
rect 8585 2533 8619 2567
rect 11253 2533 11287 2567
rect 14657 2533 14691 2567
rect 8493 2465 8527 2499
rect 9137 2465 9171 2499
rect 10149 2465 10183 2499
rect 11805 2465 11839 2499
rect 13001 2465 13035 2499
rect 13645 2465 13679 2499
rect 14381 2465 14415 2499
rect 15485 2465 15519 2499
rect 1685 2397 1719 2431
rect 2513 2397 2547 2431
rect 3525 2397 3559 2431
rect 5089 2397 5123 2431
rect 6009 2397 6043 2431
rect 6929 2397 6963 2431
rect 7757 2397 7791 2431
rect 8769 2397 8803 2431
rect 10333 2397 10367 2431
rect 11345 2397 11379 2431
rect 11989 2397 12023 2431
rect 13185 2397 13219 2431
rect 13829 2397 13863 2431
rect 15669 2397 15703 2431
rect 5457 2329 5491 2363
rect 8125 2329 8159 2363
rect 9321 2261 9355 2295
<< metal1 >>
rect 4062 15172 4068 15224
rect 4120 15212 4126 15224
rect 9950 15212 9956 15224
rect 4120 15184 9956 15212
rect 4120 15172 4126 15184
rect 9950 15172 9956 15184
rect 10008 15172 10014 15224
rect 2222 14968 2228 15020
rect 2280 15008 2286 15020
rect 6546 15008 6552 15020
rect 2280 14980 6552 15008
rect 2280 14968 2286 14980
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 9398 14968 9404 15020
rect 9456 15008 9462 15020
rect 15102 15008 15108 15020
rect 9456 14980 15108 15008
rect 9456 14968 9462 14980
rect 15102 14968 15108 14980
rect 15160 14968 15166 15020
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 10134 14940 10140 14952
rect 4120 14912 10140 14940
rect 4120 14900 4126 14912
rect 10134 14900 10140 14912
rect 10192 14900 10198 14952
rect 4154 14832 4160 14884
rect 4212 14872 4218 14884
rect 14642 14872 14648 14884
rect 4212 14844 14648 14872
rect 4212 14832 4218 14844
rect 14642 14832 14648 14844
rect 14700 14832 14706 14884
rect 3510 14764 3516 14816
rect 3568 14804 3574 14816
rect 9490 14804 9496 14816
rect 3568 14776 9496 14804
rect 3568 14764 3574 14776
rect 9490 14764 9496 14776
rect 9548 14764 9554 14816
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 14090 14804 14096 14816
rect 12860 14776 14096 14804
rect 12860 14764 12866 14776
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 1104 14714 16836 14736
rect 1104 14662 6246 14714
rect 6298 14662 6310 14714
rect 6362 14662 6374 14714
rect 6426 14662 6438 14714
rect 6490 14662 11510 14714
rect 11562 14662 11574 14714
rect 11626 14662 11638 14714
rect 11690 14662 11702 14714
rect 11754 14662 16836 14714
rect 1104 14640 16836 14662
rect 4154 14600 4160 14612
rect 4115 14572 4160 14600
rect 4154 14560 4160 14572
rect 4212 14560 4218 14612
rect 7377 14603 7435 14609
rect 7377 14569 7389 14603
rect 7423 14600 7435 14603
rect 8294 14600 8300 14612
rect 7423 14572 8300 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 10686 14600 10692 14612
rect 10599 14572 10692 14600
rect 10686 14560 10692 14572
rect 10744 14600 10750 14612
rect 11701 14603 11759 14609
rect 11701 14600 11713 14603
rect 10744 14572 11713 14600
rect 10744 14560 10750 14572
rect 11701 14569 11713 14572
rect 11747 14569 11759 14603
rect 11701 14563 11759 14569
rect 12989 14603 13047 14609
rect 12989 14569 13001 14603
rect 13035 14600 13047 14603
rect 13633 14603 13691 14609
rect 13633 14600 13645 14603
rect 13035 14572 13645 14600
rect 13035 14569 13047 14572
rect 12989 14563 13047 14569
rect 13633 14569 13645 14572
rect 13679 14569 13691 14603
rect 13633 14563 13691 14569
rect 13722 14560 13728 14612
rect 13780 14600 13786 14612
rect 15841 14603 15899 14609
rect 15841 14600 15853 14603
rect 13780 14572 15853 14600
rect 13780 14560 13786 14572
rect 15841 14569 15853 14572
rect 15887 14569 15899 14603
rect 15841 14563 15899 14569
rect 1394 14492 1400 14544
rect 1452 14532 1458 14544
rect 2501 14535 2559 14541
rect 2501 14532 2513 14535
rect 1452 14504 2513 14532
rect 1452 14492 1458 14504
rect 2501 14501 2513 14504
rect 2547 14532 2559 14535
rect 13354 14532 13360 14544
rect 2547 14504 13360 14532
rect 2547 14501 2559 14504
rect 2501 14495 2559 14501
rect 13004 14476 13032 14504
rect 13354 14492 13360 14504
rect 13412 14492 13418 14544
rect 14921 14535 14979 14541
rect 14921 14501 14933 14535
rect 14967 14532 14979 14535
rect 15746 14532 15752 14544
rect 14967 14504 15752 14532
rect 14967 14501 14979 14504
rect 14921 14495 14979 14501
rect 15746 14492 15752 14504
rect 15804 14492 15810 14544
rect 2406 14464 2412 14476
rect 2367 14436 2412 14464
rect 2406 14424 2412 14436
rect 2464 14424 2470 14476
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 4525 14467 4583 14473
rect 4525 14464 4537 14467
rect 4212 14436 4537 14464
rect 4212 14424 4218 14436
rect 4525 14433 4537 14436
rect 4571 14433 4583 14467
rect 5534 14464 5540 14476
rect 5495 14436 5540 14464
rect 4525 14427 4583 14433
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 6086 14464 6092 14476
rect 5675 14436 6092 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 7285 14467 7343 14473
rect 7285 14433 7297 14467
rect 7331 14464 7343 14467
rect 8570 14464 8576 14476
rect 7331 14436 8576 14464
rect 7331 14433 7343 14436
rect 7285 14427 7343 14433
rect 8570 14424 8576 14436
rect 8628 14424 8634 14476
rect 8662 14424 8668 14476
rect 8720 14464 8726 14476
rect 9033 14467 9091 14473
rect 9033 14464 9045 14467
rect 8720 14436 9045 14464
rect 8720 14424 8726 14436
rect 9033 14433 9045 14436
rect 9079 14433 9091 14467
rect 9033 14427 9091 14433
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 9674 14464 9680 14476
rect 9171 14436 9680 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14464 10655 14467
rect 11609 14467 11667 14473
rect 11609 14464 11621 14467
rect 10643 14436 11621 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 11609 14433 11621 14436
rect 11655 14464 11667 14467
rect 12158 14464 12164 14476
rect 11655 14436 12164 14464
rect 11655 14433 11667 14436
rect 11609 14427 11667 14433
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 12986 14424 12992 14476
rect 13044 14424 13050 14476
rect 13998 14464 14004 14476
rect 13959 14436 14004 14464
rect 13998 14424 14004 14436
rect 14056 14424 14062 14476
rect 14090 14424 14096 14476
rect 14148 14464 14154 14476
rect 14642 14464 14648 14476
rect 14148 14436 14193 14464
rect 14603 14436 14648 14464
rect 14148 14424 14154 14436
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 2590 14396 2596 14408
rect 2551 14368 2596 14396
rect 2590 14356 2596 14368
rect 2648 14356 2654 14408
rect 4614 14396 4620 14408
rect 4575 14368 4620 14396
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14365 4767 14399
rect 5718 14396 5724 14408
rect 5679 14368 5724 14396
rect 4709 14359 4767 14365
rect 4338 14288 4344 14340
rect 4396 14328 4402 14340
rect 4724 14328 4752 14359
rect 5718 14356 5724 14368
rect 5776 14356 5782 14408
rect 7098 14356 7104 14408
rect 7156 14396 7162 14408
rect 7469 14399 7527 14405
rect 7469 14396 7481 14399
rect 7156 14368 7481 14396
rect 7156 14356 7162 14368
rect 7469 14365 7481 14368
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 6638 14328 6644 14340
rect 4396 14300 4752 14328
rect 4816 14300 6644 14328
rect 4396 14288 4402 14300
rect 2041 14263 2099 14269
rect 2041 14229 2053 14263
rect 2087 14260 2099 14263
rect 3418 14260 3424 14272
rect 2087 14232 3424 14260
rect 2087 14229 2099 14232
rect 2041 14223 2099 14229
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 4816 14260 4844 14300
rect 6638 14288 6644 14300
rect 6696 14288 6702 14340
rect 7484 14328 7512 14359
rect 8754 14356 8760 14408
rect 8812 14396 8818 14408
rect 9217 14399 9275 14405
rect 9217 14396 9229 14399
rect 8812 14368 9229 14396
rect 8812 14356 8818 14368
rect 9217 14365 9229 14368
rect 9263 14365 9275 14399
rect 9217 14359 9275 14365
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 11793 14399 11851 14405
rect 10836 14368 10881 14396
rect 10836 14356 10842 14368
rect 11793 14365 11805 14399
rect 11839 14365 11851 14399
rect 13078 14396 13084 14408
rect 13039 14368 13084 14396
rect 11793 14359 11851 14365
rect 11808 14328 11836 14359
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 13265 14399 13323 14405
rect 13265 14365 13277 14399
rect 13311 14396 13323 14399
rect 13814 14396 13820 14408
rect 13311 14368 13820 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 7484 14300 11836 14328
rect 11974 14288 11980 14340
rect 12032 14328 12038 14340
rect 13280 14328 13308 14359
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 14185 14399 14243 14405
rect 14185 14365 14197 14399
rect 14231 14365 14243 14399
rect 14185 14359 14243 14365
rect 12032 14300 13308 14328
rect 12032 14288 12038 14300
rect 13630 14288 13636 14340
rect 13688 14328 13694 14340
rect 14200 14328 14228 14359
rect 15378 14356 15384 14408
rect 15436 14396 15442 14408
rect 15933 14399 15991 14405
rect 15933 14396 15945 14399
rect 15436 14368 15945 14396
rect 15436 14356 15442 14368
rect 15933 14365 15945 14368
rect 15979 14365 15991 14399
rect 16114 14396 16120 14408
rect 16075 14368 16120 14396
rect 15933 14359 15991 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 13688 14300 14228 14328
rect 13688 14288 13694 14300
rect 4120 14232 4844 14260
rect 4120 14220 4126 14232
rect 4982 14220 4988 14272
rect 5040 14260 5046 14272
rect 5169 14263 5227 14269
rect 5169 14260 5181 14263
rect 5040 14232 5181 14260
rect 5040 14220 5046 14232
rect 5169 14229 5181 14232
rect 5215 14229 5227 14263
rect 5169 14223 5227 14229
rect 6917 14263 6975 14269
rect 6917 14229 6929 14263
rect 6963 14260 6975 14263
rect 7374 14260 7380 14272
rect 6963 14232 7380 14260
rect 6963 14229 6975 14232
rect 6917 14223 6975 14229
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 8386 14220 8392 14272
rect 8444 14260 8450 14272
rect 8665 14263 8723 14269
rect 8665 14260 8677 14263
rect 8444 14232 8677 14260
rect 8444 14220 8450 14232
rect 8665 14229 8677 14232
rect 8711 14229 8723 14263
rect 8665 14223 8723 14229
rect 10042 14220 10048 14272
rect 10100 14260 10106 14272
rect 10229 14263 10287 14269
rect 10229 14260 10241 14263
rect 10100 14232 10241 14260
rect 10100 14220 10106 14232
rect 10229 14229 10241 14232
rect 10275 14229 10287 14263
rect 10229 14223 10287 14229
rect 11054 14220 11060 14272
rect 11112 14260 11118 14272
rect 11241 14263 11299 14269
rect 11241 14260 11253 14263
rect 11112 14232 11253 14260
rect 11112 14220 11118 14232
rect 11241 14229 11253 14232
rect 11287 14229 11299 14263
rect 12618 14260 12624 14272
rect 12579 14232 12624 14260
rect 11241 14223 11299 14229
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 15470 14260 15476 14272
rect 15431 14232 15476 14260
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 1104 14170 16836 14192
rect 1104 14118 3614 14170
rect 3666 14118 3678 14170
rect 3730 14118 3742 14170
rect 3794 14118 3806 14170
rect 3858 14118 8878 14170
rect 8930 14118 8942 14170
rect 8994 14118 9006 14170
rect 9058 14118 9070 14170
rect 9122 14118 14142 14170
rect 14194 14118 14206 14170
rect 14258 14118 14270 14170
rect 14322 14118 14334 14170
rect 14386 14118 16836 14170
rect 1104 14096 16836 14118
rect 4154 14056 4160 14068
rect 4115 14028 4160 14056
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 4246 14016 4252 14068
rect 4304 14056 4310 14068
rect 5718 14056 5724 14068
rect 4304 14028 5724 14056
rect 4304 14016 4310 14028
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 8205 14059 8263 14065
rect 8205 14056 8217 14059
rect 5920 14028 8217 14056
rect 2041 13991 2099 13997
rect 2041 13957 2053 13991
rect 2087 13988 2099 13991
rect 3053 13991 3111 13997
rect 2087 13960 2820 13988
rect 2087 13957 2099 13960
rect 2041 13951 2099 13957
rect 2590 13920 2596 13932
rect 2551 13892 2596 13920
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 2792 13920 2820 13960
rect 3053 13957 3065 13991
rect 3099 13988 3111 13991
rect 5534 13988 5540 14000
rect 3099 13960 5540 13988
rect 3099 13957 3111 13960
rect 3053 13951 3111 13957
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 3513 13923 3571 13929
rect 3513 13920 3525 13923
rect 2792 13892 3525 13920
rect 3513 13889 3525 13892
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13889 3663 13923
rect 4798 13920 4804 13932
rect 4759 13892 4804 13920
rect 3605 13883 3663 13889
rect 2498 13852 2504 13864
rect 2459 13824 2504 13852
rect 2498 13812 2504 13824
rect 2556 13812 2562 13864
rect 3142 13812 3148 13864
rect 3200 13852 3206 13864
rect 3620 13852 3648 13883
rect 4798 13880 4804 13892
rect 4856 13880 4862 13932
rect 5350 13880 5356 13932
rect 5408 13920 5414 13932
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5408 13892 5825 13920
rect 5408 13880 5414 13892
rect 5813 13889 5825 13892
rect 5859 13920 5871 13923
rect 5920 13920 5948 14028
rect 8205 14025 8217 14028
rect 8251 14025 8263 14059
rect 8662 14056 8668 14068
rect 8623 14028 8668 14056
rect 8205 14019 8263 14025
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 12802 14056 12808 14068
rect 8772 14028 12808 14056
rect 6822 13920 6828 13932
rect 5859 13892 5948 13920
rect 6783 13892 6828 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 6822 13880 6828 13892
rect 6880 13880 6886 13932
rect 8772 13920 8800 14028
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 14093 14059 14151 14065
rect 14093 14056 14105 14059
rect 13136 14028 14105 14056
rect 13136 14016 13142 14028
rect 14093 14025 14105 14028
rect 14139 14025 14151 14059
rect 15378 14056 15384 14068
rect 15339 14028 15384 14056
rect 14093 14019 14151 14025
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 9582 13948 9588 14000
rect 9640 13988 9646 14000
rect 9677 13991 9735 13997
rect 9677 13988 9689 13991
rect 9640 13960 9689 13988
rect 9640 13948 9646 13960
rect 9677 13957 9689 13960
rect 9723 13957 9735 13991
rect 9677 13951 9735 13957
rect 11333 13991 11391 13997
rect 11333 13957 11345 13991
rect 11379 13988 11391 13991
rect 12434 13988 12440 14000
rect 11379 13960 12440 13988
rect 11379 13957 11391 13960
rect 11333 13951 11391 13957
rect 12434 13948 12440 13960
rect 12492 13948 12498 14000
rect 13814 13988 13820 14000
rect 13775 13960 13820 13988
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 9306 13920 9312 13932
rect 7852 13892 8800 13920
rect 9267 13892 9312 13920
rect 7098 13861 7104 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 3200 13824 3648 13852
rect 5552 13824 5641 13852
rect 3200 13812 3206 13824
rect 3418 13784 3424 13796
rect 3379 13756 3424 13784
rect 3418 13744 3424 13756
rect 3476 13744 3482 13796
rect 4525 13787 4583 13793
rect 4525 13753 4537 13787
rect 4571 13784 4583 13787
rect 4571 13756 5212 13784
rect 4571 13753 4583 13756
rect 4525 13747 4583 13753
rect 2409 13719 2467 13725
rect 2409 13685 2421 13719
rect 2455 13716 2467 13719
rect 2682 13716 2688 13728
rect 2455 13688 2688 13716
rect 2455 13685 2467 13688
rect 2409 13679 2467 13685
rect 2682 13676 2688 13688
rect 2740 13676 2746 13728
rect 4614 13716 4620 13728
rect 4575 13688 4620 13716
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 5184 13725 5212 13756
rect 5258 13744 5264 13796
rect 5316 13784 5322 13796
rect 5552 13784 5580 13824
rect 5629 13821 5641 13824
rect 5675 13852 5687 13855
rect 7092 13852 7104 13861
rect 5675 13824 6960 13852
rect 7059 13824 7104 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 5316 13756 5580 13784
rect 6932 13784 6960 13824
rect 7092 13815 7104 13824
rect 7098 13812 7104 13815
rect 7156 13812 7162 13864
rect 7852 13852 7880 13892
rect 9306 13880 9312 13892
rect 9364 13880 9370 13932
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 10321 13923 10379 13929
rect 10321 13920 10333 13923
rect 9916 13892 10333 13920
rect 9916 13880 9922 13892
rect 10321 13889 10333 13892
rect 10367 13920 10379 13923
rect 10778 13920 10784 13932
rect 10367 13892 10784 13920
rect 10367 13889 10379 13892
rect 10321 13883 10379 13889
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 11974 13920 11980 13932
rect 11935 13892 11980 13920
rect 11974 13880 11980 13892
rect 12032 13880 12038 13932
rect 13630 13880 13636 13932
rect 13688 13920 13694 13932
rect 14645 13923 14703 13929
rect 14645 13920 14657 13923
rect 13688 13892 14657 13920
rect 13688 13880 13694 13892
rect 14645 13889 14657 13892
rect 14691 13889 14703 13923
rect 15930 13920 15936 13932
rect 15891 13892 15936 13920
rect 14645 13883 14703 13889
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 7668 13824 7880 13852
rect 7668 13784 7696 13824
rect 8662 13812 8668 13864
rect 8720 13852 8726 13864
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 8720 13824 9137 13852
rect 8720 13812 8726 13824
rect 9125 13821 9137 13824
rect 9171 13852 9183 13855
rect 9398 13852 9404 13864
rect 9171 13824 9404 13852
rect 9171 13821 9183 13824
rect 9125 13815 9183 13821
rect 9398 13812 9404 13824
rect 9456 13812 9462 13864
rect 11624 13824 12296 13852
rect 6932 13756 7696 13784
rect 9033 13787 9091 13793
rect 5316 13744 5322 13756
rect 9033 13753 9045 13787
rect 9079 13784 9091 13787
rect 9214 13784 9220 13796
rect 9079 13756 9220 13784
rect 9079 13753 9091 13756
rect 9033 13747 9091 13753
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 10873 13787 10931 13793
rect 10873 13753 10885 13787
rect 10919 13784 10931 13787
rect 11624 13784 11652 13824
rect 10919 13756 11652 13784
rect 11701 13787 11759 13793
rect 10919 13753 10931 13756
rect 10873 13747 10931 13753
rect 11701 13753 11713 13787
rect 11747 13784 11759 13787
rect 12268 13784 12296 13824
rect 12342 13812 12348 13864
rect 12400 13852 12406 13864
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12400 13824 12449 13852
rect 12400 13812 12406 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 12544 13824 12848 13852
rect 12544 13784 12572 13824
rect 12710 13793 12716 13796
rect 12704 13784 12716 13793
rect 11747 13756 12204 13784
rect 12268 13756 12572 13784
rect 12671 13756 12716 13784
rect 11747 13753 11759 13756
rect 11701 13747 11759 13753
rect 5169 13719 5227 13725
rect 5169 13685 5181 13719
rect 5215 13685 5227 13719
rect 5169 13679 5227 13685
rect 5537 13719 5595 13725
rect 5537 13685 5549 13719
rect 5583 13716 5595 13719
rect 6181 13719 6239 13725
rect 6181 13716 6193 13719
rect 5583 13688 6193 13716
rect 5583 13685 5595 13688
rect 5537 13679 5595 13685
rect 6181 13685 6193 13688
rect 6227 13685 6239 13719
rect 6181 13679 6239 13685
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 10045 13719 10103 13725
rect 10045 13716 10057 13719
rect 9824 13688 10057 13716
rect 9824 13676 9830 13688
rect 10045 13685 10057 13688
rect 10091 13685 10103 13719
rect 10045 13679 10103 13685
rect 10137 13719 10195 13725
rect 10137 13685 10149 13719
rect 10183 13716 10195 13719
rect 10594 13716 10600 13728
rect 10183 13688 10600 13716
rect 10183 13685 10195 13688
rect 10137 13679 10195 13685
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 11793 13719 11851 13725
rect 11793 13685 11805 13719
rect 11839 13716 11851 13719
rect 11882 13716 11888 13728
rect 11839 13688 11888 13716
rect 11839 13685 11851 13688
rect 11793 13679 11851 13685
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 12176 13716 12204 13756
rect 12704 13747 12716 13756
rect 12710 13744 12716 13747
rect 12768 13744 12774 13796
rect 12820 13784 12848 13824
rect 13262 13812 13268 13864
rect 13320 13852 13326 13864
rect 14553 13855 14611 13861
rect 13320 13824 14136 13852
rect 13320 13812 13326 13824
rect 13998 13784 14004 13796
rect 12820 13756 14004 13784
rect 13998 13744 14004 13756
rect 14056 13744 14062 13796
rect 14108 13784 14136 13824
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 14734 13852 14740 13864
rect 14599 13824 14740 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15841 13787 15899 13793
rect 15841 13784 15853 13787
rect 14108 13756 15853 13784
rect 15841 13753 15853 13756
rect 15887 13753 15899 13787
rect 15841 13747 15899 13753
rect 13446 13716 13452 13728
rect 12176 13688 13452 13716
rect 13446 13676 13452 13688
rect 13504 13676 13510 13728
rect 13538 13676 13544 13728
rect 13596 13716 13602 13728
rect 14461 13719 14519 13725
rect 14461 13716 14473 13719
rect 13596 13688 14473 13716
rect 13596 13676 13602 13688
rect 14461 13685 14473 13688
rect 14507 13685 14519 13719
rect 14461 13679 14519 13685
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 15749 13719 15807 13725
rect 15749 13716 15761 13719
rect 15712 13688 15761 13716
rect 15712 13676 15718 13688
rect 15749 13685 15761 13688
rect 15795 13685 15807 13719
rect 15749 13679 15807 13685
rect 1104 13626 16836 13648
rect 1104 13574 6246 13626
rect 6298 13574 6310 13626
rect 6362 13574 6374 13626
rect 6426 13574 6438 13626
rect 6490 13574 11510 13626
rect 11562 13574 11574 13626
rect 11626 13574 11638 13626
rect 11690 13574 11702 13626
rect 11754 13574 16836 13626
rect 1104 13552 16836 13574
rect 2599 13484 3924 13512
rect 2599 13453 2627 13484
rect 2584 13447 2642 13453
rect 2584 13413 2596 13447
rect 2630 13413 2642 13447
rect 2584 13407 2642 13413
rect 2682 13404 2688 13456
rect 2740 13444 2746 13456
rect 2740 13416 3823 13444
rect 2740 13404 2746 13416
rect 2317 13379 2375 13385
rect 2317 13345 2329 13379
rect 2363 13376 2375 13379
rect 2958 13376 2964 13388
rect 2363 13348 2964 13376
rect 2363 13345 2375 13348
rect 2317 13339 2375 13345
rect 2958 13336 2964 13348
rect 3016 13336 3022 13388
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 3697 13175 3755 13181
rect 3697 13172 3709 13175
rect 3568 13144 3709 13172
rect 3568 13132 3574 13144
rect 3697 13141 3709 13144
rect 3743 13141 3755 13175
rect 3795 13172 3823 13416
rect 3896 13376 3924 13484
rect 4614 13472 4620 13524
rect 4672 13512 4678 13524
rect 4709 13515 4767 13521
rect 4709 13512 4721 13515
rect 4672 13484 4721 13512
rect 4672 13472 4678 13484
rect 4709 13481 4721 13484
rect 4755 13481 4767 13515
rect 7098 13512 7104 13524
rect 4709 13475 4767 13481
rect 5092 13484 6960 13512
rect 7011 13484 7104 13512
rect 3970 13404 3976 13456
rect 4028 13444 4034 13456
rect 5092 13453 5120 13484
rect 5077 13447 5135 13453
rect 5077 13444 5089 13447
rect 4028 13416 5089 13444
rect 4028 13404 4034 13416
rect 5077 13413 5089 13416
rect 5123 13413 5135 13447
rect 5077 13407 5135 13413
rect 5988 13447 6046 13453
rect 5988 13413 6000 13447
rect 6034 13444 6046 13447
rect 6730 13444 6736 13456
rect 6034 13416 6736 13444
rect 6034 13413 6046 13416
rect 5988 13407 6046 13413
rect 6730 13404 6736 13416
rect 6788 13404 6794 13456
rect 6932 13444 6960 13484
rect 7098 13472 7104 13484
rect 7156 13512 7162 13524
rect 7282 13512 7288 13524
rect 7156 13484 7288 13512
rect 7156 13472 7162 13484
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7929 13515 7987 13521
rect 7929 13481 7941 13515
rect 7975 13512 7987 13515
rect 8386 13512 8392 13524
rect 7975 13484 8392 13512
rect 7975 13481 7987 13484
rect 7929 13475 7987 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 9674 13512 9680 13524
rect 9635 13484 9680 13512
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 10008 13484 10057 13512
rect 10008 13472 10014 13484
rect 10045 13481 10057 13484
rect 10091 13481 10103 13515
rect 10045 13475 10103 13481
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 10502 13512 10508 13524
rect 10183 13484 10508 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 12434 13472 12440 13524
rect 12492 13472 12498 13524
rect 12618 13472 12624 13524
rect 12676 13512 12682 13524
rect 13265 13515 13323 13521
rect 13265 13512 13277 13515
rect 12676 13484 13277 13512
rect 12676 13472 12682 13484
rect 13265 13481 13277 13484
rect 13311 13481 13323 13515
rect 13265 13475 13323 13481
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 13909 13515 13967 13521
rect 13909 13512 13921 13515
rect 13504 13484 13921 13512
rect 13504 13472 13510 13484
rect 13909 13481 13921 13484
rect 13955 13481 13967 13515
rect 13909 13475 13967 13481
rect 14458 13472 14464 13524
rect 14516 13512 14522 13524
rect 15010 13512 15016 13524
rect 14516 13484 15016 13512
rect 14516 13472 14522 13484
rect 15010 13472 15016 13484
rect 15068 13512 15074 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15068 13484 16037 13512
rect 15068 13472 15074 13484
rect 16025 13481 16037 13484
rect 16071 13481 16083 13515
rect 16025 13475 16083 13481
rect 7834 13444 7840 13456
rect 6932 13416 7840 13444
rect 7834 13404 7840 13416
rect 7892 13404 7898 13456
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 9033 13447 9091 13453
rect 9033 13444 9045 13447
rect 8352 13416 9045 13444
rect 8352 13404 8358 13416
rect 9033 13413 9045 13416
rect 9079 13444 9091 13447
rect 11508 13447 11566 13453
rect 9079 13416 11468 13444
rect 9079 13413 9091 13416
rect 9033 13407 9091 13413
rect 3896 13348 5396 13376
rect 3988 13320 4016 13348
rect 5368 13320 5396 13348
rect 5810 13336 5816 13388
rect 5868 13376 5874 13388
rect 8021 13379 8079 13385
rect 8021 13376 8033 13379
rect 5868 13348 8033 13376
rect 5868 13336 5874 13348
rect 8021 13345 8033 13348
rect 8067 13345 8079 13379
rect 8021 13339 8079 13345
rect 8570 13336 8576 13388
rect 8628 13376 8634 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8628 13348 8953 13376
rect 8628 13336 8634 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 9490 13336 9496 13388
rect 9548 13376 9554 13388
rect 10689 13379 10747 13385
rect 10689 13376 10701 13379
rect 9548 13348 9996 13376
rect 9548 13336 9554 13348
rect 3970 13268 3976 13320
rect 4028 13268 4034 13320
rect 5166 13308 5172 13320
rect 5127 13280 5172 13308
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 5350 13308 5356 13320
rect 5311 13280 5356 13308
rect 5350 13268 5356 13280
rect 5408 13268 5414 13320
rect 5626 13268 5632 13320
rect 5684 13308 5690 13320
rect 5721 13311 5779 13317
rect 5721 13308 5733 13311
rect 5684 13280 5733 13308
rect 5684 13268 5690 13280
rect 5721 13277 5733 13280
rect 5767 13277 5779 13311
rect 8202 13308 8208 13320
rect 8163 13280 8208 13308
rect 5721 13271 5779 13277
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 9674 13308 9680 13320
rect 9263 13280 9680 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 9674 13268 9680 13280
rect 9732 13308 9738 13320
rect 9858 13308 9864 13320
rect 9732 13280 9864 13308
rect 9732 13268 9738 13280
rect 9858 13268 9864 13280
rect 9916 13268 9922 13320
rect 9968 13308 9996 13348
rect 10152 13348 10701 13376
rect 10152 13308 10180 13348
rect 10689 13345 10701 13348
rect 10735 13345 10747 13379
rect 11440 13376 11468 13416
rect 11508 13413 11520 13447
rect 11554 13444 11566 13447
rect 11974 13444 11980 13456
rect 11554 13416 11980 13444
rect 11554 13413 11566 13416
rect 11508 13407 11566 13413
rect 11974 13404 11980 13416
rect 12032 13404 12038 13456
rect 12452 13444 12480 13472
rect 13357 13447 13415 13453
rect 13357 13444 13369 13447
rect 12452 13416 13369 13444
rect 13357 13413 13369 13416
rect 13403 13413 13415 13447
rect 13357 13407 13415 13413
rect 12250 13376 12256 13388
rect 11440 13348 12256 13376
rect 10689 13339 10747 13345
rect 12250 13336 12256 13348
rect 12308 13336 12314 13388
rect 12342 13336 12348 13388
rect 12400 13376 12406 13388
rect 12434 13376 12440 13388
rect 12400 13348 12440 13376
rect 12400 13336 12406 13348
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 14277 13379 14335 13385
rect 12676 13348 13584 13376
rect 12676 13336 12682 13348
rect 10318 13308 10324 13320
rect 9968 13280 10180 13308
rect 10279 13280 10324 13308
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 11238 13308 11244 13320
rect 11199 13280 11244 13308
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 13449 13311 13507 13317
rect 13449 13308 13461 13311
rect 12636 13280 13461 13308
rect 11146 13240 11152 13252
rect 6656 13212 11152 13240
rect 6656 13172 6684 13212
rect 11146 13200 11152 13212
rect 11204 13200 11210 13252
rect 12636 13249 12664 13280
rect 13449 13277 13461 13280
rect 13495 13277 13507 13311
rect 13556 13308 13584 13348
rect 14277 13345 14289 13379
rect 14323 13376 14335 13379
rect 15010 13376 15016 13388
rect 14323 13348 15016 13376
rect 14323 13345 14335 13348
rect 14277 13339 14335 13345
rect 15010 13336 15016 13348
rect 15068 13336 15074 13388
rect 15194 13336 15200 13388
rect 15252 13376 15258 13388
rect 15933 13379 15991 13385
rect 15933 13376 15945 13379
rect 15252 13348 15945 13376
rect 15252 13336 15258 13348
rect 15933 13345 15945 13348
rect 15979 13345 15991 13379
rect 15933 13339 15991 13345
rect 14369 13311 14427 13317
rect 14369 13308 14381 13311
rect 13556 13280 14381 13308
rect 13449 13271 13507 13277
rect 14369 13277 14381 13280
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 14461 13311 14519 13317
rect 14461 13277 14473 13311
rect 14507 13277 14519 13311
rect 16114 13308 16120 13320
rect 16075 13280 16120 13308
rect 14461 13271 14519 13277
rect 12621 13243 12679 13249
rect 12621 13209 12633 13243
rect 12667 13209 12679 13243
rect 12621 13203 12679 13209
rect 3795 13144 6684 13172
rect 3697 13135 3755 13141
rect 7098 13132 7104 13184
rect 7156 13172 7162 13184
rect 7561 13175 7619 13181
rect 7561 13172 7573 13175
rect 7156 13144 7573 13172
rect 7156 13132 7162 13144
rect 7561 13141 7573 13144
rect 7607 13141 7619 13175
rect 7561 13135 7619 13141
rect 8573 13175 8631 13181
rect 8573 13141 8585 13175
rect 8619 13172 8631 13175
rect 9398 13172 9404 13184
rect 8619 13144 9404 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 9858 13132 9864 13184
rect 9916 13172 9922 13184
rect 10134 13172 10140 13184
rect 9916 13144 10140 13172
rect 9916 13132 9922 13144
rect 10134 13132 10140 13144
rect 10192 13132 10198 13184
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10284 13144 10885 13172
rect 10284 13132 10290 13144
rect 10873 13141 10885 13144
rect 10919 13141 10931 13175
rect 10873 13135 10931 13141
rect 11422 13132 11428 13184
rect 11480 13172 11486 13184
rect 12636 13172 12664 13203
rect 12710 13200 12716 13252
rect 12768 13240 12774 13252
rect 13630 13240 13636 13252
rect 12768 13212 13636 13240
rect 12768 13200 12774 13212
rect 13630 13200 13636 13212
rect 13688 13240 13694 13252
rect 14476 13240 14504 13271
rect 16114 13268 16120 13280
rect 16172 13268 16178 13320
rect 13688 13212 14504 13240
rect 13688 13200 13694 13212
rect 12894 13172 12900 13184
rect 11480 13144 12664 13172
rect 12855 13144 12900 13172
rect 11480 13132 11486 13144
rect 12894 13132 12900 13144
rect 12952 13132 12958 13184
rect 15562 13172 15568 13184
rect 15523 13144 15568 13172
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 1104 13082 16836 13104
rect 1104 13030 3614 13082
rect 3666 13030 3678 13082
rect 3730 13030 3742 13082
rect 3794 13030 3806 13082
rect 3858 13030 8878 13082
rect 8930 13030 8942 13082
rect 8994 13030 9006 13082
rect 9058 13030 9070 13082
rect 9122 13030 14142 13082
rect 14194 13030 14206 13082
rect 14258 13030 14270 13082
rect 14322 13030 14334 13082
rect 14386 13030 16836 13082
rect 1104 13008 16836 13030
rect 4338 12968 4344 12980
rect 4299 12940 4344 12968
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 4706 12968 4712 12980
rect 4667 12940 4712 12968
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 4890 12928 4896 12980
rect 4948 12968 4954 12980
rect 5721 12971 5779 12977
rect 4948 12940 5396 12968
rect 4948 12928 4954 12940
rect 2590 12832 2596 12844
rect 2551 12804 2596 12832
rect 2590 12792 2596 12804
rect 2648 12792 2654 12844
rect 2958 12832 2964 12844
rect 2919 12804 2964 12832
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 4798 12832 4804 12844
rect 4264 12804 4804 12832
rect 2314 12764 2320 12776
rect 2275 12736 2320 12764
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 3228 12767 3286 12773
rect 3228 12733 3240 12767
rect 3274 12764 3286 12767
rect 3510 12764 3516 12776
rect 3274 12736 3516 12764
rect 3274 12733 3286 12736
rect 3228 12727 3286 12733
rect 3510 12724 3516 12736
rect 3568 12764 3574 12776
rect 4264 12764 4292 12804
rect 4798 12792 4804 12804
rect 4856 12832 4862 12844
rect 5261 12835 5319 12841
rect 5261 12832 5273 12835
rect 4856 12804 5273 12832
rect 4856 12792 4862 12804
rect 5261 12801 5273 12804
rect 5307 12801 5319 12835
rect 5261 12795 5319 12801
rect 3568 12736 4292 12764
rect 5169 12767 5227 12773
rect 3568 12724 3574 12736
rect 5169 12733 5181 12767
rect 5215 12764 5227 12767
rect 5368 12764 5396 12940
rect 5721 12937 5733 12971
rect 5767 12968 5779 12971
rect 5810 12968 5816 12980
rect 5767 12940 5816 12968
rect 5767 12937 5779 12940
rect 5721 12931 5779 12937
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 9677 12971 9735 12977
rect 9677 12968 9689 12971
rect 6196 12940 9689 12968
rect 6196 12841 6224 12940
rect 9677 12937 9689 12940
rect 9723 12937 9735 12971
rect 9677 12931 9735 12937
rect 11333 12971 11391 12977
rect 11333 12937 11345 12971
rect 11379 12968 11391 12971
rect 11882 12968 11888 12980
rect 11379 12940 11888 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 14550 12968 14556 12980
rect 12452 12940 14556 12968
rect 8754 12900 8760 12912
rect 8715 12872 8760 12900
rect 8754 12860 8760 12872
rect 8812 12860 8818 12912
rect 9858 12860 9864 12912
rect 9916 12900 9922 12912
rect 10965 12903 11023 12909
rect 9916 12872 10824 12900
rect 9916 12860 9922 12872
rect 6181 12835 6239 12841
rect 6181 12801 6193 12835
rect 6227 12801 6239 12835
rect 6181 12795 6239 12801
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 5215 12736 5396 12764
rect 6380 12764 6408 12795
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6972 12804 7389 12832
rect 6972 12792 6978 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 7466 12764 7472 12776
rect 6380 12736 7472 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 7466 12724 7472 12736
rect 7524 12764 7530 12776
rect 8772 12764 8800 12860
rect 9214 12832 9220 12844
rect 9175 12804 9220 12832
rect 9214 12792 9220 12804
rect 9272 12792 9278 12844
rect 9398 12792 9404 12844
rect 9456 12832 9462 12844
rect 10137 12835 10195 12841
rect 10137 12832 10149 12835
rect 9456 12804 10149 12832
rect 9456 12792 9462 12804
rect 10137 12801 10149 12804
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 10229 12835 10287 12841
rect 10229 12801 10241 12835
rect 10275 12832 10287 12835
rect 10318 12832 10324 12844
rect 10275 12804 10324 12832
rect 10275 12801 10287 12804
rect 10229 12795 10287 12801
rect 10042 12764 10048 12776
rect 7524 12736 8800 12764
rect 10003 12736 10048 12764
rect 7524 12724 7530 12736
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10244 12764 10272 12795
rect 10318 12792 10324 12804
rect 10376 12792 10382 12844
rect 10796 12773 10824 12872
rect 10965 12869 10977 12903
rect 11011 12900 11023 12903
rect 12452 12900 12480 12940
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 11011 12872 12480 12900
rect 11011 12869 11023 12872
rect 10965 12863 11023 12869
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 12584 12872 13032 12900
rect 12584 12860 12590 12872
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12832 12035 12835
rect 12710 12832 12716 12844
rect 12023 12804 12716 12832
rect 12023 12801 12035 12804
rect 11977 12795 12035 12801
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 13004 12841 13032 12872
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 13035 12804 13124 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 13096 12776 13124 12804
rect 10152 12736 10272 12764
rect 10781 12767 10839 12773
rect 2332 12696 2360 12724
rect 3418 12696 3424 12708
rect 2332 12668 3424 12696
rect 3418 12656 3424 12668
rect 3476 12656 3482 12708
rect 4430 12656 4436 12708
rect 4488 12696 4494 12708
rect 4890 12696 4896 12708
rect 4488 12668 4896 12696
rect 4488 12656 4494 12668
rect 4890 12656 4896 12668
rect 4948 12656 4954 12708
rect 7644 12699 7702 12705
rect 7644 12665 7656 12699
rect 7690 12696 7702 12699
rect 9306 12696 9312 12708
rect 7690 12668 9312 12696
rect 7690 12665 7702 12668
rect 7644 12659 7702 12665
rect 9306 12656 9312 12668
rect 9364 12696 9370 12708
rect 10152 12696 10180 12736
rect 10781 12733 10793 12767
rect 10827 12733 10839 12767
rect 10781 12727 10839 12733
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 12342 12764 12348 12776
rect 11204 12736 12348 12764
rect 11204 12724 11210 12736
rect 12342 12724 12348 12736
rect 12400 12724 12406 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12492 12736 12537 12764
rect 12492 12724 12498 12736
rect 13078 12724 13084 12776
rect 13136 12764 13142 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 13136 12736 14933 12764
rect 13136 12724 13142 12736
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 14921 12727 14979 12733
rect 9364 12668 10180 12696
rect 11701 12699 11759 12705
rect 9364 12656 9370 12668
rect 11701 12665 11713 12699
rect 11747 12696 11759 12699
rect 12710 12696 12716 12708
rect 11747 12668 12716 12696
rect 11747 12665 11759 12668
rect 11701 12659 11759 12665
rect 12710 12656 12716 12668
rect 12768 12656 12774 12708
rect 13256 12699 13314 12705
rect 13256 12665 13268 12699
rect 13302 12696 13314 12699
rect 13354 12696 13360 12708
rect 13302 12668 13360 12696
rect 13302 12665 13314 12668
rect 13256 12659 13314 12665
rect 13354 12656 13360 12668
rect 13412 12656 13418 12708
rect 15188 12699 15246 12705
rect 15188 12665 15200 12699
rect 15234 12696 15246 12699
rect 15378 12696 15384 12708
rect 15234 12668 15384 12696
rect 15234 12665 15246 12668
rect 15188 12659 15246 12665
rect 15378 12656 15384 12668
rect 15436 12656 15442 12708
rect 1949 12631 2007 12637
rect 1949 12597 1961 12631
rect 1995 12628 2007 12631
rect 2222 12628 2228 12640
rect 1995 12600 2228 12628
rect 1995 12597 2007 12600
rect 1949 12591 2007 12597
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 2409 12631 2467 12637
rect 2409 12597 2421 12631
rect 2455 12628 2467 12631
rect 3050 12628 3056 12640
rect 2455 12600 3056 12628
rect 2455 12597 2467 12600
rect 2409 12591 2467 12597
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 5074 12588 5080 12640
rect 5132 12628 5138 12640
rect 6089 12631 6147 12637
rect 5132 12600 5177 12628
rect 5132 12588 5138 12600
rect 6089 12597 6101 12631
rect 6135 12628 6147 12631
rect 8018 12628 8024 12640
rect 6135 12600 8024 12628
rect 6135 12597 6147 12600
rect 6089 12591 6147 12597
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10778 12628 10784 12640
rect 9824 12600 10784 12628
rect 9824 12588 9830 12600
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 11793 12631 11851 12637
rect 11793 12597 11805 12631
rect 11839 12628 11851 12631
rect 12526 12628 12532 12640
rect 11839 12600 12532 12628
rect 11839 12597 11851 12600
rect 11793 12591 11851 12597
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 12621 12631 12679 12637
rect 12621 12597 12633 12631
rect 12667 12628 12679 12631
rect 13078 12628 13084 12640
rect 12667 12600 13084 12628
rect 12667 12597 12679 12600
rect 12621 12591 12679 12597
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 13630 12588 13636 12640
rect 13688 12628 13694 12640
rect 14369 12631 14427 12637
rect 14369 12628 14381 12631
rect 13688 12600 14381 12628
rect 13688 12588 13694 12600
rect 14369 12597 14381 12600
rect 14415 12597 14427 12631
rect 14369 12591 14427 12597
rect 15286 12588 15292 12640
rect 15344 12628 15350 12640
rect 16301 12631 16359 12637
rect 16301 12628 16313 12631
rect 15344 12600 16313 12628
rect 15344 12588 15350 12600
rect 16301 12597 16313 12600
rect 16347 12597 16359 12631
rect 16301 12591 16359 12597
rect 1104 12538 16836 12560
rect 1104 12486 6246 12538
rect 6298 12486 6310 12538
rect 6362 12486 6374 12538
rect 6426 12486 6438 12538
rect 6490 12486 11510 12538
rect 11562 12486 11574 12538
rect 11626 12486 11638 12538
rect 11690 12486 11702 12538
rect 11754 12486 16836 12538
rect 1104 12464 16836 12486
rect 1489 12427 1547 12433
rect 1489 12393 1501 12427
rect 1535 12424 1547 12427
rect 2406 12424 2412 12436
rect 1535 12396 2412 12424
rect 1535 12393 1547 12396
rect 1489 12387 1547 12393
rect 2406 12384 2412 12396
rect 2464 12384 2470 12436
rect 2961 12427 3019 12433
rect 2961 12393 2973 12427
rect 3007 12424 3019 12427
rect 5074 12424 5080 12436
rect 3007 12396 5080 12424
rect 3007 12393 3019 12396
rect 2961 12387 3019 12393
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 6748 12396 8156 12424
rect 6748 12368 6776 12396
rect 4338 12365 4344 12368
rect 4332 12356 4344 12365
rect 4299 12328 4344 12356
rect 4332 12319 4344 12328
rect 4338 12316 4344 12319
rect 4396 12316 4402 12368
rect 4798 12316 4804 12368
rect 4856 12356 4862 12368
rect 6641 12359 6699 12365
rect 6641 12356 6653 12359
rect 4856 12328 6653 12356
rect 4856 12316 4862 12328
rect 6641 12325 6653 12328
rect 6687 12325 6699 12359
rect 6641 12319 6699 12325
rect 6730 12316 6736 12368
rect 6788 12316 6794 12368
rect 7466 12365 7472 12368
rect 7460 12356 7472 12365
rect 7427 12328 7472 12356
rect 7460 12319 7472 12328
rect 7466 12316 7472 12319
rect 7524 12316 7530 12368
rect 8128 12356 8156 12396
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8260 12396 8585 12424
rect 8260 12384 8266 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 9766 12424 9772 12436
rect 8573 12387 8631 12393
rect 8680 12396 9772 12424
rect 8680 12356 8708 12396
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10318 12424 10324 12436
rect 10100 12396 10324 12424
rect 10100 12384 10106 12396
rect 10318 12384 10324 12396
rect 10376 12424 10382 12436
rect 11793 12427 11851 12433
rect 11793 12424 11805 12427
rect 10376 12396 11805 12424
rect 10376 12384 10382 12396
rect 11793 12393 11805 12396
rect 11839 12393 11851 12427
rect 11793 12387 11851 12393
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12713 12427 12771 12433
rect 12713 12424 12725 12427
rect 12584 12396 12725 12424
rect 12584 12384 12590 12396
rect 12713 12393 12725 12396
rect 12759 12393 12771 12427
rect 12713 12387 12771 12393
rect 12894 12384 12900 12436
rect 12952 12424 12958 12436
rect 13446 12424 13452 12436
rect 12952 12396 13452 12424
rect 12952 12384 12958 12396
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 14553 12427 14611 12433
rect 14553 12393 14565 12427
rect 14599 12424 14611 12427
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 14599 12396 15301 12424
rect 14599 12393 14611 12396
rect 14553 12387 14611 12393
rect 15289 12393 15301 12396
rect 15335 12393 15347 12427
rect 15289 12387 15347 12393
rect 15562 12384 15568 12436
rect 15620 12424 15626 12436
rect 15657 12427 15715 12433
rect 15657 12424 15669 12427
rect 15620 12396 15669 12424
rect 15620 12384 15626 12396
rect 15657 12393 15669 12396
rect 15703 12393 15715 12427
rect 15657 12387 15715 12393
rect 8128 12328 8708 12356
rect 9674 12316 9680 12368
rect 9732 12356 9738 12368
rect 10658 12359 10716 12365
rect 10658 12356 10670 12359
rect 9732 12328 10670 12356
rect 9732 12316 9738 12328
rect 10658 12325 10670 12328
rect 10704 12325 10716 12359
rect 10658 12319 10716 12325
rect 10778 12316 10784 12368
rect 10836 12356 10842 12368
rect 14918 12356 14924 12368
rect 10836 12328 14924 12356
rect 10836 12316 10842 12328
rect 14918 12316 14924 12328
rect 14976 12316 14982 12368
rect 1946 12248 1952 12300
rect 2004 12288 2010 12300
rect 2317 12291 2375 12297
rect 2317 12288 2329 12291
rect 2004 12260 2329 12288
rect 2004 12248 2010 12260
rect 2317 12257 2329 12260
rect 2363 12257 2375 12291
rect 3326 12288 3332 12300
rect 3287 12260 3332 12288
rect 2317 12251 2375 12257
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 3970 12288 3976 12300
rect 3528 12260 3976 12288
rect 2406 12220 2412 12232
rect 2367 12192 2412 12220
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 2498 12180 2504 12232
rect 2556 12220 2562 12232
rect 3528 12229 3556 12260
rect 3970 12248 3976 12260
rect 4028 12248 4034 12300
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 6549 12291 6607 12297
rect 6549 12288 6561 12291
rect 4212 12260 6561 12288
rect 4212 12248 4218 12260
rect 6549 12257 6561 12260
rect 6595 12257 6607 12291
rect 9030 12288 9036 12300
rect 8991 12260 9036 12288
rect 6549 12251 6607 12257
rect 9030 12248 9036 12260
rect 9088 12248 9094 12300
rect 9769 12291 9827 12297
rect 9769 12257 9781 12291
rect 9815 12288 9827 12291
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 9815 12260 9873 12288
rect 9815 12257 9827 12260
rect 9769 12251 9827 12257
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 10413 12291 10471 12297
rect 10413 12257 10425 12291
rect 10459 12288 10471 12291
rect 11238 12288 11244 12300
rect 10459 12260 11244 12288
rect 10459 12257 10471 12260
rect 10413 12251 10471 12257
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 11514 12248 11520 12300
rect 11572 12288 11578 12300
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 11572 12260 12173 12288
rect 11572 12248 11578 12260
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 12161 12251 12219 12257
rect 12250 12248 12256 12300
rect 12308 12288 12314 12300
rect 12621 12291 12679 12297
rect 12621 12288 12633 12291
rect 12308 12260 12633 12288
rect 12308 12248 12314 12260
rect 12621 12257 12633 12260
rect 12667 12257 12679 12291
rect 12621 12251 12679 12257
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12288 13139 12291
rect 13446 12288 13452 12300
rect 13127 12260 13452 12288
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 15286 12288 15292 12300
rect 13556 12260 15292 12288
rect 3421 12223 3479 12229
rect 3421 12220 3433 12223
rect 2556 12192 2601 12220
rect 2792 12192 3433 12220
rect 2556 12180 2562 12192
rect 2682 12112 2688 12164
rect 2740 12152 2746 12164
rect 2792 12152 2820 12192
rect 3421 12189 3433 12192
rect 3467 12189 3479 12223
rect 3421 12183 3479 12189
rect 3513 12223 3571 12229
rect 3513 12189 3525 12223
rect 3559 12189 3571 12223
rect 3513 12183 3571 12189
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12189 4123 12223
rect 4065 12183 4123 12189
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 2740 12124 2820 12152
rect 2740 12112 2746 12124
rect 2958 12112 2964 12164
rect 3016 12152 3022 12164
rect 4080 12152 4108 12183
rect 3016 12124 4108 12152
rect 6748 12152 6776 12183
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 6972 12192 7205 12220
rect 6972 12180 6978 12192
rect 7193 12189 7205 12192
rect 7239 12189 7251 12223
rect 9048 12220 9076 12248
rect 10226 12220 10232 12232
rect 9048 12192 10232 12220
rect 7193 12183 7251 12189
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12189 13231 12223
rect 13354 12220 13360 12232
rect 13267 12192 13360 12220
rect 13173 12183 13231 12189
rect 7006 12152 7012 12164
rect 6748 12124 7012 12152
rect 3016 12112 3022 12124
rect 7006 12112 7012 12124
rect 7064 12112 7070 12164
rect 9769 12155 9827 12161
rect 9769 12152 9781 12155
rect 9140 12124 9781 12152
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12084 2007 12087
rect 2038 12084 2044 12096
rect 1995 12056 2044 12084
rect 1995 12053 2007 12056
rect 1949 12047 2007 12053
rect 2038 12044 2044 12056
rect 2096 12044 2102 12096
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 5445 12087 5503 12093
rect 5445 12084 5457 12087
rect 4120 12056 5457 12084
rect 4120 12044 4126 12056
rect 5445 12053 5457 12056
rect 5491 12053 5503 12087
rect 5445 12047 5503 12053
rect 6181 12087 6239 12093
rect 6181 12053 6193 12087
rect 6227 12084 6239 12087
rect 7558 12084 7564 12096
rect 6227 12056 7564 12084
rect 6227 12053 6239 12056
rect 6181 12047 6239 12053
rect 7558 12044 7564 12056
rect 7616 12044 7622 12096
rect 7926 12044 7932 12096
rect 7984 12084 7990 12096
rect 9140 12084 9168 12124
rect 9769 12121 9781 12124
rect 9815 12121 9827 12155
rect 9769 12115 9827 12121
rect 11974 12112 11980 12164
rect 12032 12152 12038 12164
rect 12345 12155 12403 12161
rect 12345 12152 12357 12155
rect 12032 12124 12357 12152
rect 12032 12112 12038 12124
rect 12345 12121 12357 12124
rect 12391 12121 12403 12155
rect 12345 12115 12403 12121
rect 12526 12112 12532 12164
rect 12584 12152 12590 12164
rect 12621 12155 12679 12161
rect 12621 12152 12633 12155
rect 12584 12124 12633 12152
rect 12584 12112 12590 12124
rect 12621 12121 12633 12124
rect 12667 12152 12679 12155
rect 13188 12152 13216 12183
rect 13354 12180 13360 12192
rect 13412 12220 13418 12232
rect 13556 12220 13584 12260
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 13722 12220 13728 12232
rect 13412 12192 13584 12220
rect 13683 12192 13728 12220
rect 13412 12180 13418 12192
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 14642 12220 14648 12232
rect 14603 12192 14648 12220
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12220 14887 12223
rect 15378 12220 15384 12232
rect 14875 12192 15384 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 15749 12223 15807 12229
rect 15749 12189 15761 12223
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 12667 12124 13216 12152
rect 12667 12121 12679 12124
rect 12621 12115 12679 12121
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 15764 12152 15792 12183
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 15896 12192 15941 12220
rect 15896 12180 15902 12192
rect 14056 12124 15792 12152
rect 14056 12112 14062 12124
rect 7984 12056 9168 12084
rect 9217 12087 9275 12093
rect 7984 12044 7990 12056
rect 9217 12053 9229 12087
rect 9263 12084 9275 12087
rect 9306 12084 9312 12096
rect 9263 12056 9312 12084
rect 9263 12053 9275 12056
rect 9217 12047 9275 12053
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 10045 12087 10103 12093
rect 10045 12053 10057 12087
rect 10091 12084 10103 12087
rect 10778 12084 10784 12096
rect 10091 12056 10784 12084
rect 10091 12053 10103 12056
rect 10045 12047 10103 12053
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 11422 12044 11428 12096
rect 11480 12084 11486 12096
rect 13814 12084 13820 12096
rect 11480 12056 13820 12084
rect 11480 12044 11486 12056
rect 13814 12044 13820 12056
rect 13872 12044 13878 12096
rect 14185 12087 14243 12093
rect 14185 12053 14197 12087
rect 14231 12084 14243 12087
rect 14734 12084 14740 12096
rect 14231 12056 14740 12084
rect 14231 12053 14243 12056
rect 14185 12047 14243 12053
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 1104 11994 16836 12016
rect 1104 11942 3614 11994
rect 3666 11942 3678 11994
rect 3730 11942 3742 11994
rect 3794 11942 3806 11994
rect 3858 11942 8878 11994
rect 8930 11942 8942 11994
rect 8994 11942 9006 11994
rect 9058 11942 9070 11994
rect 9122 11942 14142 11994
rect 14194 11942 14206 11994
rect 14258 11942 14270 11994
rect 14322 11942 14334 11994
rect 14386 11942 16836 11994
rect 1104 11920 16836 11942
rect 2866 11840 2872 11892
rect 2924 11880 2930 11892
rect 5994 11880 6000 11892
rect 2924 11852 6000 11880
rect 2924 11840 2930 11852
rect 5994 11840 6000 11852
rect 6052 11880 6058 11892
rect 6052 11852 7420 11880
rect 6052 11840 6058 11852
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 6273 11747 6331 11753
rect 6273 11744 6285 11747
rect 5684 11716 6285 11744
rect 5684 11704 5690 11716
rect 6273 11713 6285 11716
rect 6319 11713 6331 11747
rect 7392 11744 7420 11852
rect 8018 11840 8024 11892
rect 8076 11880 8082 11892
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 8076 11852 9229 11880
rect 8076 11840 8082 11852
rect 9217 11849 9229 11852
rect 9263 11849 9275 11883
rect 9217 11843 9275 11849
rect 9674 11840 9680 11892
rect 9732 11840 9738 11892
rect 10321 11883 10379 11889
rect 10321 11849 10333 11883
rect 10367 11880 10379 11883
rect 13998 11880 14004 11892
rect 10367 11852 14004 11880
rect 10367 11849 10379 11852
rect 10321 11843 10379 11849
rect 13998 11840 14004 11852
rect 14056 11840 14062 11892
rect 14108 11852 15332 11880
rect 8757 11815 8815 11821
rect 8757 11781 8769 11815
rect 8803 11812 8815 11815
rect 9692 11812 9720 11840
rect 11333 11815 11391 11821
rect 8803 11784 9720 11812
rect 10796 11784 11284 11812
rect 8803 11781 8815 11784
rect 8757 11775 8815 11781
rect 7392 11716 7512 11744
rect 6273 11707 6331 11713
rect 1486 11636 1492 11688
rect 1544 11676 1550 11688
rect 1765 11679 1823 11685
rect 1765 11676 1777 11679
rect 1544 11648 1777 11676
rect 1544 11636 1550 11648
rect 1765 11645 1777 11648
rect 1811 11676 1823 11679
rect 2958 11676 2964 11688
rect 1811 11648 2964 11676
rect 1811 11645 1823 11648
rect 1765 11639 1823 11645
rect 2958 11636 2964 11648
rect 3016 11676 3022 11688
rect 3513 11679 3571 11685
rect 3513 11676 3525 11679
rect 3016 11648 3525 11676
rect 3016 11636 3022 11648
rect 3513 11645 3525 11648
rect 3559 11645 3571 11679
rect 3513 11639 3571 11645
rect 3602 11636 3608 11688
rect 3660 11676 3666 11688
rect 3780 11679 3838 11685
rect 3780 11676 3792 11679
rect 3660 11648 3792 11676
rect 3660 11636 3666 11648
rect 3780 11645 3792 11648
rect 3826 11676 3838 11679
rect 4062 11676 4068 11688
rect 3826 11648 4068 11676
rect 3826 11645 3838 11648
rect 3780 11639 3838 11645
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 5810 11636 5816 11688
rect 5868 11676 5874 11688
rect 6914 11676 6920 11688
rect 5868 11648 6920 11676
rect 5868 11636 5874 11648
rect 6914 11636 6920 11648
rect 6972 11676 6978 11688
rect 7377 11679 7435 11685
rect 7377 11676 7389 11679
rect 6972 11648 7389 11676
rect 6972 11636 6978 11648
rect 7377 11645 7389 11648
rect 7423 11645 7435 11679
rect 7484 11676 7512 11716
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 9677 11747 9735 11753
rect 9677 11744 9689 11747
rect 9640 11716 9689 11744
rect 9640 11704 9646 11716
rect 9677 11713 9689 11716
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 9861 11747 9919 11753
rect 9861 11713 9873 11747
rect 9907 11744 9919 11747
rect 10042 11744 10048 11756
rect 9907 11716 10048 11744
rect 9907 11713 9919 11716
rect 9861 11707 9919 11713
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 10796 11685 10824 11784
rect 10962 11744 10968 11756
rect 10923 11716 10968 11744
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11256 11744 11284 11784
rect 11333 11781 11345 11815
rect 11379 11812 11391 11815
rect 12618 11812 12624 11824
rect 11379 11784 12624 11812
rect 11379 11781 11391 11784
rect 11333 11775 11391 11781
rect 12618 11772 12624 11784
rect 12676 11772 12682 11824
rect 14108 11812 14136 11852
rect 13740 11784 14136 11812
rect 15304 11812 15332 11852
rect 15378 11840 15384 11892
rect 15436 11880 15442 11892
rect 15749 11883 15807 11889
rect 15749 11880 15761 11883
rect 15436 11852 15761 11880
rect 15436 11840 15442 11852
rect 15749 11849 15761 11852
rect 15795 11849 15807 11883
rect 15749 11843 15807 11849
rect 16114 11812 16120 11824
rect 15304 11784 16120 11812
rect 11422 11744 11428 11756
rect 11256 11716 11428 11744
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 12023 11716 12848 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 7484 11648 10793 11676
rect 7377 11639 7435 11645
rect 10781 11645 10793 11648
rect 10827 11645 10839 11679
rect 11514 11676 11520 11688
rect 10781 11639 10839 11645
rect 10888 11648 11520 11676
rect 2032 11611 2090 11617
rect 2032 11577 2044 11611
rect 2078 11608 2090 11611
rect 2498 11608 2504 11620
rect 2078 11580 2504 11608
rect 2078 11577 2090 11580
rect 2032 11571 2090 11577
rect 2498 11568 2504 11580
rect 2556 11608 2562 11620
rect 2556 11580 3740 11608
rect 2556 11568 2562 11580
rect 1670 11500 1676 11552
rect 1728 11540 1734 11552
rect 2314 11540 2320 11552
rect 1728 11512 2320 11540
rect 1728 11500 1734 11512
rect 2314 11500 2320 11512
rect 2372 11540 2378 11552
rect 2866 11540 2872 11552
rect 2372 11512 2872 11540
rect 2372 11500 2378 11512
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3142 11540 3148 11552
rect 3016 11512 3148 11540
rect 3016 11500 3022 11512
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 3712 11540 3740 11580
rect 4982 11568 4988 11620
rect 5040 11608 5046 11620
rect 5350 11608 5356 11620
rect 5040 11580 5356 11608
rect 5040 11568 5046 11580
rect 5350 11568 5356 11580
rect 5408 11568 5414 11620
rect 5902 11568 5908 11620
rect 5960 11608 5966 11620
rect 6089 11611 6147 11617
rect 6089 11608 6101 11611
rect 5960 11580 6101 11608
rect 5960 11568 5966 11580
rect 6089 11577 6101 11580
rect 6135 11577 6147 11611
rect 6089 11571 6147 11577
rect 6181 11611 6239 11617
rect 6181 11577 6193 11611
rect 6227 11608 6239 11611
rect 7282 11608 7288 11620
rect 6227 11580 7288 11608
rect 6227 11577 6239 11580
rect 6181 11571 6239 11577
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 7466 11568 7472 11620
rect 7524 11608 7530 11620
rect 7622 11611 7680 11617
rect 7622 11608 7634 11611
rect 7524 11580 7634 11608
rect 7524 11568 7530 11580
rect 7622 11577 7634 11580
rect 7668 11577 7680 11611
rect 7622 11571 7680 11577
rect 7742 11568 7748 11620
rect 7800 11608 7806 11620
rect 10689 11611 10747 11617
rect 10689 11608 10701 11611
rect 7800 11580 10701 11608
rect 7800 11568 7806 11580
rect 10689 11577 10701 11580
rect 10735 11608 10747 11611
rect 10888 11608 10916 11648
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 11698 11676 11704 11688
rect 11659 11648 11704 11676
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 12158 11636 12164 11688
rect 12216 11676 12222 11688
rect 12713 11679 12771 11685
rect 12713 11676 12725 11679
rect 12216 11648 12725 11676
rect 12216 11636 12222 11648
rect 12713 11645 12725 11648
rect 12759 11645 12771 11679
rect 12820 11676 12848 11716
rect 13354 11676 13360 11688
rect 12820 11648 13360 11676
rect 12713 11639 12771 11645
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 10735 11580 10916 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 11054 11568 11060 11620
rect 11112 11568 11118 11620
rect 12250 11568 12256 11620
rect 12308 11608 12314 11620
rect 12980 11611 13038 11617
rect 12980 11608 12992 11611
rect 12308 11580 12992 11608
rect 12308 11568 12314 11580
rect 12980 11577 12992 11580
rect 13026 11608 13038 11611
rect 13740 11608 13768 11784
rect 16114 11772 16120 11784
rect 16172 11772 16178 11824
rect 13026 11580 13768 11608
rect 13832 11716 14504 11744
rect 13026 11577 13038 11580
rect 12980 11571 13038 11577
rect 4893 11543 4951 11549
rect 4893 11540 4905 11543
rect 3712 11512 4905 11540
rect 4893 11509 4905 11512
rect 4939 11509 4951 11543
rect 5718 11540 5724 11552
rect 5679 11512 5724 11540
rect 4893 11503 4951 11509
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 6822 11540 6828 11552
rect 6696 11512 6828 11540
rect 6696 11500 6702 11512
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 6917 11543 6975 11549
rect 6917 11509 6929 11543
rect 6963 11540 6975 11543
rect 8110 11540 8116 11552
rect 6963 11512 8116 11540
rect 6963 11509 6975 11512
rect 6917 11503 6975 11509
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 9548 11512 9597 11540
rect 9548 11500 9554 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 11072 11540 11100 11568
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11072 11512 11805 11540
rect 9585 11503 9643 11509
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 11882 11500 11888 11552
rect 11940 11540 11946 11552
rect 13832 11540 13860 11716
rect 14366 11676 14372 11688
rect 14327 11648 14372 11676
rect 14366 11636 14372 11648
rect 14424 11636 14430 11688
rect 14476 11676 14504 11716
rect 15194 11676 15200 11688
rect 14476 11648 15200 11676
rect 15194 11636 15200 11648
rect 15252 11636 15258 11688
rect 16022 11676 16028 11688
rect 15983 11648 16028 11676
rect 16022 11636 16028 11648
rect 16080 11636 16086 11688
rect 14636 11611 14694 11617
rect 14636 11608 14648 11611
rect 14108 11580 14648 11608
rect 14108 11549 14136 11580
rect 14636 11577 14648 11580
rect 14682 11608 14694 11611
rect 15838 11608 15844 11620
rect 14682 11580 15844 11608
rect 14682 11577 14694 11580
rect 14636 11571 14694 11577
rect 15838 11568 15844 11580
rect 15896 11568 15902 11620
rect 11940 11512 13860 11540
rect 14093 11543 14151 11549
rect 11940 11500 11946 11512
rect 14093 11509 14105 11543
rect 14139 11509 14151 11543
rect 14093 11503 14151 11509
rect 16209 11543 16267 11549
rect 16209 11509 16221 11543
rect 16255 11540 16267 11543
rect 16390 11540 16396 11552
rect 16255 11512 16396 11540
rect 16255 11509 16267 11512
rect 16209 11503 16267 11509
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 1104 11450 16836 11472
rect 1104 11398 6246 11450
rect 6298 11398 6310 11450
rect 6362 11398 6374 11450
rect 6426 11398 6438 11450
rect 6490 11398 11510 11450
rect 11562 11398 11574 11450
rect 11626 11398 11638 11450
rect 11690 11398 11702 11450
rect 11754 11398 16836 11450
rect 1104 11376 16836 11398
rect 1946 11336 1952 11348
rect 1907 11308 1952 11336
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 2406 11296 2412 11348
rect 2464 11336 2470 11348
rect 2961 11339 3019 11345
rect 2961 11336 2973 11339
rect 2464 11308 2973 11336
rect 2464 11296 2470 11308
rect 2961 11305 2973 11308
rect 3007 11305 3019 11339
rect 4246 11336 4252 11348
rect 2961 11299 3019 11305
rect 3068 11308 4252 11336
rect 2866 11228 2872 11280
rect 2924 11268 2930 11280
rect 3068 11268 3096 11308
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 4985 11339 5043 11345
rect 4985 11305 4997 11339
rect 5031 11336 5043 11339
rect 7377 11339 7435 11345
rect 5031 11308 7328 11336
rect 5031 11305 5043 11308
rect 4985 11299 5043 11305
rect 2924 11240 3096 11268
rect 3421 11271 3479 11277
rect 2924 11228 2930 11240
rect 3421 11237 3433 11271
rect 3467 11268 3479 11271
rect 3467 11240 4292 11268
rect 3467 11237 3479 11240
rect 3421 11231 3479 11237
rect 4264 11212 4292 11240
rect 4522 11228 4528 11280
rect 4580 11228 4586 11280
rect 5813 11271 5871 11277
rect 5813 11237 5825 11271
rect 5859 11268 5871 11271
rect 7300 11268 7328 11308
rect 7377 11305 7389 11339
rect 7423 11336 7435 11339
rect 7466 11336 7472 11348
rect 7423 11308 7472 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 7466 11296 7472 11308
rect 7524 11296 7530 11348
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 7742 11336 7748 11348
rect 7699 11308 7748 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 7742 11296 7748 11308
rect 7800 11336 7806 11348
rect 10137 11339 10195 11345
rect 7800 11308 7972 11336
rect 7800 11296 7806 11308
rect 7561 11271 7619 11277
rect 7561 11268 7573 11271
rect 5859 11240 7052 11268
rect 7300 11240 7573 11268
rect 5859 11237 5871 11240
rect 5813 11231 5871 11237
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 2314 11160 2320 11212
rect 2372 11200 2378 11212
rect 2372 11172 2417 11200
rect 2372 11160 2378 11172
rect 3142 11160 3148 11212
rect 3200 11200 3206 11212
rect 3329 11203 3387 11209
rect 3329 11200 3341 11203
rect 3200 11172 3341 11200
rect 3200 11160 3206 11172
rect 3329 11169 3341 11172
rect 3375 11169 3387 11203
rect 4062 11200 4068 11212
rect 4023 11172 4068 11200
rect 3329 11163 3387 11169
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4246 11160 4252 11212
rect 4304 11160 4310 11212
rect 4540 11200 4568 11228
rect 4893 11203 4951 11209
rect 4540 11172 4660 11200
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11132 2467 11135
rect 2498 11132 2504 11144
rect 2455 11104 2504 11132
rect 2455 11101 2467 11104
rect 2409 11095 2467 11101
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11101 2651 11135
rect 3602 11132 3608 11144
rect 3563 11104 3608 11132
rect 2593 11095 2651 11101
rect 1578 11064 1584 11076
rect 1539 11036 1584 11064
rect 1578 11024 1584 11036
rect 1636 11024 1642 11076
rect 2608 11064 2636 11095
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 4522 11132 4528 11144
rect 3936 11104 4528 11132
rect 3936 11092 3942 11104
rect 4522 11092 4528 11104
rect 4580 11092 4586 11144
rect 3620 11064 3648 11092
rect 2608 11036 3648 11064
rect 4338 11024 4344 11076
rect 4396 11064 4402 11076
rect 4632 11064 4660 11172
rect 4893 11169 4905 11203
rect 4939 11200 4951 11203
rect 5074 11200 5080 11212
rect 4939 11172 5080 11200
rect 4939 11169 4951 11172
rect 4893 11163 4951 11169
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 5166 11160 5172 11212
rect 5224 11200 5230 11212
rect 5353 11203 5411 11209
rect 5353 11200 5365 11203
rect 5224 11172 5365 11200
rect 5224 11160 5230 11172
rect 5353 11169 5365 11172
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 6264 11203 6322 11209
rect 6264 11169 6276 11203
rect 6310 11200 6322 11203
rect 6546 11200 6552 11212
rect 6310 11172 6552 11200
rect 6310 11169 6322 11172
rect 6264 11163 6322 11169
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 5445 11135 5503 11141
rect 5445 11132 5457 11135
rect 5092 11104 5457 11132
rect 5092 11064 5120 11104
rect 5445 11101 5457 11104
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 5537 11135 5595 11141
rect 5537 11101 5549 11135
rect 5583 11101 5595 11135
rect 5537 11095 5595 11101
rect 4396 11036 5120 11064
rect 4396 11024 4402 11036
rect 5166 11024 5172 11076
rect 5224 11064 5230 11076
rect 5552 11064 5580 11095
rect 5810 11092 5816 11144
rect 5868 11132 5874 11144
rect 5997 11135 6055 11141
rect 5997 11132 6009 11135
rect 5868 11104 6009 11132
rect 5868 11092 5874 11104
rect 5997 11101 6009 11104
rect 6043 11101 6055 11135
rect 7024 11132 7052 11240
rect 7561 11237 7573 11240
rect 7607 11237 7619 11271
rect 7561 11231 7619 11237
rect 7944 11209 7972 11308
rect 10137 11305 10149 11339
rect 10183 11336 10195 11339
rect 15657 11339 15715 11345
rect 15657 11336 15669 11339
rect 10183 11308 12020 11336
rect 10183 11305 10195 11308
rect 10137 11299 10195 11305
rect 8202 11277 8208 11280
rect 8196 11268 8208 11277
rect 8163 11240 8208 11268
rect 8196 11231 8208 11240
rect 8202 11228 8208 11231
rect 8260 11228 8266 11280
rect 9677 11271 9735 11277
rect 9677 11237 9689 11271
rect 9723 11268 9735 11271
rect 11882 11268 11888 11280
rect 9723 11240 11888 11268
rect 9723 11237 9735 11240
rect 9677 11231 9735 11237
rect 11882 11228 11888 11240
rect 11940 11228 11946 11280
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 7392 11172 7849 11200
rect 7392 11132 7420 11172
rect 7837 11169 7849 11172
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 7929 11203 7987 11209
rect 7929 11169 7941 11203
rect 7975 11169 7987 11203
rect 10134 11200 10140 11212
rect 7929 11163 7987 11169
rect 8036 11172 10140 11200
rect 7024 11104 7420 11132
rect 7561 11135 7619 11141
rect 5997 11095 6055 11101
rect 7561 11101 7573 11135
rect 7607 11132 7619 11135
rect 8036 11132 8064 11172
rect 10134 11160 10140 11172
rect 10192 11160 10198 11212
rect 10226 11160 10232 11212
rect 10284 11200 10290 11212
rect 10505 11203 10563 11209
rect 10505 11200 10517 11203
rect 10284 11172 10517 11200
rect 10284 11160 10290 11172
rect 10505 11169 10517 11172
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11200 10655 11203
rect 10870 11200 10876 11212
rect 10643 11172 10876 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 10870 11160 10876 11172
rect 10928 11160 10934 11212
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11200 11207 11203
rect 11238 11200 11244 11212
rect 11195 11172 11244 11200
rect 11195 11169 11207 11172
rect 11149 11163 11207 11169
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11416 11203 11474 11209
rect 11416 11169 11428 11203
rect 11462 11200 11474 11203
rect 11698 11200 11704 11212
rect 11462 11172 11704 11200
rect 11462 11169 11474 11172
rect 11416 11163 11474 11169
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 11992 11200 12020 11308
rect 12452 11308 15669 11336
rect 12452 11200 12480 11308
rect 15657 11305 15669 11308
rect 15703 11305 15715 11339
rect 15657 11299 15715 11305
rect 12713 11271 12771 11277
rect 12713 11237 12725 11271
rect 12759 11268 12771 11271
rect 13170 11268 13176 11280
rect 12759 11240 13176 11268
rect 12759 11237 12771 11240
rect 12713 11231 12771 11237
rect 13170 11228 13176 11240
rect 13228 11268 13234 11280
rect 14366 11268 14372 11280
rect 13228 11240 14372 11268
rect 13228 11228 13234 11240
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 15470 11228 15476 11280
rect 15528 11268 15534 11280
rect 15749 11271 15807 11277
rect 15749 11268 15761 11271
rect 15528 11240 15761 11268
rect 15528 11228 15534 11240
rect 15749 11237 15761 11240
rect 15795 11237 15807 11271
rect 15749 11231 15807 11237
rect 13072 11203 13130 11209
rect 13072 11200 13084 11203
rect 11992 11172 12480 11200
rect 12544 11172 13084 11200
rect 7607 11104 8064 11132
rect 10781 11135 10839 11141
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 10781 11101 10793 11135
rect 10827 11132 10839 11135
rect 10962 11132 10968 11144
rect 10827 11104 10968 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 10962 11092 10968 11104
rect 11020 11092 11026 11144
rect 12544 11073 12572 11172
rect 13072 11169 13084 11172
rect 13118 11200 13130 11203
rect 13814 11200 13820 11212
rect 13118 11172 13820 11200
rect 13118 11169 13130 11172
rect 13072 11163 13130 11169
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 13906 11160 13912 11212
rect 13964 11200 13970 11212
rect 14645 11203 14703 11209
rect 14645 11200 14657 11203
rect 13964 11172 14657 11200
rect 13964 11160 13970 11172
rect 14645 11169 14657 11172
rect 14691 11169 14703 11203
rect 16482 11200 16488 11212
rect 16443 11172 16488 11200
rect 14645 11163 14703 11169
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11132 12771 11135
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 12759 11104 12817 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 14366 11092 14372 11144
rect 14424 11132 14430 11144
rect 15838 11132 15844 11144
rect 14424 11104 15424 11132
rect 15799 11104 15844 11132
rect 14424 11092 14430 11104
rect 12529 11067 12587 11073
rect 5224 11036 6040 11064
rect 5224 11024 5230 11036
rect 2314 10956 2320 11008
rect 2372 10996 2378 11008
rect 2682 10996 2688 11008
rect 2372 10968 2688 10996
rect 2372 10956 2378 10968
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 4062 10956 4068 11008
rect 4120 10996 4126 11008
rect 4249 10999 4307 11005
rect 4249 10996 4261 10999
rect 4120 10968 4261 10996
rect 4120 10956 4126 10968
rect 4249 10965 4261 10968
rect 4295 10965 4307 10999
rect 4706 10996 4712 11008
rect 4619 10968 4712 10996
rect 4249 10959 4307 10965
rect 4706 10956 4712 10968
rect 4764 10996 4770 11008
rect 5813 10999 5871 11005
rect 5813 10996 5825 10999
rect 4764 10968 5825 10996
rect 4764 10956 4770 10968
rect 5813 10965 5825 10968
rect 5859 10965 5871 10999
rect 6012 10996 6040 11036
rect 7107 11036 7972 11064
rect 7107 10996 7135 11036
rect 6012 10968 7135 10996
rect 5813 10959 5871 10965
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 7742 10996 7748 11008
rect 7248 10968 7748 10996
rect 7248 10956 7254 10968
rect 7742 10956 7748 10968
rect 7800 10956 7806 11008
rect 7944 10996 7972 11036
rect 12529 11033 12541 11067
rect 12575 11033 12587 11067
rect 12529 11027 12587 11033
rect 14642 11024 14648 11076
rect 14700 11064 14706 11076
rect 15289 11067 15347 11073
rect 15289 11064 15301 11067
rect 14700 11036 15301 11064
rect 14700 11024 14706 11036
rect 15289 11033 15301 11036
rect 15335 11033 15347 11067
rect 15396 11064 15424 11104
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 16301 11067 16359 11073
rect 16301 11064 16313 11067
rect 15396 11036 16313 11064
rect 15289 11027 15347 11033
rect 16301 11033 16313 11036
rect 16347 11033 16359 11067
rect 16301 11027 16359 11033
rect 9214 10996 9220 11008
rect 7944 10968 9220 10996
rect 9214 10956 9220 10968
rect 9272 10996 9278 11008
rect 9309 10999 9367 11005
rect 9309 10996 9321 10999
rect 9272 10968 9321 10996
rect 9272 10956 9278 10968
rect 9309 10965 9321 10968
rect 9355 10965 9367 10999
rect 9309 10959 9367 10965
rect 10686 10956 10692 11008
rect 10744 10996 10750 11008
rect 11514 10996 11520 11008
rect 10744 10968 11520 10996
rect 10744 10956 10750 10968
rect 11514 10956 11520 10968
rect 11572 10956 11578 11008
rect 11790 10956 11796 11008
rect 11848 10996 11854 11008
rect 13906 10996 13912 11008
rect 11848 10968 13912 10996
rect 11848 10956 11854 10968
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 13998 10956 14004 11008
rect 14056 10996 14062 11008
rect 14185 10999 14243 11005
rect 14185 10996 14197 10999
rect 14056 10968 14197 10996
rect 14056 10956 14062 10968
rect 14185 10965 14197 10968
rect 14231 10965 14243 10999
rect 14185 10959 14243 10965
rect 14829 10999 14887 11005
rect 14829 10965 14841 10999
rect 14875 10996 14887 10999
rect 14918 10996 14924 11008
rect 14875 10968 14924 10996
rect 14875 10965 14887 10968
rect 14829 10959 14887 10965
rect 14918 10956 14924 10968
rect 14976 10956 14982 11008
rect 1104 10906 16836 10928
rect 1104 10854 3614 10906
rect 3666 10854 3678 10906
rect 3730 10854 3742 10906
rect 3794 10854 3806 10906
rect 3858 10854 8878 10906
rect 8930 10854 8942 10906
rect 8994 10854 9006 10906
rect 9058 10854 9070 10906
rect 9122 10854 14142 10906
rect 14194 10854 14206 10906
rect 14258 10854 14270 10906
rect 14322 10854 14334 10906
rect 14386 10854 16836 10906
rect 1104 10832 16836 10854
rect 2777 10795 2835 10801
rect 2777 10761 2789 10795
rect 2823 10792 2835 10795
rect 2866 10792 2872 10804
rect 2823 10764 2872 10792
rect 2823 10761 2835 10764
rect 2777 10755 2835 10761
rect 2866 10752 2872 10764
rect 2924 10752 2930 10804
rect 3050 10792 3056 10804
rect 3011 10764 3056 10792
rect 3050 10752 3056 10764
rect 3108 10752 3114 10804
rect 4065 10795 4123 10801
rect 4065 10761 4077 10795
rect 4111 10792 4123 10795
rect 4154 10792 4160 10804
rect 4111 10764 4160 10792
rect 4111 10761 4123 10764
rect 4065 10755 4123 10761
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 5810 10792 5816 10804
rect 5092 10764 5816 10792
rect 3510 10684 3516 10736
rect 3568 10724 3574 10736
rect 3568 10696 3740 10724
rect 3568 10684 3574 10696
rect 2406 10616 2412 10668
rect 2464 10656 2470 10668
rect 3712 10665 3740 10696
rect 3697 10659 3755 10665
rect 2464 10628 3648 10656
rect 2464 10616 2470 10628
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1486 10588 1492 10600
rect 1443 10560 1492 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1486 10548 1492 10560
rect 1544 10548 1550 10600
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 3234 10588 3240 10600
rect 3108 10560 3240 10588
rect 3108 10548 3114 10560
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 3326 10548 3332 10600
rect 3384 10588 3390 10600
rect 3513 10591 3571 10597
rect 3513 10588 3525 10591
rect 3384 10560 3525 10588
rect 3384 10548 3390 10560
rect 3513 10557 3525 10560
rect 3559 10557 3571 10591
rect 3620 10588 3648 10628
rect 3697 10625 3709 10659
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 5092 10665 5120 10764
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 11238 10792 11244 10804
rect 8680 10764 11244 10792
rect 6178 10684 6184 10736
rect 6236 10724 6242 10736
rect 8478 10724 8484 10736
rect 6236 10696 8484 10724
rect 6236 10684 6242 10696
rect 8478 10684 8484 10696
rect 8536 10684 8542 10736
rect 4617 10659 4675 10665
rect 4617 10656 4629 10659
rect 4396 10628 4629 10656
rect 4396 10616 4402 10628
rect 4617 10625 4629 10628
rect 4663 10625 4675 10659
rect 4617 10619 4675 10625
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10625 5135 10659
rect 7466 10656 7472 10668
rect 7427 10628 7472 10656
rect 5077 10619 5135 10625
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 8680 10665 8708 10764
rect 10045 10727 10103 10733
rect 10045 10724 10057 10727
rect 9692 10696 10057 10724
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 4433 10591 4491 10597
rect 4433 10588 4445 10591
rect 3620 10560 4445 10588
rect 3513 10551 3571 10557
rect 4433 10557 4445 10560
rect 4479 10588 4491 10591
rect 4982 10588 4988 10600
rect 4479 10560 4988 10588
rect 4479 10557 4491 10560
rect 4433 10551 4491 10557
rect 4982 10548 4988 10560
rect 5040 10548 5046 10600
rect 5344 10591 5402 10597
rect 5344 10557 5356 10591
rect 5390 10588 5402 10591
rect 5626 10588 5632 10600
rect 5390 10560 5632 10588
rect 5390 10557 5402 10560
rect 5344 10551 5402 10557
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 7006 10548 7012 10600
rect 7064 10588 7070 10600
rect 7834 10588 7840 10600
rect 7064 10560 7840 10588
rect 7064 10548 7070 10560
rect 7834 10548 7840 10560
rect 7892 10588 7898 10600
rect 7892 10560 7972 10588
rect 7892 10548 7898 10560
rect 1664 10523 1722 10529
rect 1664 10489 1676 10523
rect 1710 10520 1722 10523
rect 2958 10520 2964 10532
rect 1710 10492 2964 10520
rect 1710 10489 1722 10492
rect 1664 10483 1722 10489
rect 2958 10480 2964 10492
rect 3016 10480 3022 10532
rect 4154 10520 4160 10532
rect 3068 10492 4160 10520
rect 2498 10412 2504 10464
rect 2556 10452 2562 10464
rect 3068 10452 3096 10492
rect 4154 10480 4160 10492
rect 4212 10520 4218 10532
rect 4212 10492 4568 10520
rect 4212 10480 4218 10492
rect 3418 10452 3424 10464
rect 2556 10424 3096 10452
rect 3379 10424 3424 10452
rect 2556 10412 2562 10424
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 4540 10461 4568 10492
rect 5534 10480 5540 10532
rect 5592 10520 5598 10532
rect 7285 10523 7343 10529
rect 7285 10520 7297 10523
rect 5592 10492 7297 10520
rect 5592 10480 5598 10492
rect 7285 10489 7297 10492
rect 7331 10489 7343 10523
rect 7944 10520 7972 10560
rect 8018 10548 8024 10600
rect 8076 10588 8082 10600
rect 8113 10591 8171 10597
rect 8113 10588 8125 10591
rect 8076 10560 8125 10588
rect 8076 10548 8082 10560
rect 8113 10557 8125 10560
rect 8159 10588 8171 10591
rect 8202 10588 8208 10600
rect 8159 10560 8208 10588
rect 8159 10557 8171 10560
rect 8113 10551 8171 10557
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 8932 10591 8990 10597
rect 8932 10557 8944 10591
rect 8978 10588 8990 10591
rect 9214 10588 9220 10600
rect 8978 10560 9220 10588
rect 8978 10557 8990 10560
rect 8932 10551 8990 10557
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9692 10588 9720 10696
rect 10045 10693 10057 10696
rect 10091 10693 10103 10727
rect 10045 10687 10103 10693
rect 10336 10665 10364 10764
rect 11238 10752 11244 10764
rect 11296 10792 11302 10804
rect 12158 10792 12164 10804
rect 11296 10764 12164 10792
rect 11296 10752 11302 10764
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12268 10764 12848 10792
rect 11698 10724 11704 10736
rect 11611 10696 11704 10724
rect 11698 10684 11704 10696
rect 11756 10724 11762 10736
rect 11882 10724 11888 10736
rect 11756 10696 11888 10724
rect 11756 10684 11762 10696
rect 11882 10684 11888 10696
rect 11940 10684 11946 10736
rect 11974 10684 11980 10736
rect 12032 10724 12038 10736
rect 12032 10696 12077 10724
rect 12032 10684 12038 10696
rect 10321 10659 10379 10665
rect 10321 10625 10333 10659
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 12268 10656 12296 10764
rect 12710 10724 12716 10736
rect 12671 10696 12716 10724
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 12820 10724 12848 10764
rect 12894 10752 12900 10804
rect 12952 10792 12958 10804
rect 16482 10792 16488 10804
rect 12952 10764 16488 10792
rect 12952 10752 12958 10764
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 13354 10724 13360 10736
rect 12820 10696 13216 10724
rect 11572 10628 12296 10656
rect 11572 10616 11578 10628
rect 12342 10616 12348 10668
rect 12400 10656 12406 10668
rect 13078 10656 13084 10668
rect 12400 10628 13084 10656
rect 12400 10616 12406 10628
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 13188 10665 13216 10696
rect 13280 10696 13360 10724
rect 13280 10665 13308 10696
rect 13354 10684 13360 10696
rect 13412 10684 13418 10736
rect 13446 10684 13452 10736
rect 13504 10724 13510 10736
rect 13504 10696 14504 10724
rect 13504 10684 13510 10696
rect 14476 10668 14504 10696
rect 16114 10684 16120 10736
rect 16172 10724 16178 10736
rect 16301 10727 16359 10733
rect 16301 10724 16313 10727
rect 16172 10696 16313 10724
rect 16172 10684 16178 10696
rect 16301 10693 16313 10696
rect 16347 10693 16359 10727
rect 16301 10687 16359 10693
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 13265 10659 13323 10665
rect 13265 10625 13277 10659
rect 13311 10625 13323 10659
rect 13265 10619 13323 10625
rect 9324 10560 9720 10588
rect 10588 10591 10646 10597
rect 9324 10520 9352 10560
rect 10588 10557 10600 10591
rect 10634 10588 10646 10591
rect 10962 10588 10968 10600
rect 10634 10560 10968 10588
rect 10634 10557 10646 10560
rect 10588 10551 10646 10557
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 12158 10588 12164 10600
rect 12119 10560 12164 10588
rect 12158 10548 12164 10560
rect 12216 10548 12222 10600
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12710 10588 12716 10600
rect 12492 10560 12716 10588
rect 12492 10548 12498 10560
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 7944 10492 9352 10520
rect 7285 10483 7343 10489
rect 10042 10480 10048 10532
rect 10100 10520 10106 10532
rect 11054 10520 11060 10532
rect 10100 10492 11060 10520
rect 10100 10480 10106 10492
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 13188 10520 13216 10619
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 14277 10659 14335 10665
rect 14277 10656 14289 10659
rect 13872 10628 14289 10656
rect 13872 10616 13878 10628
rect 14277 10625 14289 10628
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 14458 10616 14464 10668
rect 14516 10616 14522 10668
rect 14642 10616 14648 10668
rect 14700 10656 14706 10668
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 14700 10628 14933 10656
rect 14700 10616 14706 10628
rect 14921 10625 14933 10628
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 13630 10548 13636 10600
rect 13688 10548 13694 10600
rect 15188 10591 15246 10597
rect 15188 10557 15200 10591
rect 15234 10588 15246 10591
rect 15930 10588 15936 10600
rect 15234 10560 15936 10588
rect 15234 10557 15246 10560
rect 15188 10551 15246 10557
rect 15930 10548 15936 10560
rect 15988 10548 15994 10600
rect 13648 10520 13676 10548
rect 13188 10492 13584 10520
rect 13648 10492 13768 10520
rect 4525 10455 4583 10461
rect 4525 10421 4537 10455
rect 4571 10452 4583 10455
rect 5902 10452 5908 10464
rect 4571 10424 5908 10452
rect 4571 10421 4583 10424
rect 4525 10415 4583 10421
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 6457 10455 6515 10461
rect 6457 10421 6469 10455
rect 6503 10452 6515 10455
rect 6546 10452 6552 10464
rect 6503 10424 6552 10452
rect 6503 10421 6515 10424
rect 6457 10415 6515 10421
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 6825 10455 6883 10461
rect 6825 10421 6837 10455
rect 6871 10452 6883 10455
rect 6914 10452 6920 10464
rect 6871 10424 6920 10452
rect 6871 10421 6883 10424
rect 6825 10415 6883 10421
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 7190 10452 7196 10464
rect 7151 10424 7196 10452
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 8297 10455 8355 10461
rect 8297 10421 8309 10455
rect 8343 10452 8355 10455
rect 12342 10452 12348 10464
rect 8343 10424 12348 10452
rect 8343 10421 8355 10424
rect 8297 10415 8355 10421
rect 12342 10412 12348 10424
rect 12400 10412 12406 10464
rect 13078 10452 13084 10464
rect 12991 10424 13084 10452
rect 13078 10412 13084 10424
rect 13136 10452 13142 10464
rect 13354 10452 13360 10464
rect 13136 10424 13360 10452
rect 13136 10412 13142 10424
rect 13354 10412 13360 10424
rect 13412 10412 13418 10464
rect 13556 10452 13584 10492
rect 13630 10452 13636 10464
rect 13556 10424 13636 10452
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 13740 10461 13768 10492
rect 13814 10480 13820 10532
rect 13872 10520 13878 10532
rect 14093 10523 14151 10529
rect 14093 10520 14105 10523
rect 13872 10492 14105 10520
rect 13872 10480 13878 10492
rect 14093 10489 14105 10492
rect 14139 10489 14151 10523
rect 14093 10483 14151 10489
rect 13725 10455 13783 10461
rect 13725 10421 13737 10455
rect 13771 10421 13783 10455
rect 14182 10452 14188 10464
rect 14143 10424 14188 10452
rect 13725 10415 13783 10421
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 14550 10412 14556 10464
rect 14608 10452 14614 10464
rect 15838 10452 15844 10464
rect 14608 10424 15844 10452
rect 14608 10412 14614 10424
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 1104 10362 16836 10384
rect 1104 10310 6246 10362
rect 6298 10310 6310 10362
rect 6362 10310 6374 10362
rect 6426 10310 6438 10362
rect 6490 10310 11510 10362
rect 11562 10310 11574 10362
rect 11626 10310 11638 10362
rect 11690 10310 11702 10362
rect 11754 10310 16836 10362
rect 1104 10288 16836 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 2682 10248 2688 10260
rect 1544 10220 2688 10248
rect 1544 10208 1550 10220
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1854 10112 1860 10124
rect 1443 10084 1860 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 1964 10121 1992 10220
rect 2682 10208 2688 10220
rect 2740 10248 2746 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 2740 10220 3617 10248
rect 2740 10208 2746 10220
rect 3605 10217 3617 10220
rect 3651 10217 3663 10251
rect 3605 10211 3663 10217
rect 4525 10251 4583 10257
rect 4525 10217 4537 10251
rect 4571 10217 4583 10251
rect 4982 10248 4988 10260
rect 4943 10220 4988 10248
rect 4525 10211 4583 10217
rect 2216 10183 2274 10189
rect 2216 10149 2228 10183
rect 2262 10180 2274 10183
rect 2866 10180 2872 10192
rect 2262 10152 2872 10180
rect 2262 10149 2274 10152
rect 2216 10143 2274 10149
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 3510 10140 3516 10192
rect 3568 10140 3574 10192
rect 4540 10180 4568 10211
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 5534 10248 5540 10260
rect 5495 10220 5540 10248
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 5718 10208 5724 10260
rect 5776 10248 5782 10260
rect 5997 10251 6055 10257
rect 5997 10248 6009 10251
rect 5776 10220 6009 10248
rect 5776 10208 5782 10220
rect 5997 10217 6009 10220
rect 6043 10217 6055 10251
rect 5997 10211 6055 10217
rect 6825 10251 6883 10257
rect 6825 10217 6837 10251
rect 6871 10217 6883 10251
rect 7190 10248 7196 10260
rect 7151 10220 7196 10248
rect 6825 10211 6883 10217
rect 5905 10183 5963 10189
rect 5905 10180 5917 10183
rect 4540 10152 5917 10180
rect 5905 10149 5917 10152
rect 5951 10149 5963 10183
rect 5905 10143 5963 10149
rect 6362 10140 6368 10192
rect 6420 10180 6426 10192
rect 6840 10180 6868 10211
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 7561 10251 7619 10257
rect 7561 10217 7573 10251
rect 7607 10248 7619 10251
rect 8205 10251 8263 10257
rect 8205 10248 8217 10251
rect 7607 10220 8217 10248
rect 7607 10217 7619 10220
rect 7561 10211 7619 10217
rect 8205 10217 8217 10220
rect 8251 10217 8263 10251
rect 8205 10211 8263 10217
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 8665 10251 8723 10257
rect 8665 10248 8677 10251
rect 8352 10220 8677 10248
rect 8352 10208 8358 10220
rect 8665 10217 8677 10220
rect 8711 10248 8723 10251
rect 9398 10248 9404 10260
rect 8711 10220 9404 10248
rect 8711 10217 8723 10220
rect 8665 10211 8723 10217
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 14182 10248 14188 10260
rect 10183 10220 14188 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 14182 10208 14188 10220
rect 14240 10208 14246 10260
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 15657 10251 15715 10257
rect 15657 10248 15669 10251
rect 14516 10220 15669 10248
rect 14516 10208 14522 10220
rect 15657 10217 15669 10220
rect 15703 10248 15715 10251
rect 16114 10248 16120 10260
rect 15703 10220 16120 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 6420 10152 6868 10180
rect 8573 10183 8631 10189
rect 6420 10140 6426 10152
rect 8573 10149 8585 10183
rect 8619 10180 8631 10183
rect 9677 10183 9735 10189
rect 9677 10180 9689 10183
rect 8619 10152 9689 10180
rect 8619 10149 8631 10152
rect 8573 10143 8631 10149
rect 9677 10149 9689 10152
rect 9723 10149 9735 10183
rect 11974 10180 11980 10192
rect 9677 10143 9735 10149
rect 10336 10152 11980 10180
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10081 2007 10115
rect 1949 10075 2007 10081
rect 2774 10072 2780 10124
rect 2832 10112 2838 10124
rect 3142 10112 3148 10124
rect 2832 10084 3148 10112
rect 2832 10072 2838 10084
rect 3142 10072 3148 10084
rect 3200 10072 3206 10124
rect 3528 10044 3556 10140
rect 3789 10115 3847 10121
rect 3789 10081 3801 10115
rect 3835 10112 3847 10115
rect 4706 10112 4712 10124
rect 3835 10084 4712 10112
rect 3835 10081 3847 10084
rect 3789 10075 3847 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 4893 10115 4951 10121
rect 4893 10081 4905 10115
rect 4939 10081 4951 10115
rect 4893 10075 4951 10081
rect 4908 10044 4936 10075
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 6641 10115 6699 10121
rect 6641 10112 6653 10115
rect 5500 10084 6653 10112
rect 5500 10072 5506 10084
rect 6641 10081 6653 10084
rect 6687 10112 6699 10115
rect 9493 10115 9551 10121
rect 6687 10084 8892 10112
rect 6687 10081 6699 10084
rect 6641 10075 6699 10081
rect 3528 10016 4936 10044
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10044 5227 10047
rect 5534 10044 5540 10056
rect 5215 10016 5540 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 3694 9936 3700 9988
rect 3752 9936 3758 9988
rect 6196 9976 6224 10007
rect 6454 10004 6460 10056
rect 6512 10044 6518 10056
rect 6730 10044 6736 10056
rect 6512 10016 6736 10044
rect 6512 10004 6518 10016
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 7006 10004 7012 10056
rect 7064 10044 7070 10056
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 7064 10016 7665 10044
rect 7064 10004 7070 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 8754 10044 8760 10056
rect 8715 10016 8760 10044
rect 7745 10007 7803 10013
rect 6546 9976 6552 9988
rect 6196 9948 6552 9976
rect 6546 9936 6552 9948
rect 6604 9976 6610 9988
rect 7760 9976 7788 10007
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 8864 10044 8892 10084
rect 9493 10081 9505 10115
rect 9539 10112 9551 10115
rect 10336 10112 10364 10152
rect 11974 10140 11980 10152
rect 12032 10140 12038 10192
rect 12526 10140 12532 10192
rect 12584 10140 12590 10192
rect 12710 10180 12716 10192
rect 12671 10152 12716 10180
rect 12710 10140 12716 10152
rect 12768 10140 12774 10192
rect 12805 10183 12863 10189
rect 12805 10149 12817 10183
rect 12851 10180 12863 10183
rect 12894 10180 12900 10192
rect 12851 10152 12900 10180
rect 12851 10149 12863 10152
rect 12805 10143 12863 10149
rect 12894 10140 12900 10152
rect 12952 10140 12958 10192
rect 13808 10183 13866 10189
rect 13096 10152 13768 10180
rect 10502 10112 10508 10124
rect 9539 10084 10364 10112
rect 10463 10084 10508 10112
rect 9539 10081 9551 10084
rect 9493 10075 9551 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 11238 10112 11244 10124
rect 10704 10084 11244 10112
rect 10226 10044 10232 10056
rect 8864 10016 10232 10044
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 10318 10004 10324 10056
rect 10376 10044 10382 10056
rect 10597 10047 10655 10053
rect 10597 10044 10609 10047
rect 10376 10016 10609 10044
rect 10376 10004 10382 10016
rect 10597 10013 10609 10016
rect 10643 10013 10655 10047
rect 10597 10007 10655 10013
rect 6604 9948 7788 9976
rect 9309 9979 9367 9985
rect 6604 9936 6610 9948
rect 9309 9945 9321 9979
rect 9355 9976 9367 9979
rect 10704 9976 10732 10084
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10112 11575 10115
rect 12544 10112 12572 10140
rect 13096 10112 13124 10152
rect 11563 10084 12480 10112
rect 12544 10084 13124 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 10781 10047 10839 10053
rect 10781 10013 10793 10047
rect 10827 10013 10839 10047
rect 10781 10007 10839 10013
rect 9355 9948 10732 9976
rect 10796 9976 10824 10007
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11609 10047 11667 10053
rect 11609 10044 11621 10047
rect 11112 10016 11621 10044
rect 11112 10004 11118 10016
rect 11609 10013 11621 10016
rect 11655 10013 11667 10047
rect 11790 10044 11796 10056
rect 11751 10016 11796 10044
rect 11609 10007 11667 10013
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 12452 10044 12480 10084
rect 13170 10072 13176 10124
rect 13228 10112 13234 10124
rect 13538 10112 13544 10124
rect 13228 10084 13544 10112
rect 13228 10072 13234 10084
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 13740 10112 13768 10152
rect 13808 10149 13820 10183
rect 13854 10180 13866 10183
rect 13906 10180 13912 10192
rect 13854 10152 13912 10180
rect 13854 10149 13866 10152
rect 13808 10143 13866 10149
rect 13906 10140 13912 10152
rect 13964 10180 13970 10192
rect 13964 10152 15884 10180
rect 13964 10140 13970 10152
rect 14090 10112 14096 10124
rect 13740 10084 14096 10112
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 15620 10084 15761 10112
rect 15620 10072 15626 10084
rect 15749 10081 15761 10084
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 12526 10044 12532 10056
rect 12452 10016 12532 10044
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 12989 10047 13047 10053
rect 12989 10013 13001 10047
rect 13035 10044 13047 10047
rect 13078 10044 13084 10056
rect 13035 10016 13084 10044
rect 13035 10013 13047 10016
rect 12989 10007 13047 10013
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 15856 10053 15884 10152
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10013 15899 10047
rect 15841 10007 15899 10013
rect 11882 9976 11888 9988
rect 10796 9948 11888 9976
rect 9355 9945 9367 9948
rect 9309 9939 9367 9945
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 12434 9976 12440 9988
rect 11992 9948 12440 9976
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 2866 9908 2872 9920
rect 1627 9880 2872 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 2866 9868 2872 9880
rect 2924 9868 2930 9920
rect 3326 9908 3332 9920
rect 3287 9880 3332 9908
rect 3326 9868 3332 9880
rect 3384 9868 3390 9920
rect 3712 9908 3740 9936
rect 6270 9908 6276 9920
rect 3712 9880 6276 9908
rect 6270 9868 6276 9880
rect 6328 9868 6334 9920
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 9214 9908 9220 9920
rect 8444 9880 9220 9908
rect 8444 9868 8450 9880
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 9582 9868 9588 9920
rect 9640 9908 9646 9920
rect 9766 9908 9772 9920
rect 9640 9880 9772 9908
rect 9640 9868 9646 9880
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 10594 9868 10600 9920
rect 10652 9908 10658 9920
rect 11149 9911 11207 9917
rect 11149 9908 11161 9911
rect 10652 9880 11161 9908
rect 10652 9868 10658 9880
rect 11149 9877 11161 9880
rect 11195 9877 11207 9911
rect 11149 9871 11207 9877
rect 11422 9868 11428 9920
rect 11480 9908 11486 9920
rect 11992 9908 12020 9948
rect 12434 9936 12440 9948
rect 12492 9976 12498 9988
rect 13170 9976 13176 9988
rect 12492 9948 13176 9976
rect 12492 9936 12498 9948
rect 13170 9936 13176 9948
rect 13228 9936 13234 9988
rect 11480 9880 12020 9908
rect 12345 9911 12403 9917
rect 11480 9868 11486 9880
rect 12345 9877 12357 9911
rect 12391 9908 12403 9911
rect 13906 9908 13912 9920
rect 12391 9880 13912 9908
rect 12391 9877 12403 9880
rect 12345 9871 12403 9877
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 14921 9911 14979 9917
rect 14921 9877 14933 9911
rect 14967 9908 14979 9911
rect 15010 9908 15016 9920
rect 14967 9880 15016 9908
rect 14967 9877 14979 9880
rect 14921 9871 14979 9877
rect 15010 9868 15016 9880
rect 15068 9868 15074 9920
rect 15286 9908 15292 9920
rect 15247 9880 15292 9908
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 1104 9818 16836 9840
rect 1104 9766 3614 9818
rect 3666 9766 3678 9818
rect 3730 9766 3742 9818
rect 3794 9766 3806 9818
rect 3858 9766 8878 9818
rect 8930 9766 8942 9818
rect 8994 9766 9006 9818
rect 9058 9766 9070 9818
rect 9122 9766 14142 9818
rect 14194 9766 14206 9818
rect 14258 9766 14270 9818
rect 14322 9766 14334 9818
rect 14386 9766 16836 9818
rect 1104 9744 16836 9766
rect 2682 9664 2688 9716
rect 2740 9704 2746 9716
rect 3053 9707 3111 9713
rect 3053 9704 3065 9707
rect 2740 9676 3065 9704
rect 2740 9664 2746 9676
rect 3053 9673 3065 9676
rect 3099 9673 3111 9707
rect 3418 9704 3424 9716
rect 3053 9667 3111 9673
rect 3160 9676 3424 9704
rect 1946 9528 1952 9580
rect 2004 9568 2010 9580
rect 2593 9571 2651 9577
rect 2593 9568 2605 9571
rect 2004 9540 2605 9568
rect 2004 9528 2010 9540
rect 2593 9537 2605 9540
rect 2639 9568 2651 9571
rect 2682 9568 2688 9580
rect 2639 9540 2688 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9537 2835 9571
rect 3160 9568 3188 9676
rect 3418 9664 3424 9676
rect 3476 9664 3482 9716
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 6730 9704 6736 9716
rect 6420 9676 6736 9704
rect 6420 9664 6426 9676
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 6840 9676 8217 9704
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 5442 9636 5448 9648
rect 4304 9608 5448 9636
rect 4304 9596 4310 9608
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 5721 9639 5779 9645
rect 5721 9605 5733 9639
rect 5767 9636 5779 9639
rect 6546 9636 6552 9648
rect 5767 9608 6552 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 6546 9596 6552 9608
rect 6604 9596 6610 9648
rect 3160 9540 3271 9568
rect 2777 9531 2835 9537
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9500 1639 9503
rect 1670 9500 1676 9512
rect 1627 9472 1676 9500
rect 1627 9469 1639 9472
rect 1581 9463 1639 9469
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 2501 9435 2559 9441
rect 2501 9401 2513 9435
rect 2547 9432 2559 9435
rect 2792 9432 2820 9531
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9500 3111 9503
rect 3145 9503 3203 9509
rect 3145 9500 3157 9503
rect 3099 9472 3157 9500
rect 3099 9469 3111 9472
rect 3053 9463 3111 9469
rect 3145 9469 3157 9472
rect 3191 9469 3203 9503
rect 3243 9500 3271 9540
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4522 9568 4528 9580
rect 4212 9540 4528 9568
rect 4212 9528 4218 9540
rect 4522 9528 4528 9540
rect 4580 9568 4586 9580
rect 4580 9540 5396 9568
rect 4580 9528 4586 9540
rect 3412 9503 3470 9509
rect 3412 9500 3424 9503
rect 3243 9472 3424 9500
rect 3145 9463 3203 9469
rect 3412 9469 3424 9472
rect 3458 9500 3470 9503
rect 3694 9500 3700 9512
rect 3458 9472 3700 9500
rect 3458 9469 3470 9472
rect 3412 9463 3470 9469
rect 3694 9460 3700 9472
rect 3752 9460 3758 9512
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9500 4859 9503
rect 5258 9500 5264 9512
rect 4847 9472 5264 9500
rect 4847 9469 4859 9472
rect 4801 9463 4859 9469
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 2547 9404 2728 9432
rect 2792 9404 3280 9432
rect 2547 9401 2559 9404
rect 2501 9395 2559 9401
rect 1762 9364 1768 9376
rect 1723 9336 1768 9364
rect 1762 9324 1768 9336
rect 1820 9324 1826 9376
rect 2130 9364 2136 9376
rect 2091 9336 2136 9364
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 2700 9364 2728 9404
rect 2774 9364 2780 9376
rect 2700 9336 2780 9364
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 3252 9364 3280 9404
rect 3326 9392 3332 9444
rect 3384 9432 3390 9444
rect 5368 9432 5396 9540
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 5592 9540 6377 9568
rect 5592 9528 5598 9540
rect 6365 9537 6377 9540
rect 6411 9568 6423 9571
rect 6840 9568 6868 9676
rect 8205 9673 8217 9676
rect 8251 9704 8263 9707
rect 8754 9704 8760 9716
rect 8251 9676 8760 9704
rect 8251 9673 8263 9676
rect 8205 9667 8263 9673
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 10137 9707 10195 9713
rect 10137 9673 10149 9707
rect 10183 9704 10195 9707
rect 10502 9704 10508 9716
rect 10183 9676 10508 9704
rect 10183 9673 10195 9676
rect 10137 9667 10195 9673
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 11422 9704 11428 9716
rect 10836 9676 11428 9704
rect 10836 9664 10842 9676
rect 11422 9664 11428 9676
rect 11480 9664 11486 9716
rect 11882 9664 11888 9716
rect 11940 9704 11946 9716
rect 11940 9676 13216 9704
rect 11940 9664 11946 9676
rect 11149 9639 11207 9645
rect 11149 9605 11161 9639
rect 11195 9605 11207 9639
rect 11149 9599 11207 9605
rect 9769 9571 9827 9577
rect 6411 9540 6868 9568
rect 8312 9540 9720 9568
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 5994 9460 6000 9512
rect 6052 9500 6058 9512
rect 6181 9503 6239 9509
rect 6181 9500 6193 9503
rect 6052 9472 6193 9500
rect 6052 9460 6058 9472
rect 6181 9469 6193 9472
rect 6227 9469 6239 9503
rect 6822 9500 6828 9512
rect 6783 9472 6828 9500
rect 6181 9463 6239 9469
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 7098 9509 7104 9512
rect 7092 9463 7104 9509
rect 7156 9500 7162 9512
rect 7156 9472 7192 9500
rect 7098 9460 7104 9463
rect 7156 9460 7162 9472
rect 7558 9460 7564 9512
rect 7616 9500 7622 9512
rect 8202 9500 8208 9512
rect 7616 9472 8208 9500
rect 7616 9460 7622 9472
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 8312 9432 8340 9540
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 9582 9500 9588 9512
rect 8619 9472 9588 9500
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 3384 9404 5028 9432
rect 5368 9404 8340 9432
rect 3384 9392 3390 9404
rect 4338 9364 4344 9376
rect 3252 9336 4344 9364
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 4614 9364 4620 9376
rect 4571 9336 4620 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 5000 9373 5028 9404
rect 4985 9367 5043 9373
rect 4985 9333 4997 9367
rect 5031 9333 5043 9367
rect 4985 9327 5043 9333
rect 6089 9367 6147 9373
rect 6089 9333 6101 9367
rect 6135 9364 6147 9367
rect 7466 9364 7472 9376
rect 6135 9336 7472 9364
rect 6135 9333 6147 9336
rect 6089 9327 6147 9333
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 7926 9324 7932 9376
rect 7984 9364 7990 9376
rect 8588 9364 8616 9463
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 8846 9392 8852 9444
rect 8904 9432 8910 9444
rect 9493 9435 9551 9441
rect 9493 9432 9505 9435
rect 8904 9404 9505 9432
rect 8904 9392 8910 9404
rect 9493 9401 9505 9404
rect 9539 9401 9551 9435
rect 9692 9432 9720 9540
rect 9769 9537 9781 9571
rect 9815 9568 9827 9571
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9815 9540 9965 9568
rect 9815 9537 9827 9540
rect 9769 9531 9827 9537
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 10594 9568 10600 9580
rect 10555 9540 10600 9568
rect 9953 9531 10011 9537
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9568 10839 9571
rect 10962 9568 10968 9580
rect 10827 9540 10968 9568
rect 10827 9537 10839 9540
rect 10781 9531 10839 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11164 9568 11192 9599
rect 11422 9568 11428 9580
rect 11164 9540 11428 9568
rect 11422 9528 11428 9540
rect 11480 9528 11486 9580
rect 11790 9568 11796 9580
rect 11751 9540 11796 9568
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 12894 9528 12900 9580
rect 12952 9568 12958 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12952 9540 13001 9568
rect 12952 9528 12958 9540
rect 12989 9537 13001 9540
rect 13035 9568 13047 9571
rect 13078 9568 13084 9580
rect 13035 9540 13084 9568
rect 13035 9537 13047 9540
rect 12989 9531 13047 9537
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 13188 9568 13216 9676
rect 13538 9664 13544 9716
rect 13596 9704 13602 9716
rect 13596 9676 14320 9704
rect 13596 9664 13602 9676
rect 13449 9639 13507 9645
rect 13449 9605 13461 9639
rect 13495 9636 13507 9639
rect 13814 9636 13820 9648
rect 13495 9608 13820 9636
rect 13495 9605 13507 9608
rect 13449 9599 13507 9605
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14001 9571 14059 9577
rect 14001 9568 14013 9571
rect 13188 9540 14013 9568
rect 14001 9537 14013 9540
rect 14047 9537 14059 9571
rect 14292 9568 14320 9676
rect 15930 9664 15936 9716
rect 15988 9704 15994 9716
rect 16209 9707 16267 9713
rect 16209 9704 16221 9707
rect 15988 9676 16221 9704
rect 15988 9664 15994 9676
rect 16209 9673 16221 9676
rect 16255 9673 16267 9707
rect 16209 9667 16267 9673
rect 14829 9571 14887 9577
rect 14829 9568 14841 9571
rect 14292 9540 14841 9568
rect 14001 9531 14059 9537
rect 14829 9537 14841 9540
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 10226 9460 10232 9512
rect 10284 9500 10290 9512
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 10284 9472 10517 9500
rect 10284 9460 10290 9472
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 10505 9463 10563 9469
rect 12805 9503 12863 9509
rect 12805 9469 12817 9503
rect 12851 9500 12863 9503
rect 13722 9500 13728 9512
rect 12851 9472 13728 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 13722 9460 13728 9472
rect 13780 9460 13786 9512
rect 13906 9500 13912 9512
rect 13867 9472 13912 9500
rect 13906 9460 13912 9472
rect 13964 9460 13970 9512
rect 11882 9432 11888 9444
rect 9692 9404 11888 9432
rect 9493 9395 9551 9401
rect 11882 9392 11888 9404
rect 11940 9392 11946 9444
rect 12897 9435 12955 9441
rect 12897 9401 12909 9435
rect 12943 9432 12955 9435
rect 12986 9432 12992 9444
rect 12943 9404 12992 9432
rect 12943 9401 12955 9404
rect 12897 9395 12955 9401
rect 12986 9392 12992 9404
rect 13044 9392 13050 9444
rect 13078 9392 13084 9444
rect 13136 9432 13142 9444
rect 14826 9432 14832 9444
rect 13136 9404 14832 9432
rect 13136 9392 13142 9404
rect 14826 9392 14832 9404
rect 14884 9392 14890 9444
rect 14918 9392 14924 9444
rect 14976 9432 14982 9444
rect 15074 9435 15132 9441
rect 15074 9432 15086 9435
rect 14976 9404 15086 9432
rect 14976 9392 14982 9404
rect 15074 9401 15086 9404
rect 15120 9401 15132 9435
rect 15074 9395 15132 9401
rect 8754 9364 8760 9376
rect 7984 9336 8616 9364
rect 8715 9336 8760 9364
rect 7984 9324 7990 9336
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 9125 9367 9183 9373
rect 9125 9333 9137 9367
rect 9171 9364 9183 9367
rect 9398 9364 9404 9376
rect 9171 9336 9404 9364
rect 9171 9333 9183 9336
rect 9125 9327 9183 9333
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9582 9364 9588 9376
rect 9543 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 9824 9336 9965 9364
rect 9824 9324 9830 9336
rect 9953 9333 9965 9336
rect 9999 9333 10011 9367
rect 9953 9327 10011 9333
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 10594 9364 10600 9376
rect 10100 9336 10600 9364
rect 10100 9324 10106 9336
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 10836 9336 11529 9364
rect 10836 9324 10842 9336
rect 11517 9333 11529 9336
rect 11563 9333 11575 9367
rect 11517 9327 11575 9333
rect 11609 9367 11667 9373
rect 11609 9333 11621 9367
rect 11655 9364 11667 9367
rect 12250 9364 12256 9376
rect 11655 9336 12256 9364
rect 11655 9333 11667 9336
rect 11609 9327 11667 9333
rect 12250 9324 12256 9336
rect 12308 9324 12314 9376
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 12483 9336 13829 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 13817 9327 13875 9333
rect 1104 9274 16836 9296
rect 1104 9222 6246 9274
rect 6298 9222 6310 9274
rect 6362 9222 6374 9274
rect 6426 9222 6438 9274
rect 6490 9222 11510 9274
rect 11562 9222 11574 9274
rect 11626 9222 11638 9274
rect 11690 9222 11702 9274
rect 11754 9222 16836 9274
rect 1104 9200 16836 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 3421 9163 3479 9169
rect 3421 9160 3433 9163
rect 1995 9132 3433 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 3421 9129 3433 9132
rect 3467 9129 3479 9163
rect 3421 9123 3479 9129
rect 3510 9120 3516 9172
rect 3568 9160 3574 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 3568 9132 4077 9160
rect 3568 9120 3574 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 4433 9163 4491 9169
rect 4433 9160 4445 9163
rect 4212 9132 4445 9160
rect 4212 9120 4218 9132
rect 4433 9129 4445 9132
rect 4479 9129 4491 9163
rect 4433 9123 4491 9129
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 4890 9160 4896 9172
rect 4571 9132 4896 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 5810 9160 5816 9172
rect 5184 9132 5816 9160
rect 2130 9052 2136 9104
rect 2188 9092 2194 9104
rect 4798 9092 4804 9104
rect 2188 9064 4804 9092
rect 2188 9052 2194 9064
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 8993 2375 9027
rect 2317 8987 2375 8993
rect 2409 9027 2467 9033
rect 2409 8993 2421 9027
rect 2455 9024 2467 9027
rect 2682 9024 2688 9036
rect 2455 8996 2688 9024
rect 2455 8993 2467 8996
rect 2409 8987 2467 8993
rect 2332 8956 2360 8987
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 3234 8984 3240 9036
rect 3292 9024 3298 9036
rect 3329 9027 3387 9033
rect 3329 9024 3341 9027
rect 3292 8996 3341 9024
rect 3292 8984 3298 8996
rect 3329 8993 3341 8996
rect 3375 8993 3387 9027
rect 3694 9024 3700 9036
rect 3329 8987 3387 8993
rect 3427 8996 3700 9024
rect 2498 8956 2504 8968
rect 2332 8928 2504 8956
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 3427 8956 3455 8996
rect 3694 8984 3700 8996
rect 3752 8984 3758 9036
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4212 8996 5120 9024
rect 4212 8984 4218 8996
rect 2639 8928 3455 8956
rect 3605 8959 3663 8965
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 3605 8925 3617 8959
rect 3651 8956 3663 8959
rect 4614 8956 4620 8968
rect 3651 8928 4620 8956
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 1670 8848 1676 8900
rect 1728 8888 1734 8900
rect 1728 8860 4200 8888
rect 1728 8848 1734 8860
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 2774 8820 2780 8832
rect 1627 8792 2780 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 2961 8823 3019 8829
rect 2961 8789 2973 8823
rect 3007 8820 3019 8823
rect 3234 8820 3240 8832
rect 3007 8792 3240 8820
rect 3007 8789 3019 8792
rect 2961 8783 3019 8789
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 4172 8820 4200 8860
rect 4338 8848 4344 8900
rect 4396 8888 4402 8900
rect 4522 8888 4528 8900
rect 4396 8860 4528 8888
rect 4396 8848 4402 8860
rect 4522 8848 4528 8860
rect 4580 8848 4586 8900
rect 5092 8888 5120 8996
rect 5184 8956 5212 9132
rect 5810 9120 5816 9132
rect 5868 9160 5874 9172
rect 6822 9160 6828 9172
rect 5868 9132 6828 9160
rect 5868 9120 5874 9132
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7190 9120 7196 9172
rect 7248 9160 7254 9172
rect 8662 9160 8668 9172
rect 7248 9132 8668 9160
rect 7248 9120 7254 9132
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 14918 9160 14924 9172
rect 9508 9132 13400 9160
rect 9508 9101 9536 9132
rect 9493 9095 9551 9101
rect 9493 9092 9505 9095
rect 5276 9064 9505 9092
rect 5276 9033 5304 9064
rect 9493 9061 9505 9064
rect 9539 9061 9551 9095
rect 9493 9055 9551 9061
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 9824 9064 11928 9092
rect 9824 9052 9830 9064
rect 5626 9033 5632 9036
rect 5261 9027 5319 9033
rect 5261 8993 5273 9027
rect 5307 8993 5319 9027
rect 5620 9024 5632 9033
rect 5587 8996 5632 9024
rect 5261 8987 5319 8993
rect 5620 8987 5632 8996
rect 5626 8984 5632 8987
rect 5684 8984 5690 9036
rect 7009 9027 7067 9033
rect 7009 8993 7021 9027
rect 7055 9024 7067 9027
rect 7190 9024 7196 9036
rect 7055 8996 7196 9024
rect 7055 8993 7067 8996
rect 7009 8987 7067 8993
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 7745 9027 7803 9033
rect 7745 8993 7757 9027
rect 7791 8993 7803 9027
rect 7745 8987 7803 8993
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 5184 8928 5365 8956
rect 5353 8925 5365 8928
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 6638 8916 6644 8968
rect 6696 8956 6702 8968
rect 7760 8956 7788 8987
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 9858 9024 9864 9036
rect 8076 8996 9864 9024
rect 8076 8984 8082 8996
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 9953 9027 10011 9033
rect 9953 8993 9965 9027
rect 9999 8993 10011 9027
rect 9953 8987 10011 8993
rect 6696 8928 7788 8956
rect 6696 8916 6702 8928
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8846 8956 8852 8968
rect 8352 8928 8852 8956
rect 8352 8916 8358 8928
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 6733 8891 6791 8897
rect 5092 8860 5212 8888
rect 4706 8820 4712 8832
rect 4172 8792 4712 8820
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 5074 8820 5080 8832
rect 5035 8792 5080 8820
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5184 8820 5212 8860
rect 6733 8857 6745 8891
rect 6779 8888 6791 8891
rect 7098 8888 7104 8900
rect 6779 8860 7104 8888
rect 6779 8857 6791 8860
rect 6733 8851 6791 8857
rect 7098 8848 7104 8860
rect 7156 8888 7162 8900
rect 7926 8888 7932 8900
rect 7156 8860 7932 8888
rect 7156 8848 7162 8860
rect 7926 8848 7932 8860
rect 7984 8848 7990 8900
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 9122 8888 9128 8900
rect 8260 8860 9128 8888
rect 8260 8848 8266 8860
rect 9122 8848 9128 8860
rect 9180 8888 9186 8900
rect 9968 8888 9996 8987
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 10870 9024 10876 9036
rect 10560 8996 10876 9024
rect 10560 8984 10566 8996
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 11790 9033 11796 9036
rect 11784 9024 11796 9033
rect 11164 8996 11796 9024
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 11164 8965 11192 8996
rect 11784 8987 11796 8996
rect 11790 8984 11796 8987
rect 11848 8984 11854 9036
rect 11900 9024 11928 9064
rect 11974 9052 11980 9104
rect 12032 9092 12038 9104
rect 12158 9092 12164 9104
rect 12032 9064 12164 9092
rect 12032 9052 12038 9064
rect 12158 9052 12164 9064
rect 12216 9092 12222 9104
rect 12989 9095 13047 9101
rect 12989 9092 13001 9095
rect 12216 9064 13001 9092
rect 12216 9052 12222 9064
rect 12989 9061 13001 9064
rect 13035 9061 13047 9095
rect 12989 9055 13047 9061
rect 13372 9033 13400 9132
rect 13464 9132 14924 9160
rect 13357 9027 13415 9033
rect 11900 8996 13308 9024
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10744 8928 10977 8956
rect 10744 8916 10750 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11517 8959 11575 8965
rect 11517 8956 11529 8959
rect 11296 8928 11529 8956
rect 11296 8916 11302 8928
rect 11517 8925 11529 8928
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13280 8956 13308 8996
rect 13357 8993 13369 9027
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 13464 8956 13492 9132
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 15654 9120 15660 9172
rect 15712 9120 15718 9172
rect 15749 9163 15807 9169
rect 15749 9129 15761 9163
rect 15795 9160 15807 9163
rect 16206 9160 16212 9172
rect 15795 9132 16212 9160
rect 15795 9129 15807 9132
rect 15749 9123 15807 9129
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 13998 9052 14004 9104
rect 14056 9092 14062 9104
rect 15194 9092 15200 9104
rect 14056 9064 15200 9092
rect 14056 9052 14062 9064
rect 15194 9052 15200 9064
rect 15252 9052 15258 9104
rect 15672 9092 15700 9120
rect 15838 9092 15844 9104
rect 15672 9064 15844 9092
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 13814 9033 13820 9036
rect 13808 9024 13820 9033
rect 13596 8996 13641 9024
rect 13775 8996 13820 9024
rect 13596 8984 13602 8996
rect 13808 8987 13820 8996
rect 13814 8984 13820 8987
rect 13872 8984 13878 9036
rect 14642 8984 14648 9036
rect 14700 9024 14706 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 14700 8996 15669 9024
rect 14700 8984 14706 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 15838 8956 15844 8968
rect 13035 8928 13216 8956
rect 13280 8928 13492 8956
rect 15799 8928 15844 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 9180 8860 9996 8888
rect 10137 8891 10195 8897
rect 9180 8848 9186 8860
rect 10137 8857 10149 8891
rect 10183 8888 10195 8891
rect 10870 8888 10876 8900
rect 10183 8860 10876 8888
rect 10183 8857 10195 8860
rect 10137 8851 10195 8857
rect 10870 8848 10876 8860
rect 10928 8848 10934 8900
rect 12526 8848 12532 8900
rect 12584 8888 12590 8900
rect 13188 8897 13216 8928
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 13173 8891 13231 8897
rect 12584 8860 13023 8888
rect 12584 8848 12590 8860
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 5184 8792 7205 8820
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 7193 8783 7251 8789
rect 10505 8823 10563 8829
rect 10505 8789 10517 8823
rect 10551 8820 10563 8823
rect 10686 8820 10692 8832
rect 10551 8792 10692 8820
rect 10551 8789 10563 8792
rect 10505 8783 10563 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 10962 8780 10968 8832
rect 11020 8820 11026 8832
rect 11238 8820 11244 8832
rect 11020 8792 11244 8820
rect 11020 8780 11026 8792
rect 11238 8780 11244 8792
rect 11296 8820 11302 8832
rect 12894 8820 12900 8832
rect 11296 8792 12900 8820
rect 11296 8780 11302 8792
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 12995 8820 13023 8860
rect 13173 8857 13185 8891
rect 13219 8857 13231 8891
rect 13173 8851 13231 8857
rect 15194 8848 15200 8900
rect 15252 8888 15258 8900
rect 16114 8888 16120 8900
rect 15252 8860 16120 8888
rect 15252 8848 15258 8860
rect 16114 8848 16120 8860
rect 16172 8848 16178 8900
rect 15289 8823 15347 8829
rect 15289 8820 15301 8823
rect 12995 8792 15301 8820
rect 15289 8789 15301 8792
rect 15335 8789 15347 8823
rect 15289 8783 15347 8789
rect 1104 8730 16836 8752
rect 1104 8678 3614 8730
rect 3666 8678 3678 8730
rect 3730 8678 3742 8730
rect 3794 8678 3806 8730
rect 3858 8678 8878 8730
rect 8930 8678 8942 8730
rect 8994 8678 9006 8730
rect 9058 8678 9070 8730
rect 9122 8678 14142 8730
rect 14194 8678 14206 8730
rect 14258 8678 14270 8730
rect 14322 8678 14334 8730
rect 14386 8678 16836 8730
rect 1104 8656 16836 8678
rect 4614 8616 4620 8628
rect 2424 8588 4620 8616
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1486 8412 1492 8424
rect 1443 8384 1492 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1486 8372 1492 8384
rect 1544 8372 1550 8424
rect 1664 8415 1722 8421
rect 1664 8381 1676 8415
rect 1710 8412 1722 8415
rect 2424 8412 2452 8588
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9582 8616 9588 8628
rect 9355 8588 9588 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 10318 8616 10324 8628
rect 10279 8588 10324 8616
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 14369 8619 14427 8625
rect 14369 8616 14381 8619
rect 10428 8588 14381 8616
rect 2777 8551 2835 8557
rect 2777 8517 2789 8551
rect 2823 8548 2835 8551
rect 2823 8520 3740 8548
rect 2823 8517 2835 8520
rect 2777 8511 2835 8517
rect 3234 8440 3240 8492
rect 3292 8480 3298 8492
rect 3712 8489 3740 8520
rect 4246 8508 4252 8560
rect 4304 8508 4310 8560
rect 5626 8508 5632 8560
rect 5684 8548 5690 8560
rect 5813 8551 5871 8557
rect 5813 8548 5825 8551
rect 5684 8520 5825 8548
rect 5684 8508 5690 8520
rect 5813 8517 5825 8520
rect 5859 8548 5871 8551
rect 7098 8548 7104 8560
rect 5859 8520 7104 8548
rect 5859 8517 5871 8520
rect 5813 8511 5871 8517
rect 7098 8508 7104 8520
rect 7156 8508 7162 8560
rect 10428 8548 10456 8588
rect 14369 8585 14381 8588
rect 14415 8585 14427 8619
rect 14369 8579 14427 8585
rect 15381 8551 15439 8557
rect 15381 8548 15393 8551
rect 9784 8520 10456 8548
rect 10520 8520 12296 8548
rect 3513 8483 3571 8489
rect 3513 8480 3525 8483
rect 3292 8452 3525 8480
rect 3292 8440 3298 8452
rect 3513 8449 3525 8452
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8480 3755 8483
rect 3786 8480 3792 8492
rect 3743 8452 3792 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 4264 8480 4292 8508
rect 4264 8452 4384 8480
rect 3418 8412 3424 8424
rect 1710 8384 2452 8412
rect 3379 8384 3424 8412
rect 1710 8381 1722 8384
rect 1664 8375 1722 8381
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 4065 8415 4123 8421
rect 4065 8381 4077 8415
rect 4111 8412 4123 8415
rect 4246 8412 4252 8424
rect 4111 8384 4252 8412
rect 4111 8381 4123 8384
rect 4065 8375 4123 8381
rect 4246 8372 4252 8384
rect 4304 8372 4310 8424
rect 1762 8304 1768 8356
rect 1820 8344 1826 8356
rect 3142 8344 3148 8356
rect 1820 8316 3148 8344
rect 1820 8304 1826 8316
rect 3142 8304 3148 8316
rect 3200 8304 3206 8356
rect 3510 8304 3516 8356
rect 3568 8344 3574 8356
rect 3568 8316 4292 8344
rect 3568 8304 3574 8316
rect 3050 8276 3056 8288
rect 3011 8248 3056 8276
rect 3050 8236 3056 8248
rect 3108 8236 3114 8288
rect 4264 8285 4292 8316
rect 4249 8279 4307 8285
rect 4249 8245 4261 8279
rect 4295 8245 4307 8279
rect 4356 8276 4384 8452
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 9784 8489 9812 8520
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 6880 8452 7573 8480
rect 6880 8440 6886 8452
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 9769 8483 9827 8489
rect 9769 8449 9781 8483
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 9953 8483 10011 8489
rect 9953 8449 9965 8483
rect 9999 8480 10011 8483
rect 10042 8480 10048 8492
rect 9999 8452 10048 8480
rect 9999 8449 10011 8452
rect 9953 8443 10011 8449
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4522 8412 4528 8424
rect 4479 8384 4528 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 8662 8412 8668 8424
rect 7760 8384 8668 8412
rect 4706 8353 4712 8356
rect 4700 8344 4712 8353
rect 4667 8316 4712 8344
rect 4700 8307 4712 8316
rect 4706 8304 4712 8307
rect 4764 8304 4770 8356
rect 4890 8304 4896 8356
rect 4948 8344 4954 8356
rect 5902 8344 5908 8356
rect 4948 8316 5908 8344
rect 4948 8304 4954 8316
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 6181 8347 6239 8353
rect 6181 8313 6193 8347
rect 6227 8344 6239 8347
rect 6273 8347 6331 8353
rect 6273 8344 6285 8347
rect 6227 8316 6285 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 6273 8313 6285 8316
rect 6319 8344 6331 8347
rect 7285 8347 7343 8353
rect 6319 8316 7236 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 6638 8276 6644 8288
rect 4356 8248 6644 8276
rect 4249 8239 4307 8245
rect 6638 8236 6644 8248
rect 6696 8236 6702 8288
rect 7208 8276 7236 8316
rect 7285 8313 7297 8347
rect 7331 8344 7343 8347
rect 7760 8344 7788 8384
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 10520 8412 10548 8520
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 11238 8480 11244 8492
rect 11011 8452 11244 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11882 8440 11888 8492
rect 11940 8480 11946 8492
rect 11940 8452 11985 8480
rect 11940 8440 11946 8452
rect 10686 8412 10692 8424
rect 9723 8384 10548 8412
rect 10647 8384 10692 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11422 8412 11428 8424
rect 10827 8384 11428 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 11422 8372 11428 8384
rect 11480 8372 11486 8424
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8412 11759 8415
rect 12158 8412 12164 8424
rect 11747 8384 12164 8412
rect 11747 8381 11759 8384
rect 11701 8375 11759 8381
rect 12158 8372 12164 8384
rect 12216 8372 12222 8424
rect 12268 8412 12296 8520
rect 13740 8520 15393 8548
rect 12710 8480 12716 8492
rect 12671 8452 12716 8480
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 13740 8412 13768 8520
rect 15381 8517 15393 8520
rect 15427 8517 15439 8551
rect 15381 8511 15439 8517
rect 14921 8483 14979 8489
rect 14921 8480 14933 8483
rect 14016 8452 14933 8480
rect 14016 8424 14044 8452
rect 14921 8449 14933 8452
rect 14967 8480 14979 8483
rect 15010 8480 15016 8492
rect 14967 8452 15016 8480
rect 14967 8449 14979 8452
rect 14921 8443 14979 8449
rect 15010 8440 15016 8452
rect 15068 8480 15074 8492
rect 15838 8480 15844 8492
rect 15068 8452 15844 8480
rect 15068 8440 15074 8452
rect 15838 8440 15844 8452
rect 15896 8480 15902 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15896 8452 15945 8480
rect 15896 8440 15902 8452
rect 15933 8449 15945 8452
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 12268 8384 13768 8412
rect 13998 8372 14004 8424
rect 14056 8372 14062 8424
rect 14090 8372 14096 8424
rect 14148 8412 14154 8424
rect 14148 8384 14228 8412
rect 14148 8372 14154 8384
rect 7834 8353 7840 8356
rect 7331 8316 7788 8344
rect 7331 8313 7343 8316
rect 7285 8307 7343 8313
rect 7828 8307 7840 8353
rect 7892 8344 7898 8356
rect 9858 8344 9864 8356
rect 7892 8316 7928 8344
rect 8036 8316 9864 8344
rect 7834 8304 7840 8307
rect 7892 8304 7898 8316
rect 8036 8276 8064 8316
rect 9858 8304 9864 8316
rect 9916 8304 9922 8356
rect 11793 8347 11851 8353
rect 11793 8313 11805 8347
rect 11839 8344 11851 8347
rect 12980 8347 13038 8353
rect 11839 8316 12940 8344
rect 11839 8313 11851 8316
rect 11793 8307 11851 8313
rect 7208 8248 8064 8276
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 8941 8279 8999 8285
rect 8941 8276 8953 8279
rect 8628 8248 8953 8276
rect 8628 8236 8634 8248
rect 8941 8245 8953 8248
rect 8987 8245 8999 8279
rect 8941 8239 8999 8245
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 9950 8276 9956 8288
rect 9088 8248 9956 8276
rect 9088 8236 9094 8248
rect 9950 8236 9956 8248
rect 10008 8236 10014 8288
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10318 8276 10324 8288
rect 10192 8248 10324 8276
rect 10192 8236 10198 8248
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 11333 8279 11391 8285
rect 11333 8245 11345 8279
rect 11379 8276 11391 8279
rect 12250 8276 12256 8288
rect 11379 8248 12256 8276
rect 11379 8245 11391 8248
rect 11333 8239 11391 8245
rect 12250 8236 12256 8248
rect 12308 8236 12314 8288
rect 12912 8276 12940 8316
rect 12980 8313 12992 8347
rect 13026 8344 13038 8347
rect 13026 8316 13768 8344
rect 13026 8313 13038 8316
rect 12980 8307 13038 8313
rect 13630 8276 13636 8288
rect 12912 8248 13636 8276
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 13740 8276 13768 8316
rect 13814 8304 13820 8356
rect 13872 8344 13878 8356
rect 14200 8344 14228 8384
rect 14458 8372 14464 8424
rect 14516 8412 14522 8424
rect 14737 8415 14795 8421
rect 14737 8412 14749 8415
rect 14516 8384 14749 8412
rect 14516 8372 14522 8384
rect 14737 8381 14749 8384
rect 14783 8381 14795 8415
rect 14737 8375 14795 8381
rect 14829 8415 14887 8421
rect 14829 8381 14841 8415
rect 14875 8412 14887 8415
rect 15286 8412 15292 8424
rect 14875 8384 15292 8412
rect 14875 8381 14887 8384
rect 14829 8375 14887 8381
rect 15286 8372 15292 8384
rect 15344 8372 15350 8424
rect 15470 8372 15476 8424
rect 15528 8412 15534 8424
rect 15528 8384 15884 8412
rect 15528 8372 15534 8384
rect 15856 8353 15884 8384
rect 15749 8347 15807 8353
rect 15749 8344 15761 8347
rect 13872 8316 14136 8344
rect 14200 8316 15761 8344
rect 13872 8304 13878 8316
rect 13998 8276 14004 8288
rect 13740 8248 14004 8276
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 14108 8285 14136 8316
rect 15749 8313 15761 8316
rect 15795 8313 15807 8347
rect 15749 8307 15807 8313
rect 15841 8347 15899 8353
rect 15841 8313 15853 8347
rect 15887 8313 15899 8347
rect 15841 8307 15899 8313
rect 14093 8279 14151 8285
rect 14093 8245 14105 8279
rect 14139 8276 14151 8279
rect 14139 8248 14173 8276
rect 14139 8245 14151 8248
rect 14093 8239 14151 8245
rect 1104 8186 16836 8208
rect 1104 8134 6246 8186
rect 6298 8134 6310 8186
rect 6362 8134 6374 8186
rect 6426 8134 6438 8186
rect 6490 8134 11510 8186
rect 11562 8134 11574 8186
rect 11626 8134 11638 8186
rect 11690 8134 11702 8186
rect 11754 8134 16836 8186
rect 1104 8112 16836 8134
rect 2222 8032 2228 8084
rect 2280 8072 2286 8084
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 2280 8044 2329 8072
rect 2280 8032 2286 8044
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 2317 8035 2375 8041
rect 2961 8075 3019 8081
rect 2961 8041 2973 8075
rect 3007 8072 3019 8075
rect 7009 8075 7067 8081
rect 7009 8072 7021 8075
rect 3007 8044 7021 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 7009 8041 7021 8044
rect 7055 8041 7067 8075
rect 7009 8035 7067 8041
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 7377 8075 7435 8081
rect 7377 8072 7389 8075
rect 7340 8044 7389 8072
rect 7340 8032 7346 8044
rect 7377 8041 7389 8044
rect 7423 8041 7435 8075
rect 8294 8072 8300 8084
rect 7377 8035 7435 8041
rect 7760 8044 8156 8072
rect 8255 8044 8300 8072
rect 2038 7964 2044 8016
rect 2096 8004 2102 8016
rect 2409 8007 2467 8013
rect 2409 8004 2421 8007
rect 2096 7976 2421 8004
rect 2096 7964 2102 7976
rect 2409 7973 2421 7976
rect 2455 7973 2467 8007
rect 2409 7967 2467 7973
rect 4982 7964 4988 8016
rect 5040 8004 5046 8016
rect 5138 8007 5196 8013
rect 5138 8004 5150 8007
rect 5040 7976 5150 8004
rect 5040 7964 5046 7976
rect 5138 7973 5150 7976
rect 5184 7973 5196 8007
rect 5718 8004 5724 8016
rect 5138 7967 5196 7973
rect 5368 7976 5724 8004
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1670 7936 1676 7948
rect 1443 7908 1676 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 3326 7936 3332 7948
rect 3287 7908 3332 7936
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 5368 7936 5396 7976
rect 5718 7964 5724 7976
rect 5776 7964 5782 8016
rect 6638 7964 6644 8016
rect 6696 8004 6702 8016
rect 7760 8013 7788 8044
rect 7745 8007 7803 8013
rect 7745 8004 7757 8007
rect 6696 7976 7757 8004
rect 6696 7964 6702 7976
rect 7745 7973 7757 7976
rect 7791 7973 7803 8007
rect 8128 8004 8156 8044
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 8665 8075 8723 8081
rect 8665 8041 8677 8075
rect 8711 8072 8723 8075
rect 12526 8072 12532 8084
rect 8711 8044 9628 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 8478 8004 8484 8016
rect 8128 7976 8484 8004
rect 7745 7967 7803 7973
rect 8478 7964 8484 7976
rect 8536 7964 8542 8016
rect 9600 8004 9628 8044
rect 9968 8044 12532 8072
rect 9968 8004 9996 8044
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 12805 8075 12863 8081
rect 12805 8072 12817 8075
rect 12676 8044 12817 8072
rect 12676 8032 12682 8044
rect 12805 8041 12817 8044
rect 12851 8041 12863 8075
rect 12805 8035 12863 8041
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 13412 8044 13461 8072
rect 13412 8032 13418 8044
rect 13449 8041 13461 8044
rect 13495 8041 13507 8075
rect 13449 8035 13507 8041
rect 13722 8032 13728 8084
rect 13780 8072 13786 8084
rect 14458 8072 14464 8084
rect 13780 8044 14464 8072
rect 13780 8032 13786 8044
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 15289 8075 15347 8081
rect 15289 8041 15301 8075
rect 15335 8041 15347 8075
rect 15289 8035 15347 8041
rect 9600 7976 9996 8004
rect 10045 8007 10103 8013
rect 10045 7973 10057 8007
rect 10091 8004 10103 8007
rect 10226 8004 10232 8016
rect 10091 7976 10232 8004
rect 10091 7973 10103 7976
rect 10045 7967 10103 7973
rect 10226 7964 10232 7976
rect 10284 7964 10290 8016
rect 10318 7964 10324 8016
rect 10376 7964 10382 8016
rect 10686 7964 10692 8016
rect 10744 8004 10750 8016
rect 15304 8004 15332 8035
rect 10744 7976 15332 8004
rect 10744 7964 10750 7976
rect 4111 7908 5396 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6880 7908 6929 7936
rect 6880 7896 6886 7908
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 8294 7936 8300 7948
rect 7883 7908 8300 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7936 10195 7939
rect 10336 7936 10364 7964
rect 10183 7908 10364 7936
rect 10772 7939 10830 7945
rect 10183 7905 10195 7908
rect 10137 7899 10195 7905
rect 10772 7905 10784 7939
rect 10818 7936 10830 7939
rect 11882 7936 11888 7948
rect 10818 7908 11888 7936
rect 10818 7905 10830 7908
rect 10772 7899 10830 7905
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2958 7868 2964 7880
rect 2639 7840 2964 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 4706 7868 4712 7880
rect 3651 7840 4712 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 3436 7800 3464 7831
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 4890 7868 4896 7880
rect 4851 7840 4896 7868
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 7098 7868 7104 7880
rect 7059 7840 7104 7868
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 7984 7840 8029 7868
rect 7984 7828 7990 7840
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 8536 7840 8769 7868
rect 8536 7828 8542 7840
rect 8757 7837 8769 7840
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7868 8999 7871
rect 9030 7868 9036 7880
rect 8987 7840 9036 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 4798 7800 4804 7812
rect 3436 7772 4804 7800
rect 4798 7760 4804 7772
rect 4856 7760 4862 7812
rect 5994 7760 6000 7812
rect 6052 7800 6058 7812
rect 6549 7803 6607 7809
rect 6549 7800 6561 7803
rect 6052 7772 6561 7800
rect 6052 7760 6058 7772
rect 6549 7769 6561 7772
rect 6595 7769 6607 7803
rect 6549 7763 6607 7769
rect 1394 7692 1400 7744
rect 1452 7732 1458 7744
rect 1581 7735 1639 7741
rect 1581 7732 1593 7735
rect 1452 7704 1593 7732
rect 1452 7692 1458 7704
rect 1581 7701 1593 7704
rect 1627 7701 1639 7735
rect 1946 7732 1952 7744
rect 1907 7704 1952 7732
rect 1581 7695 1639 7701
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 3142 7692 3148 7744
rect 3200 7732 3206 7744
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 3200 7704 4261 7732
rect 3200 7692 3206 7704
rect 4249 7701 4261 7704
rect 4295 7701 4307 7735
rect 4249 7695 4307 7701
rect 4706 7692 4712 7744
rect 4764 7732 4770 7744
rect 6270 7732 6276 7744
rect 4764 7704 6276 7732
rect 4764 7692 4770 7704
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 9309 7735 9367 7741
rect 9309 7732 9321 7735
rect 8260 7704 9321 7732
rect 8260 7692 8266 7704
rect 9309 7701 9321 7704
rect 9355 7701 9367 7735
rect 9508 7732 9536 7899
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 13814 7936 13820 7948
rect 13775 7908 13820 7936
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 13909 7939 13967 7945
rect 13909 7905 13921 7939
rect 13955 7936 13967 7939
rect 14090 7936 14096 7948
rect 13955 7908 14096 7936
rect 13955 7905 13967 7908
rect 13909 7899 13967 7905
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 14642 7936 14648 7948
rect 14603 7908 14648 7936
rect 14642 7896 14648 7908
rect 14700 7936 14706 7948
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 14700 7908 15669 7936
rect 14700 7896 14706 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 16298 7936 16304 7948
rect 15657 7899 15715 7905
rect 15764 7908 16304 7936
rect 9582 7828 9588 7880
rect 9640 7868 9646 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 9640 7840 10241 7868
rect 9640 7828 9646 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 10376 7840 10517 7868
rect 10376 7828 10382 7840
rect 10505 7837 10517 7840
rect 10551 7837 10563 7871
rect 12894 7868 12900 7880
rect 12855 7840 12900 7868
rect 10505 7831 10563 7837
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7868 13139 7871
rect 13722 7868 13728 7880
rect 13127 7840 13728 7868
rect 13127 7837 13139 7840
rect 13081 7831 13139 7837
rect 13722 7828 13728 7840
rect 13780 7868 13786 7880
rect 15764 7877 15792 7908
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 14001 7871 14059 7877
rect 14001 7868 14013 7871
rect 13780 7840 14013 7868
rect 13780 7828 13786 7840
rect 14001 7837 14013 7840
rect 14047 7837 14059 7871
rect 14001 7831 14059 7837
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 9674 7760 9680 7812
rect 9732 7800 9738 7812
rect 9732 7772 9777 7800
rect 9732 7760 9738 7772
rect 11790 7760 11796 7812
rect 11848 7800 11854 7812
rect 11885 7803 11943 7809
rect 11885 7800 11897 7803
rect 11848 7772 11897 7800
rect 11848 7760 11854 7772
rect 11885 7769 11897 7772
rect 11931 7769 11943 7803
rect 11885 7763 11943 7769
rect 11992 7772 12664 7800
rect 10226 7732 10232 7744
rect 9508 7704 10232 7732
rect 9309 7695 9367 7701
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 11698 7692 11704 7744
rect 11756 7732 11762 7744
rect 11992 7732 12020 7772
rect 11756 7704 12020 7732
rect 12437 7735 12495 7741
rect 11756 7692 11762 7704
rect 12437 7701 12449 7735
rect 12483 7732 12495 7735
rect 12526 7732 12532 7744
rect 12483 7704 12532 7732
rect 12483 7701 12495 7704
rect 12437 7695 12495 7701
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 12636 7732 12664 7772
rect 15102 7760 15108 7812
rect 15160 7800 15166 7812
rect 15764 7800 15792 7831
rect 15838 7828 15844 7880
rect 15896 7868 15902 7880
rect 15896 7840 15941 7868
rect 15896 7828 15902 7840
rect 15160 7772 15792 7800
rect 15160 7760 15166 7772
rect 13078 7732 13084 7744
rect 12636 7704 13084 7732
rect 13078 7692 13084 7704
rect 13136 7732 13142 7744
rect 13814 7732 13820 7744
rect 13136 7704 13820 7732
rect 13136 7692 13142 7704
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 14829 7735 14887 7741
rect 14829 7701 14841 7735
rect 14875 7732 14887 7735
rect 15286 7732 15292 7744
rect 14875 7704 15292 7732
rect 14875 7701 14887 7704
rect 14829 7695 14887 7701
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 1104 7642 16836 7664
rect 1104 7590 3614 7642
rect 3666 7590 3678 7642
rect 3730 7590 3742 7642
rect 3794 7590 3806 7642
rect 3858 7590 8878 7642
rect 8930 7590 8942 7642
rect 8994 7590 9006 7642
rect 9058 7590 9070 7642
rect 9122 7590 14142 7642
rect 14194 7590 14206 7642
rect 14258 7590 14270 7642
rect 14322 7590 14334 7642
rect 14386 7590 16836 7642
rect 1104 7568 16836 7590
rect 1946 7488 1952 7540
rect 2004 7528 2010 7540
rect 2004 7500 4476 7528
rect 2004 7488 2010 7500
rect 2958 7460 2964 7472
rect 2871 7432 2964 7460
rect 2958 7420 2964 7432
rect 3016 7460 3022 7472
rect 4448 7460 4476 7500
rect 4798 7488 4804 7540
rect 4856 7528 4862 7540
rect 6546 7528 6552 7540
rect 4856 7500 6552 7528
rect 4856 7488 4862 7500
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 6822 7528 6828 7540
rect 6783 7500 6828 7528
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 11238 7528 11244 7540
rect 8312 7500 11244 7528
rect 6086 7460 6092 7472
rect 3016 7432 3832 7460
rect 4448 7432 6092 7460
rect 3016 7420 3022 7432
rect 1486 7352 1492 7404
rect 1544 7392 1550 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 1544 7364 1593 7392
rect 1544 7352 1550 7364
rect 1581 7361 1593 7364
rect 1627 7361 1639 7395
rect 1581 7355 1639 7361
rect 3050 7352 3056 7404
rect 3108 7392 3114 7404
rect 3804 7401 3832 7432
rect 6086 7420 6092 7432
rect 6144 7420 6150 7472
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 3108 7364 3709 7392
rect 3108 7352 3114 7364
rect 3697 7361 3709 7364
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4801 7395 4859 7401
rect 4801 7392 4813 7395
rect 4028 7364 4813 7392
rect 4028 7352 4034 7364
rect 4801 7361 4813 7364
rect 4847 7361 4859 7395
rect 5718 7392 5724 7404
rect 5679 7364 5724 7392
rect 4801 7355 4859 7361
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 1848 7327 1906 7333
rect 1848 7293 1860 7327
rect 1894 7324 1906 7327
rect 3988 7324 4016 7352
rect 1894 7296 4016 7324
rect 1894 7293 1906 7296
rect 1848 7287 1906 7293
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 5828 7324 5856 7355
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 6328 7364 7389 7392
rect 6328 7352 6334 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8312 7392 8340 7500
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 11701 7531 11759 7537
rect 11701 7497 11713 7531
rect 11747 7528 11759 7531
rect 11882 7528 11888 7540
rect 11747 7500 11888 7528
rect 11747 7497 11759 7500
rect 11701 7491 11759 7497
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12989 7531 13047 7537
rect 12989 7497 13001 7531
rect 13035 7528 13047 7531
rect 13998 7528 14004 7540
rect 13035 7500 14004 7528
rect 13035 7497 13047 7500
rect 12989 7491 13047 7497
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 15381 7531 15439 7537
rect 15381 7528 15393 7531
rect 14516 7500 15393 7528
rect 14516 7488 14522 7500
rect 15381 7497 15393 7500
rect 15427 7497 15439 7531
rect 15381 7491 15439 7497
rect 13357 7463 13415 7469
rect 13357 7429 13369 7463
rect 13403 7460 13415 7463
rect 13403 7432 15884 7460
rect 13403 7429 13415 7432
rect 13357 7423 13415 7429
rect 9858 7392 9864 7404
rect 7883 7364 8340 7392
rect 9416 7364 9864 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 7282 7324 7288 7336
rect 4764 7296 5856 7324
rect 7243 7296 7288 7324
rect 4764 7284 4770 7296
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 7742 7284 7748 7336
rect 7800 7324 7806 7336
rect 7926 7324 7932 7336
rect 7800 7296 7932 7324
rect 7800 7284 7806 7296
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 8297 7327 8355 7333
rect 8297 7324 8309 7327
rect 8260 7296 8309 7324
rect 8260 7284 8266 7296
rect 8297 7293 8309 7296
rect 8343 7324 8355 7327
rect 9416 7324 9444 7364
rect 9858 7352 9864 7364
rect 9916 7392 9922 7404
rect 10318 7392 10324 7404
rect 9916 7364 10324 7392
rect 9916 7352 9922 7364
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 13722 7352 13728 7404
rect 13780 7392 13786 7404
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13780 7364 13921 7392
rect 13780 7352 13786 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7392 14887 7395
rect 14918 7392 14924 7404
rect 14875 7364 14924 7392
rect 14875 7361 14887 7364
rect 14829 7355 14887 7361
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7392 15071 7395
rect 15102 7392 15108 7404
rect 15059 7364 15108 7392
rect 15059 7361 15071 7364
rect 15013 7355 15071 7361
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 15856 7401 15884 7432
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7361 15899 7395
rect 15841 7355 15899 7361
rect 15930 7352 15936 7404
rect 15988 7392 15994 7404
rect 15988 7364 16033 7392
rect 15988 7352 15994 7364
rect 8343 7296 9444 7324
rect 8343 7293 8355 7296
rect 8297 7287 8355 7293
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 9548 7296 9965 7324
rect 9548 7284 9554 7296
rect 9953 7293 9965 7296
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 10588 7327 10646 7333
rect 10588 7293 10600 7327
rect 10634 7324 10646 7327
rect 12618 7324 12624 7336
rect 10634 7296 12624 7324
rect 10634 7293 10646 7296
rect 10588 7287 10646 7293
rect 2314 7216 2320 7268
rect 2372 7256 2378 7268
rect 2590 7256 2596 7268
rect 2372 7228 2596 7256
rect 2372 7216 2378 7228
rect 2590 7216 2596 7228
rect 2648 7216 2654 7268
rect 3605 7259 3663 7265
rect 3605 7225 3617 7259
rect 3651 7256 3663 7259
rect 3651 7228 4292 7256
rect 3651 7225 3663 7228
rect 3605 7219 3663 7225
rect 3142 7148 3148 7200
rect 3200 7188 3206 7200
rect 4264 7197 4292 7228
rect 6730 7216 6736 7268
rect 6788 7256 6794 7268
rect 8570 7265 8576 7268
rect 6788 7228 7328 7256
rect 6788 7216 6794 7228
rect 3237 7191 3295 7197
rect 3237 7188 3249 7191
rect 3200 7160 3249 7188
rect 3200 7148 3206 7160
rect 3237 7157 3249 7160
rect 3283 7157 3295 7191
rect 3237 7151 3295 7157
rect 4249 7191 4307 7197
rect 4249 7157 4261 7191
rect 4295 7157 4307 7191
rect 4249 7151 4307 7157
rect 4338 7148 4344 7200
rect 4396 7188 4402 7200
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 4396 7160 4629 7188
rect 4396 7148 4402 7160
rect 4617 7157 4629 7160
rect 4663 7157 4675 7191
rect 4617 7151 4675 7157
rect 4709 7191 4767 7197
rect 4709 7157 4721 7191
rect 4755 7188 4767 7191
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 4755 7160 5273 7188
rect 4755 7157 4767 7160
rect 4709 7151 4767 7157
rect 5261 7157 5273 7160
rect 5307 7157 5319 7191
rect 5626 7188 5632 7200
rect 5587 7160 5632 7188
rect 5261 7151 5319 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6273 7191 6331 7197
rect 6273 7157 6285 7191
rect 6319 7188 6331 7191
rect 6638 7188 6644 7200
rect 6319 7160 6644 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7300 7188 7328 7228
rect 8564 7219 8576 7265
rect 8628 7256 8634 7268
rect 9968 7256 9996 7287
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 11054 7256 11060 7268
rect 8628 7228 8664 7256
rect 9968 7228 11060 7256
rect 8570 7216 8576 7219
rect 8628 7216 8634 7228
rect 11054 7216 11060 7228
rect 11112 7216 11118 7268
rect 11238 7216 11244 7268
rect 11296 7256 11302 7268
rect 12820 7256 12848 7287
rect 13354 7284 13360 7336
rect 13412 7324 13418 7336
rect 15749 7327 15807 7333
rect 15749 7324 15761 7327
rect 13412 7296 15761 7324
rect 13412 7284 13418 7296
rect 15749 7293 15761 7296
rect 15795 7293 15807 7327
rect 15749 7287 15807 7293
rect 11296 7228 12848 7256
rect 13725 7259 13783 7265
rect 11296 7216 11302 7228
rect 13725 7225 13737 7259
rect 13771 7256 13783 7259
rect 13771 7228 14412 7256
rect 13771 7225 13783 7228
rect 13725 7219 13783 7225
rect 9582 7188 9588 7200
rect 7300 7160 9588 7188
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 9677 7191 9735 7197
rect 9677 7157 9689 7191
rect 9723 7188 9735 7191
rect 9766 7188 9772 7200
rect 9723 7160 9772 7188
rect 9723 7157 9735 7160
rect 9677 7151 9735 7157
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 10137 7191 10195 7197
rect 10137 7157 10149 7191
rect 10183 7188 10195 7191
rect 13630 7188 13636 7200
rect 10183 7160 13636 7188
rect 10183 7157 10195 7160
rect 10137 7151 10195 7157
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 13817 7191 13875 7197
rect 13817 7157 13829 7191
rect 13863 7188 13875 7191
rect 14182 7188 14188 7200
rect 13863 7160 14188 7188
rect 13863 7157 13875 7160
rect 13817 7151 13875 7157
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 14384 7197 14412 7228
rect 14369 7191 14427 7197
rect 14369 7157 14381 7191
rect 14415 7157 14427 7191
rect 14369 7151 14427 7157
rect 14642 7148 14648 7200
rect 14700 7188 14706 7200
rect 14737 7191 14795 7197
rect 14737 7188 14749 7191
rect 14700 7160 14749 7188
rect 14700 7148 14706 7160
rect 14737 7157 14749 7160
rect 14783 7188 14795 7191
rect 15470 7188 15476 7200
rect 14783 7160 15476 7188
rect 14783 7157 14795 7160
rect 14737 7151 14795 7157
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 1104 7098 16836 7120
rect 1104 7046 6246 7098
rect 6298 7046 6310 7098
rect 6362 7046 6374 7098
rect 6426 7046 6438 7098
rect 6490 7046 11510 7098
rect 11562 7046 11574 7098
rect 11626 7046 11638 7098
rect 11690 7046 11702 7098
rect 11754 7046 16836 7098
rect 1104 7024 16836 7046
rect 4433 6987 4491 6993
rect 4433 6953 4445 6987
rect 4479 6984 4491 6987
rect 6638 6984 6644 6996
rect 4479 6956 6644 6984
rect 4479 6953 4491 6956
rect 4433 6947 4491 6953
rect 6638 6944 6644 6956
rect 6696 6944 6702 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 8478 6984 8484 6996
rect 7340 6956 8484 6984
rect 7340 6944 7346 6956
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 11333 6987 11391 6993
rect 11333 6953 11345 6987
rect 11379 6984 11391 6987
rect 12989 6987 13047 6993
rect 11379 6956 12572 6984
rect 11379 6953 11391 6956
rect 11333 6947 11391 6953
rect 5276 6888 5672 6916
rect 1489 6851 1547 6857
rect 1489 6817 1501 6851
rect 1535 6817 1547 6851
rect 1489 6811 1547 6817
rect 1504 6712 1532 6811
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 2409 6851 2467 6857
rect 2409 6848 2421 6851
rect 1636 6820 2421 6848
rect 1636 6808 1642 6820
rect 2409 6817 2421 6820
rect 2455 6817 2467 6851
rect 2409 6811 2467 6817
rect 3053 6851 3111 6857
rect 3053 6817 3065 6851
rect 3099 6848 3111 6851
rect 3418 6848 3424 6860
rect 3099 6820 3424 6848
rect 3099 6817 3111 6820
rect 3053 6811 3111 6817
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 5074 6848 5080 6860
rect 3927 6820 5080 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 1854 6740 1860 6792
rect 1912 6780 1918 6792
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 1912 6752 2513 6780
rect 1912 6740 1918 6752
rect 2501 6749 2513 6752
rect 2547 6749 2559 6783
rect 2501 6743 2559 6749
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 2648 6752 2693 6780
rect 2648 6740 2654 6752
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3234 6780 3240 6792
rect 2832 6752 3240 6780
rect 2832 6740 2838 6752
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 4525 6783 4583 6789
rect 3988 6752 4476 6780
rect 3988 6712 4016 6752
rect 1504 6684 4016 6712
rect 4065 6715 4123 6721
rect 4065 6681 4077 6715
rect 4111 6712 4123 6715
rect 4338 6712 4344 6724
rect 4111 6684 4344 6712
rect 4111 6681 4123 6684
rect 4065 6675 4123 6681
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 842 6604 848 6656
rect 900 6644 906 6656
rect 1673 6647 1731 6653
rect 1673 6644 1685 6647
rect 900 6616 1685 6644
rect 900 6604 906 6616
rect 1673 6613 1685 6616
rect 1719 6613 1731 6647
rect 2038 6644 2044 6656
rect 1999 6616 2044 6644
rect 1673 6607 1731 6613
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 3237 6647 3295 6653
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 3418 6644 3424 6656
rect 3283 6616 3424 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3697 6647 3755 6653
rect 3697 6613 3709 6647
rect 3743 6644 3755 6647
rect 3970 6644 3976 6656
rect 3743 6616 3976 6644
rect 3743 6613 3755 6616
rect 3697 6607 3755 6613
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4448 6644 4476 6752
rect 4525 6749 4537 6783
rect 4571 6749 4583 6783
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 4525 6743 4583 6749
rect 4540 6712 4568 6743
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5276 6789 5304 6888
rect 5534 6857 5540 6860
rect 5528 6848 5540 6857
rect 5495 6820 5540 6848
rect 5528 6811 5540 6820
rect 5534 6808 5540 6811
rect 5592 6808 5598 6860
rect 5644 6848 5672 6888
rect 5718 6876 5724 6928
rect 5776 6916 5782 6928
rect 6178 6916 6184 6928
rect 5776 6888 6184 6916
rect 5776 6876 5782 6888
rect 6178 6876 6184 6888
rect 6236 6916 6242 6928
rect 8754 6916 8760 6928
rect 6236 6888 7604 6916
rect 8715 6888 8760 6916
rect 6236 6876 6242 6888
rect 6917 6851 6975 6857
rect 6917 6848 6929 6851
rect 5644 6820 6929 6848
rect 6917 6817 6929 6820
rect 6963 6817 6975 6851
rect 6917 6811 6975 6817
rect 7184 6851 7242 6857
rect 7184 6817 7196 6851
rect 7230 6848 7242 6851
rect 7466 6848 7472 6860
rect 7230 6820 7472 6848
rect 7230 6817 7242 6820
rect 7184 6811 7242 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7576 6848 7604 6888
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 9214 6876 9220 6928
rect 9272 6916 9278 6928
rect 9490 6916 9496 6928
rect 9272 6888 9496 6916
rect 9272 6876 9278 6888
rect 9490 6876 9496 6888
rect 9548 6876 9554 6928
rect 10226 6876 10232 6928
rect 10284 6916 10290 6928
rect 11348 6916 11376 6947
rect 11974 6916 11980 6928
rect 10284 6888 11376 6916
rect 11808 6888 11980 6916
rect 10284 6876 10290 6888
rect 7576 6820 8524 6848
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 4948 6752 5273 6780
rect 4948 6740 4954 6752
rect 5261 6749 5273 6752
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 4614 6712 4620 6724
rect 4540 6684 4620 6712
rect 4614 6672 4620 6684
rect 4672 6672 4678 6724
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 8389 6715 8447 6721
rect 8389 6712 8401 6715
rect 8168 6684 8401 6712
rect 8168 6672 8174 6684
rect 8389 6681 8401 6684
rect 8435 6681 8447 6715
rect 8496 6712 8524 6820
rect 8570 6808 8576 6860
rect 8628 6848 8634 6860
rect 8628 6820 8984 6848
rect 8628 6808 8634 6820
rect 8846 6780 8852 6792
rect 8807 6752 8852 6780
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 8956 6789 8984 6820
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 9933 6851 9991 6857
rect 9933 6848 9945 6851
rect 9824 6820 9945 6848
rect 9824 6808 9830 6820
rect 9933 6817 9945 6820
rect 9979 6817 9991 6851
rect 9933 6811 9991 6817
rect 11517 6851 11575 6857
rect 11517 6817 11529 6851
rect 11563 6848 11575 6851
rect 11808 6848 11836 6888
rect 11974 6876 11980 6888
rect 12032 6876 12038 6928
rect 11563 6820 11836 6848
rect 11876 6851 11934 6857
rect 11563 6817 11575 6820
rect 11517 6811 11575 6817
rect 11876 6817 11888 6851
rect 11922 6848 11934 6851
rect 12434 6848 12440 6860
rect 11922 6820 12440 6848
rect 11922 6817 11934 6820
rect 11876 6811 11934 6817
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 12544 6848 12572 6956
rect 12989 6953 13001 6987
rect 13035 6953 13047 6987
rect 14182 6984 14188 6996
rect 14143 6956 14188 6984
rect 12989 6947 13047 6953
rect 12618 6876 12624 6928
rect 12676 6916 12682 6928
rect 13004 6916 13032 6947
rect 14182 6944 14188 6956
rect 14240 6944 14246 6996
rect 14645 6987 14703 6993
rect 14645 6953 14657 6987
rect 14691 6984 14703 6987
rect 15562 6984 15568 6996
rect 14691 6956 15568 6984
rect 14691 6953 14703 6956
rect 14645 6947 14703 6953
rect 15562 6944 15568 6956
rect 15620 6944 15626 6996
rect 15657 6987 15715 6993
rect 15657 6953 15669 6987
rect 15703 6984 15715 6987
rect 15746 6984 15752 6996
rect 15703 6956 15752 6984
rect 15703 6953 15715 6956
rect 15657 6947 15715 6953
rect 15746 6944 15752 6956
rect 15804 6944 15810 6996
rect 15930 6916 15936 6928
rect 12676 6888 15936 6916
rect 12676 6876 12682 6888
rect 15930 6876 15936 6888
rect 15988 6876 15994 6928
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 12544 6820 13461 6848
rect 13449 6817 13461 6820
rect 13495 6817 13507 6851
rect 13449 6811 13507 6817
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6817 13691 6851
rect 14553 6851 14611 6857
rect 14553 6848 14565 6851
rect 13633 6811 13691 6817
rect 13740 6820 14565 6848
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6780 8999 6783
rect 9214 6780 9220 6792
rect 8987 6752 9220 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 9122 6712 9128 6724
rect 8496 6684 9128 6712
rect 8389 6675 8447 6681
rect 9122 6672 9128 6684
rect 9180 6672 9186 6724
rect 6178 6644 6184 6656
rect 4448 6616 6184 6644
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 6638 6644 6644 6656
rect 6599 6616 6644 6644
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 8297 6647 8355 6653
rect 8297 6613 8309 6647
rect 8343 6644 8355 6647
rect 9306 6644 9312 6656
rect 8343 6616 9312 6644
rect 8343 6613 8355 6616
rect 8297 6607 8355 6613
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 9692 6644 9720 6743
rect 9858 6644 9864 6656
rect 9692 6616 9864 6644
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 11054 6644 11060 6656
rect 11015 6616 11060 6644
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11624 6644 11652 6743
rect 13262 6740 13268 6792
rect 13320 6780 13326 6792
rect 13648 6780 13676 6811
rect 13320 6752 13676 6780
rect 13320 6740 13326 6752
rect 12894 6672 12900 6724
rect 12952 6712 12958 6724
rect 13740 6712 13768 6820
rect 14553 6817 14565 6820
rect 14599 6848 14611 6851
rect 15194 6848 15200 6860
rect 14599 6820 15200 6848
rect 14599 6817 14611 6820
rect 14553 6811 14611 6817
rect 15194 6808 15200 6820
rect 15252 6808 15258 6860
rect 16022 6848 16028 6860
rect 15764 6820 16028 6848
rect 15764 6792 15792 6820
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6780 14887 6783
rect 15102 6780 15108 6792
rect 14875 6752 15108 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 15102 6740 15108 6752
rect 15160 6780 15166 6792
rect 15746 6780 15752 6792
rect 15160 6752 15516 6780
rect 15707 6752 15752 6780
rect 15160 6740 15166 6752
rect 12952 6684 13768 6712
rect 12952 6672 12958 6684
rect 13906 6672 13912 6724
rect 13964 6712 13970 6724
rect 15289 6715 15347 6721
rect 15289 6712 15301 6715
rect 13964 6684 15301 6712
rect 13964 6672 13970 6684
rect 15289 6681 15301 6684
rect 15335 6681 15347 6715
rect 15488 6712 15516 6752
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 15856 6712 15884 6743
rect 15488 6684 15884 6712
rect 15289 6675 15347 6681
rect 13170 6644 13176 6656
rect 11624 6616 13176 6644
rect 13170 6604 13176 6616
rect 13228 6644 13234 6656
rect 13265 6647 13323 6653
rect 13265 6644 13277 6647
rect 13228 6616 13277 6644
rect 13228 6604 13234 6616
rect 13265 6613 13277 6616
rect 13311 6613 13323 6647
rect 13265 6607 13323 6613
rect 13817 6647 13875 6653
rect 13817 6613 13829 6647
rect 13863 6644 13875 6647
rect 14826 6644 14832 6656
rect 13863 6616 14832 6644
rect 13863 6613 13875 6616
rect 13817 6607 13875 6613
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 1104 6554 16836 6576
rect 1104 6502 3614 6554
rect 3666 6502 3678 6554
rect 3730 6502 3742 6554
rect 3794 6502 3806 6554
rect 3858 6502 8878 6554
rect 8930 6502 8942 6554
rect 8994 6502 9006 6554
rect 9058 6502 9070 6554
rect 9122 6502 14142 6554
rect 14194 6502 14206 6554
rect 14258 6502 14270 6554
rect 14322 6502 14334 6554
rect 14386 6502 16836 6554
rect 1104 6480 16836 6502
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4706 6440 4712 6452
rect 4212 6412 4712 6440
rect 4212 6400 4218 6412
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 7101 6443 7159 6449
rect 7101 6409 7113 6443
rect 7147 6440 7159 6443
rect 7282 6440 7288 6452
rect 7147 6412 7288 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 7484 6412 9505 6440
rect 4249 6375 4307 6381
rect 4249 6341 4261 6375
rect 4295 6372 4307 6375
rect 4433 6375 4491 6381
rect 4433 6372 4445 6375
rect 4295 6344 4445 6372
rect 4295 6341 4307 6344
rect 4249 6335 4307 6341
rect 4433 6341 4445 6344
rect 4479 6341 4491 6375
rect 4433 6335 4491 6341
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 7484 6372 7512 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 12342 6440 12348 6452
rect 9493 6403 9551 6409
rect 9692 6412 12348 6440
rect 5592 6344 7512 6372
rect 7576 6344 8064 6372
rect 5592 6332 5598 6344
rect 7300 6316 7328 6344
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6304 1455 6307
rect 1578 6304 1584 6316
rect 1443 6276 1584 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 1578 6264 1584 6276
rect 1636 6264 1642 6316
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6304 2559 6307
rect 2590 6304 2596 6316
rect 2547 6276 2596 6304
rect 2547 6273 2559 6276
rect 2501 6267 2559 6273
rect 2590 6264 2596 6276
rect 2648 6264 2654 6316
rect 3878 6264 3884 6316
rect 3936 6304 3942 6316
rect 4522 6304 4528 6316
rect 3936 6276 4528 6304
rect 3936 6264 3942 6276
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 6822 6304 6828 6316
rect 6104 6276 6828 6304
rect 1486 6196 1492 6248
rect 1544 6236 1550 6248
rect 2866 6236 2872 6248
rect 1544 6208 2872 6236
rect 1544 6196 1550 6208
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 3125 6239 3183 6245
rect 3125 6236 3137 6239
rect 3016 6208 3137 6236
rect 3016 6196 3022 6208
rect 3125 6205 3137 6208
rect 3171 6205 3183 6239
rect 4154 6236 4160 6248
rect 3125 6199 3183 6205
rect 3620 6208 4160 6236
rect 2225 6171 2283 6177
rect 2225 6137 2237 6171
rect 2271 6168 2283 6171
rect 3620 6168 3648 6208
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 6104 6236 6132 6276
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 7282 6264 7288 6316
rect 7340 6264 7346 6316
rect 7576 6313 7604 6344
rect 8036 6316 8064 6344
rect 9582 6332 9588 6384
rect 9640 6372 9646 6384
rect 9692 6372 9720 6412
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 13078 6440 13084 6452
rect 12492 6412 13084 6440
rect 12492 6400 12498 6412
rect 13078 6400 13084 6412
rect 13136 6440 13142 6452
rect 13722 6440 13728 6452
rect 13136 6412 13728 6440
rect 13136 6400 13142 6412
rect 13722 6400 13728 6412
rect 13780 6440 13786 6452
rect 16209 6443 16267 6449
rect 16209 6440 16221 6443
rect 13780 6412 16221 6440
rect 13780 6400 13786 6412
rect 16209 6409 16221 6412
rect 16255 6409 16267 6443
rect 16209 6403 16267 6409
rect 9640 6344 9720 6372
rect 11609 6375 11667 6381
rect 9640 6332 9646 6344
rect 11609 6341 11621 6375
rect 11655 6372 11667 6375
rect 11790 6372 11796 6384
rect 11655 6344 11796 6372
rect 11655 6341 11667 6344
rect 11609 6335 11667 6341
rect 11790 6332 11796 6344
rect 11848 6332 11854 6384
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6273 7619 6307
rect 7742 6304 7748 6316
rect 7703 6276 7748 6304
rect 7561 6267 7619 6273
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 8018 6264 8024 6316
rect 8076 6264 8082 6316
rect 11238 6264 11244 6316
rect 11296 6304 11302 6316
rect 12434 6304 12440 6316
rect 11296 6276 12440 6304
rect 11296 6264 11302 6276
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 12802 6264 12808 6316
rect 12860 6304 12866 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12860 6276 13001 6304
rect 12860 6264 12866 6276
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 13078 6264 13084 6316
rect 13136 6304 13142 6316
rect 13136 6276 13181 6304
rect 13136 6264 13142 6276
rect 13906 6264 13912 6316
rect 13964 6304 13970 6316
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 13964 6276 14197 6304
rect 13964 6264 13970 6276
rect 14185 6273 14197 6276
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 5000 6208 6132 6236
rect 6181 6239 6239 6245
rect 2271 6140 3648 6168
rect 4433 6171 4491 6177
rect 2271 6137 2283 6140
rect 2225 6131 2283 6137
rect 4433 6137 4445 6171
rect 4479 6168 4491 6171
rect 4706 6168 4712 6180
rect 4479 6140 4712 6168
rect 4479 6137 4491 6140
rect 4433 6131 4491 6137
rect 4706 6128 4712 6140
rect 4764 6177 4770 6180
rect 4764 6171 4828 6177
rect 4764 6137 4782 6171
rect 4816 6137 4828 6171
rect 4764 6131 4828 6137
rect 4764 6128 4770 6131
rect 1854 6100 1860 6112
rect 1815 6072 1860 6100
rect 1854 6060 1860 6072
rect 1912 6060 1918 6112
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 5000 6100 5028 6208
rect 6181 6205 6193 6239
rect 6227 6236 6239 6239
rect 6730 6236 6736 6248
rect 6227 6208 6736 6236
rect 6227 6205 6239 6208
rect 6181 6199 6239 6205
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6236 7527 6239
rect 7650 6236 7656 6248
rect 7515 6208 7656 6236
rect 7515 6205 7527 6208
rect 7469 6199 7527 6205
rect 7650 6196 7656 6208
rect 7708 6196 7714 6248
rect 7926 6196 7932 6248
rect 7984 6236 7990 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7984 6208 8125 6236
rect 7984 6196 7990 6208
rect 8113 6205 8125 6208
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 9858 6196 9864 6248
rect 9916 6236 9922 6248
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 9916 6208 10241 6236
rect 9916 6196 9922 6208
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 10496 6239 10554 6245
rect 10496 6205 10508 6239
rect 10542 6236 10554 6239
rect 11054 6236 11060 6248
rect 10542 6208 11060 6236
rect 10542 6205 10554 6208
rect 10496 6199 10554 6205
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 12066 6196 12072 6248
rect 12124 6236 12130 6248
rect 12124 6208 13032 6236
rect 12124 6196 12130 6208
rect 5166 6128 5172 6180
rect 5224 6168 5230 6180
rect 8380 6171 8438 6177
rect 5224 6140 6408 6168
rect 5224 6128 5230 6140
rect 2363 6072 5028 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 5074 6060 5080 6112
rect 5132 6100 5138 6112
rect 6380 6109 6408 6140
rect 8380 6137 8392 6171
rect 8426 6168 8438 6171
rect 8478 6168 8484 6180
rect 8426 6140 8484 6168
rect 8426 6137 8438 6140
rect 8380 6131 8438 6137
rect 8478 6128 8484 6140
rect 8536 6128 8542 6180
rect 12897 6171 12955 6177
rect 12897 6168 12909 6171
rect 11072 6140 12909 6168
rect 5905 6103 5963 6109
rect 5905 6100 5917 6103
rect 5132 6072 5917 6100
rect 5132 6060 5138 6072
rect 5905 6069 5917 6072
rect 5951 6069 5963 6103
rect 5905 6063 5963 6069
rect 6365 6103 6423 6109
rect 6365 6069 6377 6103
rect 6411 6069 6423 6103
rect 6365 6063 6423 6069
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 9122 6100 9128 6112
rect 8260 6072 9128 6100
rect 8260 6060 8266 6072
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9769 6103 9827 6109
rect 9769 6069 9781 6103
rect 9815 6100 9827 6103
rect 11072 6100 11100 6140
rect 12897 6137 12909 6140
rect 12943 6137 12955 6171
rect 12897 6131 12955 6137
rect 13004 6112 13032 6208
rect 13170 6196 13176 6248
rect 13228 6236 13234 6248
rect 14829 6239 14887 6245
rect 14829 6236 14841 6239
rect 13228 6208 14841 6236
rect 13228 6196 13234 6208
rect 14829 6205 14841 6208
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 14936 6208 15240 6236
rect 14001 6171 14059 6177
rect 14001 6137 14013 6171
rect 14047 6168 14059 6171
rect 14936 6168 14964 6208
rect 15212 6180 15240 6208
rect 15102 6177 15108 6180
rect 15096 6168 15108 6177
rect 14047 6140 14964 6168
rect 15063 6140 15108 6168
rect 14047 6137 14059 6140
rect 14001 6131 14059 6137
rect 15096 6131 15108 6140
rect 15102 6128 15108 6131
rect 15160 6128 15166 6180
rect 15194 6128 15200 6180
rect 15252 6128 15258 6180
rect 11882 6100 11888 6112
rect 9815 6072 11100 6100
rect 11843 6072 11888 6100
rect 9815 6069 9827 6072
rect 9769 6063 9827 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 12529 6103 12587 6109
rect 12529 6069 12541 6103
rect 12575 6100 12587 6103
rect 12802 6100 12808 6112
rect 12575 6072 12808 6100
rect 12575 6069 12587 6072
rect 12529 6063 12587 6069
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 12986 6060 12992 6112
rect 13044 6060 13050 6112
rect 13078 6060 13084 6112
rect 13136 6100 13142 6112
rect 13633 6103 13691 6109
rect 13633 6100 13645 6103
rect 13136 6072 13645 6100
rect 13136 6060 13142 6072
rect 13633 6069 13645 6072
rect 13679 6069 13691 6103
rect 13633 6063 13691 6069
rect 14093 6103 14151 6109
rect 14093 6069 14105 6103
rect 14139 6100 14151 6103
rect 15286 6100 15292 6112
rect 14139 6072 15292 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 1104 6010 16836 6032
rect 1104 5958 6246 6010
rect 6298 5958 6310 6010
rect 6362 5958 6374 6010
rect 6426 5958 6438 6010
rect 6490 5958 11510 6010
rect 11562 5958 11574 6010
rect 11626 5958 11638 6010
rect 11690 5958 11702 6010
rect 11754 5958 16836 6010
rect 1104 5936 16836 5958
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3697 5899 3755 5905
rect 3697 5896 3709 5899
rect 2924 5868 3709 5896
rect 2924 5856 2930 5868
rect 3697 5865 3709 5868
rect 3743 5896 3755 5899
rect 3878 5896 3884 5908
rect 3743 5868 3884 5896
rect 3743 5865 3755 5868
rect 3697 5859 3755 5865
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 4525 5899 4583 5905
rect 4525 5896 4537 5899
rect 4396 5868 4537 5896
rect 4396 5856 4402 5868
rect 4525 5865 4537 5868
rect 4571 5865 4583 5899
rect 4525 5859 4583 5865
rect 4617 5899 4675 5905
rect 4617 5865 4629 5899
rect 4663 5896 4675 5899
rect 4798 5896 4804 5908
rect 4663 5868 4804 5896
rect 4663 5865 4675 5868
rect 4617 5859 4675 5865
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5721 5899 5779 5905
rect 5721 5896 5733 5899
rect 4948 5868 5733 5896
rect 4948 5856 4954 5868
rect 5721 5865 5733 5868
rect 5767 5896 5779 5899
rect 5810 5896 5816 5908
rect 5767 5868 5816 5896
rect 5767 5865 5779 5868
rect 5721 5859 5779 5865
rect 5810 5856 5816 5868
rect 5868 5896 5874 5908
rect 7926 5896 7932 5908
rect 5868 5868 7932 5896
rect 5868 5856 5874 5868
rect 2308 5831 2366 5837
rect 2308 5797 2320 5831
rect 2354 5828 2366 5831
rect 2590 5828 2596 5840
rect 2354 5800 2596 5828
rect 2354 5797 2366 5800
rect 2308 5791 2366 5797
rect 2590 5788 2596 5800
rect 2648 5788 2654 5840
rect 3970 5788 3976 5840
rect 4028 5828 4034 5840
rect 4028 5800 5948 5828
rect 4028 5788 4034 5800
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5729 1547 5763
rect 1489 5723 1547 5729
rect 1504 5692 1532 5723
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 2041 5763 2099 5769
rect 2041 5760 2053 5763
rect 1636 5732 2053 5760
rect 1636 5720 1642 5732
rect 2041 5729 2053 5732
rect 2087 5729 2099 5763
rect 3881 5763 3939 5769
rect 2041 5723 2099 5729
rect 2148 5732 3832 5760
rect 2148 5692 2176 5732
rect 1504 5664 2176 5692
rect 3804 5692 3832 5732
rect 3881 5729 3893 5763
rect 3927 5760 3939 5763
rect 3988 5760 4016 5788
rect 3927 5732 4016 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4212 5732 4844 5760
rect 4212 5720 4218 5732
rect 4430 5692 4436 5704
rect 3804 5664 4436 5692
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 4706 5692 4712 5704
rect 4667 5664 4712 5692
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 4816 5692 4844 5732
rect 4890 5720 4896 5772
rect 4948 5760 4954 5772
rect 5169 5763 5227 5769
rect 5169 5760 5181 5763
rect 4948 5732 5181 5760
rect 4948 5720 4954 5732
rect 5169 5729 5181 5732
rect 5215 5760 5227 5763
rect 5258 5760 5264 5772
rect 5215 5732 5264 5760
rect 5215 5729 5227 5732
rect 5169 5723 5227 5729
rect 5258 5720 5264 5732
rect 5316 5720 5322 5772
rect 5920 5769 5948 5800
rect 6012 5769 6040 5868
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 8110 5896 8116 5908
rect 8071 5868 8116 5896
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 8205 5899 8263 5905
rect 8205 5865 8217 5899
rect 8251 5896 8263 5899
rect 8573 5899 8631 5905
rect 8573 5896 8585 5899
rect 8251 5868 8585 5896
rect 8251 5865 8263 5868
rect 8205 5859 8263 5865
rect 8573 5865 8585 5868
rect 8619 5865 8631 5899
rect 8573 5859 8631 5865
rect 8941 5899 8999 5905
rect 8941 5865 8953 5899
rect 8987 5896 8999 5899
rect 9674 5896 9680 5908
rect 8987 5868 9680 5896
rect 8987 5865 8999 5868
rect 8941 5859 8999 5865
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 10134 5856 10140 5908
rect 10192 5896 10198 5908
rect 10413 5899 10471 5905
rect 10413 5896 10425 5899
rect 10192 5868 10425 5896
rect 10192 5856 10198 5868
rect 10413 5865 10425 5868
rect 10459 5865 10471 5899
rect 10413 5859 10471 5865
rect 10505 5899 10563 5905
rect 10505 5865 10517 5899
rect 10551 5896 10563 5899
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 10551 5868 11069 5896
rect 10551 5865 10563 5868
rect 10505 5859 10563 5865
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 11146 5856 11152 5908
rect 11204 5896 11210 5908
rect 11517 5899 11575 5905
rect 11517 5896 11529 5899
rect 11204 5868 11529 5896
rect 11204 5856 11210 5868
rect 11517 5865 11529 5868
rect 11563 5896 11575 5899
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 11563 5868 11897 5896
rect 11563 5865 11575 5868
rect 11517 5859 11575 5865
rect 11885 5865 11897 5868
rect 11931 5865 11943 5899
rect 11885 5859 11943 5865
rect 12069 5899 12127 5905
rect 12069 5865 12081 5899
rect 12115 5896 12127 5899
rect 12158 5896 12164 5908
rect 12115 5868 12164 5896
rect 12115 5865 12127 5868
rect 12069 5859 12127 5865
rect 12158 5856 12164 5868
rect 12216 5856 12222 5908
rect 12437 5899 12495 5905
rect 12437 5865 12449 5899
rect 12483 5896 12495 5899
rect 12802 5896 12808 5908
rect 12483 5868 12808 5896
rect 12483 5865 12495 5868
rect 12437 5859 12495 5865
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 15286 5896 15292 5908
rect 15247 5868 15292 5896
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 15746 5896 15752 5908
rect 15707 5868 15752 5896
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 6822 5828 6828 5840
rect 6104 5800 6828 5828
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5729 5963 5763
rect 5905 5723 5963 5729
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5729 6055 5763
rect 5997 5723 6055 5729
rect 6104 5692 6132 5800
rect 6822 5788 6828 5800
rect 6880 5788 6886 5840
rect 10226 5828 10232 5840
rect 8036 5800 10232 5828
rect 6264 5763 6322 5769
rect 6264 5729 6276 5763
rect 6310 5760 6322 5763
rect 6638 5760 6644 5772
rect 6310 5732 6644 5760
rect 6310 5729 6322 5732
rect 6264 5723 6322 5729
rect 6638 5720 6644 5732
rect 6696 5760 6702 5772
rect 7650 5760 7656 5772
rect 6696 5732 7656 5760
rect 6696 5720 6702 5732
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7466 5692 7472 5704
rect 4816 5664 6132 5692
rect 7379 5664 7472 5692
rect 7392 5633 7420 5664
rect 7466 5652 7472 5664
rect 7524 5692 7530 5704
rect 8036 5692 8064 5800
rect 10226 5788 10232 5800
rect 10284 5788 10290 5840
rect 11425 5831 11483 5837
rect 11425 5828 11437 5831
rect 10612 5800 11437 5828
rect 9766 5760 9772 5772
rect 8312 5732 9772 5760
rect 8312 5701 8340 5732
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 7524 5664 8064 5692
rect 8297 5695 8355 5701
rect 7524 5652 7530 5664
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 8938 5652 8944 5704
rect 8996 5692 9002 5704
rect 9033 5695 9091 5701
rect 9033 5692 9045 5695
rect 8996 5664 9045 5692
rect 8996 5652 9002 5664
rect 9033 5661 9045 5664
rect 9079 5661 9091 5695
rect 9214 5692 9220 5704
rect 9175 5664 9220 5692
rect 9033 5655 9091 5661
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9582 5652 9588 5704
rect 9640 5692 9646 5704
rect 10612 5692 10640 5800
rect 11425 5797 11437 5800
rect 11471 5828 11483 5831
rect 12526 5828 12532 5840
rect 11471 5800 11928 5828
rect 12487 5800 12532 5828
rect 11471 5797 11483 5800
rect 11425 5791 11483 5797
rect 11054 5720 11060 5772
rect 11112 5760 11118 5772
rect 11112 5732 11468 5760
rect 11112 5720 11118 5732
rect 9640 5664 10640 5692
rect 10689 5695 10747 5701
rect 9640 5652 9646 5664
rect 10689 5661 10701 5695
rect 10735 5692 10747 5695
rect 10962 5692 10968 5704
rect 10735 5664 10968 5692
rect 10735 5661 10747 5664
rect 10689 5655 10747 5661
rect 10962 5652 10968 5664
rect 11020 5692 11026 5704
rect 11440 5692 11468 5732
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 11020 5664 11376 5692
rect 11440 5664 11621 5692
rect 11020 5652 11026 5664
rect 5353 5627 5411 5633
rect 5353 5624 5365 5627
rect 2976 5596 5365 5624
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 1946 5516 1952 5568
rect 2004 5556 2010 5568
rect 2976 5556 3004 5596
rect 5353 5593 5365 5596
rect 5399 5593 5411 5627
rect 5353 5587 5411 5593
rect 7377 5627 7435 5633
rect 7377 5593 7389 5627
rect 7423 5593 7435 5627
rect 7377 5587 7435 5593
rect 7745 5627 7803 5633
rect 7745 5593 7757 5627
rect 7791 5624 7803 5627
rect 11238 5624 11244 5636
rect 7791 5596 11244 5624
rect 7791 5593 7803 5596
rect 7745 5587 7803 5593
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 11348 5624 11376 5664
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 11790 5624 11796 5636
rect 11348 5596 11796 5624
rect 11790 5584 11796 5596
rect 11848 5584 11854 5636
rect 11900 5624 11928 5800
rect 12526 5788 12532 5800
rect 12584 5788 12590 5840
rect 15657 5831 15715 5837
rect 15657 5828 15669 5831
rect 12636 5800 15669 5828
rect 12636 5760 12664 5800
rect 15657 5797 15669 5800
rect 15703 5797 15715 5831
rect 15657 5791 15715 5797
rect 11992 5732 12664 5760
rect 13081 5763 13139 5769
rect 11992 5704 12020 5732
rect 13081 5729 13093 5763
rect 13127 5760 13139 5763
rect 13170 5760 13176 5772
rect 13127 5732 13176 5760
rect 13127 5729 13139 5732
rect 13081 5723 13139 5729
rect 13170 5720 13176 5732
rect 13228 5720 13234 5772
rect 13354 5769 13360 5772
rect 13348 5760 13360 5769
rect 13315 5732 13360 5760
rect 13348 5723 13360 5732
rect 13354 5720 13360 5723
rect 13412 5720 13418 5772
rect 11974 5652 11980 5704
rect 12032 5652 12038 5704
rect 12618 5692 12624 5704
rect 12579 5664 12624 5692
rect 12618 5652 12624 5664
rect 12676 5652 12682 5704
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5692 14795 5695
rect 15562 5692 15568 5704
rect 14783 5664 15568 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 15562 5652 15568 5664
rect 15620 5652 15626 5704
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 12894 5624 12900 5636
rect 11900 5596 12900 5624
rect 12894 5584 12900 5596
rect 12952 5584 12958 5636
rect 14461 5627 14519 5633
rect 14461 5593 14473 5627
rect 14507 5624 14519 5627
rect 15102 5624 15108 5636
rect 14507 5596 15108 5624
rect 14507 5593 14519 5596
rect 14461 5587 14519 5593
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 15286 5584 15292 5636
rect 15344 5624 15350 5636
rect 15856 5624 15884 5655
rect 15344 5596 15884 5624
rect 15344 5584 15350 5596
rect 2004 5528 3004 5556
rect 3421 5559 3479 5565
rect 2004 5516 2010 5528
rect 3421 5525 3433 5559
rect 3467 5556 3479 5559
rect 3510 5556 3516 5568
rect 3467 5528 3516 5556
rect 3467 5525 3479 5528
rect 3421 5519 3479 5525
rect 3510 5516 3516 5528
rect 3568 5516 3574 5568
rect 4154 5556 4160 5568
rect 4115 5528 4160 5556
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 5534 5556 5540 5568
rect 4672 5528 5540 5556
rect 4672 5516 4678 5528
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 5902 5516 5908 5568
rect 5960 5556 5966 5568
rect 6178 5556 6184 5568
rect 5960 5528 6184 5556
rect 5960 5516 5966 5528
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 10042 5556 10048 5568
rect 10003 5528 10048 5556
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 10134 5516 10140 5568
rect 10192 5556 10198 5568
rect 11330 5556 11336 5568
rect 10192 5528 11336 5556
rect 10192 5516 10198 5528
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 11885 5559 11943 5565
rect 11885 5525 11897 5559
rect 11931 5556 11943 5559
rect 15654 5556 15660 5568
rect 11931 5528 15660 5556
rect 11931 5525 11943 5528
rect 11885 5519 11943 5525
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 1104 5466 16836 5488
rect 1104 5414 3614 5466
rect 3666 5414 3678 5466
rect 3730 5414 3742 5466
rect 3794 5414 3806 5466
rect 3858 5414 8878 5466
rect 8930 5414 8942 5466
rect 8994 5414 9006 5466
rect 9058 5414 9070 5466
rect 9122 5414 14142 5466
rect 14194 5414 14206 5466
rect 14258 5414 14270 5466
rect 14322 5414 14334 5466
rect 14386 5414 16836 5466
rect 1104 5392 16836 5414
rect 2774 5312 2780 5364
rect 2832 5312 2838 5364
rect 5074 5352 5080 5364
rect 3896 5324 5080 5352
rect 2792 5284 2820 5312
rect 1688 5256 2820 5284
rect 1688 5225 1716 5256
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 2590 5176 2596 5228
rect 2648 5216 2654 5228
rect 2777 5219 2835 5225
rect 2777 5216 2789 5219
rect 2648 5188 2789 5216
rect 2648 5176 2654 5188
rect 2777 5185 2789 5188
rect 2823 5216 2835 5219
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 2823 5188 3801 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 3789 5185 3801 5188
rect 3835 5216 3847 5219
rect 3896 5216 3924 5324
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6825 5355 6883 5361
rect 6825 5352 6837 5355
rect 6328 5324 6837 5352
rect 6328 5312 6334 5324
rect 6825 5321 6837 5324
rect 6871 5321 6883 5355
rect 6825 5315 6883 5321
rect 7282 5312 7288 5364
rect 7340 5352 7346 5364
rect 8018 5352 8024 5364
rect 7340 5324 8024 5352
rect 7340 5312 7346 5324
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 8573 5355 8631 5361
rect 8573 5321 8585 5355
rect 8619 5352 8631 5355
rect 8754 5352 8760 5364
rect 8619 5324 8760 5352
rect 8619 5321 8631 5324
rect 8573 5315 8631 5321
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 9858 5352 9864 5364
rect 9600 5324 9864 5352
rect 4157 5287 4215 5293
rect 4157 5253 4169 5287
rect 4203 5284 4215 5287
rect 4203 5256 7328 5284
rect 4203 5253 4215 5256
rect 4157 5247 4215 5253
rect 3835 5188 3924 5216
rect 4801 5219 4859 5225
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 4890 5216 4896 5228
rect 4847 5188 4896 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 4890 5176 4896 5188
rect 4948 5216 4954 5228
rect 5718 5216 5724 5228
rect 4948 5188 5724 5216
rect 4948 5176 4954 5188
rect 5718 5176 5724 5188
rect 5776 5176 5782 5228
rect 7300 5225 7328 5256
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5185 7343 5219
rect 7466 5216 7472 5228
rect 7427 5188 7472 5216
rect 7285 5179 7343 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 7742 5176 7748 5228
rect 7800 5216 7806 5228
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 7800 5188 9137 5216
rect 7800 5176 7806 5188
rect 9125 5185 9137 5188
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 2314 5148 2320 5160
rect 1443 5120 2320 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 2314 5108 2320 5120
rect 2372 5108 2378 5160
rect 2406 5108 2412 5160
rect 2464 5148 2470 5160
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 2464 5120 2513 5148
rect 2464 5108 2470 5120
rect 2501 5117 2513 5120
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 3605 5151 3663 5157
rect 3605 5117 3617 5151
rect 3651 5148 3663 5151
rect 4154 5148 4160 5160
rect 3651 5120 4160 5148
rect 3651 5117 3663 5120
rect 3605 5111 3663 5117
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 4614 5148 4620 5160
rect 4571 5120 4620 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5148 5595 5151
rect 5902 5148 5908 5160
rect 5583 5120 5908 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 6178 5148 6184 5160
rect 6139 5120 6184 5148
rect 6178 5108 6184 5120
rect 6236 5148 6242 5160
rect 6638 5148 6644 5160
rect 6236 5120 6644 5148
rect 6236 5108 6242 5120
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 7653 5151 7711 5157
rect 7653 5148 7665 5151
rect 6972 5120 7665 5148
rect 6972 5108 6978 5120
rect 7653 5117 7665 5120
rect 7699 5117 7711 5151
rect 7653 5111 7711 5117
rect 8662 5108 8668 5160
rect 8720 5148 8726 5160
rect 9600 5157 9628 5324
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 15010 5352 15016 5364
rect 10928 5324 15016 5352
rect 10928 5312 10934 5324
rect 15010 5312 15016 5324
rect 15068 5312 15074 5364
rect 10965 5287 11023 5293
rect 10965 5253 10977 5287
rect 11011 5253 11023 5287
rect 10965 5247 11023 5253
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 10980 5216 11008 5247
rect 14090 5244 14096 5296
rect 14148 5284 14154 5296
rect 14642 5284 14648 5296
rect 14148 5256 14648 5284
rect 14148 5244 14154 5256
rect 14642 5244 14648 5256
rect 14700 5244 14706 5296
rect 11793 5219 11851 5225
rect 11793 5216 11805 5219
rect 10744 5188 11805 5216
rect 10744 5176 10750 5188
rect 11793 5185 11805 5188
rect 11839 5185 11851 5219
rect 14829 5219 14887 5225
rect 14829 5216 14841 5219
rect 11793 5179 11851 5185
rect 13464 5188 14841 5216
rect 8941 5151 8999 5157
rect 8941 5148 8953 5151
rect 8720 5120 8953 5148
rect 8720 5108 8726 5120
rect 8941 5117 8953 5120
rect 8987 5117 8999 5151
rect 8941 5111 8999 5117
rect 9585 5151 9643 5157
rect 9585 5117 9597 5151
rect 9631 5148 9643 5151
rect 9674 5148 9680 5160
rect 9631 5120 9680 5148
rect 9631 5117 9643 5120
rect 9585 5111 9643 5117
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 9852 5151 9910 5157
rect 9852 5117 9864 5151
rect 9898 5148 9910 5151
rect 10962 5148 10968 5160
rect 9898 5120 10968 5148
rect 9898 5117 9910 5120
rect 9852 5111 9910 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 13170 5148 13176 5160
rect 12483 5120 13176 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 13170 5108 13176 5120
rect 13228 5148 13234 5160
rect 13464 5148 13492 5188
rect 14829 5185 14841 5188
rect 14875 5185 14887 5219
rect 14829 5179 14887 5185
rect 13228 5120 13492 5148
rect 13228 5108 13234 5120
rect 13722 5108 13728 5160
rect 13780 5148 13786 5160
rect 14277 5151 14335 5157
rect 14277 5148 14289 5151
rect 13780 5120 14289 5148
rect 13780 5108 13786 5120
rect 14277 5117 14289 5120
rect 14323 5117 14335 5151
rect 14277 5111 14335 5117
rect 2593 5083 2651 5089
rect 2593 5049 2605 5083
rect 2639 5080 2651 5083
rect 2958 5080 2964 5092
rect 2639 5052 2964 5080
rect 2639 5049 2651 5052
rect 2593 5043 2651 5049
rect 2958 5040 2964 5052
rect 3016 5040 3022 5092
rect 4430 5080 4436 5092
rect 3160 5052 4436 5080
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 3160 5021 3188 5052
rect 4430 5040 4436 5052
rect 4488 5040 4494 5092
rect 7193 5083 7251 5089
rect 7193 5080 7205 5083
rect 5184 5052 7205 5080
rect 3145 5015 3203 5021
rect 3145 4981 3157 5015
rect 3191 4981 3203 5015
rect 3145 4975 3203 4981
rect 3513 5015 3571 5021
rect 3513 4981 3525 5015
rect 3559 5012 3571 5015
rect 3602 5012 3608 5024
rect 3559 4984 3608 5012
rect 3559 4981 3571 4984
rect 3513 4975 3571 4981
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 4614 5012 4620 5024
rect 4575 4984 4620 5012
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 5184 5021 5212 5052
rect 7193 5049 7205 5052
rect 7239 5049 7251 5083
rect 7193 5043 7251 5049
rect 7282 5040 7288 5092
rect 7340 5080 7346 5092
rect 7929 5083 7987 5089
rect 7929 5080 7941 5083
rect 7340 5052 7941 5080
rect 7340 5040 7346 5052
rect 7929 5049 7941 5052
rect 7975 5049 7987 5083
rect 7929 5043 7987 5049
rect 8110 5040 8116 5092
rect 8168 5080 8174 5092
rect 8168 5052 11100 5080
rect 8168 5040 8174 5052
rect 11072 5024 11100 5052
rect 11146 5040 11152 5092
rect 11204 5080 11210 5092
rect 11701 5083 11759 5089
rect 11701 5080 11713 5083
rect 11204 5052 11713 5080
rect 11204 5040 11210 5052
rect 11701 5049 11713 5052
rect 11747 5049 11759 5083
rect 11701 5043 11759 5049
rect 12704 5083 12762 5089
rect 12704 5049 12716 5083
rect 12750 5080 12762 5083
rect 13906 5080 13912 5092
rect 12750 5052 13912 5080
rect 12750 5049 12762 5052
rect 12704 5043 12762 5049
rect 13906 5040 13912 5052
rect 13964 5080 13970 5092
rect 15096 5083 15154 5089
rect 13964 5052 15056 5080
rect 13964 5040 13970 5052
rect 5169 5015 5227 5021
rect 5169 4981 5181 5015
rect 5215 4981 5227 5015
rect 5169 4975 5227 4981
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 5629 5015 5687 5021
rect 5629 5012 5641 5015
rect 5592 4984 5641 5012
rect 5592 4972 5598 4984
rect 5629 4981 5641 4984
rect 5675 4981 5687 5015
rect 5629 4975 5687 4981
rect 5718 4972 5724 5024
rect 5776 5012 5782 5024
rect 6365 5015 6423 5021
rect 6365 5012 6377 5015
rect 5776 4984 6377 5012
rect 5776 4972 5782 4984
rect 6365 4981 6377 4984
rect 6411 4981 6423 5015
rect 6365 4975 6423 4981
rect 8386 4972 8392 5024
rect 8444 5012 8450 5024
rect 9033 5015 9091 5021
rect 9033 5012 9045 5015
rect 8444 4984 9045 5012
rect 8444 4972 8450 4984
rect 9033 4981 9045 4984
rect 9079 4981 9091 5015
rect 9033 4975 9091 4981
rect 9766 4972 9772 5024
rect 9824 5012 9830 5024
rect 10502 5012 10508 5024
rect 9824 4984 10508 5012
rect 9824 4972 9830 4984
rect 10502 4972 10508 4984
rect 10560 5012 10566 5024
rect 10962 5012 10968 5024
rect 10560 4984 10968 5012
rect 10560 4972 10566 4984
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11054 4972 11060 5024
rect 11112 4972 11118 5024
rect 11238 5012 11244 5024
rect 11199 4984 11244 5012
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 11330 4972 11336 5024
rect 11388 5012 11394 5024
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 11388 4984 11621 5012
rect 11388 4972 11394 4984
rect 11609 4981 11621 4984
rect 11655 4981 11667 5015
rect 11609 4975 11667 4981
rect 12802 4972 12808 5024
rect 12860 5012 12866 5024
rect 13354 5012 13360 5024
rect 12860 4984 13360 5012
rect 12860 4972 12866 4984
rect 13354 4972 13360 4984
rect 13412 5012 13418 5024
rect 13817 5015 13875 5021
rect 13817 5012 13829 5015
rect 13412 4984 13829 5012
rect 13412 4972 13418 4984
rect 13817 4981 13829 4984
rect 13863 4981 13875 5015
rect 13817 4975 13875 4981
rect 14461 5015 14519 5021
rect 14461 4981 14473 5015
rect 14507 5012 14519 5015
rect 14918 5012 14924 5024
rect 14507 4984 14924 5012
rect 14507 4981 14519 4984
rect 14461 4975 14519 4981
rect 14918 4972 14924 4984
rect 14976 4972 14982 5024
rect 15028 5012 15056 5052
rect 15096 5049 15108 5083
rect 15142 5080 15154 5083
rect 15286 5080 15292 5092
rect 15142 5052 15292 5080
rect 15142 5049 15154 5052
rect 15096 5043 15154 5049
rect 15286 5040 15292 5052
rect 15344 5040 15350 5092
rect 16209 5015 16267 5021
rect 16209 5012 16221 5015
rect 15028 4984 16221 5012
rect 16209 4981 16221 4984
rect 16255 4981 16267 5015
rect 16209 4975 16267 4981
rect 1104 4922 16836 4944
rect 1104 4870 6246 4922
rect 6298 4870 6310 4922
rect 6362 4870 6374 4922
rect 6426 4870 6438 4922
rect 6490 4870 11510 4922
rect 11562 4870 11574 4922
rect 11626 4870 11638 4922
rect 11690 4870 11702 4922
rect 11754 4870 16836 4922
rect 1104 4848 16836 4870
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 5718 4808 5724 4820
rect 2556 4780 5724 4808
rect 2556 4768 2562 4780
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 5960 4780 6500 4808
rect 5960 4768 5966 4780
rect 6472 4752 6500 4780
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 6696 4780 8432 4808
rect 6696 4768 6702 4780
rect 2406 4740 2412 4752
rect 1504 4712 2412 4740
rect 1504 4684 1532 4712
rect 2406 4700 2412 4712
rect 2464 4700 2470 4752
rect 4154 4740 4160 4752
rect 3252 4712 4160 4740
rect 1486 4672 1492 4684
rect 1447 4644 1492 4672
rect 1486 4632 1492 4644
rect 1544 4632 1550 4684
rect 1762 4681 1768 4684
rect 1756 4635 1768 4681
rect 1820 4672 1826 4684
rect 3252 4681 3280 4712
rect 4154 4700 4160 4712
rect 4212 4700 4218 4752
rect 4614 4700 4620 4752
rect 4672 4740 4678 4752
rect 6086 4740 6092 4752
rect 4672 4712 6092 4740
rect 4672 4700 4678 4712
rect 6086 4700 6092 4712
rect 6144 4700 6150 4752
rect 6454 4700 6460 4752
rect 6512 4700 6518 4752
rect 7006 4700 7012 4752
rect 7064 4740 7070 4752
rect 7644 4743 7702 4749
rect 7064 4712 7604 4740
rect 7064 4700 7070 4712
rect 3237 4675 3295 4681
rect 1820 4644 1856 4672
rect 1762 4632 1768 4635
rect 1820 4632 1826 4644
rect 3237 4641 3249 4675
rect 3283 4641 3295 4675
rect 3237 4635 3295 4641
rect 3878 4632 3884 4684
rect 3936 4672 3942 4684
rect 4065 4675 4123 4681
rect 4065 4672 4077 4675
rect 3936 4644 4077 4672
rect 3936 4632 3942 4644
rect 4065 4641 4077 4644
rect 4111 4641 4123 4675
rect 4065 4635 4123 4641
rect 4332 4675 4390 4681
rect 4332 4641 4344 4675
rect 4378 4672 4390 4675
rect 4890 4672 4896 4684
rect 4378 4644 4896 4672
rect 4378 4641 4390 4644
rect 4332 4635 4390 4641
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5977 4675 6035 4681
rect 5977 4672 5989 4675
rect 5644 4644 5989 4672
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4604 3571 4607
rect 3970 4604 3976 4616
rect 3559 4576 3976 4604
rect 3559 4573 3571 4576
rect 3513 4567 3571 4573
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 5644 4536 5672 4644
rect 5977 4641 5989 4644
rect 6023 4672 6035 4675
rect 7466 4672 7472 4684
rect 6023 4644 7472 4672
rect 6023 4641 6035 4644
rect 5977 4635 6035 4641
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 7576 4672 7604 4712
rect 7644 4709 7656 4743
rect 7690 4740 7702 4743
rect 8110 4740 8116 4752
rect 7690 4712 8116 4740
rect 7690 4709 7702 4712
rect 7644 4703 7702 4709
rect 8110 4700 8116 4712
rect 8168 4700 8174 4752
rect 8404 4740 8432 4780
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 10505 4811 10563 4817
rect 10505 4808 10517 4811
rect 10100 4780 10517 4808
rect 10100 4768 10106 4780
rect 10505 4777 10517 4780
rect 10551 4777 10563 4811
rect 10505 4771 10563 4777
rect 11425 4811 11483 4817
rect 11425 4777 11437 4811
rect 11471 4808 11483 4811
rect 11974 4808 11980 4820
rect 11471 4780 11980 4808
rect 11471 4777 11483 4780
rect 11425 4771 11483 4777
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 12621 4811 12679 4817
rect 12621 4777 12633 4811
rect 12667 4808 12679 4811
rect 13173 4811 13231 4817
rect 13173 4808 13185 4811
rect 12667 4780 13185 4808
rect 12667 4777 12679 4780
rect 12621 4771 12679 4777
rect 13173 4777 13185 4780
rect 13219 4777 13231 4811
rect 13173 4771 13231 4777
rect 13541 4811 13599 4817
rect 13541 4777 13553 4811
rect 13587 4808 13599 4811
rect 14185 4811 14243 4817
rect 14185 4808 14197 4811
rect 13587 4780 14197 4808
rect 13587 4777 13599 4780
rect 13541 4771 13599 4777
rect 14185 4777 14197 4780
rect 14231 4777 14243 4811
rect 14185 4771 14243 4777
rect 14458 4768 14464 4820
rect 14516 4808 14522 4820
rect 14553 4811 14611 4817
rect 14553 4808 14565 4811
rect 14516 4780 14565 4808
rect 14516 4768 14522 4780
rect 14553 4777 14565 4780
rect 14599 4777 14611 4811
rect 14553 4771 14611 4777
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15289 4811 15347 4817
rect 15289 4808 15301 4811
rect 15252 4780 15301 4808
rect 15252 4768 15258 4780
rect 15289 4777 15301 4780
rect 15335 4777 15347 4811
rect 15289 4771 15347 4777
rect 15562 4768 15568 4820
rect 15620 4808 15626 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15620 4780 15669 4808
rect 15620 4768 15626 4780
rect 15657 4777 15669 4780
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 10413 4743 10471 4749
rect 8404 4712 9812 4740
rect 8849 4675 8907 4681
rect 8849 4672 8861 4675
rect 7576 4644 8861 4672
rect 8849 4641 8861 4644
rect 8895 4641 8907 4675
rect 8849 4635 8907 4641
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 9784 4672 9812 4712
rect 10413 4709 10425 4743
rect 10459 4740 10471 4743
rect 10873 4743 10931 4749
rect 10873 4740 10885 4743
rect 10459 4712 10885 4740
rect 10459 4709 10471 4712
rect 10413 4703 10471 4709
rect 10873 4709 10885 4712
rect 10919 4709 10931 4743
rect 10873 4703 10931 4709
rect 10962 4700 10968 4752
rect 11020 4740 11026 4752
rect 14645 4743 14703 4749
rect 14645 4740 14657 4743
rect 11020 4712 14657 4740
rect 11020 4700 11026 4712
rect 14645 4709 14657 4712
rect 14691 4709 14703 4743
rect 14645 4703 14703 4709
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 9784 4644 11529 4672
rect 9677 4635 9735 4641
rect 11517 4641 11529 4644
rect 11563 4672 11575 4675
rect 12342 4672 12348 4684
rect 11563 4644 12348 4672
rect 11563 4641 11575 4644
rect 11517 4635 11575 4641
rect 5718 4564 5724 4616
rect 5776 4604 5782 4616
rect 7377 4607 7435 4613
rect 7377 4604 7389 4607
rect 5776 4576 5821 4604
rect 6748 4576 7389 4604
rect 5776 4564 5782 4576
rect 5460 4508 5672 4536
rect 2866 4468 2872 4480
rect 2827 4440 2872 4468
rect 2866 4428 2872 4440
rect 2924 4428 2930 4480
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 4062 4468 4068 4480
rect 3292 4440 4068 4468
rect 3292 4428 3298 4440
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 5460 4477 5488 4508
rect 5445 4471 5503 4477
rect 5445 4468 5457 4471
rect 5316 4440 5457 4468
rect 5316 4428 5322 4440
rect 5445 4437 5457 4440
rect 5491 4437 5503 4471
rect 5736 4468 5764 4564
rect 6748 4468 6776 4576
rect 7377 4573 7389 4576
rect 7423 4573 7435 4607
rect 7377 4567 7435 4573
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 9033 4607 9091 4613
rect 9033 4604 9045 4607
rect 8444 4576 9045 4604
rect 8444 4564 8450 4576
rect 9033 4573 9045 4576
rect 9079 4573 9091 4607
rect 9033 4567 9091 4573
rect 9692 4604 9720 4635
rect 12342 4632 12348 4644
rect 12400 4632 12406 4684
rect 12529 4675 12587 4681
rect 12529 4641 12541 4675
rect 12575 4672 12587 4675
rect 13078 4672 13084 4684
rect 12575 4644 13084 4672
rect 12575 4641 12587 4644
rect 12529 4635 12587 4641
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13633 4675 13691 4681
rect 13633 4641 13645 4675
rect 13679 4672 13691 4675
rect 13814 4672 13820 4684
rect 13679 4644 13820 4672
rect 13679 4641 13691 4644
rect 13633 4635 13691 4641
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 10410 4604 10416 4616
rect 9692 4576 10416 4604
rect 9692 4536 9720 4576
rect 10410 4564 10416 4576
rect 10468 4564 10474 4616
rect 10686 4604 10692 4616
rect 10647 4576 10692 4604
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4604 11759 4607
rect 11790 4604 11796 4616
rect 11747 4576 11796 4604
rect 11747 4573 11759 4576
rect 11701 4567 11759 4573
rect 11790 4564 11796 4576
rect 11848 4604 11854 4616
rect 11974 4604 11980 4616
rect 11848 4576 11980 4604
rect 11848 4564 11854 4576
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 12802 4604 12808 4616
rect 12763 4576 12808 4604
rect 12802 4564 12808 4576
rect 12860 4564 12866 4616
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4604 13783 4607
rect 13906 4604 13912 4616
rect 13771 4576 13912 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 13906 4564 13912 4576
rect 13964 4564 13970 4616
rect 14829 4607 14887 4613
rect 14829 4573 14841 4607
rect 14875 4604 14887 4607
rect 15194 4604 15200 4616
rect 14875 4576 15200 4604
rect 14875 4573 14887 4576
rect 14829 4567 14887 4573
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 15746 4604 15752 4616
rect 15707 4576 15752 4604
rect 15746 4564 15752 4576
rect 15804 4564 15810 4616
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 8312 4508 9720 4536
rect 9861 4539 9919 4545
rect 6822 4468 6828 4480
rect 5736 4440 6828 4468
rect 5445 4431 5503 4437
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 7064 4440 7113 4468
rect 7064 4428 7070 4440
rect 7101 4437 7113 4440
rect 7147 4437 7159 4471
rect 7101 4431 7159 4437
rect 7650 4428 7656 4480
rect 7708 4468 7714 4480
rect 8312 4468 8340 4508
rect 9861 4505 9873 4539
rect 9907 4536 9919 4539
rect 14734 4536 14740 4548
rect 9907 4508 14740 4536
rect 9907 4505 9919 4508
rect 9861 4499 9919 4505
rect 14734 4496 14740 4508
rect 14792 4496 14798 4548
rect 15212 4536 15240 4564
rect 15856 4536 15884 4567
rect 15212 4508 15884 4536
rect 7708 4440 8340 4468
rect 7708 4428 7714 4440
rect 8478 4428 8484 4480
rect 8536 4468 8542 4480
rect 8757 4471 8815 4477
rect 8757 4468 8769 4471
rect 8536 4440 8769 4468
rect 8536 4428 8542 4440
rect 8757 4437 8769 4440
rect 8803 4468 8815 4471
rect 9398 4468 9404 4480
rect 8803 4440 9404 4468
rect 8803 4437 8815 4440
rect 8757 4431 8815 4437
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 10045 4471 10103 4477
rect 10045 4437 10057 4471
rect 10091 4468 10103 4471
rect 10502 4468 10508 4480
rect 10091 4440 10508 4468
rect 10091 4437 10103 4440
rect 10045 4431 10103 4437
rect 10502 4428 10508 4440
rect 10560 4428 10566 4480
rect 10873 4471 10931 4477
rect 10873 4437 10885 4471
rect 10919 4468 10931 4471
rect 11057 4471 11115 4477
rect 11057 4468 11069 4471
rect 10919 4440 11069 4468
rect 10919 4437 10931 4440
rect 10873 4431 10931 4437
rect 11057 4437 11069 4440
rect 11103 4437 11115 4471
rect 11057 4431 11115 4437
rect 12161 4471 12219 4477
rect 12161 4437 12173 4471
rect 12207 4468 12219 4471
rect 13906 4468 13912 4480
rect 12207 4440 13912 4468
rect 12207 4437 12219 4440
rect 12161 4431 12219 4437
rect 13906 4428 13912 4440
rect 13964 4428 13970 4480
rect 1104 4378 16836 4400
rect 1104 4326 3614 4378
rect 3666 4326 3678 4378
rect 3730 4326 3742 4378
rect 3794 4326 3806 4378
rect 3858 4326 8878 4378
rect 8930 4326 8942 4378
rect 8994 4326 9006 4378
rect 9058 4326 9070 4378
rect 9122 4326 14142 4378
rect 14194 4326 14206 4378
rect 14258 4326 14270 4378
rect 14322 4326 14334 4378
rect 14386 4326 16836 4378
rect 1104 4304 16836 4326
rect 3510 4264 3516 4276
rect 1964 4236 3516 4264
rect 1762 4156 1768 4208
rect 1820 4196 1826 4208
rect 1964 4196 1992 4236
rect 3510 4224 3516 4236
rect 3568 4264 3574 4276
rect 3568 4236 4660 4264
rect 3568 4224 3574 4236
rect 1820 4168 1992 4196
rect 1820 4156 1826 4168
rect 1854 4128 1860 4140
rect 1815 4100 1860 4128
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 1964 4137 1992 4168
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 2406 4128 2412 4140
rect 2367 4100 2412 4128
rect 1949 4091 2007 4097
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 4632 4137 4660 4236
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 5592 4236 7788 4264
rect 5592 4224 5598 4236
rect 5074 4196 5080 4208
rect 5035 4168 5080 4196
rect 5074 4156 5080 4168
rect 5132 4156 5138 4208
rect 5902 4156 5908 4208
rect 5960 4196 5966 4208
rect 6638 4196 6644 4208
rect 5960 4168 6644 4196
rect 5960 4156 5966 4168
rect 6638 4156 6644 4168
rect 6696 4156 6702 4208
rect 7760 4196 7788 4236
rect 8110 4224 8116 4276
rect 8168 4264 8174 4276
rect 8205 4267 8263 4273
rect 8205 4264 8217 4267
rect 8168 4236 8217 4264
rect 8168 4224 8174 4236
rect 8205 4233 8217 4236
rect 8251 4233 8263 4267
rect 10778 4264 10784 4276
rect 8205 4227 8263 4233
rect 8404 4236 10784 4264
rect 8404 4196 8432 4236
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 12250 4224 12256 4276
rect 12308 4264 12314 4276
rect 12434 4264 12440 4276
rect 12308 4236 12440 4264
rect 12308 4224 12314 4236
rect 12434 4224 12440 4236
rect 12492 4224 12498 4276
rect 15194 4224 15200 4276
rect 15252 4264 15258 4276
rect 15473 4267 15531 4273
rect 15473 4264 15485 4267
rect 15252 4236 15485 4264
rect 15252 4224 15258 4236
rect 15473 4233 15485 4236
rect 15519 4233 15531 4267
rect 15473 4227 15531 4233
rect 7760 4168 8432 4196
rect 8481 4199 8539 4205
rect 8481 4165 8493 4199
rect 8527 4165 8539 4199
rect 8481 4159 8539 4165
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 4488 4100 4537 4128
rect 4488 4088 4494 4100
rect 4525 4097 4537 4100
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 5626 4128 5632 4140
rect 5587 4100 5632 4128
rect 4617 4091 4675 4097
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 6822 4128 6828 4140
rect 6783 4100 6828 4128
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 1765 4063 1823 4069
rect 1765 4029 1777 4063
rect 1811 4060 1823 4063
rect 2038 4060 2044 4072
rect 1811 4032 2044 4060
rect 1811 4029 1823 4032
rect 1765 4023 1823 4029
rect 2038 4020 2044 4032
rect 2096 4020 2102 4072
rect 2130 4020 2136 4072
rect 2188 4060 2194 4072
rect 4338 4060 4344 4072
rect 2188 4032 4344 4060
rect 2188 4020 2194 4032
rect 4338 4020 4344 4032
rect 4396 4020 4402 4072
rect 6086 4060 6092 4072
rect 6047 4032 6092 4060
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 2676 3995 2734 4001
rect 2676 3961 2688 3995
rect 2722 3992 2734 3995
rect 2866 3992 2872 4004
rect 2722 3964 2872 3992
rect 2722 3961 2734 3964
rect 2676 3955 2734 3961
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 3878 3952 3884 4004
rect 3936 3992 3942 4004
rect 3936 3964 6316 3992
rect 3936 3952 3942 3964
rect 1394 3924 1400 3936
rect 1355 3896 1400 3924
rect 1394 3884 1400 3896
rect 1452 3884 1458 3936
rect 2406 3884 2412 3936
rect 2464 3924 2470 3936
rect 3510 3924 3516 3936
rect 2464 3896 3516 3924
rect 2464 3884 2470 3896
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 3786 3924 3792 3936
rect 3747 3896 3792 3924
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4062 3924 4068 3936
rect 4023 3896 4068 3924
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 4433 3927 4491 3933
rect 4433 3924 4445 3927
rect 4396 3896 4445 3924
rect 4396 3884 4402 3896
rect 4433 3893 4445 3896
rect 4479 3893 4491 3927
rect 4433 3887 4491 3893
rect 4522 3884 4528 3936
rect 4580 3924 4586 3936
rect 5445 3927 5503 3933
rect 5445 3924 5457 3927
rect 4580 3896 5457 3924
rect 4580 3884 4586 3896
rect 5445 3893 5457 3896
rect 5491 3893 5503 3927
rect 5445 3887 5503 3893
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 6288 3933 6316 3964
rect 6454 3952 6460 4004
rect 6512 3992 6518 4004
rect 6638 3992 6644 4004
rect 6512 3964 6644 3992
rect 6512 3952 6518 3964
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 7006 3952 7012 4004
rect 7064 4001 7070 4004
rect 7064 3995 7128 4001
rect 7064 3961 7082 3995
rect 7116 3961 7128 3995
rect 8496 3992 8524 4159
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8996 4100 9045 4128
rect 8996 4088 9002 4100
rect 9033 4097 9045 4100
rect 9079 4128 9091 4131
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9079 4100 10057 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 9490 4060 9496 4072
rect 8720 4032 9496 4060
rect 8720 4020 8726 4032
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 9732 4032 10609 4060
rect 9732 4020 9738 4032
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 10597 4023 10655 4029
rect 10686 4020 10692 4072
rect 10744 4060 10750 4072
rect 10853 4063 10911 4069
rect 10853 4060 10865 4063
rect 10744 4032 10865 4060
rect 10744 4020 10750 4032
rect 10853 4029 10865 4032
rect 10899 4029 10911 4063
rect 10853 4023 10911 4029
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 13170 4060 13176 4072
rect 12483 4032 13176 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 13170 4020 13176 4032
rect 13228 4060 13234 4072
rect 14093 4063 14151 4069
rect 14093 4060 14105 4063
rect 13228 4032 14105 4060
rect 13228 4020 13234 4032
rect 14093 4029 14105 4032
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 15749 4063 15807 4069
rect 15749 4029 15761 4063
rect 15795 4029 15807 4063
rect 15749 4023 15807 4029
rect 11054 3992 11060 4004
rect 8496 3964 11060 3992
rect 7064 3955 7128 3961
rect 7064 3952 7070 3955
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 12682 3995 12740 4001
rect 12682 3992 12694 3995
rect 11992 3964 12694 3992
rect 6273 3927 6331 3933
rect 5592 3896 5637 3924
rect 5592 3884 5598 3896
rect 6273 3893 6285 3927
rect 6319 3893 6331 3927
rect 6273 3887 6331 3893
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 8846 3924 8852 3936
rect 7984 3896 8852 3924
rect 7984 3884 7990 3896
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9490 3924 9496 3936
rect 8996 3896 9041 3924
rect 9451 3896 9496 3924
rect 8996 3884 9002 3896
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9824 3896 9873 3924
rect 9824 3884 9830 3896
rect 9861 3893 9873 3896
rect 9907 3893 9919 3927
rect 9861 3887 9919 3893
rect 9950 3884 9956 3936
rect 10008 3924 10014 3936
rect 10008 3896 10053 3924
rect 10008 3884 10014 3896
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 11992 3933 12020 3964
rect 12682 3961 12694 3964
rect 12728 3961 12740 3995
rect 14338 3995 14396 4001
rect 14338 3992 14350 3995
rect 12682 3955 12740 3961
rect 13832 3964 14350 3992
rect 13832 3933 13860 3964
rect 14338 3961 14350 3964
rect 14384 3992 14396 3995
rect 14458 3992 14464 4004
rect 14384 3964 14464 3992
rect 14384 3961 14396 3964
rect 14338 3955 14396 3961
rect 14458 3952 14464 3964
rect 14516 3952 14522 4004
rect 15764 3992 15792 4023
rect 16022 3992 16028 4004
rect 14568 3964 15792 3992
rect 15983 3964 16028 3992
rect 11977 3927 12035 3933
rect 11977 3924 11989 3927
rect 10928 3896 11989 3924
rect 10928 3884 10934 3896
rect 11977 3893 11989 3896
rect 12023 3893 12035 3927
rect 11977 3887 12035 3893
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3893 13875 3927
rect 13817 3887 13875 3893
rect 13906 3884 13912 3936
rect 13964 3924 13970 3936
rect 14568 3924 14596 3964
rect 16022 3952 16028 3964
rect 16080 3952 16086 4004
rect 13964 3896 14596 3924
rect 13964 3884 13970 3896
rect 1104 3834 16836 3856
rect 1104 3782 6246 3834
rect 6298 3782 6310 3834
rect 6362 3782 6374 3834
rect 6426 3782 6438 3834
rect 6490 3782 11510 3834
rect 11562 3782 11574 3834
rect 11626 3782 11638 3834
rect 11690 3782 11702 3834
rect 11754 3782 16836 3834
rect 1104 3760 16836 3782
rect 1394 3680 1400 3732
rect 1452 3720 1458 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 1452 3692 2697 3720
rect 1452 3680 1458 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 4062 3720 4068 3732
rect 2823 3692 4068 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 5445 3723 5503 3729
rect 5445 3689 5457 3723
rect 5491 3689 5503 3723
rect 5445 3683 5503 3689
rect 1504 3624 3740 3652
rect 1504 3593 1532 3624
rect 1489 3587 1547 3593
rect 1489 3553 1501 3587
rect 1535 3553 1547 3587
rect 3329 3587 3387 3593
rect 3329 3584 3341 3587
rect 1489 3547 1547 3553
rect 3252 3556 3341 3584
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1673 3519 1731 3525
rect 1673 3516 1685 3519
rect 624 3488 1685 3516
rect 624 3476 630 3488
rect 1673 3485 1685 3488
rect 1719 3485 1731 3519
rect 2866 3516 2872 3528
rect 2827 3488 2872 3516
rect 1673 3479 1731 3485
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 2314 3448 2320 3460
rect 2275 3420 2320 3448
rect 2314 3408 2320 3420
rect 2372 3408 2378 3460
rect 2590 3408 2596 3460
rect 2648 3448 2654 3460
rect 3252 3448 3280 3556
rect 3329 3553 3341 3556
rect 3375 3553 3387 3587
rect 3712 3584 3740 3624
rect 3786 3612 3792 3664
rect 3844 3652 3850 3664
rect 4310 3655 4368 3661
rect 4310 3652 4322 3655
rect 3844 3624 4322 3652
rect 3844 3612 3850 3624
rect 4310 3621 4322 3624
rect 4356 3652 4368 3655
rect 5460 3652 5488 3683
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 6733 3723 6791 3729
rect 6733 3720 6745 3723
rect 5592 3692 6745 3720
rect 5592 3680 5598 3692
rect 6733 3689 6745 3692
rect 6779 3689 6791 3723
rect 8389 3723 8447 3729
rect 6733 3683 6791 3689
rect 7484 3692 8340 3720
rect 5626 3652 5632 3664
rect 4356 3624 5396 3652
rect 5460 3624 5632 3652
rect 4356 3621 4368 3624
rect 4310 3615 4368 3621
rect 5368 3584 5396 3624
rect 5626 3612 5632 3624
rect 5684 3652 5690 3664
rect 5684 3624 6316 3652
rect 5684 3612 5690 3624
rect 5810 3584 5816 3596
rect 3712 3556 5304 3584
rect 5368 3556 5816 3584
rect 3329 3547 3387 3553
rect 3510 3476 3516 3528
rect 3568 3516 3574 3528
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 3568 3488 4077 3516
rect 3568 3476 3574 3488
rect 4065 3485 4077 3488
rect 4111 3485 4123 3519
rect 5276 3516 5304 3556
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 6086 3584 6092 3596
rect 6047 3556 6092 3584
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 5350 3516 5356 3528
rect 5276 3488 5356 3516
rect 4065 3479 4123 3485
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 6288 3525 6316 3624
rect 6362 3612 6368 3664
rect 6420 3652 6426 3664
rect 7484 3652 7512 3692
rect 6420 3624 7512 3652
rect 6420 3612 6426 3624
rect 7558 3612 7564 3664
rect 7616 3652 7622 3664
rect 7616 3624 7788 3652
rect 7616 3612 7622 3624
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6880 3556 7113 3584
rect 6880 3544 6886 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 7650 3584 7656 3596
rect 7101 3547 7159 3553
rect 7208 3556 7656 3584
rect 6181 3519 6239 3525
rect 6181 3516 6193 3519
rect 5500 3488 6193 3516
rect 5500 3476 5506 3488
rect 6181 3485 6193 3488
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 7208 3525 7236 3556
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 7760 3593 7788 3624
rect 8312 3596 8340 3692
rect 8389 3689 8401 3723
rect 8435 3689 8447 3723
rect 8846 3720 8852 3732
rect 8807 3692 8852 3720
rect 8389 3683 8447 3689
rect 8404 3652 8432 3683
rect 8846 3680 8852 3692
rect 8904 3680 8910 3732
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 12250 3720 12256 3732
rect 9548 3692 12256 3720
rect 9548 3680 9554 3692
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 12713 3723 12771 3729
rect 12713 3720 12725 3723
rect 12360 3692 12725 3720
rect 12158 3652 12164 3664
rect 8404 3624 11652 3652
rect 12119 3624 12164 3652
rect 7745 3587 7803 3593
rect 7745 3553 7757 3587
rect 7791 3553 7803 3587
rect 7745 3547 7803 3553
rect 8294 3544 8300 3596
rect 8352 3544 8358 3596
rect 8757 3587 8815 3593
rect 8757 3553 8769 3587
rect 8803 3553 8815 3587
rect 8757 3547 8815 3553
rect 7193 3519 7251 3525
rect 7193 3516 7205 3519
rect 6972 3488 7205 3516
rect 6972 3476 6978 3488
rect 7193 3485 7205 3488
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3516 7435 3519
rect 7561 3519 7619 3525
rect 7561 3516 7573 3519
rect 7423 3488 7573 3516
rect 7423 3485 7435 3488
rect 7377 3479 7435 3485
rect 7561 3485 7573 3488
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 8772 3516 8800 3547
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 9582 3584 9588 3596
rect 9180 3556 9588 3584
rect 9180 3544 9186 3556
rect 9582 3544 9588 3556
rect 9640 3584 9646 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 9640 3556 10057 3584
rect 9640 3544 9646 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3584 10195 3587
rect 10318 3584 10324 3596
rect 10183 3556 10324 3584
rect 10183 3553 10195 3556
rect 10137 3547 10195 3553
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 10781 3587 10839 3593
rect 10781 3584 10793 3587
rect 10744 3556 10793 3584
rect 10744 3544 10750 3556
rect 10781 3553 10793 3556
rect 10827 3553 10839 3587
rect 10781 3547 10839 3553
rect 10962 3544 10968 3596
rect 11020 3584 11026 3596
rect 11517 3587 11575 3593
rect 11517 3584 11529 3587
rect 11020 3556 11529 3584
rect 11020 3544 11026 3556
rect 11517 3553 11529 3556
rect 11563 3553 11575 3587
rect 11624 3584 11652 3624
rect 12158 3612 12164 3624
rect 12216 3652 12222 3664
rect 12360 3652 12388 3692
rect 12713 3689 12725 3692
rect 12759 3689 12771 3723
rect 12713 3683 12771 3689
rect 12802 3680 12808 3732
rect 12860 3720 12866 3732
rect 13814 3720 13820 3732
rect 12860 3692 12905 3720
rect 13775 3692 13820 3720
rect 12860 3680 12866 3692
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 12216 3624 12388 3652
rect 12216 3612 12222 3624
rect 12434 3612 12440 3664
rect 12492 3652 12498 3664
rect 12492 3624 15332 3652
rect 12492 3612 12498 3624
rect 12618 3584 12624 3596
rect 11624 3556 12624 3584
rect 11517 3547 11575 3553
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 13262 3584 13268 3596
rect 12728 3556 13268 3584
rect 8938 3516 8944 3528
rect 8720 3488 8800 3516
rect 8899 3488 8944 3516
rect 8720 3476 8726 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 11609 3519 11667 3525
rect 10284 3488 10329 3516
rect 11072 3488 11560 3516
rect 10284 3476 10290 3488
rect 3878 3448 3884 3460
rect 2648 3420 3884 3448
rect 2648 3408 2654 3420
rect 3878 3408 3884 3420
rect 3936 3408 3942 3460
rect 7929 3451 7987 3457
rect 7929 3448 7941 3451
rect 5000 3420 7941 3448
rect 3050 3340 3056 3392
rect 3108 3380 3114 3392
rect 3513 3383 3571 3389
rect 3513 3380 3525 3383
rect 3108 3352 3525 3380
rect 3108 3340 3114 3352
rect 3513 3349 3525 3352
rect 3559 3349 3571 3383
rect 3513 3343 3571 3349
rect 4062 3340 4068 3392
rect 4120 3380 4126 3392
rect 5000 3380 5028 3420
rect 7929 3417 7941 3420
rect 7975 3417 7987 3451
rect 7929 3411 7987 3417
rect 9950 3408 9956 3460
rect 10008 3448 10014 3460
rect 11072 3448 11100 3488
rect 10008 3420 11100 3448
rect 11532 3448 11560 3488
rect 11609 3485 11621 3519
rect 11655 3516 11667 3519
rect 11698 3516 11704 3528
rect 11655 3488 11704 3516
rect 11655 3485 11667 3488
rect 11609 3479 11667 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 11793 3519 11851 3525
rect 11793 3485 11805 3519
rect 11839 3516 11851 3519
rect 11974 3516 11980 3528
rect 11839 3488 11980 3516
rect 11839 3485 11851 3488
rect 11793 3479 11851 3485
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12728 3448 12756 3556
rect 13262 3544 13268 3556
rect 13320 3584 13326 3596
rect 15304 3593 15332 3624
rect 14185 3587 14243 3593
rect 14185 3584 14197 3587
rect 13320 3556 14197 3584
rect 13320 3544 13326 3556
rect 14185 3553 14197 3556
rect 14231 3553 14243 3587
rect 14185 3547 14243 3553
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 15654 3544 15660 3596
rect 15712 3584 15718 3596
rect 16025 3587 16083 3593
rect 16025 3584 16037 3587
rect 15712 3556 16037 3584
rect 15712 3544 15718 3556
rect 16025 3553 16037 3556
rect 16071 3553 16083 3587
rect 16025 3547 16083 3553
rect 12894 3476 12900 3528
rect 12952 3516 12958 3528
rect 12952 3488 12997 3516
rect 12952 3476 12958 3488
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13780 3488 14289 3516
rect 13780 3476 13786 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 15194 3516 15200 3528
rect 14507 3488 15200 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 15473 3519 15531 3525
rect 15473 3485 15485 3519
rect 15519 3485 15531 3519
rect 15473 3479 15531 3485
rect 11532 3420 12756 3448
rect 10008 3408 10014 3420
rect 13078 3408 13084 3460
rect 13136 3448 13142 3460
rect 15488 3448 15516 3479
rect 13136 3420 15516 3448
rect 13136 3408 13142 3420
rect 5718 3380 5724 3392
rect 4120 3352 5028 3380
rect 5679 3352 5724 3380
rect 4120 3340 4126 3352
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 7561 3383 7619 3389
rect 7561 3380 7573 3383
rect 5868 3352 7573 3380
rect 5868 3340 5874 3352
rect 7561 3349 7573 3352
rect 7607 3349 7619 3383
rect 7561 3343 7619 3349
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 9306 3380 9312 3392
rect 7708 3352 9312 3380
rect 7708 3340 7714 3352
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9674 3380 9680 3392
rect 9635 3352 9680 3380
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 10962 3380 10968 3392
rect 10923 3352 10968 3380
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 12342 3380 12348 3392
rect 11204 3352 11249 3380
rect 12303 3352 12348 3380
rect 11204 3340 11210 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 15102 3340 15108 3392
rect 15160 3380 15166 3392
rect 16209 3383 16267 3389
rect 16209 3380 16221 3383
rect 15160 3352 16221 3380
rect 15160 3340 15166 3352
rect 16209 3349 16221 3352
rect 16255 3349 16267 3383
rect 16209 3343 16267 3349
rect 1104 3290 16836 3312
rect 1104 3238 3614 3290
rect 3666 3238 3678 3290
rect 3730 3238 3742 3290
rect 3794 3238 3806 3290
rect 3858 3238 8878 3290
rect 8930 3238 8942 3290
rect 8994 3238 9006 3290
rect 9058 3238 9070 3290
rect 9122 3238 14142 3290
rect 14194 3238 14206 3290
rect 14258 3238 14270 3290
rect 14322 3238 14334 3290
rect 14386 3238 16836 3290
rect 1104 3216 16836 3238
rect 2222 3176 2228 3188
rect 2183 3148 2228 3176
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 3237 3179 3295 3185
rect 3237 3145 3249 3179
rect 3283 3176 3295 3179
rect 3326 3176 3332 3188
rect 3283 3148 3332 3176
rect 3283 3145 3295 3148
rect 3237 3139 3295 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 4249 3179 4307 3185
rect 4249 3176 4261 3179
rect 4212 3148 4261 3176
rect 4212 3136 4218 3148
rect 4249 3145 4261 3148
rect 4295 3145 4307 3179
rect 4249 3139 4307 3145
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 4982 3176 4988 3188
rect 4672 3148 4988 3176
rect 4672 3136 4678 3148
rect 4982 3136 4988 3148
rect 5040 3176 5046 3188
rect 7193 3179 7251 3185
rect 7193 3176 7205 3179
rect 5040 3148 7205 3176
rect 5040 3136 5046 3148
rect 7193 3145 7205 3148
rect 7239 3145 7251 3179
rect 7193 3139 7251 3145
rect 7742 3136 7748 3188
rect 7800 3176 7806 3188
rect 9125 3179 9183 3185
rect 9125 3176 9137 3179
rect 7800 3148 9137 3176
rect 7800 3136 7806 3148
rect 9125 3145 9137 3148
rect 9171 3145 9183 3179
rect 9306 3176 9312 3188
rect 9267 3148 9312 3176
rect 9125 3139 9183 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9582 3136 9588 3188
rect 9640 3176 9646 3188
rect 9858 3176 9864 3188
rect 9640 3148 9864 3176
rect 9640 3136 9646 3148
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 10870 3176 10876 3188
rect 10796 3148 10876 3176
rect 5442 3068 5448 3120
rect 5500 3108 5506 3120
rect 7006 3108 7012 3120
rect 5500 3080 5545 3108
rect 5736 3080 7012 3108
rect 5500 3068 5506 3080
rect 2682 3000 2688 3052
rect 2740 3040 2746 3052
rect 2777 3043 2835 3049
rect 2777 3040 2789 3043
rect 2740 3012 2789 3040
rect 2740 3000 2746 3012
rect 2777 3009 2789 3012
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 2958 3000 2964 3052
rect 3016 3040 3022 3052
rect 3881 3043 3939 3049
rect 3016 3012 3648 3040
rect 3016 3000 3022 3012
rect 3620 2981 3648 3012
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 4614 3040 4620 3052
rect 3927 3012 4620 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3040 4951 3043
rect 5736 3040 5764 3080
rect 7006 3068 7012 3080
rect 7064 3068 7070 3120
rect 10594 3108 10600 3120
rect 7668 3080 10600 3108
rect 4939 3012 5764 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 5994 3040 6000 3052
rect 5868 3012 6000 3040
rect 5868 3000 5874 3012
rect 5994 3000 6000 3012
rect 6052 3000 6058 3052
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3040 7251 3043
rect 7558 3040 7564 3052
rect 7239 3012 7564 3040
rect 7239 3009 7251 3012
rect 7193 3003 7251 3009
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 1489 2975 1547 2981
rect 1489 2941 1501 2975
rect 1535 2972 1547 2975
rect 3605 2975 3663 2981
rect 1535 2944 3464 2972
rect 1535 2941 1547 2944
rect 1489 2935 1547 2941
rect 1762 2904 1768 2916
rect 1723 2876 1768 2904
rect 1762 2864 1768 2876
rect 1820 2864 1826 2916
rect 2593 2907 2651 2913
rect 2593 2873 2605 2907
rect 2639 2904 2651 2907
rect 3326 2904 3332 2916
rect 2639 2876 3332 2904
rect 2639 2873 2651 2876
rect 2593 2867 2651 2873
rect 3326 2864 3332 2876
rect 3384 2864 3390 2916
rect 2682 2836 2688 2848
rect 2643 2808 2688 2836
rect 2682 2796 2688 2808
rect 2740 2796 2746 2848
rect 3436 2836 3464 2944
rect 3605 2941 3617 2975
rect 3651 2941 3663 2975
rect 3605 2935 3663 2941
rect 3697 2975 3755 2981
rect 3697 2941 3709 2975
rect 3743 2972 3755 2975
rect 5534 2972 5540 2984
rect 3743 2944 5540 2972
rect 3743 2941 3755 2944
rect 3697 2935 3755 2941
rect 5534 2932 5540 2944
rect 5592 2932 5598 2984
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6696 2944 6837 2972
rect 6696 2932 6702 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 7374 2972 7380 2984
rect 6825 2935 6883 2941
rect 7199 2944 7380 2972
rect 4430 2864 4436 2916
rect 4488 2904 4494 2916
rect 4709 2907 4767 2913
rect 4709 2904 4721 2907
rect 4488 2876 4721 2904
rect 4488 2864 4494 2876
rect 4709 2873 4721 2876
rect 4755 2873 4767 2907
rect 4709 2867 4767 2873
rect 5442 2864 5448 2916
rect 5500 2904 5506 2916
rect 5905 2907 5963 2913
rect 5905 2904 5917 2907
rect 5500 2876 5917 2904
rect 5500 2864 5506 2876
rect 5905 2873 5917 2876
rect 5951 2904 5963 2907
rect 6362 2904 6368 2916
rect 5951 2876 6368 2904
rect 5951 2873 5963 2876
rect 5905 2867 5963 2873
rect 6362 2864 6368 2876
rect 6420 2864 6426 2916
rect 4338 2836 4344 2848
rect 3436 2808 4344 2836
rect 4338 2796 4344 2808
rect 4396 2796 4402 2848
rect 4614 2836 4620 2848
rect 4575 2808 4620 2836
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 5350 2796 5356 2848
rect 5408 2836 5414 2848
rect 5813 2839 5871 2845
rect 5813 2836 5825 2839
rect 5408 2808 5825 2836
rect 5408 2796 5414 2808
rect 5813 2805 5825 2808
rect 5859 2805 5871 2839
rect 5813 2799 5871 2805
rect 6638 2796 6644 2848
rect 6696 2836 6702 2848
rect 7199 2836 7227 2944
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 7668 2981 7696 3080
rect 10594 3068 10600 3080
rect 10652 3068 10658 3120
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3040 7987 3043
rect 8018 3040 8024 3052
rect 7975 3012 8024 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 8754 3040 8760 3052
rect 8715 3012 8760 3040
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3040 8999 3043
rect 9030 3040 9036 3052
rect 8987 3012 9036 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9171 3012 9873 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 10796 3040 10824 3148
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11330 3176 11336 3188
rect 11291 3148 11336 3176
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 11514 3136 11520 3188
rect 11572 3176 11578 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 11572 3148 12449 3176
rect 11572 3136 11578 3148
rect 12437 3145 12449 3148
rect 12483 3145 12495 3179
rect 13722 3176 13728 3188
rect 13683 3148 13728 3176
rect 12437 3139 12495 3145
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 10796 3012 10885 3040
rect 9861 3003 9919 3009
rect 10873 3009 10885 3012
rect 10919 3009 10931 3043
rect 11790 3040 11796 3052
rect 11751 3012 11796 3040
rect 10873 3003 10931 3009
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 11974 3040 11980 3052
rect 11935 3012 11980 3040
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 12894 3000 12900 3052
rect 12952 3040 12958 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12952 3012 13001 3040
rect 12952 3000 12958 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 14185 3043 14243 3049
rect 14185 3040 14197 3043
rect 13872 3012 14197 3040
rect 13872 3000 13878 3012
rect 14185 3009 14197 3012
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3040 14427 3043
rect 14458 3040 14464 3052
rect 14415 3012 14464 3040
rect 14415 3009 14427 3012
rect 14369 3003 14427 3009
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 14642 3000 14648 3052
rect 14700 3040 14706 3052
rect 14700 3012 15516 3040
rect 14700 3000 14706 3012
rect 7653 2975 7711 2981
rect 7653 2941 7665 2975
rect 7699 2941 7711 2975
rect 7653 2935 7711 2941
rect 7745 2975 7803 2981
rect 7745 2941 7757 2975
rect 7791 2972 7803 2975
rect 10594 2972 10600 2984
rect 7791 2944 10600 2972
rect 7791 2941 7803 2944
rect 7745 2935 7803 2941
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 10689 2975 10747 2981
rect 10689 2941 10701 2975
rect 10735 2972 10747 2975
rect 11238 2972 11244 2984
rect 10735 2944 11244 2972
rect 10735 2941 10747 2944
rect 10689 2935 10747 2941
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 11348 2944 12296 2972
rect 9769 2907 9827 2913
rect 9769 2904 9781 2907
rect 7300 2876 9781 2904
rect 7300 2845 7328 2876
rect 9769 2873 9781 2876
rect 9815 2873 9827 2907
rect 9769 2867 9827 2873
rect 10042 2864 10048 2916
rect 10100 2904 10106 2916
rect 10410 2904 10416 2916
rect 10100 2876 10416 2904
rect 10100 2864 10106 2876
rect 10410 2864 10416 2876
rect 10468 2904 10474 2916
rect 11348 2904 11376 2944
rect 10468 2876 11376 2904
rect 11701 2907 11759 2913
rect 10468 2864 10474 2876
rect 11701 2873 11713 2907
rect 11747 2904 11759 2907
rect 11882 2904 11888 2916
rect 11747 2876 11888 2904
rect 11747 2873 11759 2876
rect 11701 2867 11759 2873
rect 11882 2864 11888 2876
rect 11940 2864 11946 2916
rect 6696 2808 7227 2836
rect 7285 2839 7343 2845
rect 6696 2796 6702 2808
rect 7285 2805 7297 2839
rect 7331 2805 7343 2839
rect 7285 2799 7343 2805
rect 8297 2839 8355 2845
rect 8297 2805 8309 2839
rect 8343 2836 8355 2839
rect 8570 2836 8576 2848
rect 8343 2808 8576 2836
rect 8343 2805 8355 2808
rect 8297 2799 8355 2805
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 8665 2839 8723 2845
rect 8665 2805 8677 2839
rect 8711 2836 8723 2839
rect 9582 2836 9588 2848
rect 8711 2808 9588 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 9677 2839 9735 2845
rect 9677 2805 9689 2839
rect 9723 2836 9735 2839
rect 9950 2836 9956 2848
rect 9723 2808 9956 2836
rect 9723 2805 9735 2808
rect 9677 2799 9735 2805
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 10318 2836 10324 2848
rect 10279 2808 10324 2836
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 10502 2796 10508 2848
rect 10560 2836 10566 2848
rect 10781 2839 10839 2845
rect 10781 2836 10793 2839
rect 10560 2808 10793 2836
rect 10560 2796 10566 2808
rect 10781 2805 10793 2808
rect 10827 2805 10839 2839
rect 12268 2836 12296 2944
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 12492 2944 12817 2972
rect 12492 2932 12498 2944
rect 12805 2941 12817 2944
rect 12851 2941 12863 2975
rect 12805 2935 12863 2941
rect 13170 2932 13176 2984
rect 13228 2972 13234 2984
rect 15488 2981 15516 3012
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 13228 2944 14749 2972
rect 13228 2932 13234 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 15473 2975 15531 2981
rect 15473 2941 15485 2975
rect 15519 2941 15531 2975
rect 15473 2935 15531 2941
rect 12618 2864 12624 2916
rect 12676 2904 12682 2916
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 12676 2876 12909 2904
rect 12676 2864 12682 2876
rect 12897 2873 12909 2876
rect 12943 2873 12955 2907
rect 12897 2867 12955 2873
rect 15013 2907 15071 2913
rect 15013 2873 15025 2907
rect 15059 2904 15071 2907
rect 15194 2904 15200 2916
rect 15059 2876 15200 2904
rect 15059 2873 15071 2876
rect 15013 2867 15071 2873
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 15749 2907 15807 2913
rect 15749 2873 15761 2907
rect 15795 2904 15807 2907
rect 16298 2904 16304 2916
rect 15795 2876 16304 2904
rect 15795 2873 15807 2876
rect 15749 2867 15807 2873
rect 16298 2864 16304 2876
rect 16356 2864 16362 2916
rect 14093 2839 14151 2845
rect 14093 2836 14105 2839
rect 12268 2808 14105 2836
rect 10781 2799 10839 2805
rect 14093 2805 14105 2808
rect 14139 2805 14151 2839
rect 14093 2799 14151 2805
rect 1104 2746 16836 2768
rect 1104 2694 6246 2746
rect 6298 2694 6310 2746
rect 6362 2694 6374 2746
rect 6426 2694 6438 2746
rect 6490 2694 11510 2746
rect 11562 2694 11574 2746
rect 11626 2694 11638 2746
rect 11690 2694 11702 2746
rect 11754 2694 16836 2746
rect 1104 2672 16836 2694
rect 2961 2635 3019 2641
rect 2961 2601 2973 2635
rect 3007 2632 3019 2635
rect 4246 2632 4252 2644
rect 3007 2604 4252 2632
rect 3007 2601 3019 2604
rect 2961 2595 3019 2601
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4430 2632 4436 2644
rect 4391 2604 4436 2632
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 4801 2635 4859 2641
rect 4801 2601 4813 2635
rect 4847 2632 4859 2635
rect 5074 2632 5080 2644
rect 4847 2604 5080 2632
rect 4847 2601 4859 2604
rect 4801 2595 4859 2601
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 5905 2635 5963 2641
rect 5905 2632 5917 2635
rect 5684 2604 5917 2632
rect 5684 2592 5690 2604
rect 5905 2601 5917 2604
rect 5951 2632 5963 2635
rect 6917 2635 6975 2641
rect 6917 2632 6929 2635
rect 5951 2604 6929 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 6917 2601 6929 2604
rect 6963 2601 6975 2635
rect 6917 2595 6975 2601
rect 7101 2635 7159 2641
rect 7101 2601 7113 2635
rect 7147 2632 7159 2635
rect 7190 2632 7196 2644
rect 7147 2604 7196 2632
rect 7147 2601 7159 2604
rect 7101 2595 7159 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 7466 2632 7472 2644
rect 7427 2604 7472 2632
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 9950 2632 9956 2644
rect 9815 2604 9956 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10781 2635 10839 2641
rect 10781 2632 10793 2635
rect 10275 2604 10793 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10781 2601 10793 2604
rect 10827 2601 10839 2635
rect 10781 2595 10839 2601
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 11112 2604 11161 2632
rect 11112 2592 11118 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 11149 2595 11207 2601
rect 11330 2592 11336 2644
rect 11388 2632 11394 2644
rect 12621 2635 12679 2641
rect 12621 2632 12633 2635
rect 11388 2604 12633 2632
rect 11388 2592 11394 2604
rect 12621 2601 12633 2604
rect 12667 2601 12679 2635
rect 12621 2595 12679 2601
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 13081 2635 13139 2641
rect 13081 2632 13093 2635
rect 12768 2604 13093 2632
rect 12768 2592 12774 2604
rect 13081 2601 13093 2604
rect 13127 2601 13139 2635
rect 13081 2595 13139 2601
rect 3142 2564 3148 2576
rect 1504 2536 3148 2564
rect 1504 2505 1532 2536
rect 3142 2524 3148 2536
rect 3200 2524 3206 2576
rect 4893 2567 4951 2573
rect 4893 2533 4905 2567
rect 4939 2564 4951 2567
rect 5718 2564 5724 2576
rect 4939 2536 5724 2564
rect 4939 2533 4951 2536
rect 4893 2527 4951 2533
rect 5718 2524 5724 2536
rect 5776 2524 5782 2576
rect 5810 2524 5816 2576
rect 5868 2564 5874 2576
rect 7561 2567 7619 2573
rect 7561 2564 7573 2567
rect 5868 2536 5913 2564
rect 7116 2536 7573 2564
rect 5868 2524 5874 2536
rect 7116 2508 7144 2536
rect 7561 2533 7573 2536
rect 7607 2533 7619 2567
rect 7561 2527 7619 2533
rect 8573 2567 8631 2573
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 9674 2564 9680 2576
rect 8619 2536 9680 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 11241 2567 11299 2573
rect 11241 2533 11253 2567
rect 11287 2564 11299 2567
rect 11974 2564 11980 2576
rect 11287 2536 11980 2564
rect 11287 2533 11299 2536
rect 11241 2527 11299 2533
rect 11974 2524 11980 2536
rect 12032 2524 12038 2576
rect 12342 2564 12348 2576
rect 12084 2536 12348 2564
rect 1489 2499 1547 2505
rect 1489 2465 1501 2499
rect 1535 2465 1547 2499
rect 1489 2459 1547 2465
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2465 2283 2499
rect 3326 2496 3332 2508
rect 3287 2468 3332 2496
rect 2225 2459 2283 2465
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 2240 2292 2268 2459
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 6638 2496 6644 2508
rect 3467 2468 6644 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 6638 2456 6644 2468
rect 6696 2456 6702 2508
rect 7098 2456 7104 2508
rect 7156 2456 7162 2508
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 7484 2468 8493 2496
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 2516 2360 2544 2391
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 3292 2400 3525 2428
rect 3292 2388 3298 2400
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 5258 2428 5264 2440
rect 5123 2400 5264 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5994 2428 6000 2440
rect 5955 2400 6000 2428
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7484 2428 7512 2468
rect 8481 2465 8493 2468
rect 8527 2496 8539 2499
rect 9125 2499 9183 2505
rect 8527 2468 8984 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 6963 2400 7512 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 7616 2400 7757 2428
rect 7616 2388 7622 2400
rect 7745 2397 7757 2400
rect 7791 2428 7803 2431
rect 8757 2431 8815 2437
rect 8757 2428 8769 2431
rect 7791 2400 8769 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 8757 2397 8769 2400
rect 8803 2428 8815 2431
rect 8846 2428 8852 2440
rect 8803 2400 8852 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 8956 2428 8984 2468
rect 9125 2465 9137 2499
rect 9171 2496 9183 2499
rect 9950 2496 9956 2508
rect 9171 2468 9956 2496
rect 9171 2465 9183 2468
rect 9125 2459 9183 2465
rect 9950 2456 9956 2468
rect 10008 2456 10014 2508
rect 10137 2499 10195 2505
rect 10137 2465 10149 2499
rect 10183 2496 10195 2499
rect 11790 2496 11796 2508
rect 10183 2468 11468 2496
rect 11751 2468 11796 2496
rect 10183 2465 10195 2468
rect 10137 2459 10195 2465
rect 9766 2428 9772 2440
rect 8956 2400 9772 2428
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 11330 2428 11336 2440
rect 10321 2391 10379 2397
rect 10612 2400 11336 2428
rect 3142 2360 3148 2372
rect 2516 2332 3148 2360
rect 3142 2320 3148 2332
rect 3200 2320 3206 2372
rect 5445 2363 5503 2369
rect 5445 2329 5457 2363
rect 5491 2360 5503 2363
rect 6086 2360 6092 2372
rect 5491 2332 6092 2360
rect 5491 2329 5503 2332
rect 5445 2323 5503 2329
rect 6086 2320 6092 2332
rect 6144 2320 6150 2372
rect 6546 2320 6552 2372
rect 6604 2360 6610 2372
rect 8113 2363 8171 2369
rect 8113 2360 8125 2363
rect 6604 2332 8125 2360
rect 6604 2320 6610 2332
rect 8113 2329 8125 2332
rect 8159 2329 8171 2363
rect 8113 2323 8171 2329
rect 8202 2320 8208 2372
rect 8260 2360 8266 2372
rect 10336 2360 10364 2391
rect 8260 2332 10364 2360
rect 8260 2320 8266 2332
rect 4890 2292 4896 2304
rect 2240 2264 4896 2292
rect 4890 2252 4896 2264
rect 4948 2252 4954 2304
rect 6914 2252 6920 2304
rect 6972 2292 6978 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 6972 2264 9321 2292
rect 6972 2252 6978 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 9398 2252 9404 2304
rect 9456 2292 9462 2304
rect 10612 2292 10640 2400
rect 11330 2388 11336 2400
rect 11388 2388 11394 2440
rect 11440 2428 11468 2468
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 12084 2496 12112 2536
rect 12342 2524 12348 2536
rect 12400 2524 12406 2576
rect 12526 2524 12532 2576
rect 12584 2564 12590 2576
rect 14645 2567 14703 2573
rect 12584 2536 13676 2564
rect 12584 2524 12590 2536
rect 11900 2468 12112 2496
rect 11900 2428 11928 2468
rect 12250 2456 12256 2508
rect 12308 2496 12314 2508
rect 13648 2505 13676 2536
rect 14645 2533 14657 2567
rect 14691 2564 14703 2567
rect 17402 2564 17408 2576
rect 14691 2536 17408 2564
rect 14691 2533 14703 2536
rect 14645 2527 14703 2533
rect 17402 2524 17408 2536
rect 17460 2524 17466 2576
rect 12989 2499 13047 2505
rect 12989 2496 13001 2499
rect 12308 2468 13001 2496
rect 12308 2456 12314 2468
rect 12989 2465 13001 2468
rect 13035 2465 13047 2499
rect 12989 2459 13047 2465
rect 13633 2499 13691 2505
rect 13633 2465 13645 2499
rect 13679 2465 13691 2499
rect 13633 2459 13691 2465
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2496 14427 2499
rect 14550 2496 14556 2508
rect 14415 2468 14556 2496
rect 14415 2465 14427 2468
rect 14369 2459 14427 2465
rect 14550 2456 14556 2468
rect 14608 2456 14614 2508
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15436 2468 15485 2496
rect 15436 2456 15442 2468
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 11440 2400 11928 2428
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2397 13231 2431
rect 13814 2428 13820 2440
rect 13775 2400 13820 2428
rect 13173 2391 13231 2397
rect 10686 2320 10692 2372
rect 10744 2360 10750 2372
rect 11992 2360 12020 2391
rect 10744 2332 12020 2360
rect 10744 2320 10750 2332
rect 12802 2320 12808 2372
rect 12860 2360 12866 2372
rect 13188 2360 13216 2391
rect 13814 2388 13820 2400
rect 13872 2388 13878 2440
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 12860 2332 13216 2360
rect 12860 2320 12866 2332
rect 14458 2320 14464 2372
rect 14516 2360 14522 2372
rect 15672 2360 15700 2391
rect 14516 2332 15700 2360
rect 14516 2320 14522 2332
rect 9456 2264 10640 2292
rect 9456 2252 9462 2264
rect 1104 2202 16836 2224
rect 1104 2150 3614 2202
rect 3666 2150 3678 2202
rect 3730 2150 3742 2202
rect 3794 2150 3806 2202
rect 3858 2150 8878 2202
rect 8930 2150 8942 2202
rect 8994 2150 9006 2202
rect 9058 2150 9070 2202
rect 9122 2150 14142 2202
rect 14194 2150 14206 2202
rect 14258 2150 14270 2202
rect 14322 2150 14334 2202
rect 14386 2150 16836 2202
rect 1104 2128 16836 2150
rect 3234 2048 3240 2100
rect 3292 2088 3298 2100
rect 5166 2088 5172 2100
rect 3292 2060 5172 2088
rect 3292 2048 3298 2060
rect 5166 2048 5172 2060
rect 5224 2048 5230 2100
rect 10134 2088 10140 2100
rect 6104 2060 10140 2088
rect 3326 1980 3332 2032
rect 3384 2020 3390 2032
rect 6104 2020 6132 2060
rect 10134 2048 10140 2060
rect 10192 2048 10198 2100
rect 11330 2048 11336 2100
rect 11388 2088 11394 2100
rect 12802 2088 12808 2100
rect 11388 2060 12808 2088
rect 11388 2048 11394 2060
rect 12802 2048 12808 2060
rect 12860 2048 12866 2100
rect 3384 1992 6132 2020
rect 3384 1980 3390 1992
rect 3142 1912 3148 1964
rect 3200 1952 3206 1964
rect 6178 1952 6184 1964
rect 3200 1924 6184 1952
rect 3200 1912 3206 1924
rect 6178 1912 6184 1924
rect 6236 1912 6242 1964
rect 9582 1368 9588 1420
rect 9640 1408 9646 1420
rect 13814 1408 13820 1420
rect 9640 1380 13820 1408
rect 9640 1368 9646 1380
rect 13814 1368 13820 1380
rect 13872 1368 13878 1420
rect 3418 1300 3424 1352
rect 3476 1340 3482 1352
rect 6914 1340 6920 1352
rect 3476 1312 6920 1340
rect 3476 1300 3482 1312
rect 6914 1300 6920 1312
rect 6972 1300 6978 1352
rect 11790 1096 11796 1148
rect 11848 1136 11854 1148
rect 16022 1136 16028 1148
rect 11848 1108 16028 1136
rect 11848 1096 11854 1108
rect 16022 1096 16028 1108
rect 16080 1096 16086 1148
rect 1762 620 1768 672
rect 1820 660 1826 672
rect 5074 660 5080 672
rect 1820 632 5080 660
rect 1820 620 1826 632
rect 5074 620 5080 632
rect 5132 620 5138 672
<< via1 >>
rect 4068 15172 4120 15224
rect 9956 15172 10008 15224
rect 2228 14968 2280 15020
rect 6552 14968 6604 15020
rect 9404 14968 9456 15020
rect 15108 14968 15160 15020
rect 4068 14900 4120 14952
rect 10140 14900 10192 14952
rect 4160 14832 4212 14884
rect 14648 14832 14700 14884
rect 3516 14764 3568 14816
rect 9496 14764 9548 14816
rect 12808 14764 12860 14816
rect 14096 14764 14148 14816
rect 6246 14662 6298 14714
rect 6310 14662 6362 14714
rect 6374 14662 6426 14714
rect 6438 14662 6490 14714
rect 11510 14662 11562 14714
rect 11574 14662 11626 14714
rect 11638 14662 11690 14714
rect 11702 14662 11754 14714
rect 4160 14603 4212 14612
rect 4160 14569 4169 14603
rect 4169 14569 4203 14603
rect 4203 14569 4212 14603
rect 4160 14560 4212 14569
rect 8300 14560 8352 14612
rect 10692 14603 10744 14612
rect 10692 14569 10701 14603
rect 10701 14569 10735 14603
rect 10735 14569 10744 14603
rect 10692 14560 10744 14569
rect 13728 14560 13780 14612
rect 1400 14492 1452 14544
rect 13360 14492 13412 14544
rect 15752 14492 15804 14544
rect 2412 14467 2464 14476
rect 2412 14433 2421 14467
rect 2421 14433 2455 14467
rect 2455 14433 2464 14467
rect 2412 14424 2464 14433
rect 4160 14424 4212 14476
rect 5540 14467 5592 14476
rect 5540 14433 5549 14467
rect 5549 14433 5583 14467
rect 5583 14433 5592 14467
rect 5540 14424 5592 14433
rect 6092 14424 6144 14476
rect 8576 14424 8628 14476
rect 8668 14424 8720 14476
rect 9680 14424 9732 14476
rect 12164 14424 12216 14476
rect 12992 14424 13044 14476
rect 14004 14467 14056 14476
rect 14004 14433 14013 14467
rect 14013 14433 14047 14467
rect 14047 14433 14056 14467
rect 14004 14424 14056 14433
rect 14096 14467 14148 14476
rect 14096 14433 14105 14467
rect 14105 14433 14139 14467
rect 14139 14433 14148 14467
rect 14648 14467 14700 14476
rect 14096 14424 14148 14433
rect 14648 14433 14657 14467
rect 14657 14433 14691 14467
rect 14691 14433 14700 14467
rect 14648 14424 14700 14433
rect 2596 14399 2648 14408
rect 2596 14365 2605 14399
rect 2605 14365 2639 14399
rect 2639 14365 2648 14399
rect 2596 14356 2648 14365
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 5724 14399 5776 14408
rect 4344 14288 4396 14340
rect 5724 14365 5733 14399
rect 5733 14365 5767 14399
rect 5767 14365 5776 14399
rect 5724 14356 5776 14365
rect 7104 14356 7156 14408
rect 3424 14220 3476 14272
rect 4068 14220 4120 14272
rect 6644 14288 6696 14340
rect 8760 14356 8812 14408
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 11980 14288 12032 14340
rect 13820 14356 13872 14408
rect 13636 14288 13688 14340
rect 15384 14356 15436 14408
rect 16120 14399 16172 14408
rect 16120 14365 16129 14399
rect 16129 14365 16163 14399
rect 16163 14365 16172 14399
rect 16120 14356 16172 14365
rect 4988 14220 5040 14272
rect 7380 14220 7432 14272
rect 8392 14220 8444 14272
rect 10048 14220 10100 14272
rect 11060 14220 11112 14272
rect 12624 14263 12676 14272
rect 12624 14229 12633 14263
rect 12633 14229 12667 14263
rect 12667 14229 12676 14263
rect 12624 14220 12676 14229
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 3614 14118 3666 14170
rect 3678 14118 3730 14170
rect 3742 14118 3794 14170
rect 3806 14118 3858 14170
rect 8878 14118 8930 14170
rect 8942 14118 8994 14170
rect 9006 14118 9058 14170
rect 9070 14118 9122 14170
rect 14142 14118 14194 14170
rect 14206 14118 14258 14170
rect 14270 14118 14322 14170
rect 14334 14118 14386 14170
rect 4160 14059 4212 14068
rect 4160 14025 4169 14059
rect 4169 14025 4203 14059
rect 4203 14025 4212 14059
rect 4160 14016 4212 14025
rect 4252 14016 4304 14068
rect 5724 14016 5776 14068
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 5540 13948 5592 14000
rect 4804 13923 4856 13932
rect 2504 13855 2556 13864
rect 2504 13821 2513 13855
rect 2513 13821 2547 13855
rect 2547 13821 2556 13855
rect 2504 13812 2556 13821
rect 3148 13812 3200 13864
rect 4804 13889 4813 13923
rect 4813 13889 4847 13923
rect 4847 13889 4856 13923
rect 4804 13880 4856 13889
rect 5356 13880 5408 13932
rect 8668 14059 8720 14068
rect 8668 14025 8677 14059
rect 8677 14025 8711 14059
rect 8711 14025 8720 14059
rect 8668 14016 8720 14025
rect 6828 13923 6880 13932
rect 6828 13889 6837 13923
rect 6837 13889 6871 13923
rect 6871 13889 6880 13923
rect 6828 13880 6880 13889
rect 12808 14016 12860 14068
rect 13084 14016 13136 14068
rect 15384 14059 15436 14068
rect 15384 14025 15393 14059
rect 15393 14025 15427 14059
rect 15427 14025 15436 14059
rect 15384 14016 15436 14025
rect 9588 13948 9640 14000
rect 12440 13948 12492 14000
rect 13820 13991 13872 14000
rect 13820 13957 13829 13991
rect 13829 13957 13863 13991
rect 13863 13957 13872 13991
rect 13820 13948 13872 13957
rect 9312 13923 9364 13932
rect 3424 13787 3476 13796
rect 3424 13753 3433 13787
rect 3433 13753 3467 13787
rect 3467 13753 3476 13787
rect 3424 13744 3476 13753
rect 2688 13676 2740 13728
rect 4620 13719 4672 13728
rect 4620 13685 4629 13719
rect 4629 13685 4663 13719
rect 4663 13685 4672 13719
rect 4620 13676 4672 13685
rect 5264 13744 5316 13796
rect 7104 13855 7156 13864
rect 7104 13821 7138 13855
rect 7138 13821 7156 13855
rect 7104 13812 7156 13821
rect 9312 13889 9321 13923
rect 9321 13889 9355 13923
rect 9355 13889 9364 13923
rect 9312 13880 9364 13889
rect 9864 13880 9916 13932
rect 10784 13880 10836 13932
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 13636 13880 13688 13932
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 8668 13812 8720 13864
rect 9404 13812 9456 13864
rect 9220 13744 9272 13796
rect 12348 13812 12400 13864
rect 12716 13787 12768 13796
rect 9772 13676 9824 13728
rect 10600 13676 10652 13728
rect 11888 13676 11940 13728
rect 12716 13753 12750 13787
rect 12750 13753 12768 13787
rect 12716 13744 12768 13753
rect 13268 13812 13320 13864
rect 14004 13744 14056 13796
rect 14740 13812 14792 13864
rect 13452 13676 13504 13728
rect 13544 13676 13596 13728
rect 15660 13676 15712 13728
rect 6246 13574 6298 13626
rect 6310 13574 6362 13626
rect 6374 13574 6426 13626
rect 6438 13574 6490 13626
rect 11510 13574 11562 13626
rect 11574 13574 11626 13626
rect 11638 13574 11690 13626
rect 11702 13574 11754 13626
rect 2688 13404 2740 13456
rect 2964 13336 3016 13388
rect 3516 13132 3568 13184
rect 4620 13472 4672 13524
rect 7104 13515 7156 13524
rect 3976 13404 4028 13456
rect 6736 13404 6788 13456
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 7288 13472 7340 13524
rect 8392 13472 8444 13524
rect 9680 13515 9732 13524
rect 9680 13481 9689 13515
rect 9689 13481 9723 13515
rect 9723 13481 9732 13515
rect 9680 13472 9732 13481
rect 9956 13472 10008 13524
rect 10508 13472 10560 13524
rect 12440 13472 12492 13524
rect 12624 13472 12676 13524
rect 13452 13472 13504 13524
rect 14464 13472 14516 13524
rect 15016 13472 15068 13524
rect 7840 13404 7892 13456
rect 8300 13404 8352 13456
rect 5816 13336 5868 13388
rect 8576 13336 8628 13388
rect 9496 13336 9548 13388
rect 3976 13268 4028 13320
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 5356 13311 5408 13320
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 5632 13268 5684 13320
rect 8208 13311 8260 13320
rect 8208 13277 8217 13311
rect 8217 13277 8251 13311
rect 8251 13277 8260 13311
rect 8208 13268 8260 13277
rect 9680 13268 9732 13320
rect 9864 13268 9916 13320
rect 11980 13404 12032 13456
rect 12256 13336 12308 13388
rect 12348 13336 12400 13388
rect 12440 13336 12492 13388
rect 12624 13336 12676 13388
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 11152 13200 11204 13252
rect 15016 13336 15068 13388
rect 15200 13336 15252 13388
rect 16120 13311 16172 13320
rect 7104 13132 7156 13184
rect 9404 13132 9456 13184
rect 9864 13132 9916 13184
rect 10140 13132 10192 13184
rect 10232 13132 10284 13184
rect 11428 13132 11480 13184
rect 12716 13200 12768 13252
rect 13636 13200 13688 13252
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 12900 13175 12952 13184
rect 12900 13141 12909 13175
rect 12909 13141 12943 13175
rect 12943 13141 12952 13175
rect 12900 13132 12952 13141
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 3614 13030 3666 13082
rect 3678 13030 3730 13082
rect 3742 13030 3794 13082
rect 3806 13030 3858 13082
rect 8878 13030 8930 13082
rect 8942 13030 8994 13082
rect 9006 13030 9058 13082
rect 9070 13030 9122 13082
rect 14142 13030 14194 13082
rect 14206 13030 14258 13082
rect 14270 13030 14322 13082
rect 14334 13030 14386 13082
rect 4344 12971 4396 12980
rect 4344 12937 4353 12971
rect 4353 12937 4387 12971
rect 4387 12937 4396 12971
rect 4344 12928 4396 12937
rect 4712 12971 4764 12980
rect 4712 12937 4721 12971
rect 4721 12937 4755 12971
rect 4755 12937 4764 12971
rect 4712 12928 4764 12937
rect 4896 12928 4948 12980
rect 2596 12835 2648 12844
rect 2596 12801 2605 12835
rect 2605 12801 2639 12835
rect 2639 12801 2648 12835
rect 2596 12792 2648 12801
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 2320 12767 2372 12776
rect 2320 12733 2329 12767
rect 2329 12733 2363 12767
rect 2363 12733 2372 12767
rect 2320 12724 2372 12733
rect 3516 12724 3568 12776
rect 4804 12792 4856 12844
rect 5816 12928 5868 12980
rect 11888 12928 11940 12980
rect 8760 12903 8812 12912
rect 8760 12869 8769 12903
rect 8769 12869 8803 12903
rect 8803 12869 8812 12903
rect 8760 12860 8812 12869
rect 9864 12860 9916 12912
rect 6920 12792 6972 12844
rect 7472 12724 7524 12776
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 9404 12792 9456 12844
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 10324 12792 10376 12844
rect 14556 12928 14608 12980
rect 12532 12860 12584 12912
rect 12716 12792 12768 12844
rect 3424 12656 3476 12708
rect 4436 12656 4488 12708
rect 4896 12656 4948 12708
rect 9312 12656 9364 12708
rect 11152 12724 11204 12776
rect 12348 12724 12400 12776
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 13084 12724 13136 12776
rect 12716 12656 12768 12708
rect 13360 12656 13412 12708
rect 15384 12656 15436 12708
rect 2228 12588 2280 12640
rect 3056 12588 3108 12640
rect 5080 12631 5132 12640
rect 5080 12597 5089 12631
rect 5089 12597 5123 12631
rect 5123 12597 5132 12631
rect 5080 12588 5132 12597
rect 8024 12588 8076 12640
rect 9772 12588 9824 12640
rect 10784 12588 10836 12640
rect 12532 12588 12584 12640
rect 13084 12588 13136 12640
rect 13636 12588 13688 12640
rect 15292 12588 15344 12640
rect 6246 12486 6298 12538
rect 6310 12486 6362 12538
rect 6374 12486 6426 12538
rect 6438 12486 6490 12538
rect 11510 12486 11562 12538
rect 11574 12486 11626 12538
rect 11638 12486 11690 12538
rect 11702 12486 11754 12538
rect 2412 12384 2464 12436
rect 5080 12384 5132 12436
rect 4344 12359 4396 12368
rect 4344 12325 4378 12359
rect 4378 12325 4396 12359
rect 4344 12316 4396 12325
rect 4804 12316 4856 12368
rect 6736 12316 6788 12368
rect 7472 12359 7524 12368
rect 7472 12325 7506 12359
rect 7506 12325 7524 12359
rect 7472 12316 7524 12325
rect 8208 12384 8260 12436
rect 9772 12384 9824 12436
rect 10048 12384 10100 12436
rect 10324 12384 10376 12436
rect 12532 12384 12584 12436
rect 12900 12384 12952 12436
rect 13452 12384 13504 12436
rect 15568 12384 15620 12436
rect 9680 12316 9732 12368
rect 10784 12316 10836 12368
rect 14924 12316 14976 12368
rect 1952 12248 2004 12300
rect 3332 12291 3384 12300
rect 3332 12257 3341 12291
rect 3341 12257 3375 12291
rect 3375 12257 3384 12291
rect 3332 12248 3384 12257
rect 2412 12223 2464 12232
rect 2412 12189 2421 12223
rect 2421 12189 2455 12223
rect 2455 12189 2464 12223
rect 2412 12180 2464 12189
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 3976 12248 4028 12300
rect 4160 12248 4212 12300
rect 9036 12291 9088 12300
rect 9036 12257 9045 12291
rect 9045 12257 9079 12291
rect 9079 12257 9088 12291
rect 9036 12248 9088 12257
rect 11244 12248 11296 12300
rect 11520 12248 11572 12300
rect 12256 12248 12308 12300
rect 13452 12248 13504 12300
rect 2504 12180 2556 12189
rect 2688 12112 2740 12164
rect 2964 12112 3016 12164
rect 6920 12180 6972 12232
rect 10232 12180 10284 12232
rect 13360 12223 13412 12232
rect 7012 12112 7064 12164
rect 2044 12044 2096 12096
rect 4068 12044 4120 12096
rect 7564 12044 7616 12096
rect 7932 12044 7984 12096
rect 11980 12112 12032 12164
rect 12532 12112 12584 12164
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 15292 12248 15344 12300
rect 13728 12223 13780 12232
rect 13360 12180 13412 12189
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 15384 12180 15436 12232
rect 14004 12112 14056 12164
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 9312 12044 9364 12096
rect 10784 12044 10836 12096
rect 11428 12044 11480 12096
rect 13820 12044 13872 12096
rect 14740 12044 14792 12096
rect 3614 11942 3666 11994
rect 3678 11942 3730 11994
rect 3742 11942 3794 11994
rect 3806 11942 3858 11994
rect 8878 11942 8930 11994
rect 8942 11942 8994 11994
rect 9006 11942 9058 11994
rect 9070 11942 9122 11994
rect 14142 11942 14194 11994
rect 14206 11942 14258 11994
rect 14270 11942 14322 11994
rect 14334 11942 14386 11994
rect 2872 11840 2924 11892
rect 6000 11840 6052 11892
rect 5632 11704 5684 11756
rect 8024 11840 8076 11892
rect 9680 11840 9732 11892
rect 14004 11840 14056 11892
rect 1492 11636 1544 11688
rect 2964 11636 3016 11688
rect 3608 11636 3660 11688
rect 4068 11636 4120 11688
rect 5816 11636 5868 11688
rect 6920 11636 6972 11688
rect 9588 11704 9640 11756
rect 10048 11704 10100 11756
rect 10968 11747 11020 11756
rect 10968 11713 10977 11747
rect 10977 11713 11011 11747
rect 11011 11713 11020 11747
rect 10968 11704 11020 11713
rect 12624 11772 12676 11824
rect 15384 11840 15436 11892
rect 11428 11704 11480 11756
rect 2504 11568 2556 11620
rect 1676 11500 1728 11552
rect 2320 11500 2372 11552
rect 2872 11500 2924 11552
rect 2964 11500 3016 11552
rect 3148 11543 3200 11552
rect 3148 11509 3157 11543
rect 3157 11509 3191 11543
rect 3191 11509 3200 11543
rect 3148 11500 3200 11509
rect 4988 11568 5040 11620
rect 5356 11568 5408 11620
rect 5908 11568 5960 11620
rect 7288 11568 7340 11620
rect 7472 11568 7524 11620
rect 7748 11568 7800 11620
rect 11520 11636 11572 11688
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 12164 11636 12216 11688
rect 13360 11636 13412 11688
rect 11060 11568 11112 11620
rect 12256 11568 12308 11620
rect 16120 11772 16172 11824
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 6644 11500 6696 11552
rect 6828 11500 6880 11552
rect 8116 11500 8168 11552
rect 9496 11500 9548 11552
rect 11888 11500 11940 11552
rect 14372 11679 14424 11688
rect 14372 11645 14381 11679
rect 14381 11645 14415 11679
rect 14415 11645 14424 11679
rect 14372 11636 14424 11645
rect 15200 11636 15252 11688
rect 16028 11679 16080 11688
rect 16028 11645 16037 11679
rect 16037 11645 16071 11679
rect 16071 11645 16080 11679
rect 16028 11636 16080 11645
rect 15844 11568 15896 11620
rect 16396 11500 16448 11552
rect 6246 11398 6298 11450
rect 6310 11398 6362 11450
rect 6374 11398 6426 11450
rect 6438 11398 6490 11450
rect 11510 11398 11562 11450
rect 11574 11398 11626 11450
rect 11638 11398 11690 11450
rect 11702 11398 11754 11450
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 2412 11296 2464 11348
rect 2872 11228 2924 11280
rect 4252 11296 4304 11348
rect 4528 11228 4580 11280
rect 7472 11296 7524 11348
rect 7748 11296 7800 11348
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 2320 11203 2372 11212
rect 2320 11169 2329 11203
rect 2329 11169 2363 11203
rect 2363 11169 2372 11203
rect 2320 11160 2372 11169
rect 3148 11160 3200 11212
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 4252 11160 4304 11212
rect 2504 11092 2556 11144
rect 3608 11135 3660 11144
rect 1584 11067 1636 11076
rect 1584 11033 1593 11067
rect 1593 11033 1627 11067
rect 1627 11033 1636 11067
rect 1584 11024 1636 11033
rect 3608 11101 3617 11135
rect 3617 11101 3651 11135
rect 3651 11101 3660 11135
rect 3608 11092 3660 11101
rect 3884 11092 3936 11144
rect 4528 11092 4580 11144
rect 4344 11024 4396 11076
rect 5080 11160 5132 11212
rect 5172 11160 5224 11212
rect 6552 11160 6604 11212
rect 5172 11024 5224 11076
rect 5816 11092 5868 11144
rect 8208 11271 8260 11280
rect 8208 11237 8242 11271
rect 8242 11237 8260 11271
rect 8208 11228 8260 11237
rect 11888 11228 11940 11280
rect 10140 11160 10192 11212
rect 10232 11160 10284 11212
rect 10876 11160 10928 11212
rect 11244 11160 11296 11212
rect 11704 11160 11756 11212
rect 13176 11228 13228 11280
rect 14372 11228 14424 11280
rect 15476 11228 15528 11280
rect 10968 11092 11020 11144
rect 13820 11160 13872 11212
rect 13912 11160 13964 11212
rect 16488 11203 16540 11212
rect 16488 11169 16497 11203
rect 16497 11169 16531 11203
rect 16531 11169 16540 11203
rect 16488 11160 16540 11169
rect 14372 11092 14424 11144
rect 15844 11135 15896 11144
rect 2320 10956 2372 11008
rect 2688 10956 2740 11008
rect 4068 10956 4120 11008
rect 4712 10999 4764 11008
rect 4712 10965 4721 10999
rect 4721 10965 4755 10999
rect 4755 10965 4764 10999
rect 4712 10956 4764 10965
rect 7196 10956 7248 11008
rect 7748 10956 7800 11008
rect 14648 11024 14700 11076
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 9220 10956 9272 11008
rect 10692 10956 10744 11008
rect 11520 10956 11572 11008
rect 11796 10956 11848 11008
rect 13912 10956 13964 11008
rect 14004 10956 14056 11008
rect 14924 10956 14976 11008
rect 3614 10854 3666 10906
rect 3678 10854 3730 10906
rect 3742 10854 3794 10906
rect 3806 10854 3858 10906
rect 8878 10854 8930 10906
rect 8942 10854 8994 10906
rect 9006 10854 9058 10906
rect 9070 10854 9122 10906
rect 14142 10854 14194 10906
rect 14206 10854 14258 10906
rect 14270 10854 14322 10906
rect 14334 10854 14386 10906
rect 2872 10752 2924 10804
rect 3056 10795 3108 10804
rect 3056 10761 3065 10795
rect 3065 10761 3099 10795
rect 3099 10761 3108 10795
rect 3056 10752 3108 10761
rect 4160 10752 4212 10804
rect 3516 10684 3568 10736
rect 2412 10616 2464 10668
rect 1492 10548 1544 10600
rect 3056 10548 3108 10600
rect 3240 10548 3292 10600
rect 3332 10548 3384 10600
rect 4344 10616 4396 10668
rect 5816 10752 5868 10804
rect 6184 10684 6236 10736
rect 8484 10684 8536 10736
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 4988 10548 5040 10600
rect 5632 10548 5684 10600
rect 7012 10548 7064 10600
rect 7840 10548 7892 10600
rect 2964 10480 3016 10532
rect 2504 10412 2556 10464
rect 4160 10480 4212 10532
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 5540 10480 5592 10532
rect 8024 10548 8076 10600
rect 8208 10548 8260 10600
rect 9220 10548 9272 10600
rect 11244 10752 11296 10804
rect 12164 10752 12216 10804
rect 11704 10727 11756 10736
rect 11704 10693 11713 10727
rect 11713 10693 11747 10727
rect 11747 10693 11756 10727
rect 11704 10684 11756 10693
rect 11888 10684 11940 10736
rect 11980 10727 12032 10736
rect 11980 10693 11989 10727
rect 11989 10693 12023 10727
rect 12023 10693 12032 10727
rect 11980 10684 12032 10693
rect 11520 10616 11572 10668
rect 12716 10727 12768 10736
rect 12716 10693 12725 10727
rect 12725 10693 12759 10727
rect 12759 10693 12768 10727
rect 12716 10684 12768 10693
rect 12900 10752 12952 10804
rect 16488 10752 16540 10804
rect 12348 10616 12400 10668
rect 13084 10616 13136 10668
rect 13360 10684 13412 10736
rect 13452 10684 13504 10736
rect 16120 10684 16172 10736
rect 10968 10548 11020 10600
rect 12164 10591 12216 10600
rect 12164 10557 12173 10591
rect 12173 10557 12207 10591
rect 12207 10557 12216 10591
rect 12164 10548 12216 10557
rect 12440 10548 12492 10600
rect 12716 10548 12768 10600
rect 10048 10480 10100 10532
rect 11060 10480 11112 10532
rect 13820 10616 13872 10668
rect 14464 10616 14516 10668
rect 14648 10616 14700 10668
rect 13636 10548 13688 10600
rect 15936 10548 15988 10600
rect 5908 10412 5960 10464
rect 6552 10412 6604 10464
rect 6920 10412 6972 10464
rect 7196 10455 7248 10464
rect 7196 10421 7205 10455
rect 7205 10421 7239 10455
rect 7239 10421 7248 10455
rect 7196 10412 7248 10421
rect 12348 10412 12400 10464
rect 13084 10455 13136 10464
rect 13084 10421 13093 10455
rect 13093 10421 13127 10455
rect 13127 10421 13136 10455
rect 13084 10412 13136 10421
rect 13360 10412 13412 10464
rect 13636 10412 13688 10464
rect 13820 10480 13872 10532
rect 14188 10455 14240 10464
rect 14188 10421 14197 10455
rect 14197 10421 14231 10455
rect 14231 10421 14240 10455
rect 14188 10412 14240 10421
rect 14556 10412 14608 10464
rect 15844 10412 15896 10464
rect 6246 10310 6298 10362
rect 6310 10310 6362 10362
rect 6374 10310 6426 10362
rect 6438 10310 6490 10362
rect 11510 10310 11562 10362
rect 11574 10310 11626 10362
rect 11638 10310 11690 10362
rect 11702 10310 11754 10362
rect 1492 10208 1544 10260
rect 1860 10072 1912 10124
rect 2688 10208 2740 10260
rect 4988 10251 5040 10260
rect 2872 10140 2924 10192
rect 3516 10140 3568 10192
rect 4988 10217 4997 10251
rect 4997 10217 5031 10251
rect 5031 10217 5040 10251
rect 4988 10208 5040 10217
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 5724 10208 5776 10260
rect 7196 10251 7248 10260
rect 6368 10140 6420 10192
rect 7196 10217 7205 10251
rect 7205 10217 7239 10251
rect 7239 10217 7248 10251
rect 7196 10208 7248 10217
rect 8300 10208 8352 10260
rect 9404 10208 9456 10260
rect 14188 10208 14240 10260
rect 14464 10208 14516 10260
rect 16120 10208 16172 10260
rect 2780 10072 2832 10124
rect 3148 10072 3200 10124
rect 4712 10072 4764 10124
rect 5448 10072 5500 10124
rect 5540 10004 5592 10056
rect 3700 9936 3752 9988
rect 6460 10004 6512 10056
rect 6736 10004 6788 10056
rect 7012 10004 7064 10056
rect 8760 10047 8812 10056
rect 6552 9936 6604 9988
rect 8760 10013 8769 10047
rect 8769 10013 8803 10047
rect 8803 10013 8812 10047
rect 8760 10004 8812 10013
rect 11980 10140 12032 10192
rect 12532 10140 12584 10192
rect 12716 10183 12768 10192
rect 12716 10149 12725 10183
rect 12725 10149 12759 10183
rect 12759 10149 12768 10183
rect 12716 10140 12768 10149
rect 12900 10140 12952 10192
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 10232 10004 10284 10056
rect 10324 10004 10376 10056
rect 11244 10072 11296 10124
rect 11060 10004 11112 10056
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 13176 10072 13228 10124
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 13912 10140 13964 10192
rect 14096 10072 14148 10124
rect 15568 10072 15620 10124
rect 12532 10004 12584 10056
rect 13084 10004 13136 10056
rect 11888 9936 11940 9988
rect 2872 9868 2924 9920
rect 3332 9911 3384 9920
rect 3332 9877 3341 9911
rect 3341 9877 3375 9911
rect 3375 9877 3384 9911
rect 3332 9868 3384 9877
rect 6276 9868 6328 9920
rect 8392 9868 8444 9920
rect 9220 9868 9272 9920
rect 9588 9868 9640 9920
rect 9772 9868 9824 9920
rect 10600 9868 10652 9920
rect 11428 9868 11480 9920
rect 12440 9936 12492 9988
rect 13176 9936 13228 9988
rect 13912 9868 13964 9920
rect 15016 9868 15068 9920
rect 15292 9911 15344 9920
rect 15292 9877 15301 9911
rect 15301 9877 15335 9911
rect 15335 9877 15344 9911
rect 15292 9868 15344 9877
rect 3614 9766 3666 9818
rect 3678 9766 3730 9818
rect 3742 9766 3794 9818
rect 3806 9766 3858 9818
rect 8878 9766 8930 9818
rect 8942 9766 8994 9818
rect 9006 9766 9058 9818
rect 9070 9766 9122 9818
rect 14142 9766 14194 9818
rect 14206 9766 14258 9818
rect 14270 9766 14322 9818
rect 14334 9766 14386 9818
rect 2688 9664 2740 9716
rect 1952 9528 2004 9580
rect 2688 9528 2740 9580
rect 3424 9664 3476 9716
rect 6368 9664 6420 9716
rect 6736 9664 6788 9716
rect 4252 9596 4304 9648
rect 5448 9596 5500 9648
rect 6552 9596 6604 9648
rect 1676 9460 1728 9512
rect 4160 9528 4212 9580
rect 4528 9528 4580 9580
rect 3700 9460 3752 9512
rect 5264 9460 5316 9512
rect 1768 9367 1820 9376
rect 1768 9333 1777 9367
rect 1777 9333 1811 9367
rect 1811 9333 1820 9367
rect 1768 9324 1820 9333
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 2780 9324 2832 9376
rect 3332 9392 3384 9444
rect 5540 9528 5592 9580
rect 8760 9664 8812 9716
rect 10508 9664 10560 9716
rect 10784 9664 10836 9716
rect 11428 9664 11480 9716
rect 11888 9664 11940 9716
rect 6000 9460 6052 9512
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 7104 9503 7156 9512
rect 7104 9469 7138 9503
rect 7138 9469 7156 9503
rect 7104 9460 7156 9469
rect 7564 9460 7616 9512
rect 8208 9460 8260 9512
rect 4344 9324 4396 9376
rect 4620 9324 4672 9376
rect 7472 9324 7524 9376
rect 7932 9324 7984 9376
rect 9588 9460 9640 9512
rect 8852 9392 8904 9444
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 10968 9528 11020 9580
rect 11428 9528 11480 9580
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 12900 9528 12952 9580
rect 13084 9528 13136 9580
rect 13544 9664 13596 9716
rect 13820 9596 13872 9648
rect 15936 9664 15988 9716
rect 10232 9460 10284 9512
rect 13728 9460 13780 9512
rect 13912 9503 13964 9512
rect 13912 9469 13921 9503
rect 13921 9469 13955 9503
rect 13955 9469 13964 9503
rect 13912 9460 13964 9469
rect 11888 9392 11940 9444
rect 12992 9392 13044 9444
rect 13084 9392 13136 9444
rect 14832 9392 14884 9444
rect 14924 9392 14976 9444
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 9404 9324 9456 9376
rect 9588 9367 9640 9376
rect 9588 9333 9597 9367
rect 9597 9333 9631 9367
rect 9631 9333 9640 9367
rect 9588 9324 9640 9333
rect 9772 9324 9824 9376
rect 10048 9324 10100 9376
rect 10600 9324 10652 9376
rect 10784 9324 10836 9376
rect 12256 9324 12308 9376
rect 6246 9222 6298 9274
rect 6310 9222 6362 9274
rect 6374 9222 6426 9274
rect 6438 9222 6490 9274
rect 11510 9222 11562 9274
rect 11574 9222 11626 9274
rect 11638 9222 11690 9274
rect 11702 9222 11754 9274
rect 3516 9120 3568 9172
rect 4160 9120 4212 9172
rect 4896 9120 4948 9172
rect 2136 9052 2188 9104
rect 4804 9052 4856 9104
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 2688 8984 2740 9036
rect 3240 8984 3292 9036
rect 2504 8916 2556 8968
rect 3700 8984 3752 9036
rect 4160 8984 4212 9036
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 1676 8848 1728 8900
rect 2780 8780 2832 8832
rect 3240 8780 3292 8832
rect 4344 8848 4396 8900
rect 4528 8848 4580 8900
rect 5816 9120 5868 9172
rect 6828 9120 6880 9172
rect 7196 9120 7248 9172
rect 8668 9120 8720 9172
rect 14924 9163 14976 9172
rect 9772 9052 9824 9104
rect 5632 9027 5684 9036
rect 5632 8993 5666 9027
rect 5666 8993 5684 9027
rect 5632 8984 5684 8993
rect 7196 8984 7248 9036
rect 6644 8916 6696 8968
rect 8024 8984 8076 9036
rect 9864 8984 9916 9036
rect 8300 8916 8352 8968
rect 8852 8916 8904 8968
rect 4712 8780 4764 8832
rect 5080 8823 5132 8832
rect 5080 8789 5089 8823
rect 5089 8789 5123 8823
rect 5123 8789 5132 8823
rect 5080 8780 5132 8789
rect 7104 8848 7156 8900
rect 7932 8848 7984 8900
rect 8208 8848 8260 8900
rect 9128 8848 9180 8900
rect 10508 8984 10560 9036
rect 10876 9027 10928 9036
rect 10876 8993 10885 9027
rect 10885 8993 10919 9027
rect 10919 8993 10928 9027
rect 10876 8984 10928 8993
rect 11796 9027 11848 9036
rect 10692 8916 10744 8968
rect 11796 8993 11830 9027
rect 11830 8993 11848 9027
rect 11796 8984 11848 8993
rect 11980 9052 12032 9104
rect 12164 9052 12216 9104
rect 11244 8916 11296 8968
rect 14924 9129 14933 9163
rect 14933 9129 14967 9163
rect 14967 9129 14976 9163
rect 14924 9120 14976 9129
rect 15660 9120 15712 9172
rect 16212 9120 16264 9172
rect 14004 9052 14056 9104
rect 15200 9052 15252 9104
rect 15844 9052 15896 9104
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13820 9027 13872 9036
rect 13544 8984 13596 8993
rect 13820 8993 13854 9027
rect 13854 8993 13872 9027
rect 13820 8984 13872 8993
rect 14648 8984 14700 9036
rect 15844 8959 15896 8968
rect 10876 8848 10928 8900
rect 12532 8848 12584 8900
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 10692 8780 10744 8832
rect 10968 8780 11020 8832
rect 11244 8780 11296 8832
rect 12900 8823 12952 8832
rect 12900 8789 12909 8823
rect 12909 8789 12943 8823
rect 12943 8789 12952 8823
rect 12900 8780 12952 8789
rect 15200 8848 15252 8900
rect 16120 8848 16172 8900
rect 3614 8678 3666 8730
rect 3678 8678 3730 8730
rect 3742 8678 3794 8730
rect 3806 8678 3858 8730
rect 8878 8678 8930 8730
rect 8942 8678 8994 8730
rect 9006 8678 9058 8730
rect 9070 8678 9122 8730
rect 14142 8678 14194 8730
rect 14206 8678 14258 8730
rect 14270 8678 14322 8730
rect 14334 8678 14386 8730
rect 1492 8372 1544 8424
rect 4620 8576 4672 8628
rect 9588 8576 9640 8628
rect 10324 8619 10376 8628
rect 10324 8585 10333 8619
rect 10333 8585 10367 8619
rect 10367 8585 10376 8619
rect 10324 8576 10376 8585
rect 3240 8440 3292 8492
rect 4252 8508 4304 8560
rect 5632 8508 5684 8560
rect 7104 8508 7156 8560
rect 3792 8440 3844 8492
rect 3424 8415 3476 8424
rect 3424 8381 3433 8415
rect 3433 8381 3467 8415
rect 3467 8381 3476 8415
rect 3424 8372 3476 8381
rect 4252 8372 4304 8424
rect 1768 8304 1820 8356
rect 3148 8304 3200 8356
rect 3516 8304 3568 8356
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 3056 8236 3108 8245
rect 6828 8440 6880 8492
rect 10048 8440 10100 8492
rect 4528 8372 4580 8424
rect 4712 8347 4764 8356
rect 4712 8313 4746 8347
rect 4746 8313 4764 8347
rect 4712 8304 4764 8313
rect 4896 8304 4948 8356
rect 5908 8304 5960 8356
rect 6644 8236 6696 8288
rect 8668 8372 8720 8424
rect 11244 8440 11296 8492
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 10692 8415 10744 8424
rect 10692 8381 10701 8415
rect 10701 8381 10735 8415
rect 10735 8381 10744 8415
rect 10692 8372 10744 8381
rect 11428 8372 11480 8424
rect 12164 8372 12216 8424
rect 12716 8483 12768 8492
rect 12716 8449 12725 8483
rect 12725 8449 12759 8483
rect 12759 8449 12768 8483
rect 12716 8440 12768 8449
rect 15016 8440 15068 8492
rect 15844 8440 15896 8492
rect 14004 8372 14056 8424
rect 14096 8372 14148 8424
rect 7840 8347 7892 8356
rect 7840 8313 7874 8347
rect 7874 8313 7892 8347
rect 7840 8304 7892 8313
rect 9864 8304 9916 8356
rect 8576 8236 8628 8288
rect 9036 8236 9088 8288
rect 9956 8236 10008 8288
rect 10140 8236 10192 8288
rect 10324 8236 10376 8288
rect 12256 8236 12308 8288
rect 13636 8236 13688 8288
rect 13820 8304 13872 8356
rect 14464 8372 14516 8424
rect 15292 8372 15344 8424
rect 15476 8372 15528 8424
rect 14004 8236 14056 8288
rect 6246 8134 6298 8186
rect 6310 8134 6362 8186
rect 6374 8134 6426 8186
rect 6438 8134 6490 8186
rect 11510 8134 11562 8186
rect 11574 8134 11626 8186
rect 11638 8134 11690 8186
rect 11702 8134 11754 8186
rect 2228 8032 2280 8084
rect 7288 8032 7340 8084
rect 8300 8075 8352 8084
rect 2044 7964 2096 8016
rect 4988 7964 5040 8016
rect 1676 7896 1728 7948
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 5724 7964 5776 8016
rect 6644 7964 6696 8016
rect 8300 8041 8309 8075
rect 8309 8041 8343 8075
rect 8343 8041 8352 8075
rect 8300 8032 8352 8041
rect 8484 7964 8536 8016
rect 12532 8032 12584 8084
rect 12624 8032 12676 8084
rect 13360 8032 13412 8084
rect 13728 8032 13780 8084
rect 14464 8032 14516 8084
rect 10232 7964 10284 8016
rect 10324 7964 10376 8016
rect 10692 7964 10744 8016
rect 6828 7896 6880 7948
rect 8300 7896 8352 7948
rect 2964 7828 3016 7880
rect 4712 7828 4764 7880
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 8484 7828 8536 7880
rect 9036 7828 9088 7880
rect 4804 7760 4856 7812
rect 6000 7760 6052 7812
rect 1400 7692 1452 7744
rect 1952 7735 2004 7744
rect 1952 7701 1961 7735
rect 1961 7701 1995 7735
rect 1995 7701 2004 7735
rect 1952 7692 2004 7701
rect 3148 7692 3200 7744
rect 4712 7692 4764 7744
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6276 7692 6328 7701
rect 8208 7692 8260 7744
rect 11888 7896 11940 7948
rect 13820 7939 13872 7948
rect 13820 7905 13829 7939
rect 13829 7905 13863 7939
rect 13863 7905 13872 7939
rect 13820 7896 13872 7905
rect 14096 7896 14148 7948
rect 14648 7939 14700 7948
rect 14648 7905 14657 7939
rect 14657 7905 14691 7939
rect 14691 7905 14700 7939
rect 14648 7896 14700 7905
rect 9588 7828 9640 7880
rect 10324 7828 10376 7880
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 13728 7828 13780 7880
rect 16304 7896 16356 7948
rect 9680 7803 9732 7812
rect 9680 7769 9689 7803
rect 9689 7769 9723 7803
rect 9723 7769 9732 7803
rect 9680 7760 9732 7769
rect 11796 7760 11848 7812
rect 10232 7692 10284 7744
rect 11704 7692 11756 7744
rect 12532 7692 12584 7744
rect 15108 7760 15160 7812
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 13084 7692 13136 7744
rect 13820 7692 13872 7744
rect 15292 7692 15344 7744
rect 3614 7590 3666 7642
rect 3678 7590 3730 7642
rect 3742 7590 3794 7642
rect 3806 7590 3858 7642
rect 8878 7590 8930 7642
rect 8942 7590 8994 7642
rect 9006 7590 9058 7642
rect 9070 7590 9122 7642
rect 14142 7590 14194 7642
rect 14206 7590 14258 7642
rect 14270 7590 14322 7642
rect 14334 7590 14386 7642
rect 1952 7488 2004 7540
rect 2964 7463 3016 7472
rect 2964 7429 2973 7463
rect 2973 7429 3007 7463
rect 3007 7429 3016 7463
rect 4804 7488 4856 7540
rect 6552 7488 6604 7540
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 2964 7420 3016 7429
rect 1492 7352 1544 7404
rect 3056 7352 3108 7404
rect 6092 7420 6144 7472
rect 3976 7352 4028 7404
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 4712 7284 4764 7336
rect 6276 7352 6328 7404
rect 11244 7488 11296 7540
rect 11888 7488 11940 7540
rect 14004 7488 14056 7540
rect 14464 7488 14516 7540
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 7748 7284 7800 7336
rect 7932 7284 7984 7336
rect 8208 7284 8260 7336
rect 9864 7352 9916 7404
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 13728 7352 13780 7404
rect 14924 7352 14976 7404
rect 15108 7352 15160 7404
rect 15936 7395 15988 7404
rect 15936 7361 15945 7395
rect 15945 7361 15979 7395
rect 15979 7361 15988 7395
rect 15936 7352 15988 7361
rect 9496 7284 9548 7336
rect 2320 7216 2372 7268
rect 2596 7216 2648 7268
rect 3148 7148 3200 7200
rect 6736 7216 6788 7268
rect 4344 7148 4396 7200
rect 5632 7191 5684 7200
rect 5632 7157 5641 7191
rect 5641 7157 5675 7191
rect 5675 7157 5684 7191
rect 5632 7148 5684 7157
rect 6644 7148 6696 7200
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 8576 7259 8628 7268
rect 8576 7225 8610 7259
rect 8610 7225 8628 7259
rect 12624 7284 12676 7336
rect 8576 7216 8628 7225
rect 11060 7216 11112 7268
rect 11244 7216 11296 7268
rect 13360 7284 13412 7336
rect 9588 7148 9640 7200
rect 9772 7148 9824 7200
rect 13636 7148 13688 7200
rect 14188 7148 14240 7200
rect 14648 7148 14700 7200
rect 15476 7148 15528 7200
rect 6246 7046 6298 7098
rect 6310 7046 6362 7098
rect 6374 7046 6426 7098
rect 6438 7046 6490 7098
rect 11510 7046 11562 7098
rect 11574 7046 11626 7098
rect 11638 7046 11690 7098
rect 11702 7046 11754 7098
rect 6644 6944 6696 6996
rect 7288 6944 7340 6996
rect 8484 6944 8536 6996
rect 1584 6808 1636 6860
rect 3424 6808 3476 6860
rect 5080 6808 5132 6860
rect 1860 6740 1912 6792
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2639 6783
rect 2639 6749 2648 6783
rect 2596 6740 2648 6749
rect 2780 6740 2832 6792
rect 3240 6740 3292 6792
rect 4344 6672 4396 6724
rect 848 6604 900 6656
rect 2044 6647 2096 6656
rect 2044 6613 2053 6647
rect 2053 6613 2087 6647
rect 2087 6613 2096 6647
rect 2044 6604 2096 6613
rect 3424 6604 3476 6656
rect 3976 6604 4028 6656
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 4896 6740 4948 6792
rect 5540 6851 5592 6860
rect 5540 6817 5574 6851
rect 5574 6817 5592 6851
rect 5540 6808 5592 6817
rect 5724 6876 5776 6928
rect 6184 6876 6236 6928
rect 8760 6919 8812 6928
rect 7472 6808 7524 6860
rect 8760 6885 8769 6919
rect 8769 6885 8803 6919
rect 8803 6885 8812 6919
rect 8760 6876 8812 6885
rect 9220 6876 9272 6928
rect 9496 6876 9548 6928
rect 10232 6876 10284 6928
rect 4620 6672 4672 6724
rect 8116 6672 8168 6724
rect 8576 6808 8628 6860
rect 8852 6783 8904 6792
rect 8852 6749 8861 6783
rect 8861 6749 8895 6783
rect 8895 6749 8904 6783
rect 8852 6740 8904 6749
rect 9772 6808 9824 6860
rect 11980 6876 12032 6928
rect 12440 6808 12492 6860
rect 14188 6987 14240 6996
rect 12624 6876 12676 6928
rect 14188 6953 14197 6987
rect 14197 6953 14231 6987
rect 14231 6953 14240 6987
rect 14188 6944 14240 6953
rect 15568 6944 15620 6996
rect 15752 6944 15804 6996
rect 15936 6876 15988 6928
rect 9220 6740 9272 6792
rect 9128 6672 9180 6724
rect 6184 6604 6236 6656
rect 6644 6647 6696 6656
rect 6644 6613 6653 6647
rect 6653 6613 6687 6647
rect 6687 6613 6696 6647
rect 6644 6604 6696 6613
rect 9312 6604 9364 6656
rect 9864 6604 9916 6656
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 13268 6740 13320 6792
rect 12900 6672 12952 6724
rect 15200 6808 15252 6860
rect 16028 6808 16080 6860
rect 15108 6740 15160 6792
rect 15752 6783 15804 6792
rect 13912 6672 13964 6724
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 13176 6604 13228 6656
rect 14832 6604 14884 6656
rect 3614 6502 3666 6554
rect 3678 6502 3730 6554
rect 3742 6502 3794 6554
rect 3806 6502 3858 6554
rect 8878 6502 8930 6554
rect 8942 6502 8994 6554
rect 9006 6502 9058 6554
rect 9070 6502 9122 6554
rect 14142 6502 14194 6554
rect 14206 6502 14258 6554
rect 14270 6502 14322 6554
rect 14334 6502 14386 6554
rect 4160 6400 4212 6452
rect 4712 6400 4764 6452
rect 7288 6400 7340 6452
rect 5540 6332 5592 6384
rect 1584 6264 1636 6316
rect 2596 6264 2648 6316
rect 3884 6264 3936 6316
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 1492 6196 1544 6248
rect 2872 6239 2924 6248
rect 2872 6205 2881 6239
rect 2881 6205 2915 6239
rect 2915 6205 2924 6239
rect 2872 6196 2924 6205
rect 2964 6196 3016 6248
rect 4160 6196 4212 6248
rect 6828 6264 6880 6316
rect 7288 6264 7340 6316
rect 9588 6332 9640 6384
rect 12348 6400 12400 6452
rect 12440 6400 12492 6452
rect 13084 6400 13136 6452
rect 13728 6400 13780 6452
rect 11796 6332 11848 6384
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 8024 6264 8076 6316
rect 11244 6264 11296 6316
rect 12440 6264 12492 6316
rect 12808 6264 12860 6316
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 13912 6264 13964 6316
rect 4712 6128 4764 6180
rect 1860 6103 1912 6112
rect 1860 6069 1869 6103
rect 1869 6069 1903 6103
rect 1903 6069 1912 6103
rect 1860 6060 1912 6069
rect 6736 6196 6788 6248
rect 7656 6196 7708 6248
rect 7932 6196 7984 6248
rect 9864 6196 9916 6248
rect 11060 6196 11112 6248
rect 12072 6196 12124 6248
rect 5172 6128 5224 6180
rect 5080 6060 5132 6112
rect 8484 6128 8536 6180
rect 8208 6060 8260 6112
rect 9128 6060 9180 6112
rect 13176 6196 13228 6248
rect 15108 6171 15160 6180
rect 15108 6137 15142 6171
rect 15142 6137 15160 6171
rect 15108 6128 15160 6137
rect 15200 6128 15252 6180
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 12808 6060 12860 6112
rect 12992 6060 13044 6112
rect 13084 6060 13136 6112
rect 15292 6060 15344 6112
rect 6246 5958 6298 6010
rect 6310 5958 6362 6010
rect 6374 5958 6426 6010
rect 6438 5958 6490 6010
rect 11510 5958 11562 6010
rect 11574 5958 11626 6010
rect 11638 5958 11690 6010
rect 11702 5958 11754 6010
rect 2872 5856 2924 5908
rect 3884 5856 3936 5908
rect 4344 5856 4396 5908
rect 4804 5856 4856 5908
rect 4896 5856 4948 5908
rect 5816 5856 5868 5908
rect 2596 5788 2648 5840
rect 3976 5788 4028 5840
rect 1584 5720 1636 5772
rect 4160 5720 4212 5772
rect 4436 5652 4488 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 4896 5720 4948 5772
rect 5264 5720 5316 5772
rect 7932 5856 7984 5908
rect 8116 5899 8168 5908
rect 8116 5865 8125 5899
rect 8125 5865 8159 5899
rect 8159 5865 8168 5899
rect 8116 5856 8168 5865
rect 9680 5856 9732 5908
rect 10140 5856 10192 5908
rect 11152 5856 11204 5908
rect 12164 5856 12216 5908
rect 12808 5856 12860 5908
rect 15292 5899 15344 5908
rect 15292 5865 15301 5899
rect 15301 5865 15335 5899
rect 15335 5865 15344 5899
rect 15292 5856 15344 5865
rect 15752 5899 15804 5908
rect 15752 5865 15761 5899
rect 15761 5865 15795 5899
rect 15795 5865 15804 5899
rect 15752 5856 15804 5865
rect 6828 5788 6880 5840
rect 6644 5720 6696 5772
rect 7656 5720 7708 5772
rect 7472 5652 7524 5704
rect 10232 5788 10284 5840
rect 9772 5720 9824 5772
rect 8944 5652 8996 5704
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 9588 5652 9640 5704
rect 12532 5831 12584 5840
rect 11060 5720 11112 5772
rect 10968 5652 11020 5704
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 1952 5516 2004 5568
rect 11244 5584 11296 5636
rect 11796 5584 11848 5636
rect 12532 5797 12541 5831
rect 12541 5797 12575 5831
rect 12575 5797 12584 5831
rect 12532 5788 12584 5797
rect 13176 5720 13228 5772
rect 13360 5763 13412 5772
rect 13360 5729 13394 5763
rect 13394 5729 13412 5763
rect 13360 5720 13412 5729
rect 11980 5652 12032 5704
rect 12624 5695 12676 5704
rect 12624 5661 12633 5695
rect 12633 5661 12667 5695
rect 12667 5661 12676 5695
rect 12624 5652 12676 5661
rect 15568 5652 15620 5704
rect 12900 5584 12952 5636
rect 15108 5584 15160 5636
rect 15292 5584 15344 5636
rect 3516 5516 3568 5568
rect 4160 5559 4212 5568
rect 4160 5525 4169 5559
rect 4169 5525 4203 5559
rect 4203 5525 4212 5559
rect 4160 5516 4212 5525
rect 4620 5516 4672 5568
rect 5540 5516 5592 5568
rect 5908 5516 5960 5568
rect 6184 5516 6236 5568
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 10140 5516 10192 5568
rect 11336 5516 11388 5568
rect 15660 5516 15712 5568
rect 3614 5414 3666 5466
rect 3678 5414 3730 5466
rect 3742 5414 3794 5466
rect 3806 5414 3858 5466
rect 8878 5414 8930 5466
rect 8942 5414 8994 5466
rect 9006 5414 9058 5466
rect 9070 5414 9122 5466
rect 14142 5414 14194 5466
rect 14206 5414 14258 5466
rect 14270 5414 14322 5466
rect 14334 5414 14386 5466
rect 2780 5312 2832 5364
rect 2596 5176 2648 5228
rect 5080 5312 5132 5364
rect 6276 5312 6328 5364
rect 7288 5312 7340 5364
rect 8024 5312 8076 5364
rect 8760 5312 8812 5364
rect 4896 5176 4948 5228
rect 5724 5219 5776 5228
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 7748 5176 7800 5228
rect 2320 5108 2372 5160
rect 2412 5108 2464 5160
rect 4160 5108 4212 5160
rect 4620 5108 4672 5160
rect 5908 5108 5960 5160
rect 6184 5151 6236 5160
rect 6184 5117 6193 5151
rect 6193 5117 6227 5151
rect 6227 5117 6236 5151
rect 6184 5108 6236 5117
rect 6644 5108 6696 5160
rect 6920 5108 6972 5160
rect 8668 5108 8720 5160
rect 9864 5312 9916 5364
rect 10876 5312 10928 5364
rect 15016 5312 15068 5364
rect 10692 5176 10744 5228
rect 14096 5244 14148 5296
rect 14648 5244 14700 5296
rect 9680 5108 9732 5160
rect 10968 5108 11020 5160
rect 13176 5108 13228 5160
rect 13728 5108 13780 5160
rect 2964 5040 3016 5092
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 4436 5040 4488 5092
rect 3608 4972 3660 5024
rect 4620 5015 4672 5024
rect 4620 4981 4629 5015
rect 4629 4981 4663 5015
rect 4663 4981 4672 5015
rect 4620 4972 4672 4981
rect 7288 5040 7340 5092
rect 8116 5040 8168 5092
rect 11152 5040 11204 5092
rect 13912 5040 13964 5092
rect 5540 4972 5592 5024
rect 5724 4972 5776 5024
rect 8392 4972 8444 5024
rect 9772 4972 9824 5024
rect 10508 4972 10560 5024
rect 10968 4972 11020 5024
rect 11060 4972 11112 5024
rect 11244 5015 11296 5024
rect 11244 4981 11253 5015
rect 11253 4981 11287 5015
rect 11287 4981 11296 5015
rect 11244 4972 11296 4981
rect 11336 4972 11388 5024
rect 12808 4972 12860 5024
rect 13360 4972 13412 5024
rect 14924 4972 14976 5024
rect 15292 5040 15344 5092
rect 6246 4870 6298 4922
rect 6310 4870 6362 4922
rect 6374 4870 6426 4922
rect 6438 4870 6490 4922
rect 11510 4870 11562 4922
rect 11574 4870 11626 4922
rect 11638 4870 11690 4922
rect 11702 4870 11754 4922
rect 2504 4768 2556 4820
rect 5724 4768 5776 4820
rect 5908 4768 5960 4820
rect 6644 4768 6696 4820
rect 2412 4700 2464 4752
rect 1492 4675 1544 4684
rect 1492 4641 1501 4675
rect 1501 4641 1535 4675
rect 1535 4641 1544 4675
rect 1492 4632 1544 4641
rect 1768 4675 1820 4684
rect 1768 4641 1802 4675
rect 1802 4641 1820 4675
rect 4160 4700 4212 4752
rect 4620 4700 4672 4752
rect 6092 4700 6144 4752
rect 6460 4700 6512 4752
rect 7012 4700 7064 4752
rect 1768 4632 1820 4641
rect 3884 4632 3936 4684
rect 4896 4632 4948 4684
rect 3976 4564 4028 4616
rect 7472 4632 7524 4684
rect 8116 4700 8168 4752
rect 10048 4768 10100 4820
rect 11980 4768 12032 4820
rect 14464 4768 14516 4820
rect 15200 4768 15252 4820
rect 15568 4768 15620 4820
rect 10968 4700 11020 4752
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 2872 4471 2924 4480
rect 2872 4437 2881 4471
rect 2881 4437 2915 4471
rect 2915 4437 2924 4471
rect 2872 4428 2924 4437
rect 3240 4428 3292 4480
rect 4068 4428 4120 4480
rect 5264 4428 5316 4480
rect 8392 4564 8444 4616
rect 12348 4632 12400 4684
rect 13084 4632 13136 4684
rect 13820 4632 13872 4684
rect 10416 4564 10468 4616
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 11796 4564 11848 4616
rect 11980 4564 12032 4616
rect 12808 4607 12860 4616
rect 12808 4573 12817 4607
rect 12817 4573 12851 4607
rect 12851 4573 12860 4607
rect 12808 4564 12860 4573
rect 13912 4564 13964 4616
rect 15200 4564 15252 4616
rect 15752 4607 15804 4616
rect 15752 4573 15761 4607
rect 15761 4573 15795 4607
rect 15795 4573 15804 4607
rect 15752 4564 15804 4573
rect 6828 4428 6880 4480
rect 7012 4428 7064 4480
rect 7656 4428 7708 4480
rect 14740 4496 14792 4548
rect 8484 4428 8536 4480
rect 9404 4428 9456 4480
rect 10508 4428 10560 4480
rect 13912 4428 13964 4480
rect 3614 4326 3666 4378
rect 3678 4326 3730 4378
rect 3742 4326 3794 4378
rect 3806 4326 3858 4378
rect 8878 4326 8930 4378
rect 8942 4326 8994 4378
rect 9006 4326 9058 4378
rect 9070 4326 9122 4378
rect 14142 4326 14194 4378
rect 14206 4326 14258 4378
rect 14270 4326 14322 4378
rect 14334 4326 14386 4378
rect 1768 4156 1820 4208
rect 3516 4224 3568 4276
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 4436 4088 4488 4140
rect 5540 4224 5592 4276
rect 5080 4199 5132 4208
rect 5080 4165 5089 4199
rect 5089 4165 5123 4199
rect 5123 4165 5132 4199
rect 5080 4156 5132 4165
rect 5908 4156 5960 4208
rect 6644 4156 6696 4208
rect 8116 4224 8168 4276
rect 10784 4224 10836 4276
rect 12256 4224 12308 4276
rect 12440 4224 12492 4276
rect 15200 4224 15252 4276
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 2044 4020 2096 4072
rect 2136 4020 2188 4072
rect 4344 4020 4396 4072
rect 6092 4063 6144 4072
rect 6092 4029 6101 4063
rect 6101 4029 6135 4063
rect 6135 4029 6144 4063
rect 6092 4020 6144 4029
rect 2872 3952 2924 4004
rect 3884 3952 3936 4004
rect 1400 3927 1452 3936
rect 1400 3893 1409 3927
rect 1409 3893 1443 3927
rect 1443 3893 1452 3927
rect 1400 3884 1452 3893
rect 2412 3884 2464 3936
rect 3516 3884 3568 3936
rect 3792 3927 3844 3936
rect 3792 3893 3801 3927
rect 3801 3893 3835 3927
rect 3835 3893 3844 3927
rect 3792 3884 3844 3893
rect 4068 3927 4120 3936
rect 4068 3893 4077 3927
rect 4077 3893 4111 3927
rect 4111 3893 4120 3927
rect 4068 3884 4120 3893
rect 4344 3884 4396 3936
rect 4528 3884 4580 3936
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 6460 3952 6512 4004
rect 6644 3952 6696 4004
rect 7012 3952 7064 4004
rect 8944 4088 8996 4140
rect 8668 4020 8720 4072
rect 9496 4020 9548 4072
rect 9680 4020 9732 4072
rect 10692 4020 10744 4072
rect 13176 4020 13228 4072
rect 11060 3952 11112 4004
rect 5540 3884 5592 3893
rect 7932 3884 7984 3936
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 8852 3884 8904 3893
rect 8944 3927 8996 3936
rect 8944 3893 8953 3927
rect 8953 3893 8987 3927
rect 8987 3893 8996 3927
rect 9496 3927 9548 3936
rect 8944 3884 8996 3893
rect 9496 3893 9505 3927
rect 9505 3893 9539 3927
rect 9539 3893 9548 3927
rect 9496 3884 9548 3893
rect 9772 3884 9824 3936
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 10876 3884 10928 3936
rect 14464 3952 14516 4004
rect 16028 3995 16080 4004
rect 13912 3884 13964 3936
rect 16028 3961 16037 3995
rect 16037 3961 16071 3995
rect 16071 3961 16080 3995
rect 16028 3952 16080 3961
rect 6246 3782 6298 3834
rect 6310 3782 6362 3834
rect 6374 3782 6426 3834
rect 6438 3782 6490 3834
rect 11510 3782 11562 3834
rect 11574 3782 11626 3834
rect 11638 3782 11690 3834
rect 11702 3782 11754 3834
rect 1400 3680 1452 3732
rect 4068 3680 4120 3732
rect 572 3476 624 3528
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 2320 3451 2372 3460
rect 2320 3417 2329 3451
rect 2329 3417 2363 3451
rect 2363 3417 2372 3451
rect 2320 3408 2372 3417
rect 2596 3408 2648 3460
rect 3792 3612 3844 3664
rect 5540 3680 5592 3732
rect 5632 3612 5684 3664
rect 3516 3476 3568 3528
rect 5816 3544 5868 3596
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 5356 3476 5408 3528
rect 5448 3476 5500 3528
rect 6368 3612 6420 3664
rect 7564 3612 7616 3664
rect 6828 3544 6880 3596
rect 6920 3476 6972 3528
rect 7656 3544 7708 3596
rect 8852 3723 8904 3732
rect 8852 3689 8861 3723
rect 8861 3689 8895 3723
rect 8895 3689 8904 3723
rect 8852 3680 8904 3689
rect 9496 3680 9548 3732
rect 12256 3680 12308 3732
rect 12164 3655 12216 3664
rect 8300 3544 8352 3596
rect 8668 3476 8720 3528
rect 9128 3544 9180 3596
rect 9588 3544 9640 3596
rect 10324 3544 10376 3596
rect 10692 3544 10744 3596
rect 10968 3544 11020 3596
rect 12164 3621 12173 3655
rect 12173 3621 12207 3655
rect 12207 3621 12216 3655
rect 12808 3723 12860 3732
rect 12808 3689 12817 3723
rect 12817 3689 12851 3723
rect 12851 3689 12860 3723
rect 13820 3723 13872 3732
rect 12808 3680 12860 3689
rect 13820 3689 13829 3723
rect 13829 3689 13863 3723
rect 13863 3689 13872 3723
rect 13820 3680 13872 3689
rect 12164 3612 12216 3621
rect 12440 3612 12492 3664
rect 12624 3544 12676 3596
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 3884 3408 3936 3460
rect 3056 3340 3108 3392
rect 4068 3340 4120 3392
rect 9956 3408 10008 3460
rect 11704 3476 11756 3528
rect 11980 3476 12032 3528
rect 13268 3544 13320 3596
rect 15660 3544 15712 3596
rect 12900 3519 12952 3528
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 13728 3476 13780 3528
rect 15200 3476 15252 3528
rect 13084 3408 13136 3460
rect 5724 3383 5776 3392
rect 5724 3349 5733 3383
rect 5733 3349 5767 3383
rect 5767 3349 5776 3383
rect 5724 3340 5776 3349
rect 5816 3340 5868 3392
rect 7656 3340 7708 3392
rect 9312 3340 9364 3392
rect 9680 3383 9732 3392
rect 9680 3349 9689 3383
rect 9689 3349 9723 3383
rect 9723 3349 9732 3383
rect 9680 3340 9732 3349
rect 10968 3383 11020 3392
rect 10968 3349 10977 3383
rect 10977 3349 11011 3383
rect 11011 3349 11020 3383
rect 10968 3340 11020 3349
rect 11152 3383 11204 3392
rect 11152 3349 11161 3383
rect 11161 3349 11195 3383
rect 11195 3349 11204 3383
rect 12348 3383 12400 3392
rect 11152 3340 11204 3349
rect 12348 3349 12357 3383
rect 12357 3349 12391 3383
rect 12391 3349 12400 3383
rect 12348 3340 12400 3349
rect 15108 3340 15160 3392
rect 3614 3238 3666 3290
rect 3678 3238 3730 3290
rect 3742 3238 3794 3290
rect 3806 3238 3858 3290
rect 8878 3238 8930 3290
rect 8942 3238 8994 3290
rect 9006 3238 9058 3290
rect 9070 3238 9122 3290
rect 14142 3238 14194 3290
rect 14206 3238 14258 3290
rect 14270 3238 14322 3290
rect 14334 3238 14386 3290
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 3332 3136 3384 3188
rect 4160 3136 4212 3188
rect 4620 3136 4672 3188
rect 4988 3136 5040 3188
rect 7748 3136 7800 3188
rect 9312 3179 9364 3188
rect 9312 3145 9321 3179
rect 9321 3145 9355 3179
rect 9355 3145 9364 3179
rect 9312 3136 9364 3145
rect 9588 3136 9640 3188
rect 9864 3136 9916 3188
rect 5448 3111 5500 3120
rect 5448 3077 5457 3111
rect 5457 3077 5491 3111
rect 5491 3077 5500 3111
rect 5448 3068 5500 3077
rect 2688 3000 2740 3052
rect 2964 3000 3016 3052
rect 4620 3000 4672 3052
rect 7012 3068 7064 3120
rect 5816 3000 5868 3052
rect 6000 3043 6052 3052
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 6000 3000 6052 3009
rect 7564 3000 7616 3052
rect 1768 2907 1820 2916
rect 1768 2873 1777 2907
rect 1777 2873 1811 2907
rect 1811 2873 1820 2907
rect 1768 2864 1820 2873
rect 3332 2864 3384 2916
rect 2688 2839 2740 2848
rect 2688 2805 2697 2839
rect 2697 2805 2731 2839
rect 2731 2805 2740 2839
rect 2688 2796 2740 2805
rect 5540 2932 5592 2984
rect 6644 2932 6696 2984
rect 4436 2864 4488 2916
rect 5448 2864 5500 2916
rect 6368 2864 6420 2916
rect 4344 2796 4396 2848
rect 4620 2839 4672 2848
rect 4620 2805 4629 2839
rect 4629 2805 4663 2839
rect 4663 2805 4672 2839
rect 4620 2796 4672 2805
rect 5356 2796 5408 2848
rect 6644 2796 6696 2848
rect 7380 2932 7432 2984
rect 10600 3068 10652 3120
rect 8024 3000 8076 3052
rect 8760 3043 8812 3052
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 9036 3000 9088 3052
rect 10876 3136 10928 3188
rect 11336 3179 11388 3188
rect 11336 3145 11345 3179
rect 11345 3145 11379 3179
rect 11379 3145 11388 3179
rect 11336 3136 11388 3145
rect 11520 3136 11572 3188
rect 13728 3179 13780 3188
rect 13728 3145 13737 3179
rect 13737 3145 13771 3179
rect 13771 3145 13780 3179
rect 13728 3136 13780 3145
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 12900 3000 12952 3052
rect 13820 3000 13872 3052
rect 14464 3000 14516 3052
rect 14648 3000 14700 3052
rect 10600 2932 10652 2984
rect 11244 2932 11296 2984
rect 10048 2864 10100 2916
rect 10416 2864 10468 2916
rect 11888 2864 11940 2916
rect 8576 2796 8628 2848
rect 9588 2796 9640 2848
rect 9956 2796 10008 2848
rect 10324 2839 10376 2848
rect 10324 2805 10333 2839
rect 10333 2805 10367 2839
rect 10367 2805 10376 2839
rect 10324 2796 10376 2805
rect 10508 2796 10560 2848
rect 12440 2932 12492 2984
rect 13176 2932 13228 2984
rect 12624 2864 12676 2916
rect 15200 2864 15252 2916
rect 16304 2864 16356 2916
rect 6246 2694 6298 2746
rect 6310 2694 6362 2746
rect 6374 2694 6426 2746
rect 6438 2694 6490 2746
rect 11510 2694 11562 2746
rect 11574 2694 11626 2746
rect 11638 2694 11690 2746
rect 11702 2694 11754 2746
rect 4252 2592 4304 2644
rect 4436 2635 4488 2644
rect 4436 2601 4445 2635
rect 4445 2601 4479 2635
rect 4479 2601 4488 2635
rect 4436 2592 4488 2601
rect 5080 2592 5132 2644
rect 5632 2592 5684 2644
rect 7196 2592 7248 2644
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 9956 2592 10008 2644
rect 11060 2592 11112 2644
rect 11336 2592 11388 2644
rect 12716 2592 12768 2644
rect 3148 2524 3200 2576
rect 5724 2524 5776 2576
rect 5816 2567 5868 2576
rect 5816 2533 5825 2567
rect 5825 2533 5859 2567
rect 5859 2533 5868 2567
rect 5816 2524 5868 2533
rect 9680 2524 9732 2576
rect 11980 2524 12032 2576
rect 3332 2499 3384 2508
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 3332 2465 3341 2499
rect 3341 2465 3375 2499
rect 3375 2465 3384 2499
rect 3332 2456 3384 2465
rect 6644 2456 6696 2508
rect 7104 2456 7156 2508
rect 3240 2388 3292 2440
rect 5264 2388 5316 2440
rect 6000 2431 6052 2440
rect 6000 2397 6009 2431
rect 6009 2397 6043 2431
rect 6043 2397 6052 2431
rect 6000 2388 6052 2397
rect 7564 2388 7616 2440
rect 8852 2388 8904 2440
rect 9956 2456 10008 2508
rect 11796 2499 11848 2508
rect 9772 2388 9824 2440
rect 11336 2431 11388 2440
rect 3148 2320 3200 2372
rect 6092 2320 6144 2372
rect 6552 2320 6604 2372
rect 8208 2320 8260 2372
rect 4896 2252 4948 2304
rect 6920 2252 6972 2304
rect 9404 2252 9456 2304
rect 11336 2397 11345 2431
rect 11345 2397 11379 2431
rect 11379 2397 11388 2431
rect 11336 2388 11388 2397
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 12348 2524 12400 2576
rect 12532 2524 12584 2576
rect 12256 2456 12308 2508
rect 17408 2524 17460 2576
rect 14556 2456 14608 2508
rect 15384 2456 15436 2508
rect 13820 2431 13872 2440
rect 10692 2320 10744 2372
rect 12808 2320 12860 2372
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 13820 2388 13872 2397
rect 14464 2320 14516 2372
rect 3614 2150 3666 2202
rect 3678 2150 3730 2202
rect 3742 2150 3794 2202
rect 3806 2150 3858 2202
rect 8878 2150 8930 2202
rect 8942 2150 8994 2202
rect 9006 2150 9058 2202
rect 9070 2150 9122 2202
rect 14142 2150 14194 2202
rect 14206 2150 14258 2202
rect 14270 2150 14322 2202
rect 14334 2150 14386 2202
rect 3240 2048 3292 2100
rect 5172 2048 5224 2100
rect 3332 1980 3384 2032
rect 10140 2048 10192 2100
rect 11336 2048 11388 2100
rect 12808 2048 12860 2100
rect 3148 1912 3200 1964
rect 6184 1912 6236 1964
rect 9588 1368 9640 1420
rect 13820 1368 13872 1420
rect 3424 1300 3476 1352
rect 6920 1300 6972 1352
rect 11796 1096 11848 1148
rect 16028 1096 16080 1148
rect 1768 620 1820 672
rect 5080 620 5132 672
<< metal2 >>
rect 2226 16520 2282 17000
rect 6734 16520 6790 17000
rect 7654 16688 7710 16697
rect 7654 16623 7710 16632
rect 2240 15026 2268 16520
rect 4066 16280 4122 16289
rect 4066 16215 4122 16224
rect 2686 15872 2742 15881
rect 2686 15807 2742 15816
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 1400 14544 1452 14550
rect 1400 14486 1452 14492
rect 1412 11218 1440 14486
rect 2412 14476 2464 14482
rect 2412 14418 2464 14424
rect 2318 13288 2374 13297
rect 2318 13223 2374 13232
rect 2332 12782 2360 13223
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1504 10606 1532 11630
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1504 10266 1532 10542
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1412 8809 1440 8978
rect 1398 8800 1454 8809
rect 1398 8735 1454 8744
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 1400 7744 1452 7750
rect 1400 7686 1452 7692
rect 1306 6896 1362 6905
rect 1306 6831 1362 6840
rect 848 6656 900 6662
rect 848 6598 900 6604
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 860 2689 888 6598
rect 1320 5681 1348 6831
rect 1306 5672 1362 5681
rect 1306 5607 1362 5616
rect 1412 4457 1440 7686
rect 1504 7410 1532 8366
rect 1596 7449 1624 11018
rect 1688 9518 1716 11494
rect 1964 11354 1992 12242
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1872 10033 1900 10066
rect 1858 10024 1914 10033
rect 1858 9959 1914 9968
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1676 8900 1728 8906
rect 1676 8842 1728 8848
rect 1688 7954 1716 8842
rect 1780 8362 1808 9318
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1582 7440 1638 7449
rect 1492 7404 1544 7410
rect 1582 7375 1638 7384
rect 1492 7346 1544 7352
rect 1504 6254 1532 7346
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1596 6322 1624 6802
rect 1872 6798 1900 9959
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1964 9081 1992 9522
rect 1950 9072 2006 9081
rect 1950 9007 2006 9016
rect 2056 8022 2084 12038
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2148 9110 2176 9318
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 2240 8090 2268 12582
rect 2424 12442 2452 14418
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2608 13938 2636 14350
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2516 12322 2544 13806
rect 2608 12850 2636 13874
rect 2700 13734 2728 15807
rect 3974 15464 4030 15473
rect 3974 15399 4030 15408
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 2688 13728 2740 13734
rect 2688 13670 2740 13676
rect 2700 13462 2728 13670
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 2976 12850 3004 13330
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2332 12294 2544 12322
rect 2332 11558 2360 12294
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2504 12232 2556 12238
rect 2608 12220 2636 12786
rect 2556 12192 2636 12220
rect 2504 12174 2556 12180
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2424 11354 2452 12174
rect 2516 11626 2544 12174
rect 2976 12170 3004 12786
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 2594 11656 2650 11665
rect 2504 11620 2556 11626
rect 2594 11591 2650 11600
rect 2504 11562 2556 11568
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2320 11212 2372 11218
rect 2372 11172 2452 11200
rect 2320 11154 2372 11160
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2044 8016 2096 8022
rect 2044 7958 2096 7964
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1964 7546 1992 7686
rect 2332 7562 2360 10950
rect 2424 10674 2452 11172
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 2240 7534 2360 7562
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 1504 5760 1532 6190
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1584 5772 1636 5778
rect 1504 5732 1584 5760
rect 1504 4690 1532 5732
rect 1584 5714 1636 5720
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1398 4448 1454 4457
rect 1398 4383 1454 4392
rect 1688 4049 1716 5510
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1780 4214 1808 4626
rect 1768 4208 1820 4214
rect 1768 4150 1820 4156
rect 1872 4146 1900 6054
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1674 4040 1730 4049
rect 1674 3975 1730 3984
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1412 3738 1440 3878
rect 1400 3732 1452 3738
rect 1400 3674 1452 3680
rect 1768 2916 1820 2922
rect 1768 2858 1820 2864
rect 846 2680 902 2689
rect 846 2615 902 2624
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1688 480 1716 2382
rect 1780 678 1808 2858
rect 1964 1873 1992 5510
rect 2056 4078 2084 6598
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2148 4078 2176 4966
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 2240 3194 2268 7534
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2332 5692 2360 7210
rect 2424 5817 2452 10610
rect 2516 10470 2544 11086
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 9897 2544 10406
rect 2502 9888 2558 9897
rect 2502 9823 2558 9832
rect 2504 8968 2556 8974
rect 2502 8936 2504 8945
rect 2556 8936 2558 8945
rect 2502 8871 2558 8880
rect 2516 6882 2544 8871
rect 2608 7313 2636 11591
rect 2700 11014 2728 12106
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2884 11558 2912 11834
rect 2976 11694 3004 12106
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2884 10810 2912 11222
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2700 9722 2728 10202
rect 2884 10198 2912 10746
rect 2976 10538 3004 11494
rect 3068 10810 3096 12582
rect 3160 11558 3188 13806
rect 3436 13802 3464 14214
rect 3528 13841 3556 14758
rect 3588 14172 3884 14192
rect 3644 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3666 14118 3668 14170
rect 3730 14118 3742 14170
rect 3804 14118 3806 14170
rect 3644 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3588 14096 3884 14116
rect 3514 13832 3570 13841
rect 3424 13796 3476 13802
rect 3514 13767 3570 13776
rect 3424 13738 3476 13744
rect 3988 13462 4016 15399
rect 4080 15230 4108 16215
rect 4068 15224 4120 15230
rect 4068 15166 4120 15172
rect 4066 15056 4122 15065
rect 4066 14991 4122 15000
rect 6552 15020 6604 15026
rect 4080 14958 4108 14991
rect 6552 14962 6604 14968
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 4066 14648 4122 14657
rect 4172 14618 4200 14826
rect 6220 14716 6516 14736
rect 6276 14714 6300 14716
rect 6356 14714 6380 14716
rect 6436 14714 6460 14716
rect 6298 14662 6300 14714
rect 6362 14662 6374 14714
rect 6436 14662 6438 14714
rect 6276 14660 6300 14662
rect 6356 14660 6380 14662
rect 6436 14660 6460 14662
rect 6220 14640 6516 14660
rect 4066 14583 4122 14592
rect 4160 14612 4212 14618
rect 4080 14278 4108 14583
rect 4160 14554 4212 14560
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 4172 14074 4200 14418
rect 4620 14408 4672 14414
rect 4672 14368 4752 14396
rect 4620 14350 4672 14356
rect 4344 14340 4396 14346
rect 4344 14282 4396 14288
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3330 12880 3386 12889
rect 3330 12815 3386 12824
rect 3344 12306 3372 12815
rect 3528 12782 3556 13126
rect 3588 13084 3884 13104
rect 3644 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3666 13030 3668 13082
rect 3730 13030 3742 13082
rect 3804 13030 3806 13082
rect 3644 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3588 13008 3884 13028
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3436 12345 3464 12650
rect 3422 12336 3478 12345
rect 3332 12300 3384 12306
rect 3252 12260 3332 12288
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2686 9616 2742 9625
rect 2686 9551 2688 9560
rect 2740 9551 2742 9560
rect 2688 9522 2740 9528
rect 2792 9382 2820 10066
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 9217 2820 9318
rect 2778 9208 2834 9217
rect 2778 9143 2834 9152
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2700 8673 2728 8978
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2686 8664 2742 8673
rect 2686 8599 2742 8608
rect 2594 7304 2650 7313
rect 2594 7239 2596 7248
rect 2648 7239 2650 7248
rect 2596 7210 2648 7216
rect 2608 7179 2636 7210
rect 2792 6905 2820 8774
rect 2778 6896 2834 6905
rect 2516 6854 2728 6882
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2608 6322 2636 6734
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2608 5846 2636 6258
rect 2596 5840 2648 5846
rect 2410 5808 2466 5817
rect 2596 5782 2648 5788
rect 2410 5743 2466 5752
rect 2332 5664 2452 5692
rect 2424 5166 2452 5664
rect 2608 5234 2636 5782
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2332 3466 2360 5102
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2424 4146 2452 4694
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2424 3942 2452 4082
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2320 3460 2372 3466
rect 2320 3402 2372 3408
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 1950 1864 2006 1873
rect 1950 1799 2006 1808
rect 2516 1057 2544 4762
rect 2700 3618 2728 6854
rect 2778 6831 2834 6840
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2792 5522 2820 6734
rect 2884 6497 2912 9862
rect 2976 7886 3004 10474
rect 3068 8401 3096 10542
rect 3160 10130 3188 11154
rect 3252 10606 3280 12260
rect 3988 12306 4016 13262
rect 3422 12271 3478 12280
rect 3976 12300 4028 12306
rect 3332 12242 3384 12248
rect 3330 10840 3386 10849
rect 3330 10775 3386 10784
rect 3344 10606 3372 10775
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3436 10554 3464 12271
rect 3976 12242 4028 12248
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 3588 11996 3884 12016
rect 3644 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3666 11942 3668 11994
rect 3730 11942 3742 11994
rect 3804 11942 3806 11994
rect 3644 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3588 11920 3884 11940
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3620 11150 3648 11630
rect 3882 11248 3938 11257
rect 3882 11183 3938 11192
rect 3896 11150 3924 11183
rect 3608 11144 3660 11150
rect 3528 11092 3608 11098
rect 3528 11086 3660 11092
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3528 11070 3648 11086
rect 3528 10742 3556 11070
rect 3588 10908 3884 10928
rect 3644 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3666 10854 3668 10906
rect 3730 10854 3742 10906
rect 3804 10854 3806 10906
rect 3644 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3588 10832 3884 10852
rect 3516 10736 3568 10742
rect 3516 10678 3568 10684
rect 3436 10526 3556 10554
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 10305 3464 10406
rect 3422 10296 3478 10305
rect 3422 10231 3478 10240
rect 3528 10198 3556 10526
rect 3698 10432 3754 10441
rect 3698 10367 3754 10376
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3712 9994 3740 10367
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3344 9738 3372 9862
rect 3588 9820 3884 9840
rect 3644 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3666 9766 3668 9818
rect 3730 9766 3742 9818
rect 3804 9766 3806 9818
rect 3644 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3588 9744 3884 9764
rect 3344 9722 3455 9738
rect 3344 9716 3476 9722
rect 3344 9710 3424 9716
rect 3424 9658 3476 9664
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3238 9344 3294 9353
rect 3238 9279 3294 9288
rect 3252 9042 3280 9279
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 8498 3280 8774
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3054 8392 3110 8401
rect 3054 8327 3110 8336
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2870 6488 2926 6497
rect 2870 6423 2926 6432
rect 2976 6254 3004 7414
rect 3068 7410 3096 8230
rect 3160 7834 3188 8298
rect 3344 8072 3372 9386
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3528 8820 3556 9114
rect 3712 9042 3740 9454
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3436 8792 3556 8820
rect 3436 8430 3464 8792
rect 3588 8732 3884 8752
rect 3644 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3666 8678 3668 8730
rect 3730 8678 3742 8730
rect 3804 8678 3806 8730
rect 3644 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3588 8656 3884 8676
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 3344 8044 3464 8072
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3160 7806 3280 7834
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3160 7290 3188 7686
rect 3068 7262 3188 7290
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2884 5914 2912 6190
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2962 5808 3018 5817
rect 2962 5743 3018 5752
rect 2792 5494 2912 5522
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2608 3590 2728 3618
rect 2608 3466 2636 3590
rect 2686 3496 2742 3505
rect 2596 3460 2648 3466
rect 2686 3431 2742 3440
rect 2596 3402 2648 3408
rect 2700 3058 2728 3431
rect 2792 3346 2820 5306
rect 2884 4865 2912 5494
rect 2976 5098 3004 5743
rect 3068 5409 3096 7262
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3054 5400 3110 5409
rect 3054 5335 3110 5344
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2870 4856 2926 4865
rect 2870 4791 2926 4800
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2884 4010 2912 4422
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2884 3534 2912 3946
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3056 3392 3108 3398
rect 2792 3318 2912 3346
rect 3056 3334 3108 3340
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 2700 2553 2728 2790
rect 2686 2544 2742 2553
rect 2686 2479 2742 2488
rect 2884 1306 2912 3318
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2976 2961 3004 2994
rect 2962 2952 3018 2961
rect 2962 2887 3018 2896
rect 2792 1278 2912 1306
rect 2502 1048 2558 1057
rect 2502 983 2558 992
rect 1768 672 1820 678
rect 1768 614 1820 620
rect 2792 480 2820 1278
rect 570 0 626 480
rect 1674 0 1730 480
rect 2778 0 2834 480
rect 3068 241 3096 3334
rect 3160 2582 3188 7142
rect 3252 6798 3280 7806
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 3252 2446 3280 4422
rect 3344 3194 3372 7890
rect 3436 7041 3464 8044
rect 3422 7032 3478 7041
rect 3422 6967 3478 6976
rect 3422 6896 3478 6905
rect 3422 6831 3424 6840
rect 3476 6831 3478 6840
rect 3424 6802 3476 6808
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3330 2952 3386 2961
rect 3330 2887 3332 2896
rect 3384 2887 3386 2896
rect 3332 2858 3384 2864
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3148 2372 3200 2378
rect 3148 2314 3200 2320
rect 3160 1970 3188 2314
rect 3240 2100 3292 2106
rect 3240 2042 3292 2048
rect 3148 1964 3200 1970
rect 3148 1906 3200 1912
rect 3252 1465 3280 2042
rect 3344 2038 3372 2450
rect 3436 2281 3464 6598
rect 3528 6089 3556 8298
rect 3804 8004 3832 8434
rect 3988 8072 4016 12242
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4080 11694 4108 12038
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4066 11248 4122 11257
rect 4066 11183 4068 11192
rect 4120 11183 4122 11192
rect 4068 11154 4120 11160
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 8265 4108 10950
rect 4172 10810 4200 12242
rect 4264 11354 4292 14010
rect 4356 12986 4384 14282
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4632 13530 4660 13670
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4724 12986 4752 14368
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4356 12374 4384 12922
rect 4816 12850 4844 13874
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4908 12714 4936 12922
rect 4436 12708 4488 12714
rect 4436 12650 4488 12656
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 4172 9897 4200 10474
rect 4158 9888 4214 9897
rect 4158 9823 4214 9832
rect 4264 9654 4292 11154
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4356 10985 4384 11018
rect 4342 10976 4398 10985
rect 4342 10911 4398 10920
rect 4342 10840 4398 10849
rect 4342 10775 4398 10784
rect 4356 10674 4384 10775
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4252 9648 4304 9654
rect 4250 9616 4252 9625
rect 4304 9616 4306 9625
rect 4160 9580 4212 9586
rect 4250 9551 4306 9560
rect 4160 9522 4212 9528
rect 4172 9178 4200 9522
rect 4356 9382 4384 10610
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4250 9208 4306 9217
rect 4160 9172 4212 9178
rect 4250 9143 4306 9152
rect 4160 9114 4212 9120
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4066 8256 4122 8265
rect 4066 8191 4122 8200
rect 3988 8044 4108 8072
rect 3804 7976 4016 8004
rect 3588 7644 3884 7664
rect 3644 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3666 7590 3668 7642
rect 3730 7590 3742 7642
rect 3804 7590 3806 7642
rect 3644 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3588 7568 3884 7588
rect 3988 7410 4016 7976
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3588 6556 3884 6576
rect 3644 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3666 6502 3668 6554
rect 3730 6502 3742 6554
rect 3804 6502 3806 6554
rect 3644 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3588 6480 3884 6500
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3514 6080 3570 6089
rect 3514 6015 3570 6024
rect 3896 5914 3924 6258
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3516 5568 3568 5574
rect 3896 5556 3924 5850
rect 3988 5846 4016 6598
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 3896 5528 4016 5556
rect 3516 5510 3568 5516
rect 3528 4282 3556 5510
rect 3588 5468 3884 5488
rect 3644 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3666 5414 3668 5466
rect 3730 5414 3742 5466
rect 3804 5414 3806 5466
rect 3644 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3588 5392 3884 5412
rect 3606 5128 3662 5137
rect 3606 5063 3662 5072
rect 3620 5030 3648 5063
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3988 4706 4016 5528
rect 3896 4690 4016 4706
rect 3884 4684 4016 4690
rect 3936 4678 4016 4684
rect 3884 4626 3936 4632
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3588 4380 3884 4400
rect 3644 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3666 4326 3668 4378
rect 3730 4326 3742 4378
rect 3804 4326 3806 4378
rect 3644 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3588 4304 3884 4324
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3528 3534 3556 3878
rect 3606 3768 3662 3777
rect 3606 3703 3662 3712
rect 3516 3528 3568 3534
rect 3620 3505 3648 3703
rect 3804 3670 3832 3878
rect 3792 3664 3844 3670
rect 3896 3641 3924 3946
rect 3792 3606 3844 3612
rect 3882 3632 3938 3641
rect 3882 3567 3938 3576
rect 3516 3470 3568 3476
rect 3606 3496 3662 3505
rect 3606 3431 3662 3440
rect 3882 3496 3938 3505
rect 3882 3431 3884 3440
rect 3936 3431 3938 3440
rect 3884 3402 3936 3408
rect 3588 3292 3884 3312
rect 3644 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3666 3238 3668 3290
rect 3730 3238 3742 3290
rect 3804 3238 3806 3290
rect 3644 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3588 3216 3884 3236
rect 3422 2272 3478 2281
rect 3422 2207 3478 2216
rect 3588 2204 3884 2224
rect 3644 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3666 2150 3668 2202
rect 3730 2150 3742 2202
rect 3804 2150 3806 2202
rect 3644 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3588 2128 3884 2148
rect 3988 2088 4016 4558
rect 4080 4486 4108 8044
rect 4172 7857 4200 8978
rect 4264 8566 4292 9143
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4158 7848 4214 7857
rect 4158 7783 4214 7792
rect 4264 7732 4292 8366
rect 4172 7704 4292 7732
rect 4172 6458 4200 7704
rect 4250 7576 4306 7585
rect 4250 7511 4306 7520
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4172 5778 4200 6190
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4172 5166 4200 5510
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3738 4108 3878
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4080 3097 4108 3334
rect 4172 3194 4200 4694
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4066 3088 4122 3097
rect 4066 3023 4122 3032
rect 4264 2650 4292 7511
rect 4356 7426 4384 8842
rect 4448 7857 4476 12650
rect 4526 12472 4582 12481
rect 4526 12407 4582 12416
rect 4540 11286 4568 12407
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 4618 11792 4674 11801
rect 4618 11727 4674 11736
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4540 9586 4568 11086
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4632 9466 4660 11727
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4724 10130 4752 10950
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4710 9888 4766 9897
rect 4710 9823 4766 9832
rect 4724 9489 4752 9823
rect 4540 9438 4660 9466
rect 4710 9480 4766 9489
rect 4540 8906 4568 9438
rect 4710 9415 4766 9424
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 8974 4660 9318
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4632 8634 4660 8910
rect 4724 8838 4752 9415
rect 4816 9110 4844 12310
rect 5000 11626 5028 14214
rect 5552 14006 5580 14418
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5736 14074 5764 14350
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5540 14000 5592 14006
rect 5446 13968 5502 13977
rect 5356 13932 5408 13938
rect 5540 13942 5592 13948
rect 5446 13903 5502 13912
rect 5356 13874 5408 13880
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 5092 12442 5120 12582
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 5184 11393 5212 13262
rect 5170 11384 5226 11393
rect 5170 11319 5226 11328
rect 5170 11248 5226 11257
rect 5080 11212 5132 11218
rect 5170 11183 5172 11192
rect 5080 11154 5132 11160
rect 5224 11183 5226 11192
rect 5172 11154 5224 11160
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 5000 10266 5028 10542
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4434 7848 4490 7857
rect 4434 7783 4490 7792
rect 4356 7398 4476 7426
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4356 6730 4384 7142
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4342 6624 4398 6633
rect 4342 6559 4398 6568
rect 4356 5914 4384 6559
rect 4448 6202 4476 7398
rect 4540 6322 4568 8366
rect 4632 7324 4660 8570
rect 4908 8362 4936 9114
rect 5092 8838 5120 11154
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5184 10849 5212 11018
rect 5170 10840 5226 10849
rect 5170 10775 5226 10784
rect 5170 10568 5226 10577
rect 5170 10503 5226 10512
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4724 7886 4752 8298
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4724 7750 4752 7822
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4816 7546 4844 7754
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4712 7336 4764 7342
rect 4632 7296 4712 7324
rect 4712 7278 4764 7284
rect 4724 6798 4752 7278
rect 4908 6798 4936 7822
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4632 6440 4660 6666
rect 4712 6452 4764 6458
rect 4632 6412 4712 6440
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4448 6174 4568 6202
rect 4434 6080 4490 6089
rect 4434 6015 4490 6024
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4356 5409 4384 5850
rect 4448 5710 4476 6015
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4342 5400 4398 5409
rect 4342 5335 4398 5344
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4448 4146 4476 5034
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4356 3942 4384 4014
rect 4540 3942 4568 6174
rect 4632 5574 4660 6412
rect 4712 6394 4764 6400
rect 4802 6216 4858 6225
rect 4712 6180 4764 6186
rect 4802 6151 4858 6160
rect 4712 6122 4764 6128
rect 4724 5710 4752 6122
rect 4816 5914 4844 6151
rect 4908 5914 4936 6734
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4896 5772 4948 5778
rect 4816 5732 4896 5760
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4618 5264 4674 5273
rect 4618 5199 4674 5208
rect 4632 5166 4660 5199
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4710 5128 4766 5137
rect 4710 5063 4766 5072
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4632 4758 4660 4966
rect 4620 4752 4672 4758
rect 4620 4694 4672 4700
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4528 3936 4580 3942
rect 4724 3924 4752 5063
rect 4528 3878 4580 3884
rect 4632 3896 4752 3924
rect 4632 3346 4660 3896
rect 4540 3318 4660 3346
rect 4342 3088 4398 3097
rect 4342 3023 4398 3032
rect 4356 2854 4384 3023
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4448 2650 4476 2858
rect 4540 2836 4568 3318
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4632 3058 4660 3130
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4816 2961 4844 5732
rect 4896 5714 4948 5720
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4908 4690 4936 5170
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4894 3224 4950 3233
rect 5000 3194 5028 7958
rect 5092 6866 5120 8774
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5184 6304 5212 10503
rect 5276 9518 5304 13738
rect 5368 13326 5396 13874
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5184 6276 5304 6304
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5092 5370 5120 6054
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 4894 3159 4950 3168
rect 4988 3188 5040 3194
rect 4802 2952 4858 2961
rect 4802 2887 4858 2896
rect 4620 2848 4672 2854
rect 4540 2808 4620 2836
rect 4620 2790 4672 2796
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4908 2310 4936 3159
rect 4988 3130 5040 3136
rect 5092 2650 5120 4150
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 5184 2106 5212 6122
rect 5276 5778 5304 6276
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5276 2446 5304 4422
rect 5368 3534 5396 11562
rect 5460 10130 5488 13903
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5644 12424 5672 13262
rect 5828 12986 5856 13330
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5644 12396 5764 12424
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5644 10606 5672 11698
rect 5736 11676 5764 12396
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5816 11688 5868 11694
rect 5736 11648 5816 11676
rect 5816 11630 5868 11636
rect 5906 11656 5962 11665
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5552 10266 5580 10474
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5540 10056 5592 10062
rect 5644 10044 5672 10542
rect 5736 10266 5764 11494
rect 5828 11150 5856 11630
rect 5906 11591 5908 11600
rect 5960 11591 5962 11600
rect 5908 11562 5960 11568
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5828 10810 5856 11086
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5722 10160 5778 10169
rect 5722 10095 5778 10104
rect 5592 10016 5672 10044
rect 5540 9998 5592 10004
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5460 6225 5488 9590
rect 5552 9586 5580 9998
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5644 8566 5672 8978
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5736 8412 5764 10095
rect 5828 9178 5856 10746
rect 5920 10470 5948 11562
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5906 10296 5962 10305
rect 5906 10231 5962 10240
rect 5920 9897 5948 10231
rect 5906 9888 5962 9897
rect 5906 9823 5962 9832
rect 6012 9518 6040 11834
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5644 8384 5764 8412
rect 5644 7206 5672 8384
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 5736 7857 5764 7958
rect 5722 7848 5778 7857
rect 5722 7783 5778 7792
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5552 6390 5580 6802
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5446 6216 5502 6225
rect 5446 6151 5502 6160
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 5030 5580 5510
rect 5644 5273 5672 7142
rect 5736 6934 5764 7346
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5630 5264 5686 5273
rect 5630 5199 5686 5208
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5736 5114 5764 5170
rect 5644 5086 5764 5114
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 4282 5580 4966
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5644 4146 5672 5086
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4826 5764 4966
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5828 4706 5856 5850
rect 5920 5574 5948 8298
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5920 4826 5948 5102
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5736 4678 5856 4706
rect 5736 4622 5764 4678
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5908 4208 5960 4214
rect 5908 4150 5960 4156
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3738 5580 3878
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5644 3670 5672 4082
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5354 3360 5410 3369
rect 5354 3295 5410 3304
rect 5368 2854 5396 3295
rect 5460 3126 5488 3470
rect 5828 3398 5856 3538
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 5356 2848 5408 2854
rect 5460 2825 5488 2858
rect 5356 2790 5408 2796
rect 5446 2816 5502 2825
rect 5446 2751 5502 2760
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5552 2394 5580 2926
rect 5630 2816 5686 2825
rect 5630 2751 5686 2760
rect 5644 2650 5672 2751
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5736 2582 5764 3334
rect 5828 3058 5856 3334
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5920 2938 5948 4150
rect 6012 3233 6040 7754
rect 6104 7478 6132 14418
rect 6220 13628 6516 13648
rect 6276 13626 6300 13628
rect 6356 13626 6380 13628
rect 6436 13626 6460 13628
rect 6298 13574 6300 13626
rect 6362 13574 6374 13626
rect 6436 13574 6438 13626
rect 6276 13572 6300 13574
rect 6356 13572 6380 13574
rect 6436 13572 6460 13574
rect 6220 13552 6516 13572
rect 6220 12540 6516 12560
rect 6276 12538 6300 12540
rect 6356 12538 6380 12540
rect 6436 12538 6460 12540
rect 6298 12486 6300 12538
rect 6362 12486 6374 12538
rect 6436 12486 6438 12538
rect 6276 12484 6300 12486
rect 6356 12484 6380 12486
rect 6436 12484 6460 12486
rect 6220 12464 6516 12484
rect 6220 11452 6516 11472
rect 6276 11450 6300 11452
rect 6356 11450 6380 11452
rect 6436 11450 6460 11452
rect 6298 11398 6300 11450
rect 6362 11398 6374 11450
rect 6436 11398 6438 11450
rect 6276 11396 6300 11398
rect 6356 11396 6380 11398
rect 6436 11396 6460 11398
rect 6220 11376 6516 11396
rect 6564 11370 6592 14962
rect 6644 14340 6696 14346
rect 6644 14282 6696 14288
rect 6656 12073 6684 14282
rect 6748 13462 6776 16520
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6840 12832 6868 13874
rect 7116 13870 7144 14350
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7116 13530 7144 13806
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 6920 12844 6972 12850
rect 6840 12804 6920 12832
rect 6920 12786 6972 12792
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6642 12064 6698 12073
rect 6642 11999 6698 12008
rect 6656 11558 6684 11999
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6564 11342 6684 11370
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6184 10736 6236 10742
rect 6182 10704 6184 10713
rect 6236 10704 6238 10713
rect 6182 10639 6238 10648
rect 6564 10470 6592 11154
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6220 10364 6516 10384
rect 6276 10362 6300 10364
rect 6356 10362 6380 10364
rect 6436 10362 6460 10364
rect 6298 10310 6300 10362
rect 6362 10310 6374 10362
rect 6436 10310 6438 10362
rect 6276 10308 6300 10310
rect 6356 10308 6380 10310
rect 6436 10308 6460 10310
rect 6220 10288 6516 10308
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6288 9625 6316 9862
rect 6380 9722 6408 10134
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6274 9616 6330 9625
rect 6274 9551 6330 9560
rect 6472 9466 6500 9998
rect 6564 9994 6592 10406
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6550 9752 6606 9761
rect 6550 9687 6606 9696
rect 6564 9654 6592 9687
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6472 9438 6592 9466
rect 6220 9276 6516 9296
rect 6276 9274 6300 9276
rect 6356 9274 6380 9276
rect 6436 9274 6460 9276
rect 6298 9222 6300 9274
rect 6362 9222 6374 9274
rect 6436 9222 6438 9274
rect 6276 9220 6300 9222
rect 6356 9220 6380 9222
rect 6436 9220 6460 9222
rect 6220 9200 6516 9220
rect 6220 8188 6516 8208
rect 6276 8186 6300 8188
rect 6356 8186 6380 8188
rect 6436 8186 6460 8188
rect 6298 8134 6300 8186
rect 6362 8134 6374 8186
rect 6436 8134 6438 8186
rect 6276 8132 6300 8134
rect 6356 8132 6380 8134
rect 6436 8132 6460 8134
rect 6220 8112 6516 8132
rect 6564 7834 6592 9438
rect 6656 8974 6684 11342
rect 6748 10062 6776 12310
rect 6932 12238 6960 12786
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6932 11694 6960 12174
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 10169 6868 11494
rect 6932 11393 6960 11630
rect 6918 11384 6974 11393
rect 6918 11319 6974 11328
rect 7024 10606 7052 12106
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6826 10160 6882 10169
rect 6826 10095 6882 10104
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 8022 6684 8230
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6196 7806 6592 7834
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 6196 7290 6224 7806
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 7410 6316 7686
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6104 7262 6224 7290
rect 6104 4758 6132 7262
rect 6220 7100 6516 7120
rect 6276 7098 6300 7100
rect 6356 7098 6380 7100
rect 6436 7098 6460 7100
rect 6298 7046 6300 7098
rect 6362 7046 6374 7098
rect 6436 7046 6438 7098
rect 6276 7044 6300 7046
rect 6356 7044 6380 7046
rect 6436 7044 6460 7046
rect 6220 7024 6516 7044
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 6196 6662 6224 6870
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6220 6012 6516 6032
rect 6276 6010 6300 6012
rect 6356 6010 6380 6012
rect 6436 6010 6460 6012
rect 6298 5958 6300 6010
rect 6362 5958 6374 6010
rect 6436 5958 6438 6010
rect 6276 5956 6300 5958
rect 6356 5956 6380 5958
rect 6436 5956 6460 5958
rect 6220 5936 6516 5956
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6196 5166 6224 5510
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6184 5160 6236 5166
rect 6288 5137 6316 5306
rect 6184 5102 6236 5108
rect 6274 5128 6330 5137
rect 6274 5063 6330 5072
rect 6220 4924 6516 4944
rect 6276 4922 6300 4924
rect 6356 4922 6380 4924
rect 6436 4922 6460 4924
rect 6298 4870 6300 4922
rect 6362 4870 6374 4922
rect 6436 4870 6438 4922
rect 6276 4868 6300 4870
rect 6356 4868 6380 4870
rect 6436 4868 6460 4870
rect 6220 4848 6516 4868
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6104 4078 6132 4694
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6472 4010 6500 4694
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6220 3836 6516 3856
rect 6276 3834 6300 3836
rect 6356 3834 6380 3836
rect 6436 3834 6460 3836
rect 6298 3782 6300 3834
rect 6362 3782 6374 3834
rect 6436 3782 6438 3834
rect 6276 3780 6300 3782
rect 6356 3780 6380 3782
rect 6436 3780 6460 3782
rect 6220 3760 6516 3780
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 5998 3224 6054 3233
rect 5998 3159 6054 3168
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 5828 2910 5948 2938
rect 5828 2582 5856 2910
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 5828 2394 5856 2518
rect 6012 2446 6040 2994
rect 5552 2366 5856 2394
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 6104 2378 6132 3538
rect 6380 2922 6408 3606
rect 6368 2916 6420 2922
rect 6368 2858 6420 2864
rect 6220 2748 6516 2768
rect 6276 2746 6300 2748
rect 6356 2746 6380 2748
rect 6436 2746 6460 2748
rect 6298 2694 6300 2746
rect 6362 2694 6374 2746
rect 6436 2694 6438 2746
rect 6276 2692 6300 2694
rect 6356 2692 6380 2694
rect 6436 2692 6460 2694
rect 6220 2672 6516 2692
rect 6564 2378 6592 7482
rect 6748 7274 6776 9658
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 9178 6868 9454
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6840 8498 6868 9114
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6840 7546 6868 7890
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6656 7002 6684 7142
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6656 5778 6684 6598
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6748 5817 6776 6190
rect 6840 6089 6868 6258
rect 6826 6080 6882 6089
rect 6826 6015 6882 6024
rect 6828 5840 6880 5846
rect 6734 5808 6790 5817
rect 6644 5772 6696 5778
rect 6828 5782 6880 5788
rect 6734 5743 6790 5752
rect 6644 5714 6696 5720
rect 6840 5681 6868 5782
rect 6826 5672 6882 5681
rect 6826 5607 6882 5616
rect 6932 5166 6960 10406
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 7024 9761 7052 9998
rect 7010 9752 7066 9761
rect 7010 9687 7066 9696
rect 7116 9602 7144 13126
rect 7300 12356 7328 13466
rect 7208 12328 7328 12356
rect 7208 11014 7236 12328
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7208 10266 7236 10406
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7024 9574 7144 9602
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6656 4826 6684 5102
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6656 4214 6684 4762
rect 7024 4758 7052 9574
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7116 8906 7144 9454
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7208 9042 7236 9114
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 7116 7886 7144 8502
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7208 7732 7236 8978
rect 7300 8090 7328 11562
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7116 7704 7236 7732
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6840 4146 6868 4422
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 7024 4010 7052 4422
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6656 2990 6684 3946
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6644 2984 6696 2990
rect 6840 2961 6868 3538
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6644 2926 6696 2932
rect 6826 2952 6882 2961
rect 6826 2887 6882 2896
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6656 2514 6684 2790
rect 6932 2553 6960 3470
rect 7024 3126 7052 3946
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 6918 2544 6974 2553
rect 6644 2508 6696 2514
rect 7116 2514 7144 7704
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 2650 7236 7142
rect 7300 7002 7328 7278
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7286 6760 7342 6769
rect 7286 6695 7342 6704
rect 7300 6458 7328 6695
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7300 5370 7328 6258
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 6918 2479 6974 2488
rect 7104 2508 7156 2514
rect 6644 2450 6696 2456
rect 7104 2450 7156 2456
rect 6092 2372 6144 2378
rect 6092 2314 6144 2320
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 3896 2060 4016 2088
rect 5172 2100 5224 2106
rect 3332 2032 3384 2038
rect 3332 1974 3384 1980
rect 3238 1456 3294 1465
rect 3238 1391 3294 1400
rect 3424 1352 3476 1358
rect 3424 1294 3476 1300
rect 3436 649 3464 1294
rect 3422 640 3478 649
rect 3422 575 3478 584
rect 3896 480 3924 2060
rect 5172 2042 5224 2048
rect 6184 1964 6236 1970
rect 6184 1906 6236 1912
rect 5080 672 5132 678
rect 5080 614 5132 620
rect 5092 480 5120 614
rect 6196 480 6224 1906
rect 6932 1358 6960 2246
rect 6920 1352 6972 1358
rect 6920 1294 6972 1300
rect 7300 480 7328 5034
rect 7392 2990 7420 14214
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7484 12374 7512 12718
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7484 11354 7512 11562
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7484 10674 7512 11290
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7576 9518 7604 12038
rect 7668 11608 7696 16623
rect 11242 16520 11298 17000
rect 15014 16688 15070 16697
rect 15014 16623 15070 16632
rect 9956 15224 10008 15230
rect 9956 15166 10008 15172
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8312 13462 8340 14554
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8404 13530 8432 14214
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 7840 13456 7892 13462
rect 7840 13398 7892 13404
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 7748 11620 7800 11626
rect 7668 11580 7748 11608
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7472 9376 7524 9382
rect 7668 9364 7696 11580
rect 7852 11608 7880 13398
rect 8588 13394 8616 14418
rect 8680 14074 8708 14418
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7932 12096 7984 12102
rect 7930 12064 7932 12073
rect 7984 12064 7986 12073
rect 7930 11999 7986 12008
rect 8036 11898 8064 12582
rect 8220 12442 8248 13262
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7852 11580 7972 11608
rect 7748 11562 7800 11568
rect 7746 11384 7802 11393
rect 7944 11370 7972 11580
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 7944 11342 8064 11370
rect 7746 11319 7748 11328
rect 7800 11319 7802 11328
rect 7748 11290 7800 11296
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7930 10976 7986 10985
rect 7524 9336 7696 9364
rect 7472 9318 7524 9324
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7484 5710 7512 6802
rect 7668 6254 7696 9336
rect 7760 7426 7788 10950
rect 7930 10911 7986 10920
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7852 8362 7880 10542
rect 7944 9382 7972 10911
rect 8036 10606 8064 11342
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8036 8945 8064 8978
rect 8022 8936 8078 8945
rect 7932 8900 7984 8906
rect 8022 8871 8078 8880
rect 7932 8842 7984 8848
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7852 8265 7880 8298
rect 7838 8256 7894 8265
rect 7838 8191 7894 8200
rect 7852 7732 7880 8191
rect 7944 7886 7972 8842
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7852 7704 7972 7732
rect 7760 7398 7880 7426
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7760 6322 7788 7278
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7562 6080 7618 6089
rect 7562 6015 7618 6024
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 4690 7512 5170
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7576 3670 7604 6015
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7668 5114 7696 5714
rect 7760 5234 7788 6258
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7668 5086 7788 5114
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7668 3602 7696 4422
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7656 3392 7708 3398
rect 7576 3340 7656 3346
rect 7576 3334 7708 3340
rect 7576 3318 7696 3334
rect 7576 3058 7604 3318
rect 7760 3194 7788 5086
rect 7852 4049 7880 7398
rect 7944 7342 7972 7704
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8036 6322 8064 8871
rect 8128 6905 8156 11494
rect 8220 11286 8248 12378
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8298 11112 8354 11121
rect 8298 11047 8354 11056
rect 8208 10600 8260 10606
rect 8206 10568 8208 10577
rect 8260 10568 8262 10577
rect 8206 10503 8262 10512
rect 8312 10266 8340 11047
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8220 9217 8248 9454
rect 8206 9208 8262 9217
rect 8206 9143 8262 9152
rect 8312 9058 8340 10202
rect 8392 9920 8444 9926
rect 8390 9888 8392 9897
rect 8444 9888 8446 9897
rect 8390 9823 8446 9832
rect 8312 9030 8432 9058
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8220 8401 8248 8842
rect 8206 8392 8262 8401
rect 8206 8327 8262 8336
rect 8312 8090 8340 8910
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7342 8248 7686
rect 8312 7449 8340 7890
rect 8298 7440 8354 7449
rect 8298 7375 8354 7384
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8114 6896 8170 6905
rect 8114 6831 8170 6840
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7944 5914 7972 6190
rect 8128 5914 8156 6666
rect 8312 6225 8340 7375
rect 8298 6216 8354 6225
rect 8298 6151 8354 6160
rect 8208 6112 8260 6118
rect 8206 6080 8208 6089
rect 8260 6080 8262 6089
rect 8206 6015 8262 6024
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 7930 5400 7986 5409
rect 7930 5335 7986 5344
rect 8024 5364 8076 5370
rect 7838 4040 7894 4049
rect 7838 3975 7894 3984
rect 7944 3942 7972 5335
rect 8024 5306 8076 5312
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 8036 3058 8064 5306
rect 8114 5264 8170 5273
rect 8114 5199 8170 5208
rect 8128 5098 8156 5199
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8128 4282 8156 4694
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8128 4185 8156 4218
rect 8114 4176 8170 4185
rect 8114 4111 8170 4120
rect 8312 4049 8340 6151
rect 8404 5030 8432 9030
rect 8496 8514 8524 10678
rect 8588 9081 8616 13330
rect 8680 9178 8708 13806
rect 8772 12918 8800 14350
rect 8852 14172 9148 14192
rect 8908 14170 8932 14172
rect 8988 14170 9012 14172
rect 9068 14170 9092 14172
rect 8930 14118 8932 14170
rect 8994 14118 9006 14170
rect 9068 14118 9070 14170
rect 8908 14116 8932 14118
rect 8988 14116 9012 14118
rect 9068 14116 9092 14118
rect 8852 14096 9148 14116
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 8852 13084 9148 13104
rect 8908 13082 8932 13084
rect 8988 13082 9012 13084
rect 9068 13082 9092 13084
rect 8930 13030 8932 13082
rect 8994 13030 9006 13082
rect 9068 13030 9070 13082
rect 8908 13028 8932 13030
rect 8988 13028 9012 13030
rect 9068 13028 9092 13030
rect 8852 13008 9148 13028
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 9232 12850 9260 13738
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9324 12714 9352 13874
rect 9416 13870 9444 14962
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9508 13394 9536 14758
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9588 14000 9640 14006
rect 9588 13942 9640 13948
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 12850 9444 13126
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9034 12336 9090 12345
rect 9034 12271 9036 12280
rect 9088 12271 9090 12280
rect 9036 12242 9088 12248
rect 9402 12200 9458 12209
rect 9402 12135 9458 12144
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 8852 11996 9148 12016
rect 8908 11994 8932 11996
rect 8988 11994 9012 11996
rect 9068 11994 9092 11996
rect 8930 11942 8932 11994
rect 8994 11942 9006 11994
rect 9068 11942 9070 11994
rect 8908 11940 8932 11942
rect 8988 11940 9012 11942
rect 9068 11940 9092 11942
rect 8852 11920 9148 11940
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 8852 10908 9148 10928
rect 8908 10906 8932 10908
rect 8988 10906 9012 10908
rect 9068 10906 9092 10908
rect 8930 10854 8932 10906
rect 8994 10854 9006 10906
rect 9068 10854 9070 10906
rect 8908 10852 8932 10854
rect 8988 10852 9012 10854
rect 9068 10852 9092 10854
rect 8852 10832 9148 10852
rect 9232 10606 9260 10950
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9218 10160 9274 10169
rect 9218 10095 9274 10104
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8772 9722 8800 9998
rect 9232 9926 9260 10095
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 8852 9820 9148 9840
rect 8908 9818 8932 9820
rect 8988 9818 9012 9820
rect 9068 9818 9092 9820
rect 8930 9766 8932 9818
rect 8994 9766 9006 9818
rect 9068 9766 9070 9818
rect 8908 9764 8932 9766
rect 8988 9764 9012 9766
rect 9068 9764 9092 9766
rect 8852 9744 9148 9764
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8574 9072 8630 9081
rect 8574 9007 8630 9016
rect 8772 8945 8800 9318
rect 8864 8974 8892 9386
rect 9126 9072 9182 9081
rect 9126 9007 9182 9016
rect 8852 8968 8904 8974
rect 8758 8936 8814 8945
rect 8852 8910 8904 8916
rect 9140 8906 9168 9007
rect 8758 8871 8814 8880
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 8852 8732 9148 8752
rect 8908 8730 8932 8732
rect 8988 8730 9012 8732
rect 9068 8730 9092 8732
rect 8930 8678 8932 8730
rect 8994 8678 9006 8730
rect 9068 8678 9070 8730
rect 8908 8676 8932 8678
rect 8988 8676 9012 8678
rect 9068 8676 9092 8678
rect 8852 8656 9148 8676
rect 8496 8486 8800 8514
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8482 8120 8538 8129
rect 8482 8055 8538 8064
rect 8496 8022 8524 8055
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8496 7177 8524 7822
rect 8588 7274 8616 8230
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8482 7168 8538 7177
rect 8482 7103 8538 7112
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8496 6304 8524 6938
rect 8588 6866 8616 7210
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8496 6276 8616 6304
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8298 4040 8354 4049
rect 8298 3975 8354 3984
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7470 2680 7526 2689
rect 7470 2615 7472 2624
rect 7524 2615 7526 2624
rect 7472 2586 7524 2592
rect 7576 2446 7604 2994
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 8036 2360 8064 2994
rect 8312 2961 8340 3538
rect 8298 2952 8354 2961
rect 8298 2887 8354 2896
rect 8208 2372 8260 2378
rect 8036 2332 8208 2360
rect 8208 2314 8260 2320
rect 8404 480 8432 4558
rect 8496 4486 8524 6122
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8588 2854 8616 6276
rect 8680 5166 8708 8366
rect 8772 7041 8800 8486
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 7886 9076 8230
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8852 7644 9148 7664
rect 8908 7642 8932 7644
rect 8988 7642 9012 7644
rect 9068 7642 9092 7644
rect 8930 7590 8932 7642
rect 8994 7590 9006 7642
rect 9068 7590 9070 7642
rect 8908 7588 8932 7590
rect 8988 7588 9012 7590
rect 9068 7588 9092 7590
rect 8852 7568 9148 7588
rect 8758 7032 8814 7041
rect 8758 6967 8814 6976
rect 9232 6934 9260 9862
rect 9324 7392 9352 12038
rect 9416 10266 9444 12135
rect 9508 11558 9536 13330
rect 9600 11762 9628 13942
rect 9692 13530 9720 14418
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9692 12374 9720 13262
rect 9784 12646 9812 13670
rect 9876 13326 9904 13874
rect 9968 13530 9996 15166
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9876 12918 9904 13126
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9784 12442 9812 12582
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9692 11898 9720 12310
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9586 11656 9642 11665
rect 9586 11591 9642 11600
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9416 8537 9444 9318
rect 9508 8809 9536 11494
rect 9600 9926 9628 11591
rect 9876 10305 9904 12854
rect 9862 10296 9918 10305
rect 9862 10231 9918 10240
rect 9862 10024 9918 10033
rect 9862 9959 9918 9968
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9588 9512 9640 9518
rect 9640 9472 9720 9500
rect 9784 9489 9812 9862
rect 9588 9454 9640 9460
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9494 8800 9550 8809
rect 9494 8735 9550 8744
rect 9600 8634 9628 9318
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9402 8528 9458 8537
rect 9402 8463 9458 8472
rect 9692 8265 9720 9472
rect 9770 9480 9826 9489
rect 9770 9415 9826 9424
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9784 9110 9812 9318
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9876 9042 9904 9959
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9968 8809 9996 13466
rect 10060 12782 10088 14214
rect 10152 13190 10180 14894
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10506 13832 10562 13841
rect 10506 13767 10562 13776
rect 10520 13530 10548 13767
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10060 11762 10088 12378
rect 10244 12322 10272 13126
rect 10336 12850 10364 13262
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10336 12442 10364 12786
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10244 12294 10456 12322
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10244 11218 10272 12174
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 10060 9625 10088 10474
rect 10046 9616 10102 9625
rect 10046 9551 10102 9560
rect 10060 9382 10088 9551
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9954 8800 10010 8809
rect 9954 8735 10010 8744
rect 10046 8664 10102 8673
rect 10046 8599 10102 8608
rect 10060 8498 10088 8599
rect 10048 8492 10100 8498
rect 9968 8452 10048 8480
rect 9862 8392 9918 8401
rect 9862 8327 9864 8336
rect 9916 8327 9918 8336
rect 9864 8298 9916 8304
rect 9968 8294 9996 8452
rect 10048 8434 10100 8440
rect 10046 8392 10102 8401
rect 10046 8327 10102 8336
rect 9956 8288 10008 8294
rect 9494 8256 9550 8265
rect 9678 8256 9734 8265
rect 9550 8214 9628 8242
rect 9494 8191 9550 8200
rect 9600 7886 9628 8214
rect 9956 8230 10008 8236
rect 9678 8191 9734 8200
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9324 7364 9444 7392
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 8772 5370 8800 6870
rect 8852 6792 8904 6798
rect 8850 6760 8852 6769
rect 9220 6792 9272 6798
rect 8904 6760 8906 6769
rect 8850 6695 8906 6704
rect 9126 6760 9182 6769
rect 9220 6734 9272 6740
rect 9126 6695 9128 6704
rect 9180 6695 9182 6704
rect 9128 6666 9180 6672
rect 8852 6556 9148 6576
rect 8908 6554 8932 6556
rect 8988 6554 9012 6556
rect 9068 6554 9092 6556
rect 8930 6502 8932 6554
rect 8994 6502 9006 6554
rect 9068 6502 9070 6554
rect 8908 6500 8932 6502
rect 8988 6500 9012 6502
rect 9068 6500 9092 6502
rect 8852 6480 9148 6500
rect 9126 6216 9182 6225
rect 9126 6151 9182 6160
rect 9140 6118 9168 6151
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 8942 5944 8998 5953
rect 8942 5879 8998 5888
rect 8956 5710 8984 5879
rect 9232 5710 9260 6734
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 8852 5468 9148 5488
rect 8908 5466 8932 5468
rect 8988 5466 9012 5468
rect 9068 5466 9092 5468
rect 8930 5414 8932 5466
rect 8994 5414 9006 5466
rect 9068 5414 9070 5466
rect 8908 5412 8932 5414
rect 8988 5412 9012 5414
rect 9068 5412 9092 5414
rect 8852 5392 9148 5412
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8852 4380 9148 4400
rect 8908 4378 8932 4380
rect 8988 4378 9012 4380
rect 9068 4378 9092 4380
rect 8930 4326 8932 4378
rect 8994 4326 9006 4378
rect 9068 4326 9070 4378
rect 8908 4324 8932 4326
rect 8988 4324 9012 4326
rect 9068 4324 9092 4326
rect 8852 4304 9148 4324
rect 8942 4176 8998 4185
rect 8998 4120 9076 4128
rect 8942 4111 8944 4120
rect 8996 4100 9076 4120
rect 8944 4082 8996 4088
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8942 4040 8998 4049
rect 8680 3534 8708 4014
rect 8942 3975 8998 3984
rect 8956 3942 8984 3975
rect 8852 3936 8904 3942
rect 8850 3904 8852 3913
rect 8944 3936 8996 3942
rect 8904 3904 8906 3913
rect 8944 3878 8996 3884
rect 8850 3839 8906 3848
rect 8850 3768 8906 3777
rect 8850 3703 8852 3712
rect 8904 3703 8906 3712
rect 8852 3674 8904 3680
rect 8758 3632 8814 3641
rect 8758 3567 8814 3576
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8772 3058 8800 3567
rect 8944 3528 8996 3534
rect 9048 3516 9076 4100
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 8996 3488 9076 3516
rect 9140 3505 9168 3538
rect 9126 3496 9182 3505
rect 8944 3470 8996 3476
rect 9126 3431 9182 3440
rect 9324 3398 9352 6598
rect 9416 5137 9444 7364
rect 9496 7336 9548 7342
rect 9494 7304 9496 7313
rect 9548 7304 9550 7313
rect 9494 7239 9550 7248
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9402 5128 9458 5137
rect 9402 5063 9458 5072
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 8852 3292 9148 3312
rect 8908 3290 8932 3292
rect 8988 3290 9012 3292
rect 9068 3290 9092 3292
rect 8930 3238 8932 3290
rect 8994 3238 9006 3290
rect 9068 3238 9070 3290
rect 8908 3236 8932 3238
rect 8988 3236 9012 3238
rect 9068 3236 9092 3238
rect 8852 3216 9148 3236
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9324 3097 9352 3130
rect 9310 3088 9366 3097
rect 8864 3058 9076 3074
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8864 3052 9088 3058
rect 8864 3046 9036 3052
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8864 2446 8892 3046
rect 9310 3023 9366 3032
rect 9036 2994 9088 3000
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 9416 2310 9444 4422
rect 9508 4078 9536 6870
rect 9600 6390 9628 7142
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9692 5914 9720 7754
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 6866 9812 7142
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9678 5808 9734 5817
rect 9784 5778 9812 6802
rect 9876 6662 9904 7346
rect 9954 6760 10010 6769
rect 9954 6695 10010 6704
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9876 6254 9904 6598
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9678 5743 9734 5752
rect 9772 5772 9824 5778
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9508 3738 9536 3878
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9600 3602 9628 5646
rect 9692 5250 9720 5743
rect 9772 5714 9824 5720
rect 9876 5370 9904 6190
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9862 5264 9918 5273
rect 9692 5222 9812 5250
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9692 4078 9720 5102
rect 9784 5030 9812 5222
rect 9862 5199 9918 5208
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9784 3942 9812 4966
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9770 3632 9826 3641
rect 9588 3596 9640 3602
rect 9770 3567 9826 3576
rect 9588 3538 9640 3544
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9600 2854 9628 3130
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9692 2582 9720 3334
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9784 2446 9812 3567
rect 9876 3194 9904 5199
rect 9968 4185 9996 6695
rect 10060 5817 10088 8327
rect 10152 8294 10180 11154
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10244 9518 10272 9998
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10244 8022 10272 9454
rect 10336 8634 10364 9998
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10336 8022 10364 8230
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10324 8016 10376 8022
rect 10324 7958 10376 7964
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 6934 10272 7686
rect 10336 7410 10364 7822
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 10138 5944 10194 5953
rect 10138 5879 10140 5888
rect 10192 5879 10194 5888
rect 10140 5850 10192 5856
rect 10232 5840 10284 5846
rect 10046 5808 10102 5817
rect 10232 5782 10284 5788
rect 10046 5743 10102 5752
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10060 4826 10088 5510
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9954 4176 10010 4185
rect 9954 4111 10010 4120
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9968 3466 9996 3878
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10048 2916 10100 2922
rect 10048 2858 10100 2864
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9968 2650 9996 2790
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9956 2508 10008 2514
rect 10060 2496 10088 2858
rect 10008 2468 10088 2496
rect 9956 2450 10008 2456
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 8852 2204 9148 2224
rect 8908 2202 8932 2204
rect 8988 2202 9012 2204
rect 9068 2202 9092 2204
rect 8930 2150 8932 2202
rect 8994 2150 9006 2202
rect 9068 2150 9070 2202
rect 8908 2148 8932 2150
rect 8988 2148 9012 2150
rect 9068 2148 9092 2150
rect 8852 2128 9148 2148
rect 10152 2106 10180 5510
rect 10244 3534 10272 5782
rect 10322 5536 10378 5545
rect 10322 5471 10378 5480
rect 10336 3602 10364 5471
rect 10428 5409 10456 12294
rect 10612 11801 10640 13670
rect 10598 11792 10654 11801
rect 10598 11727 10654 11736
rect 10704 11014 10732 14554
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10796 13938 10824 14350
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10796 12374 10824 12582
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10849 10732 10950
rect 10690 10840 10746 10849
rect 10690 10775 10746 10784
rect 10796 10305 10824 12038
rect 11072 11914 11100 14214
rect 11256 13410 11284 16520
rect 13358 15872 13414 15881
rect 13358 15807 13414 15816
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 11484 14716 11780 14736
rect 11540 14714 11564 14716
rect 11620 14714 11644 14716
rect 11700 14714 11724 14716
rect 11562 14662 11564 14714
rect 11626 14662 11638 14714
rect 11700 14662 11702 14714
rect 11540 14660 11564 14662
rect 11620 14660 11644 14662
rect 11700 14660 11724 14662
rect 11484 14640 11780 14660
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 11992 13938 12020 14282
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11484 13628 11780 13648
rect 11540 13626 11564 13628
rect 11620 13626 11644 13628
rect 11700 13626 11724 13628
rect 11562 13574 11564 13626
rect 11626 13574 11638 13626
rect 11700 13574 11702 13626
rect 11540 13572 11564 13574
rect 11620 13572 11644 13574
rect 11700 13572 11724 13574
rect 11484 13552 11780 13572
rect 11256 13382 11468 13410
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11164 12782 11192 13194
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11256 12306 11284 13262
rect 11440 13190 11468 13382
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11900 12986 11928 13670
rect 11992 13462 12020 13874
rect 12070 13832 12126 13841
rect 12070 13767 12126 13776
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11484 12540 11780 12560
rect 11540 12538 11564 12540
rect 11620 12538 11644 12540
rect 11700 12538 11724 12540
rect 11562 12486 11564 12538
rect 11626 12486 11638 12538
rect 11700 12486 11702 12538
rect 11540 12484 11564 12486
rect 11620 12484 11644 12486
rect 11700 12484 11724 12486
rect 11484 12464 11780 12484
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11072 11886 11192 11914
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10980 11665 11008 11698
rect 10966 11656 11022 11665
rect 10966 11591 11022 11600
rect 11060 11620 11112 11626
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10782 10296 10838 10305
rect 10782 10231 10838 10240
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10520 9722 10548 10066
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10603 9846 10640 9862
rect 10603 9738 10631 9846
rect 10888 9761 10916 11154
rect 10980 11150 11008 11591
rect 11060 11562 11112 11568
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10874 9752 10930 9761
rect 10508 9716 10560 9722
rect 10603 9710 10640 9738
rect 10508 9658 10560 9664
rect 10612 9586 10640 9710
rect 10784 9716 10836 9722
rect 10874 9687 10930 9696
rect 10784 9658 10836 9664
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10690 9480 10746 9489
rect 10796 9466 10824 9658
rect 10746 9438 10824 9466
rect 10690 9415 10746 9424
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10414 5400 10470 5409
rect 10414 5335 10470 5344
rect 10414 5264 10470 5273
rect 10414 5199 10470 5208
rect 10428 4622 10456 5199
rect 10520 5030 10548 8978
rect 10612 5658 10640 9318
rect 10704 8974 10732 9415
rect 10784 9376 10836 9382
rect 10782 9344 10784 9353
rect 10836 9344 10838 9353
rect 10782 9279 10838 9288
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8430 10732 8774
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10796 8129 10824 9279
rect 10888 9042 10916 9687
rect 10980 9586 11008 10542
rect 11072 10538 11100 11562
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10782 8120 10838 8129
rect 10782 8055 10838 8064
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10704 7177 10732 7958
rect 10690 7168 10746 7177
rect 10690 7103 10746 7112
rect 10612 5630 10824 5658
rect 10796 5273 10824 5630
rect 10888 5370 10916 8842
rect 10980 8838 11008 9522
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 11072 8480 11100 9998
rect 10980 8452 11100 8480
rect 10980 7426 11008 8452
rect 10980 7398 11100 7426
rect 11072 7313 11100 7398
rect 11164 7392 11192 11886
rect 11256 11218 11284 12242
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11440 11762 11468 12038
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11532 11694 11560 12242
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11704 11688 11756 11694
rect 11756 11648 11836 11676
rect 11704 11630 11756 11636
rect 11484 11452 11780 11472
rect 11540 11450 11564 11452
rect 11620 11450 11644 11452
rect 11700 11450 11724 11452
rect 11562 11398 11564 11450
rect 11626 11398 11638 11450
rect 11700 11398 11702 11450
rect 11540 11396 11564 11398
rect 11620 11396 11644 11398
rect 11700 11396 11724 11398
rect 11484 11376 11780 11396
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11256 10810 11284 11154
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11256 10130 11284 10746
rect 11532 10674 11560 10950
rect 11716 10742 11744 11154
rect 11808 11014 11836 11648
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11900 11286 11928 11494
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11704 10736 11756 10742
rect 11808 10713 11836 10950
rect 11992 10849 12020 12106
rect 11978 10840 12034 10849
rect 11978 10775 12034 10784
rect 11888 10736 11940 10742
rect 11704 10678 11756 10684
rect 11794 10704 11850 10713
rect 11520 10668 11572 10674
rect 11980 10736 12032 10742
rect 11888 10678 11940 10684
rect 11978 10704 11980 10713
rect 12032 10704 12034 10713
rect 11794 10639 11850 10648
rect 11520 10610 11572 10616
rect 11484 10364 11780 10384
rect 11540 10362 11564 10364
rect 11620 10362 11644 10364
rect 11700 10362 11724 10364
rect 11562 10310 11564 10362
rect 11626 10310 11638 10362
rect 11700 10310 11702 10362
rect 11540 10308 11564 10310
rect 11620 10308 11644 10310
rect 11700 10308 11724 10310
rect 11484 10288 11780 10308
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11256 8974 11284 10066
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11440 9722 11468 9862
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11808 9586 11836 9998
rect 11900 9994 11928 10678
rect 11978 10639 12034 10648
rect 11992 10198 12020 10639
rect 11980 10192 12032 10198
rect 11980 10134 12032 10140
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11900 9722 11928 9930
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11440 9364 11468 9522
rect 11348 9336 11468 9364
rect 11348 9160 11376 9336
rect 11484 9276 11780 9296
rect 11540 9274 11564 9276
rect 11620 9274 11644 9276
rect 11700 9274 11724 9276
rect 11562 9222 11564 9274
rect 11626 9222 11638 9274
rect 11700 9222 11702 9274
rect 11540 9220 11564 9222
rect 11620 9220 11644 9222
rect 11700 9220 11724 9222
rect 11484 9200 11780 9220
rect 11348 9132 11468 9160
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11334 8800 11390 8809
rect 11256 8498 11284 8774
rect 11334 8735 11390 8744
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11242 8392 11298 8401
rect 11242 8327 11298 8336
rect 11256 7546 11284 8327
rect 11348 7970 11376 8735
rect 11440 8430 11468 9132
rect 11808 9042 11836 9522
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11484 8188 11780 8208
rect 11540 8186 11564 8188
rect 11620 8186 11644 8188
rect 11700 8186 11724 8188
rect 11562 8134 11564 8186
rect 11626 8134 11638 8186
rect 11700 8134 11702 8186
rect 11540 8132 11564 8134
rect 11620 8132 11644 8134
rect 11700 8132 11724 8134
rect 11484 8112 11780 8132
rect 11348 7942 11560 7970
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11164 7364 11376 7392
rect 11058 7304 11114 7313
rect 11058 7239 11060 7248
rect 11112 7239 11114 7248
rect 11244 7268 11296 7274
rect 11060 7210 11112 7216
rect 11244 7210 11296 7216
rect 11256 7041 11284 7210
rect 11242 7032 11298 7041
rect 11242 6967 11298 6976
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6254 11100 6598
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11072 5778 11100 6190
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10782 5264 10838 5273
rect 10692 5228 10744 5234
rect 10782 5199 10838 5208
rect 10692 5170 10744 5176
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10704 4622 10732 5170
rect 10980 5166 11008 5646
rect 11164 5545 11192 5850
rect 11256 5642 11284 6258
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11348 5574 11376 7364
rect 11532 7290 11560 7942
rect 11702 7848 11758 7857
rect 11808 7818 11836 8978
rect 11900 8809 11928 9386
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 11886 8800 11942 8809
rect 11886 8735 11942 8744
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11900 7954 11928 8434
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11702 7783 11758 7792
rect 11796 7812 11848 7818
rect 11716 7750 11744 7783
rect 11796 7754 11848 7760
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11900 7546 11928 7890
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11532 7262 11836 7290
rect 11484 7100 11780 7120
rect 11540 7098 11564 7100
rect 11620 7098 11644 7100
rect 11700 7098 11724 7100
rect 11562 7046 11564 7098
rect 11626 7046 11638 7098
rect 11700 7046 11702 7098
rect 11540 7044 11564 7046
rect 11620 7044 11644 7046
rect 11700 7044 11724 7046
rect 11484 7024 11780 7044
rect 11808 6769 11836 7262
rect 11992 6934 12020 9046
rect 12084 8616 12112 13767
rect 12176 12186 12204 14418
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12360 14062 12572 14090
rect 12360 13870 12388 14062
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12452 13530 12480 13942
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12268 12306 12296 13330
rect 12360 12782 12388 13330
rect 12452 12782 12480 13330
rect 12544 12918 12572 14062
rect 12636 13530 12664 14214
rect 12820 14074 12848 14758
rect 13372 14550 13400 15807
rect 14094 15464 14150 15473
rect 14094 15399 14150 15408
rect 13910 15056 13966 15065
rect 13910 14991 13966 15000
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12176 12158 12388 12186
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12254 11656 12310 11665
rect 12176 10810 12204 11630
rect 12254 11591 12256 11600
rect 12308 11591 12310 11600
rect 12256 11562 12308 11568
rect 12254 11112 12310 11121
rect 12254 11047 12310 11056
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12176 9110 12204 10542
rect 12268 9382 12296 11047
rect 12360 10674 12388 12158
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12452 10606 12480 12718
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12544 12442 12572 12582
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12544 11801 12572 12106
rect 12636 11830 12664 13330
rect 12728 13258 12756 13738
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12728 12850 12756 13194
rect 12820 13025 12848 14010
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12806 13016 12862 13025
rect 12806 12951 12862 12960
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12624 11824 12676 11830
rect 12530 11792 12586 11801
rect 12624 11766 12676 11772
rect 12530 11727 12586 11736
rect 12622 11384 12678 11393
rect 12622 11319 12678 11328
rect 12530 10840 12586 10849
rect 12530 10775 12586 10784
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12438 10432 12494 10441
rect 12256 9376 12308 9382
rect 12360 9353 12388 10406
rect 12438 10367 12494 10376
rect 12452 9994 12480 10367
rect 12544 10198 12572 10775
rect 12636 10577 12664 11319
rect 12728 10742 12756 12650
rect 12912 12617 12940 13126
rect 12898 12608 12954 12617
rect 12898 12543 12954 12552
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12806 12336 12862 12345
rect 12806 12271 12862 12280
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12716 10600 12768 10606
rect 12622 10568 12678 10577
rect 12716 10542 12768 10548
rect 12622 10503 12678 10512
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12438 9888 12494 9897
rect 12438 9823 12494 9832
rect 12256 9318 12308 9324
rect 12346 9344 12402 9353
rect 12268 9217 12296 9318
rect 12346 9279 12402 9288
rect 12254 9208 12310 9217
rect 12254 9143 12310 9152
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12084 8588 12388 8616
rect 12070 8528 12126 8537
rect 12070 8463 12126 8472
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 11794 6760 11850 6769
rect 11794 6695 11850 6704
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 11484 6012 11780 6032
rect 11540 6010 11564 6012
rect 11620 6010 11644 6012
rect 11700 6010 11724 6012
rect 11562 5958 11564 6010
rect 11626 5958 11638 6010
rect 11700 5958 11702 6010
rect 11540 5956 11564 5958
rect 11620 5956 11644 5958
rect 11700 5956 11724 5958
rect 11484 5936 11780 5956
rect 11808 5642 11836 6326
rect 12084 6254 12112 8463
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11336 5568 11388 5574
rect 11150 5536 11206 5545
rect 11336 5510 11388 5516
rect 11150 5471 11206 5480
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10980 4758 11008 4966
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10414 3904 10470 3913
rect 10414 3839 10470 3848
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10336 2961 10364 3538
rect 10322 2952 10378 2961
rect 10428 2922 10456 3839
rect 10322 2887 10378 2896
rect 10416 2916 10468 2922
rect 10416 2858 10468 2864
rect 10520 2854 10548 4422
rect 10704 4078 10732 4558
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10690 3632 10746 3641
rect 10690 3567 10692 3576
rect 10744 3567 10746 3576
rect 10692 3538 10744 3544
rect 10796 3505 10824 4218
rect 11072 4162 11100 4966
rect 10980 4134 11100 4162
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10782 3496 10838 3505
rect 10782 3431 10838 3440
rect 10888 3194 10916 3878
rect 10980 3602 11008 4134
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 11072 3641 11100 3946
rect 11058 3632 11114 3641
rect 10968 3596 11020 3602
rect 11058 3567 11114 3576
rect 10968 3538 11020 3544
rect 11164 3398 11192 5034
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10600 3120 10652 3126
rect 10598 3088 10600 3097
rect 10652 3088 10654 3097
rect 10598 3023 10654 3032
rect 10600 2984 10652 2990
rect 10598 2952 10600 2961
rect 10652 2952 10654 2961
rect 10598 2887 10654 2896
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10336 2553 10364 2790
rect 10322 2544 10378 2553
rect 10322 2479 10378 2488
rect 10692 2372 10744 2378
rect 10692 2314 10744 2320
rect 10140 2100 10192 2106
rect 10140 2042 10192 2048
rect 9588 1420 9640 1426
rect 9588 1362 9640 1368
rect 9600 480 9628 1362
rect 10704 480 10732 2314
rect 10980 1057 11008 3334
rect 11256 2990 11284 4966
rect 11348 3194 11376 4966
rect 11484 4924 11780 4944
rect 11540 4922 11564 4924
rect 11620 4922 11644 4924
rect 11700 4922 11724 4924
rect 11562 4870 11564 4922
rect 11626 4870 11638 4922
rect 11700 4870 11702 4922
rect 11540 4868 11564 4870
rect 11620 4868 11644 4870
rect 11700 4868 11724 4870
rect 11484 4848 11780 4868
rect 11808 4622 11836 5578
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11794 4176 11850 4185
rect 11794 4111 11850 4120
rect 11484 3836 11780 3856
rect 11540 3834 11564 3836
rect 11620 3834 11644 3836
rect 11700 3834 11724 3836
rect 11562 3782 11564 3834
rect 11626 3782 11638 3834
rect 11700 3782 11702 3834
rect 11540 3780 11564 3782
rect 11620 3780 11644 3782
rect 11700 3780 11724 3782
rect 11484 3760 11780 3780
rect 11808 3652 11836 4111
rect 11716 3624 11836 3652
rect 11716 3534 11744 3624
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11794 3496 11850 3505
rect 11794 3431 11850 3440
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11532 3097 11560 3130
rect 11518 3088 11574 3097
rect 11808 3058 11836 3431
rect 11518 3023 11574 3032
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11334 2952 11390 2961
rect 11900 2922 11928 6054
rect 12176 5914 12204 8366
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 12162 5808 12218 5817
rect 12162 5743 12218 5752
rect 11980 5704 12032 5710
rect 11978 5672 11980 5681
rect 12032 5672 12034 5681
rect 11978 5607 12034 5616
rect 11978 4856 12034 4865
rect 11978 4791 11980 4800
rect 12032 4791 12034 4800
rect 11980 4762 12032 4768
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11992 3534 12020 4558
rect 12176 3670 12204 5743
rect 12268 4282 12296 8230
rect 12360 7721 12388 8588
rect 12452 7834 12480 9823
rect 12544 9761 12572 9998
rect 12530 9752 12586 9761
rect 12530 9687 12586 9696
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12544 8090 12572 8842
rect 12636 8090 12664 10503
rect 12728 10198 12756 10542
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12714 8936 12770 8945
rect 12714 8871 12770 8880
rect 12728 8498 12756 8871
rect 12820 8650 12848 12271
rect 12912 11393 12940 12378
rect 12898 11384 12954 11393
rect 12898 11319 12954 11328
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12912 10713 12940 10746
rect 12898 10704 12954 10713
rect 12898 10639 12954 10648
rect 12898 10296 12954 10305
rect 12898 10231 12954 10240
rect 12912 10198 12940 10231
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 12912 10033 12940 10134
rect 12898 10024 12954 10033
rect 12898 9959 12954 9968
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12912 8838 12940 9522
rect 13004 9450 13032 14418
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13096 14074 13124 14350
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13648 13938 13676 14282
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13084 12776 13136 12782
rect 13136 12736 13216 12764
rect 13084 12718 13136 12724
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13096 10985 13124 12582
rect 13188 11286 13216 12736
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 13082 10976 13138 10985
rect 13082 10911 13138 10920
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 13096 10470 13124 10610
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13188 10130 13216 11222
rect 13280 11121 13308 13806
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13464 13530 13492 13670
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13372 12238 13400 12650
rect 13556 12594 13584 13670
rect 13648 13258 13676 13874
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 13648 12646 13676 13194
rect 13464 12566 13584 12594
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13464 12442 13492 12566
rect 13740 12458 13768 14554
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13832 14006 13860 14350
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13818 13288 13874 13297
rect 13818 13223 13874 13232
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13556 12430 13768 12458
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13372 11694 13400 12174
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13266 11112 13322 11121
rect 13266 11047 13322 11056
rect 13266 10976 13322 10985
rect 13266 10911 13322 10920
rect 13280 10588 13308 10911
rect 13372 10742 13400 11630
rect 13464 10742 13492 12242
rect 13556 10849 13584 12430
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13542 10840 13598 10849
rect 13542 10775 13598 10784
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13634 10704 13690 10713
rect 13634 10639 13690 10648
rect 13648 10606 13676 10639
rect 13636 10600 13688 10606
rect 13280 10560 13584 10588
rect 13360 10464 13412 10470
rect 13556 10418 13584 10560
rect 13636 10542 13688 10548
rect 13360 10406 13412 10412
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13096 9586 13124 9998
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 13188 9874 13216 9930
rect 13188 9846 13308 9874
rect 13174 9752 13230 9761
rect 13174 9687 13230 9696
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 12990 9344 13046 9353
rect 13096 9330 13124 9386
rect 13046 9302 13124 9330
rect 12990 9279 13046 9288
rect 13082 9208 13138 9217
rect 13082 9143 13138 9152
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12820 8622 13032 8650
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 13004 7970 13032 8622
rect 12820 7942 13032 7970
rect 12452 7806 12756 7834
rect 12532 7744 12584 7750
rect 12346 7712 12402 7721
rect 12532 7686 12584 7692
rect 12346 7647 12402 7656
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12452 6458 12480 6802
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12360 5681 12388 6394
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12346 5672 12402 5681
rect 12452 5658 12480 6258
rect 12544 5846 12572 7686
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12636 6934 12664 7278
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12636 5710 12664 6870
rect 12624 5704 12676 5710
rect 12452 5630 12572 5658
rect 12624 5646 12676 5652
rect 12346 5607 12402 5616
rect 12346 4720 12402 4729
rect 12346 4655 12348 4664
rect 12400 4655 12402 4664
rect 12348 4626 12400 4632
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12164 3664 12216 3670
rect 12164 3606 12216 3612
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11992 3058 12020 3470
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11978 2952 12034 2961
rect 11334 2887 11390 2896
rect 11888 2916 11940 2922
rect 11058 2680 11114 2689
rect 11348 2650 11376 2887
rect 11978 2887 12034 2896
rect 11888 2858 11940 2864
rect 11484 2748 11780 2768
rect 11540 2746 11564 2748
rect 11620 2746 11644 2748
rect 11700 2746 11724 2748
rect 11562 2694 11564 2746
rect 11626 2694 11638 2746
rect 11700 2694 11702 2746
rect 11540 2692 11564 2694
rect 11620 2692 11644 2694
rect 11700 2692 11724 2694
rect 11484 2672 11780 2692
rect 11058 2615 11060 2624
rect 11112 2615 11114 2624
rect 11336 2644 11388 2650
rect 11060 2586 11112 2592
rect 11336 2586 11388 2592
rect 11992 2582 12020 2887
rect 11980 2576 12032 2582
rect 11794 2544 11850 2553
rect 11980 2518 12032 2524
rect 12268 2514 12296 3674
rect 12452 3670 12480 4218
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12438 3360 12494 3369
rect 12360 2582 12388 3334
rect 12438 3295 12494 3304
rect 12452 2990 12480 3295
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12544 2582 12572 5630
rect 12728 4593 12756 7806
rect 12820 6322 12848 7942
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12912 7721 12940 7822
rect 13096 7750 13124 9143
rect 13084 7744 13136 7750
rect 12898 7712 12954 7721
rect 13084 7686 13136 7692
rect 12898 7647 12954 7656
rect 13188 6746 13216 9687
rect 13280 6798 13308 9846
rect 13372 9489 13400 10406
rect 13464 10390 13584 10418
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13358 9480 13414 9489
rect 13358 9415 13414 9424
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13372 7342 13400 8026
rect 13464 7857 13492 10390
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13556 9722 13584 10066
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13556 9042 13584 9658
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13556 8945 13584 8978
rect 13542 8936 13598 8945
rect 13542 8871 13598 8880
rect 13542 8800 13598 8809
rect 13542 8735 13598 8744
rect 13450 7848 13506 7857
rect 13450 7783 13506 7792
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 13004 6718 13216 6746
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12820 5914 12848 6054
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12912 5642 12940 6666
rect 13004 6225 13032 6718
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13096 6322 13124 6394
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13188 6254 13216 6598
rect 13176 6248 13228 6254
rect 12990 6216 13046 6225
rect 13176 6190 13228 6196
rect 12990 6151 13046 6160
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12820 4622 12848 4966
rect 12808 4616 12860 4622
rect 12714 4584 12770 4593
rect 12808 4558 12860 4564
rect 12714 4519 12770 4528
rect 12728 3720 12756 4519
rect 13004 3924 13032 6054
rect 13096 4690 13124 6054
rect 13188 5778 13216 6190
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13188 5166 13216 5714
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13188 4078 13216 5102
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13004 3896 13216 3924
rect 12808 3732 12860 3738
rect 12728 3692 12808 3720
rect 12808 3674 12860 3680
rect 12714 3632 12770 3641
rect 12624 3596 12676 3602
rect 12714 3567 12770 3576
rect 12624 3538 12676 3544
rect 12636 2922 12664 3538
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 12728 2650 12756 3567
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12912 3058 12940 3470
rect 13084 3460 13136 3466
rect 13084 3402 13136 3408
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 12912 2938 12940 2994
rect 12820 2910 12940 2938
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 11794 2479 11796 2488
rect 11848 2479 11850 2488
rect 12256 2508 12308 2514
rect 11796 2450 11848 2456
rect 12256 2450 12308 2456
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11348 2106 11376 2382
rect 12820 2378 12848 2910
rect 12808 2372 12860 2378
rect 12808 2314 12860 2320
rect 12820 2106 12848 2314
rect 11336 2100 11388 2106
rect 11336 2042 11388 2048
rect 12808 2100 12860 2106
rect 12808 2042 12860 2048
rect 13096 1850 13124 3402
rect 13188 2990 13216 3896
rect 13280 3602 13308 6734
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13372 5030 13400 5714
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13556 4049 13584 8735
rect 13648 8537 13676 10406
rect 13740 9518 13768 12174
rect 13832 12102 13860 13223
rect 13924 12345 13952 14991
rect 14108 14822 14136 15399
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 14482 14136 14758
rect 14660 14482 14688 14826
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14016 13802 14044 14418
rect 14830 14240 14886 14249
rect 14116 14172 14412 14192
rect 14830 14175 14886 14184
rect 14172 14170 14196 14172
rect 14252 14170 14276 14172
rect 14332 14170 14356 14172
rect 14194 14118 14196 14170
rect 14258 14118 14270 14170
rect 14332 14118 14334 14170
rect 14172 14116 14196 14118
rect 14252 14116 14276 14118
rect 14332 14116 14356 14118
rect 14116 14096 14412 14116
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14004 13796 14056 13802
rect 14004 13738 14056 13744
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14116 13084 14412 13104
rect 14172 13082 14196 13084
rect 14252 13082 14276 13084
rect 14332 13082 14356 13084
rect 14194 13030 14196 13082
rect 14258 13030 14270 13082
rect 14332 13030 14334 13082
rect 14172 13028 14196 13030
rect 14252 13028 14276 13030
rect 14332 13028 14356 13030
rect 14116 13008 14412 13028
rect 13910 12336 13966 12345
rect 13910 12271 13966 12280
rect 14476 12209 14504 13466
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14462 12200 14518 12209
rect 14004 12164 14056 12170
rect 14462 12135 14518 12144
rect 14004 12106 14056 12112
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13910 11928 13966 11937
rect 14016 11898 14044 12106
rect 14116 11996 14412 12016
rect 14172 11994 14196 11996
rect 14252 11994 14276 11996
rect 14332 11994 14356 11996
rect 14194 11942 14196 11994
rect 14258 11942 14270 11994
rect 14332 11942 14334 11994
rect 14172 11940 14196 11942
rect 14252 11940 14276 11942
rect 14332 11940 14356 11942
rect 14116 11920 14412 11940
rect 13910 11863 13966 11872
rect 14004 11892 14056 11898
rect 13924 11218 13952 11863
rect 14004 11834 14056 11840
rect 14372 11688 14424 11694
rect 14372 11630 14424 11636
rect 14384 11286 14412 11630
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13832 10674 13860 11154
rect 14384 11150 14412 11222
rect 14372 11144 14424 11150
rect 14370 11112 14372 11121
rect 14424 11112 14426 11121
rect 14370 11047 14426 11056
rect 14384 11021 14412 11047
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 13832 9654 13860 10474
rect 13924 10441 13952 10950
rect 13910 10432 13966 10441
rect 13910 10367 13966 10376
rect 13912 10192 13964 10198
rect 14016 10180 14044 10950
rect 14116 10908 14412 10928
rect 14172 10906 14196 10908
rect 14252 10906 14276 10908
rect 14332 10906 14356 10908
rect 14194 10854 14196 10906
rect 14258 10854 14270 10906
rect 14332 10854 14334 10906
rect 14172 10852 14196 10854
rect 14252 10852 14276 10854
rect 14332 10852 14356 10854
rect 14116 10832 14412 10852
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 10266 14228 10406
rect 14476 10266 14504 10610
rect 14568 10470 14596 12922
rect 14752 12617 14780 13806
rect 14738 12608 14794 12617
rect 14738 12543 14794 12552
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14660 11082 14688 12174
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14646 10976 14702 10985
rect 14646 10911 14702 10920
rect 14660 10674 14688 10911
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 13964 10152 14044 10180
rect 14752 10180 14780 12038
rect 14844 10305 14872 14175
rect 15028 13530 15056 16623
rect 15750 16520 15806 17000
rect 15106 15328 15162 15337
rect 15106 15263 15162 15272
rect 15120 15026 15148 15263
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15106 14648 15162 14657
rect 15106 14583 15162 14592
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 14924 12368 14976 12374
rect 14924 12310 14976 12316
rect 14936 12073 14964 12310
rect 14922 12064 14978 12073
rect 14922 11999 14978 12008
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14830 10296 14886 10305
rect 14936 10282 14964 10950
rect 15028 10690 15056 13330
rect 15120 11121 15148 14583
rect 15764 14550 15792 16520
rect 16210 16280 16266 16289
rect 16210 16215 16266 16224
rect 16224 15337 16252 16215
rect 16210 15328 16266 15337
rect 16210 15263 16266 15272
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 15396 14074 15424 14350
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15212 11694 15240 13330
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15304 12306 15332 12582
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15396 12238 15424 12650
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15396 11898 15424 12174
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15488 11286 15516 14214
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15580 12442 15608 13126
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15566 11792 15622 11801
rect 15566 11727 15622 11736
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15106 11112 15162 11121
rect 15106 11047 15162 11056
rect 15382 10976 15438 10985
rect 15382 10911 15438 10920
rect 15290 10840 15346 10849
rect 15290 10775 15346 10784
rect 15028 10662 15148 10690
rect 15120 10554 15148 10662
rect 15120 10526 15240 10554
rect 14936 10254 15148 10282
rect 14830 10231 14886 10240
rect 14752 10152 14872 10180
rect 13912 10134 13964 10140
rect 14096 10124 14148 10130
rect 14016 10084 14096 10112
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13924 9518 13952 9862
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 14016 9364 14044 10084
rect 14096 10066 14148 10072
rect 14844 10044 14872 10152
rect 14752 10016 14872 10044
rect 14116 9820 14412 9840
rect 14172 9818 14196 9820
rect 14252 9818 14276 9820
rect 14332 9818 14356 9820
rect 14194 9766 14196 9818
rect 14258 9766 14270 9818
rect 14332 9766 14334 9818
rect 14172 9764 14196 9766
rect 14252 9764 14276 9766
rect 14332 9764 14356 9766
rect 14116 9744 14412 9764
rect 14554 9616 14610 9625
rect 14554 9551 14610 9560
rect 13924 9336 14044 9364
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13832 8673 13860 8978
rect 13818 8664 13874 8673
rect 13818 8599 13874 8608
rect 13634 8528 13690 8537
rect 13634 8463 13690 8472
rect 13832 8362 13860 8599
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13636 8288 13688 8294
rect 13688 8248 13768 8276
rect 13924 8265 13952 9336
rect 14016 9110 14044 9141
rect 14004 9104 14056 9110
rect 14002 9072 14004 9081
rect 14056 9072 14058 9081
rect 14002 9007 14058 9016
rect 14016 8548 14044 9007
rect 14116 8732 14412 8752
rect 14172 8730 14196 8732
rect 14252 8730 14276 8732
rect 14332 8730 14356 8732
rect 14194 8678 14196 8730
rect 14258 8678 14270 8730
rect 14332 8678 14334 8730
rect 14172 8676 14196 8678
rect 14252 8676 14276 8678
rect 14332 8676 14356 8678
rect 14116 8656 14412 8676
rect 14016 8520 14136 8548
rect 14108 8430 14136 8520
rect 14462 8528 14518 8537
rect 14462 8463 14518 8472
rect 14476 8430 14504 8463
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14016 8294 14044 8366
rect 14004 8288 14056 8294
rect 13636 8230 13688 8236
rect 13634 8120 13690 8129
rect 13740 8090 13768 8248
rect 13910 8256 13966 8265
rect 14004 8230 14056 8236
rect 13910 8191 13966 8200
rect 13634 8055 13690 8064
rect 13728 8084 13780 8090
rect 13648 7585 13676 8055
rect 13728 8026 13780 8032
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 13818 7984 13874 7993
rect 13818 7919 13820 7928
rect 13872 7919 13874 7928
rect 14096 7948 14148 7954
rect 13820 7890 13872 7896
rect 14096 7890 14148 7896
rect 13728 7880 13780 7886
rect 14108 7834 14136 7890
rect 13728 7822 13780 7828
rect 13634 7576 13690 7585
rect 13634 7511 13690 7520
rect 13740 7410 13768 7822
rect 13924 7806 14136 7834
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13542 4040 13598 4049
rect 13542 3975 13598 3984
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 13648 3097 13676 7142
rect 13740 6458 13768 7346
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13728 5160 13780 5166
rect 13832 5148 13860 7686
rect 13924 6730 13952 7806
rect 14116 7644 14412 7664
rect 14172 7642 14196 7644
rect 14252 7642 14276 7644
rect 14332 7642 14356 7644
rect 14194 7590 14196 7642
rect 14258 7590 14270 7642
rect 14332 7590 14334 7642
rect 14172 7588 14196 7590
rect 14252 7588 14276 7590
rect 14332 7588 14356 7590
rect 14116 7568 14412 7588
rect 14476 7546 14504 8026
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13780 5120 13860 5148
rect 13728 5102 13780 5108
rect 13740 3618 13768 5102
rect 13924 5098 13952 6258
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13832 3738 13860 4626
rect 13924 4622 13952 5034
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13924 3942 13952 4422
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13740 3590 13860 3618
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13740 3194 13768 3470
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13634 3088 13690 3097
rect 13832 3058 13860 3590
rect 13634 3023 13690 3032
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 13820 2440 13872 2446
rect 14016 2417 14044 7482
rect 14462 7304 14518 7313
rect 14462 7239 14518 7248
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14200 7002 14228 7142
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14116 6556 14412 6576
rect 14172 6554 14196 6556
rect 14252 6554 14276 6556
rect 14332 6554 14356 6556
rect 14194 6502 14196 6554
rect 14258 6502 14270 6554
rect 14332 6502 14334 6554
rect 14172 6500 14196 6502
rect 14252 6500 14276 6502
rect 14332 6500 14356 6502
rect 14116 6480 14412 6500
rect 14116 5468 14412 5488
rect 14172 5466 14196 5468
rect 14252 5466 14276 5468
rect 14332 5466 14356 5468
rect 14194 5414 14196 5466
rect 14258 5414 14270 5466
rect 14332 5414 14334 5466
rect 14172 5412 14196 5414
rect 14252 5412 14276 5414
rect 14332 5412 14356 5414
rect 14116 5392 14412 5412
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14108 4729 14136 5238
rect 14476 4826 14504 7239
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14094 4720 14150 4729
rect 14094 4655 14150 4664
rect 14116 4380 14412 4400
rect 14172 4378 14196 4380
rect 14252 4378 14276 4380
rect 14332 4378 14356 4380
rect 14194 4326 14196 4378
rect 14258 4326 14270 4378
rect 14332 4326 14334 4378
rect 14172 4324 14196 4326
rect 14252 4324 14276 4326
rect 14332 4324 14356 4326
rect 14116 4304 14412 4324
rect 14464 4004 14516 4010
rect 14464 3946 14516 3952
rect 14116 3292 14412 3312
rect 14172 3290 14196 3292
rect 14252 3290 14276 3292
rect 14332 3290 14356 3292
rect 14194 3238 14196 3290
rect 14258 3238 14270 3290
rect 14332 3238 14334 3290
rect 14172 3236 14196 3238
rect 14252 3236 14276 3238
rect 14332 3236 14356 3238
rect 14116 3216 14412 3236
rect 14476 3058 14504 3946
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14568 2514 14596 9551
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14660 8401 14688 8978
rect 14646 8392 14702 8401
rect 14646 8327 14702 8336
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14660 7449 14688 7890
rect 14646 7440 14702 7449
rect 14646 7375 14702 7384
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14660 5302 14688 7142
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14752 4706 14780 10016
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14844 7041 14872 9386
rect 14936 9178 14964 9386
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14922 8528 14978 8537
rect 15028 8498 15056 9862
rect 14922 8463 14978 8472
rect 15016 8492 15068 8498
rect 14936 7410 14964 8463
rect 15016 8434 15068 8440
rect 15120 8378 15148 10254
rect 15212 9110 15240 10526
rect 15304 10169 15332 10775
rect 15290 10160 15346 10169
rect 15290 10095 15346 10104
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15028 8350 15148 8378
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14830 7032 14886 7041
rect 14830 6967 14886 6976
rect 14922 6760 14978 6769
rect 14922 6695 14978 6704
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14660 4678 14780 4706
rect 14660 3058 14688 4678
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 13820 2382 13872 2388
rect 14002 2408 14058 2417
rect 12912 1822 13124 1850
rect 11796 1148 11848 1154
rect 11796 1090 11848 1096
rect 10966 1048 11022 1057
rect 10966 983 11022 992
rect 11808 480 11836 1090
rect 12912 480 12940 1822
rect 13832 1426 13860 2382
rect 14002 2343 14058 2352
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 14116 2204 14412 2224
rect 14172 2202 14196 2204
rect 14252 2202 14276 2204
rect 14332 2202 14356 2204
rect 14194 2150 14196 2202
rect 14258 2150 14270 2202
rect 14332 2150 14334 2202
rect 14172 2148 14196 2150
rect 14252 2148 14276 2150
rect 14332 2148 14356 2150
rect 14116 2128 14412 2148
rect 13820 1420 13872 1426
rect 13820 1362 13872 1368
rect 14476 1306 14504 2314
rect 14752 1873 14780 4490
rect 14738 1864 14794 1873
rect 14738 1799 14794 1808
rect 14844 1465 14872 6598
rect 14936 6089 14964 6695
rect 14922 6080 14978 6089
rect 14922 6015 14978 6024
rect 15028 5522 15056 8350
rect 15106 8120 15162 8129
rect 15106 8055 15162 8064
rect 15120 7818 15148 8055
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15120 6798 15148 7346
rect 15212 6866 15240 8842
rect 15304 8430 15332 9862
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15290 7848 15346 7857
rect 15290 7783 15346 7792
rect 15304 7750 15332 7783
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15120 6186 15148 6734
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15120 5642 15148 6122
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15028 5494 15148 5522
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14936 3890 14964 4966
rect 15028 4457 15056 5306
rect 15014 4448 15070 4457
rect 15014 4383 15070 4392
rect 14936 3862 15056 3890
rect 14830 1456 14886 1465
rect 14830 1391 14886 1400
rect 14108 1278 14504 1306
rect 14108 480 14136 1278
rect 15028 649 15056 3862
rect 15120 3641 15148 5494
rect 15212 4826 15240 6122
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15304 5914 15332 6054
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15304 5098 15332 5578
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15304 4706 15332 5034
rect 15212 4678 15332 4706
rect 15212 4622 15240 4678
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15212 4282 15240 4558
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15106 3632 15162 3641
rect 15106 3567 15162 3576
rect 15212 3534 15240 4218
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15014 640 15070 649
rect 15014 575 15070 584
rect 3054 232 3110 241
rect 3054 167 3110 176
rect 3882 0 3938 480
rect 5078 0 5134 480
rect 6182 0 6238 480
rect 7286 0 7342 480
rect 8390 0 8446 480
rect 9586 0 9642 480
rect 10690 0 10746 480
rect 11794 0 11850 480
rect 12898 0 12954 480
rect 14094 0 14150 480
rect 15120 241 15148 3334
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 15212 480 15240 2858
rect 15396 2514 15424 10911
rect 15580 10130 15608 11727
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15474 9480 15530 9489
rect 15474 9415 15530 9424
rect 15488 8430 15516 9415
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15488 7206 15516 8366
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15580 7002 15608 10066
rect 15672 9353 15700 13670
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15856 11626 15884 12174
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15750 11248 15806 11257
rect 15750 11183 15806 11192
rect 15658 9344 15714 9353
rect 15658 9279 15714 9288
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15580 5794 15608 6938
rect 15672 6497 15700 9114
rect 15764 7002 15792 11183
rect 15856 11150 15884 11562
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15948 10606 15976 13874
rect 16132 13326 16160 14350
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16132 11830 16160 13262
rect 16120 11824 16172 11830
rect 16120 11766 16172 11772
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15856 9110 15884 10406
rect 15948 9722 15976 10542
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8498 15884 8910
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15856 7886 15884 8434
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 15752 6996 15804 7002
rect 15804 6956 15884 6984
rect 15752 6938 15804 6944
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15658 6488 15714 6497
rect 15658 6423 15714 6432
rect 15764 6361 15792 6734
rect 15750 6352 15806 6361
rect 15750 6287 15806 6296
rect 15750 6216 15806 6225
rect 15750 6151 15806 6160
rect 15764 5914 15792 6151
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15580 5766 15700 5794
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15580 4826 15608 5646
rect 15672 5574 15700 5766
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15672 3602 15700 5510
rect 15752 4616 15804 4622
rect 15750 4584 15752 4593
rect 15804 4584 15806 4593
rect 15750 4519 15806 4528
rect 15856 4185 15884 6956
rect 15948 6934 15976 7346
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 16040 6866 16068 11630
rect 16132 10742 16160 11766
rect 16120 10736 16172 10742
rect 16120 10678 16172 10684
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16132 8906 16160 10202
rect 16224 9178 16252 15263
rect 16302 12608 16358 12617
rect 16302 12543 16358 12552
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16120 8900 16172 8906
rect 16120 8842 16172 8848
rect 16132 8673 16160 8842
rect 16118 8664 16174 8673
rect 16118 8599 16174 8608
rect 16316 7954 16344 12543
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 15842 4176 15898 4185
rect 15842 4111 15898 4120
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 16040 1154 16068 3946
rect 16304 2916 16356 2922
rect 16304 2858 16356 2864
rect 16028 1148 16080 1154
rect 16028 1090 16080 1096
rect 16316 480 16344 2858
rect 16408 2689 16436 11494
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16500 10810 16528 11154
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16394 2680 16450 2689
rect 16394 2615 16450 2624
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17420 480 17448 2518
rect 15106 232 15162 241
rect 15106 167 15162 176
rect 15198 0 15254 480
rect 16302 0 16358 480
rect 17406 0 17462 480
<< via2 >>
rect 7654 16632 7710 16688
rect 4066 16224 4122 16280
rect 2686 15816 2742 15872
rect 2318 13232 2374 13288
rect 1398 8744 1454 8800
rect 1306 6840 1362 6896
rect 1306 5616 1362 5672
rect 1858 9968 1914 10024
rect 1582 7384 1638 7440
rect 1950 9016 2006 9072
rect 3974 15408 4030 15464
rect 2594 11600 2650 11656
rect 1398 4392 1454 4448
rect 1674 3984 1730 4040
rect 846 2624 902 2680
rect 2502 9832 2558 9888
rect 2502 8916 2504 8936
rect 2504 8916 2556 8936
rect 2556 8916 2558 8936
rect 2502 8880 2558 8916
rect 3588 14170 3644 14172
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3588 14118 3614 14170
rect 3614 14118 3644 14170
rect 3668 14118 3678 14170
rect 3678 14118 3724 14170
rect 3748 14118 3794 14170
rect 3794 14118 3804 14170
rect 3828 14118 3858 14170
rect 3858 14118 3884 14170
rect 3588 14116 3644 14118
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3514 13776 3570 13832
rect 4066 15000 4122 15056
rect 4066 14592 4122 14648
rect 6220 14714 6276 14716
rect 6300 14714 6356 14716
rect 6380 14714 6436 14716
rect 6460 14714 6516 14716
rect 6220 14662 6246 14714
rect 6246 14662 6276 14714
rect 6300 14662 6310 14714
rect 6310 14662 6356 14714
rect 6380 14662 6426 14714
rect 6426 14662 6436 14714
rect 6460 14662 6490 14714
rect 6490 14662 6516 14714
rect 6220 14660 6276 14662
rect 6300 14660 6356 14662
rect 6380 14660 6436 14662
rect 6460 14660 6516 14662
rect 3330 12824 3386 12880
rect 3588 13082 3644 13084
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3588 13030 3614 13082
rect 3614 13030 3644 13082
rect 3668 13030 3678 13082
rect 3678 13030 3724 13082
rect 3748 13030 3794 13082
rect 3794 13030 3804 13082
rect 3828 13030 3858 13082
rect 3858 13030 3884 13082
rect 3588 13028 3644 13030
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 2686 9580 2742 9616
rect 2686 9560 2688 9580
rect 2688 9560 2740 9580
rect 2740 9560 2742 9580
rect 2778 9152 2834 9208
rect 2686 8608 2742 8664
rect 2594 7268 2650 7304
rect 2594 7248 2596 7268
rect 2596 7248 2648 7268
rect 2648 7248 2650 7268
rect 2410 5752 2466 5808
rect 1950 1808 2006 1864
rect 2778 6840 2834 6896
rect 3422 12280 3478 12336
rect 3330 10784 3386 10840
rect 3588 11994 3644 11996
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3588 11942 3614 11994
rect 3614 11942 3644 11994
rect 3668 11942 3678 11994
rect 3678 11942 3724 11994
rect 3748 11942 3794 11994
rect 3794 11942 3804 11994
rect 3828 11942 3858 11994
rect 3858 11942 3884 11994
rect 3588 11940 3644 11942
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3882 11192 3938 11248
rect 3588 10906 3644 10908
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3588 10854 3614 10906
rect 3614 10854 3644 10906
rect 3668 10854 3678 10906
rect 3678 10854 3724 10906
rect 3748 10854 3794 10906
rect 3794 10854 3804 10906
rect 3828 10854 3858 10906
rect 3858 10854 3884 10906
rect 3588 10852 3644 10854
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3422 10240 3478 10296
rect 3698 10376 3754 10432
rect 3588 9818 3644 9820
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3588 9766 3614 9818
rect 3614 9766 3644 9818
rect 3668 9766 3678 9818
rect 3678 9766 3724 9818
rect 3748 9766 3794 9818
rect 3794 9766 3804 9818
rect 3828 9766 3858 9818
rect 3858 9766 3884 9818
rect 3588 9764 3644 9766
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3238 9288 3294 9344
rect 3054 8336 3110 8392
rect 2870 6432 2926 6488
rect 3588 8730 3644 8732
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3588 8678 3614 8730
rect 3614 8678 3644 8730
rect 3668 8678 3678 8730
rect 3678 8678 3724 8730
rect 3748 8678 3794 8730
rect 3794 8678 3804 8730
rect 3828 8678 3858 8730
rect 3858 8678 3884 8730
rect 3588 8676 3644 8678
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 2962 5752 3018 5808
rect 2686 3440 2742 3496
rect 3054 5344 3110 5400
rect 2870 4800 2926 4856
rect 2686 2488 2742 2544
rect 2962 2896 3018 2952
rect 2502 992 2558 1048
rect 3422 6976 3478 7032
rect 3422 6860 3478 6896
rect 3422 6840 3424 6860
rect 3424 6840 3476 6860
rect 3476 6840 3478 6860
rect 3330 2916 3386 2952
rect 3330 2896 3332 2916
rect 3332 2896 3384 2916
rect 3384 2896 3386 2916
rect 4066 11212 4122 11248
rect 4066 11192 4068 11212
rect 4068 11192 4120 11212
rect 4120 11192 4122 11212
rect 4158 9832 4214 9888
rect 4342 10920 4398 10976
rect 4342 10784 4398 10840
rect 4250 9596 4252 9616
rect 4252 9596 4304 9616
rect 4304 9596 4306 9616
rect 4250 9560 4306 9596
rect 4250 9152 4306 9208
rect 4066 8200 4122 8256
rect 3588 7642 3644 7644
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3588 7590 3614 7642
rect 3614 7590 3644 7642
rect 3668 7590 3678 7642
rect 3678 7590 3724 7642
rect 3748 7590 3794 7642
rect 3794 7590 3804 7642
rect 3828 7590 3858 7642
rect 3858 7590 3884 7642
rect 3588 7588 3644 7590
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3588 6554 3644 6556
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3588 6502 3614 6554
rect 3614 6502 3644 6554
rect 3668 6502 3678 6554
rect 3678 6502 3724 6554
rect 3748 6502 3794 6554
rect 3794 6502 3804 6554
rect 3828 6502 3858 6554
rect 3858 6502 3884 6554
rect 3588 6500 3644 6502
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3514 6024 3570 6080
rect 3588 5466 3644 5468
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3588 5414 3614 5466
rect 3614 5414 3644 5466
rect 3668 5414 3678 5466
rect 3678 5414 3724 5466
rect 3748 5414 3794 5466
rect 3794 5414 3804 5466
rect 3828 5414 3858 5466
rect 3858 5414 3884 5466
rect 3588 5412 3644 5414
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3606 5072 3662 5128
rect 3588 4378 3644 4380
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3588 4326 3614 4378
rect 3614 4326 3644 4378
rect 3668 4326 3678 4378
rect 3678 4326 3724 4378
rect 3748 4326 3794 4378
rect 3794 4326 3804 4378
rect 3828 4326 3858 4378
rect 3858 4326 3884 4378
rect 3588 4324 3644 4326
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3606 3712 3662 3768
rect 3882 3576 3938 3632
rect 3606 3440 3662 3496
rect 3882 3460 3938 3496
rect 3882 3440 3884 3460
rect 3884 3440 3936 3460
rect 3936 3440 3938 3460
rect 3588 3290 3644 3292
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3588 3238 3614 3290
rect 3614 3238 3644 3290
rect 3668 3238 3678 3290
rect 3678 3238 3724 3290
rect 3748 3238 3794 3290
rect 3794 3238 3804 3290
rect 3828 3238 3858 3290
rect 3858 3238 3884 3290
rect 3588 3236 3644 3238
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3422 2216 3478 2272
rect 3588 2202 3644 2204
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3588 2150 3614 2202
rect 3614 2150 3644 2202
rect 3668 2150 3678 2202
rect 3678 2150 3724 2202
rect 3748 2150 3794 2202
rect 3794 2150 3804 2202
rect 3828 2150 3858 2202
rect 3858 2150 3884 2202
rect 3588 2148 3644 2150
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 4158 7792 4214 7848
rect 4250 7520 4306 7576
rect 4066 3032 4122 3088
rect 4526 12416 4582 12472
rect 4618 11736 4674 11792
rect 4710 9832 4766 9888
rect 4710 9424 4766 9480
rect 5446 13912 5502 13968
rect 5170 11328 5226 11384
rect 5170 11212 5226 11248
rect 5170 11192 5172 11212
rect 5172 11192 5224 11212
rect 5224 11192 5226 11212
rect 4434 7792 4490 7848
rect 4342 6568 4398 6624
rect 5170 10784 5226 10840
rect 5170 10512 5226 10568
rect 4434 6024 4490 6080
rect 4342 5344 4398 5400
rect 4802 6160 4858 6216
rect 4618 5208 4674 5264
rect 4710 5072 4766 5128
rect 4342 3032 4398 3088
rect 4894 3168 4950 3224
rect 4802 2896 4858 2952
rect 5906 11620 5962 11656
rect 5906 11600 5908 11620
rect 5908 11600 5960 11620
rect 5960 11600 5962 11620
rect 5722 10104 5778 10160
rect 5906 10240 5962 10296
rect 5906 9832 5962 9888
rect 5722 7792 5778 7848
rect 5446 6160 5502 6216
rect 5630 5208 5686 5264
rect 5354 3304 5410 3360
rect 5446 2760 5502 2816
rect 5630 2760 5686 2816
rect 6220 13626 6276 13628
rect 6300 13626 6356 13628
rect 6380 13626 6436 13628
rect 6460 13626 6516 13628
rect 6220 13574 6246 13626
rect 6246 13574 6276 13626
rect 6300 13574 6310 13626
rect 6310 13574 6356 13626
rect 6380 13574 6426 13626
rect 6426 13574 6436 13626
rect 6460 13574 6490 13626
rect 6490 13574 6516 13626
rect 6220 13572 6276 13574
rect 6300 13572 6356 13574
rect 6380 13572 6436 13574
rect 6460 13572 6516 13574
rect 6220 12538 6276 12540
rect 6300 12538 6356 12540
rect 6380 12538 6436 12540
rect 6460 12538 6516 12540
rect 6220 12486 6246 12538
rect 6246 12486 6276 12538
rect 6300 12486 6310 12538
rect 6310 12486 6356 12538
rect 6380 12486 6426 12538
rect 6426 12486 6436 12538
rect 6460 12486 6490 12538
rect 6490 12486 6516 12538
rect 6220 12484 6276 12486
rect 6300 12484 6356 12486
rect 6380 12484 6436 12486
rect 6460 12484 6516 12486
rect 6220 11450 6276 11452
rect 6300 11450 6356 11452
rect 6380 11450 6436 11452
rect 6460 11450 6516 11452
rect 6220 11398 6246 11450
rect 6246 11398 6276 11450
rect 6300 11398 6310 11450
rect 6310 11398 6356 11450
rect 6380 11398 6426 11450
rect 6426 11398 6436 11450
rect 6460 11398 6490 11450
rect 6490 11398 6516 11450
rect 6220 11396 6276 11398
rect 6300 11396 6356 11398
rect 6380 11396 6436 11398
rect 6460 11396 6516 11398
rect 6642 12008 6698 12064
rect 6182 10684 6184 10704
rect 6184 10684 6236 10704
rect 6236 10684 6238 10704
rect 6182 10648 6238 10684
rect 6220 10362 6276 10364
rect 6300 10362 6356 10364
rect 6380 10362 6436 10364
rect 6460 10362 6516 10364
rect 6220 10310 6246 10362
rect 6246 10310 6276 10362
rect 6300 10310 6310 10362
rect 6310 10310 6356 10362
rect 6380 10310 6426 10362
rect 6426 10310 6436 10362
rect 6460 10310 6490 10362
rect 6490 10310 6516 10362
rect 6220 10308 6276 10310
rect 6300 10308 6356 10310
rect 6380 10308 6436 10310
rect 6460 10308 6516 10310
rect 6274 9560 6330 9616
rect 6550 9696 6606 9752
rect 6220 9274 6276 9276
rect 6300 9274 6356 9276
rect 6380 9274 6436 9276
rect 6460 9274 6516 9276
rect 6220 9222 6246 9274
rect 6246 9222 6276 9274
rect 6300 9222 6310 9274
rect 6310 9222 6356 9274
rect 6380 9222 6426 9274
rect 6426 9222 6436 9274
rect 6460 9222 6490 9274
rect 6490 9222 6516 9274
rect 6220 9220 6276 9222
rect 6300 9220 6356 9222
rect 6380 9220 6436 9222
rect 6460 9220 6516 9222
rect 6220 8186 6276 8188
rect 6300 8186 6356 8188
rect 6380 8186 6436 8188
rect 6460 8186 6516 8188
rect 6220 8134 6246 8186
rect 6246 8134 6276 8186
rect 6300 8134 6310 8186
rect 6310 8134 6356 8186
rect 6380 8134 6426 8186
rect 6426 8134 6436 8186
rect 6460 8134 6490 8186
rect 6490 8134 6516 8186
rect 6220 8132 6276 8134
rect 6300 8132 6356 8134
rect 6380 8132 6436 8134
rect 6460 8132 6516 8134
rect 6918 11328 6974 11384
rect 6826 10104 6882 10160
rect 6220 7098 6276 7100
rect 6300 7098 6356 7100
rect 6380 7098 6436 7100
rect 6460 7098 6516 7100
rect 6220 7046 6246 7098
rect 6246 7046 6276 7098
rect 6300 7046 6310 7098
rect 6310 7046 6356 7098
rect 6380 7046 6426 7098
rect 6426 7046 6436 7098
rect 6460 7046 6490 7098
rect 6490 7046 6516 7098
rect 6220 7044 6276 7046
rect 6300 7044 6356 7046
rect 6380 7044 6436 7046
rect 6460 7044 6516 7046
rect 6220 6010 6276 6012
rect 6300 6010 6356 6012
rect 6380 6010 6436 6012
rect 6460 6010 6516 6012
rect 6220 5958 6246 6010
rect 6246 5958 6276 6010
rect 6300 5958 6310 6010
rect 6310 5958 6356 6010
rect 6380 5958 6426 6010
rect 6426 5958 6436 6010
rect 6460 5958 6490 6010
rect 6490 5958 6516 6010
rect 6220 5956 6276 5958
rect 6300 5956 6356 5958
rect 6380 5956 6436 5958
rect 6460 5956 6516 5958
rect 6274 5072 6330 5128
rect 6220 4922 6276 4924
rect 6300 4922 6356 4924
rect 6380 4922 6436 4924
rect 6460 4922 6516 4924
rect 6220 4870 6246 4922
rect 6246 4870 6276 4922
rect 6300 4870 6310 4922
rect 6310 4870 6356 4922
rect 6380 4870 6426 4922
rect 6426 4870 6436 4922
rect 6460 4870 6490 4922
rect 6490 4870 6516 4922
rect 6220 4868 6276 4870
rect 6300 4868 6356 4870
rect 6380 4868 6436 4870
rect 6460 4868 6516 4870
rect 6220 3834 6276 3836
rect 6300 3834 6356 3836
rect 6380 3834 6436 3836
rect 6460 3834 6516 3836
rect 6220 3782 6246 3834
rect 6246 3782 6276 3834
rect 6300 3782 6310 3834
rect 6310 3782 6356 3834
rect 6380 3782 6426 3834
rect 6426 3782 6436 3834
rect 6460 3782 6490 3834
rect 6490 3782 6516 3834
rect 6220 3780 6276 3782
rect 6300 3780 6356 3782
rect 6380 3780 6436 3782
rect 6460 3780 6516 3782
rect 5998 3168 6054 3224
rect 6220 2746 6276 2748
rect 6300 2746 6356 2748
rect 6380 2746 6436 2748
rect 6460 2746 6516 2748
rect 6220 2694 6246 2746
rect 6246 2694 6276 2746
rect 6300 2694 6310 2746
rect 6310 2694 6356 2746
rect 6380 2694 6426 2746
rect 6426 2694 6436 2746
rect 6460 2694 6490 2746
rect 6490 2694 6516 2746
rect 6220 2692 6276 2694
rect 6300 2692 6356 2694
rect 6380 2692 6436 2694
rect 6460 2692 6516 2694
rect 6826 6024 6882 6080
rect 6734 5752 6790 5808
rect 6826 5616 6882 5672
rect 7010 9696 7066 9752
rect 6826 2896 6882 2952
rect 6918 2488 6974 2544
rect 7286 6704 7342 6760
rect 3238 1400 3294 1456
rect 3422 584 3478 640
rect 15014 16632 15070 16688
rect 7930 12044 7932 12064
rect 7932 12044 7984 12064
rect 7984 12044 7986 12064
rect 7930 12008 7986 12044
rect 7746 11348 7802 11384
rect 7746 11328 7748 11348
rect 7748 11328 7800 11348
rect 7800 11328 7802 11348
rect 7930 10920 7986 10976
rect 8022 8880 8078 8936
rect 7838 8200 7894 8256
rect 7562 6024 7618 6080
rect 8298 11056 8354 11112
rect 8206 10548 8208 10568
rect 8208 10548 8260 10568
rect 8260 10548 8262 10568
rect 8206 10512 8262 10548
rect 8206 9152 8262 9208
rect 8390 9868 8392 9888
rect 8392 9868 8444 9888
rect 8444 9868 8446 9888
rect 8390 9832 8446 9868
rect 8206 8336 8262 8392
rect 8298 7384 8354 7440
rect 8114 6840 8170 6896
rect 8298 6160 8354 6216
rect 8206 6060 8208 6080
rect 8208 6060 8260 6080
rect 8260 6060 8262 6080
rect 8206 6024 8262 6060
rect 7930 5344 7986 5400
rect 7838 3984 7894 4040
rect 8114 5208 8170 5264
rect 8114 4120 8170 4176
rect 8852 14170 8908 14172
rect 8932 14170 8988 14172
rect 9012 14170 9068 14172
rect 9092 14170 9148 14172
rect 8852 14118 8878 14170
rect 8878 14118 8908 14170
rect 8932 14118 8942 14170
rect 8942 14118 8988 14170
rect 9012 14118 9058 14170
rect 9058 14118 9068 14170
rect 9092 14118 9122 14170
rect 9122 14118 9148 14170
rect 8852 14116 8908 14118
rect 8932 14116 8988 14118
rect 9012 14116 9068 14118
rect 9092 14116 9148 14118
rect 8852 13082 8908 13084
rect 8932 13082 8988 13084
rect 9012 13082 9068 13084
rect 9092 13082 9148 13084
rect 8852 13030 8878 13082
rect 8878 13030 8908 13082
rect 8932 13030 8942 13082
rect 8942 13030 8988 13082
rect 9012 13030 9058 13082
rect 9058 13030 9068 13082
rect 9092 13030 9122 13082
rect 9122 13030 9148 13082
rect 8852 13028 8908 13030
rect 8932 13028 8988 13030
rect 9012 13028 9068 13030
rect 9092 13028 9148 13030
rect 9034 12300 9090 12336
rect 9034 12280 9036 12300
rect 9036 12280 9088 12300
rect 9088 12280 9090 12300
rect 9402 12144 9458 12200
rect 8852 11994 8908 11996
rect 8932 11994 8988 11996
rect 9012 11994 9068 11996
rect 9092 11994 9148 11996
rect 8852 11942 8878 11994
rect 8878 11942 8908 11994
rect 8932 11942 8942 11994
rect 8942 11942 8988 11994
rect 9012 11942 9058 11994
rect 9058 11942 9068 11994
rect 9092 11942 9122 11994
rect 9122 11942 9148 11994
rect 8852 11940 8908 11942
rect 8932 11940 8988 11942
rect 9012 11940 9068 11942
rect 9092 11940 9148 11942
rect 8852 10906 8908 10908
rect 8932 10906 8988 10908
rect 9012 10906 9068 10908
rect 9092 10906 9148 10908
rect 8852 10854 8878 10906
rect 8878 10854 8908 10906
rect 8932 10854 8942 10906
rect 8942 10854 8988 10906
rect 9012 10854 9058 10906
rect 9058 10854 9068 10906
rect 9092 10854 9122 10906
rect 9122 10854 9148 10906
rect 8852 10852 8908 10854
rect 8932 10852 8988 10854
rect 9012 10852 9068 10854
rect 9092 10852 9148 10854
rect 9218 10104 9274 10160
rect 8852 9818 8908 9820
rect 8932 9818 8988 9820
rect 9012 9818 9068 9820
rect 9092 9818 9148 9820
rect 8852 9766 8878 9818
rect 8878 9766 8908 9818
rect 8932 9766 8942 9818
rect 8942 9766 8988 9818
rect 9012 9766 9058 9818
rect 9058 9766 9068 9818
rect 9092 9766 9122 9818
rect 9122 9766 9148 9818
rect 8852 9764 8908 9766
rect 8932 9764 8988 9766
rect 9012 9764 9068 9766
rect 9092 9764 9148 9766
rect 8574 9016 8630 9072
rect 9126 9016 9182 9072
rect 8758 8880 8814 8936
rect 8852 8730 8908 8732
rect 8932 8730 8988 8732
rect 9012 8730 9068 8732
rect 9092 8730 9148 8732
rect 8852 8678 8878 8730
rect 8878 8678 8908 8730
rect 8932 8678 8942 8730
rect 8942 8678 8988 8730
rect 9012 8678 9058 8730
rect 9058 8678 9068 8730
rect 9092 8678 9122 8730
rect 9122 8678 9148 8730
rect 8852 8676 8908 8678
rect 8932 8676 8988 8678
rect 9012 8676 9068 8678
rect 9092 8676 9148 8678
rect 8482 8064 8538 8120
rect 8482 7112 8538 7168
rect 8298 3984 8354 4040
rect 7470 2644 7526 2680
rect 7470 2624 7472 2644
rect 7472 2624 7524 2644
rect 7524 2624 7526 2644
rect 8298 2896 8354 2952
rect 8852 7642 8908 7644
rect 8932 7642 8988 7644
rect 9012 7642 9068 7644
rect 9092 7642 9148 7644
rect 8852 7590 8878 7642
rect 8878 7590 8908 7642
rect 8932 7590 8942 7642
rect 8942 7590 8988 7642
rect 9012 7590 9058 7642
rect 9058 7590 9068 7642
rect 9092 7590 9122 7642
rect 9122 7590 9148 7642
rect 8852 7588 8908 7590
rect 8932 7588 8988 7590
rect 9012 7588 9068 7590
rect 9092 7588 9148 7590
rect 8758 6976 8814 7032
rect 9586 11600 9642 11656
rect 9862 10240 9918 10296
rect 9862 9968 9918 10024
rect 9494 8744 9550 8800
rect 9402 8472 9458 8528
rect 9770 9424 9826 9480
rect 10506 13776 10562 13832
rect 10046 9560 10102 9616
rect 9954 8744 10010 8800
rect 10046 8608 10102 8664
rect 9862 8356 9918 8392
rect 9862 8336 9864 8356
rect 9864 8336 9916 8356
rect 9916 8336 9918 8356
rect 10046 8336 10102 8392
rect 9494 8200 9550 8256
rect 9678 8200 9734 8256
rect 8850 6740 8852 6760
rect 8852 6740 8904 6760
rect 8904 6740 8906 6760
rect 8850 6704 8906 6740
rect 9126 6724 9182 6760
rect 9126 6704 9128 6724
rect 9128 6704 9180 6724
rect 9180 6704 9182 6724
rect 8852 6554 8908 6556
rect 8932 6554 8988 6556
rect 9012 6554 9068 6556
rect 9092 6554 9148 6556
rect 8852 6502 8878 6554
rect 8878 6502 8908 6554
rect 8932 6502 8942 6554
rect 8942 6502 8988 6554
rect 9012 6502 9058 6554
rect 9058 6502 9068 6554
rect 9092 6502 9122 6554
rect 9122 6502 9148 6554
rect 8852 6500 8908 6502
rect 8932 6500 8988 6502
rect 9012 6500 9068 6502
rect 9092 6500 9148 6502
rect 9126 6160 9182 6216
rect 8942 5888 8998 5944
rect 8852 5466 8908 5468
rect 8932 5466 8988 5468
rect 9012 5466 9068 5468
rect 9092 5466 9148 5468
rect 8852 5414 8878 5466
rect 8878 5414 8908 5466
rect 8932 5414 8942 5466
rect 8942 5414 8988 5466
rect 9012 5414 9058 5466
rect 9058 5414 9068 5466
rect 9092 5414 9122 5466
rect 9122 5414 9148 5466
rect 8852 5412 8908 5414
rect 8932 5412 8988 5414
rect 9012 5412 9068 5414
rect 9092 5412 9148 5414
rect 8852 4378 8908 4380
rect 8932 4378 8988 4380
rect 9012 4378 9068 4380
rect 9092 4378 9148 4380
rect 8852 4326 8878 4378
rect 8878 4326 8908 4378
rect 8932 4326 8942 4378
rect 8942 4326 8988 4378
rect 9012 4326 9058 4378
rect 9058 4326 9068 4378
rect 9092 4326 9122 4378
rect 9122 4326 9148 4378
rect 8852 4324 8908 4326
rect 8932 4324 8988 4326
rect 9012 4324 9068 4326
rect 9092 4324 9148 4326
rect 8942 4140 8998 4176
rect 8942 4120 8944 4140
rect 8944 4120 8996 4140
rect 8996 4120 8998 4140
rect 8942 3984 8998 4040
rect 8850 3884 8852 3904
rect 8852 3884 8904 3904
rect 8904 3884 8906 3904
rect 8850 3848 8906 3884
rect 8850 3732 8906 3768
rect 8850 3712 8852 3732
rect 8852 3712 8904 3732
rect 8904 3712 8906 3732
rect 8758 3576 8814 3632
rect 9126 3440 9182 3496
rect 9494 7284 9496 7304
rect 9496 7284 9548 7304
rect 9548 7284 9550 7304
rect 9494 7248 9550 7284
rect 9402 5072 9458 5128
rect 8852 3290 8908 3292
rect 8932 3290 8988 3292
rect 9012 3290 9068 3292
rect 9092 3290 9148 3292
rect 8852 3238 8878 3290
rect 8878 3238 8908 3290
rect 8932 3238 8942 3290
rect 8942 3238 8988 3290
rect 9012 3238 9058 3290
rect 9058 3238 9068 3290
rect 9092 3238 9122 3290
rect 9122 3238 9148 3290
rect 8852 3236 8908 3238
rect 8932 3236 8988 3238
rect 9012 3236 9068 3238
rect 9092 3236 9148 3238
rect 9310 3032 9366 3088
rect 9678 5752 9734 5808
rect 9954 6704 10010 6760
rect 9862 5208 9918 5264
rect 9770 3576 9826 3632
rect 10138 5908 10194 5944
rect 10138 5888 10140 5908
rect 10140 5888 10192 5908
rect 10192 5888 10194 5908
rect 10046 5752 10102 5808
rect 9954 4120 10010 4176
rect 8852 2202 8908 2204
rect 8932 2202 8988 2204
rect 9012 2202 9068 2204
rect 9092 2202 9148 2204
rect 8852 2150 8878 2202
rect 8878 2150 8908 2202
rect 8932 2150 8942 2202
rect 8942 2150 8988 2202
rect 9012 2150 9058 2202
rect 9058 2150 9068 2202
rect 9092 2150 9122 2202
rect 9122 2150 9148 2202
rect 8852 2148 8908 2150
rect 8932 2148 8988 2150
rect 9012 2148 9068 2150
rect 9092 2148 9148 2150
rect 10322 5480 10378 5536
rect 10598 11736 10654 11792
rect 10690 10784 10746 10840
rect 13358 15816 13414 15872
rect 11484 14714 11540 14716
rect 11564 14714 11620 14716
rect 11644 14714 11700 14716
rect 11724 14714 11780 14716
rect 11484 14662 11510 14714
rect 11510 14662 11540 14714
rect 11564 14662 11574 14714
rect 11574 14662 11620 14714
rect 11644 14662 11690 14714
rect 11690 14662 11700 14714
rect 11724 14662 11754 14714
rect 11754 14662 11780 14714
rect 11484 14660 11540 14662
rect 11564 14660 11620 14662
rect 11644 14660 11700 14662
rect 11724 14660 11780 14662
rect 11484 13626 11540 13628
rect 11564 13626 11620 13628
rect 11644 13626 11700 13628
rect 11724 13626 11780 13628
rect 11484 13574 11510 13626
rect 11510 13574 11540 13626
rect 11564 13574 11574 13626
rect 11574 13574 11620 13626
rect 11644 13574 11690 13626
rect 11690 13574 11700 13626
rect 11724 13574 11754 13626
rect 11754 13574 11780 13626
rect 11484 13572 11540 13574
rect 11564 13572 11620 13574
rect 11644 13572 11700 13574
rect 11724 13572 11780 13574
rect 12070 13776 12126 13832
rect 11484 12538 11540 12540
rect 11564 12538 11620 12540
rect 11644 12538 11700 12540
rect 11724 12538 11780 12540
rect 11484 12486 11510 12538
rect 11510 12486 11540 12538
rect 11564 12486 11574 12538
rect 11574 12486 11620 12538
rect 11644 12486 11690 12538
rect 11690 12486 11700 12538
rect 11724 12486 11754 12538
rect 11754 12486 11780 12538
rect 11484 12484 11540 12486
rect 11564 12484 11620 12486
rect 11644 12484 11700 12486
rect 11724 12484 11780 12486
rect 10966 11600 11022 11656
rect 10782 10240 10838 10296
rect 10874 9696 10930 9752
rect 10690 9424 10746 9480
rect 10414 5344 10470 5400
rect 10414 5208 10470 5264
rect 10782 9324 10784 9344
rect 10784 9324 10836 9344
rect 10836 9324 10838 9344
rect 10782 9288 10838 9324
rect 10782 8064 10838 8120
rect 10690 7112 10746 7168
rect 11484 11450 11540 11452
rect 11564 11450 11620 11452
rect 11644 11450 11700 11452
rect 11724 11450 11780 11452
rect 11484 11398 11510 11450
rect 11510 11398 11540 11450
rect 11564 11398 11574 11450
rect 11574 11398 11620 11450
rect 11644 11398 11690 11450
rect 11690 11398 11700 11450
rect 11724 11398 11754 11450
rect 11754 11398 11780 11450
rect 11484 11396 11540 11398
rect 11564 11396 11620 11398
rect 11644 11396 11700 11398
rect 11724 11396 11780 11398
rect 11978 10784 12034 10840
rect 11794 10648 11850 10704
rect 11978 10684 11980 10704
rect 11980 10684 12032 10704
rect 12032 10684 12034 10704
rect 11484 10362 11540 10364
rect 11564 10362 11620 10364
rect 11644 10362 11700 10364
rect 11724 10362 11780 10364
rect 11484 10310 11510 10362
rect 11510 10310 11540 10362
rect 11564 10310 11574 10362
rect 11574 10310 11620 10362
rect 11644 10310 11690 10362
rect 11690 10310 11700 10362
rect 11724 10310 11754 10362
rect 11754 10310 11780 10362
rect 11484 10308 11540 10310
rect 11564 10308 11620 10310
rect 11644 10308 11700 10310
rect 11724 10308 11780 10310
rect 11978 10648 12034 10684
rect 11484 9274 11540 9276
rect 11564 9274 11620 9276
rect 11644 9274 11700 9276
rect 11724 9274 11780 9276
rect 11484 9222 11510 9274
rect 11510 9222 11540 9274
rect 11564 9222 11574 9274
rect 11574 9222 11620 9274
rect 11644 9222 11690 9274
rect 11690 9222 11700 9274
rect 11724 9222 11754 9274
rect 11754 9222 11780 9274
rect 11484 9220 11540 9222
rect 11564 9220 11620 9222
rect 11644 9220 11700 9222
rect 11724 9220 11780 9222
rect 11334 8744 11390 8800
rect 11242 8336 11298 8392
rect 11484 8186 11540 8188
rect 11564 8186 11620 8188
rect 11644 8186 11700 8188
rect 11724 8186 11780 8188
rect 11484 8134 11510 8186
rect 11510 8134 11540 8186
rect 11564 8134 11574 8186
rect 11574 8134 11620 8186
rect 11644 8134 11690 8186
rect 11690 8134 11700 8186
rect 11724 8134 11754 8186
rect 11754 8134 11780 8186
rect 11484 8132 11540 8134
rect 11564 8132 11620 8134
rect 11644 8132 11700 8134
rect 11724 8132 11780 8134
rect 11058 7268 11114 7304
rect 11058 7248 11060 7268
rect 11060 7248 11112 7268
rect 11112 7248 11114 7268
rect 11242 6976 11298 7032
rect 10782 5208 10838 5264
rect 11702 7792 11758 7848
rect 11886 8744 11942 8800
rect 11484 7098 11540 7100
rect 11564 7098 11620 7100
rect 11644 7098 11700 7100
rect 11724 7098 11780 7100
rect 11484 7046 11510 7098
rect 11510 7046 11540 7098
rect 11564 7046 11574 7098
rect 11574 7046 11620 7098
rect 11644 7046 11690 7098
rect 11690 7046 11700 7098
rect 11724 7046 11754 7098
rect 11754 7046 11780 7098
rect 11484 7044 11540 7046
rect 11564 7044 11620 7046
rect 11644 7044 11700 7046
rect 11724 7044 11780 7046
rect 14094 15408 14150 15464
rect 13910 15000 13966 15056
rect 12254 11620 12310 11656
rect 12254 11600 12256 11620
rect 12256 11600 12308 11620
rect 12308 11600 12310 11620
rect 12254 11056 12310 11112
rect 12806 12960 12862 13016
rect 12530 11736 12586 11792
rect 12622 11328 12678 11384
rect 12530 10784 12586 10840
rect 12438 10376 12494 10432
rect 12898 12552 12954 12608
rect 12806 12280 12862 12336
rect 12622 10512 12678 10568
rect 12438 9832 12494 9888
rect 12346 9288 12402 9344
rect 12254 9152 12310 9208
rect 12070 8472 12126 8528
rect 11794 6704 11850 6760
rect 11484 6010 11540 6012
rect 11564 6010 11620 6012
rect 11644 6010 11700 6012
rect 11724 6010 11780 6012
rect 11484 5958 11510 6010
rect 11510 5958 11540 6010
rect 11564 5958 11574 6010
rect 11574 5958 11620 6010
rect 11644 5958 11690 6010
rect 11690 5958 11700 6010
rect 11724 5958 11754 6010
rect 11754 5958 11780 6010
rect 11484 5956 11540 5958
rect 11564 5956 11620 5958
rect 11644 5956 11700 5958
rect 11724 5956 11780 5958
rect 11150 5480 11206 5536
rect 10414 3848 10470 3904
rect 10322 2896 10378 2952
rect 10690 3596 10746 3632
rect 10690 3576 10692 3596
rect 10692 3576 10744 3596
rect 10744 3576 10746 3596
rect 10782 3440 10838 3496
rect 11058 3576 11114 3632
rect 10598 3068 10600 3088
rect 10600 3068 10652 3088
rect 10652 3068 10654 3088
rect 10598 3032 10654 3068
rect 10598 2932 10600 2952
rect 10600 2932 10652 2952
rect 10652 2932 10654 2952
rect 10598 2896 10654 2932
rect 10322 2488 10378 2544
rect 11484 4922 11540 4924
rect 11564 4922 11620 4924
rect 11644 4922 11700 4924
rect 11724 4922 11780 4924
rect 11484 4870 11510 4922
rect 11510 4870 11540 4922
rect 11564 4870 11574 4922
rect 11574 4870 11620 4922
rect 11644 4870 11690 4922
rect 11690 4870 11700 4922
rect 11724 4870 11754 4922
rect 11754 4870 11780 4922
rect 11484 4868 11540 4870
rect 11564 4868 11620 4870
rect 11644 4868 11700 4870
rect 11724 4868 11780 4870
rect 11794 4120 11850 4176
rect 11484 3834 11540 3836
rect 11564 3834 11620 3836
rect 11644 3834 11700 3836
rect 11724 3834 11780 3836
rect 11484 3782 11510 3834
rect 11510 3782 11540 3834
rect 11564 3782 11574 3834
rect 11574 3782 11620 3834
rect 11644 3782 11690 3834
rect 11690 3782 11700 3834
rect 11724 3782 11754 3834
rect 11754 3782 11780 3834
rect 11484 3780 11540 3782
rect 11564 3780 11620 3782
rect 11644 3780 11700 3782
rect 11724 3780 11780 3782
rect 11794 3440 11850 3496
rect 11518 3032 11574 3088
rect 11334 2896 11390 2952
rect 12162 5752 12218 5808
rect 11978 5652 11980 5672
rect 11980 5652 12032 5672
rect 12032 5652 12034 5672
rect 11978 5616 12034 5652
rect 11978 4820 12034 4856
rect 11978 4800 11980 4820
rect 11980 4800 12032 4820
rect 12032 4800 12034 4820
rect 12530 9696 12586 9752
rect 12714 8880 12770 8936
rect 12898 11328 12954 11384
rect 12898 10648 12954 10704
rect 12898 10240 12954 10296
rect 12898 9968 12954 10024
rect 13082 10920 13138 10976
rect 13818 13232 13874 13288
rect 13266 11056 13322 11112
rect 13266 10920 13322 10976
rect 13542 10784 13598 10840
rect 13634 10648 13690 10704
rect 13174 9696 13230 9752
rect 12990 9288 13046 9344
rect 13082 9152 13138 9208
rect 12346 7656 12402 7712
rect 12346 5616 12402 5672
rect 12346 4684 12402 4720
rect 12346 4664 12348 4684
rect 12348 4664 12400 4684
rect 12400 4664 12402 4684
rect 11058 2644 11114 2680
rect 11978 2896 12034 2952
rect 11484 2746 11540 2748
rect 11564 2746 11620 2748
rect 11644 2746 11700 2748
rect 11724 2746 11780 2748
rect 11484 2694 11510 2746
rect 11510 2694 11540 2746
rect 11564 2694 11574 2746
rect 11574 2694 11620 2746
rect 11644 2694 11690 2746
rect 11690 2694 11700 2746
rect 11724 2694 11754 2746
rect 11754 2694 11780 2746
rect 11484 2692 11540 2694
rect 11564 2692 11620 2694
rect 11644 2692 11700 2694
rect 11724 2692 11780 2694
rect 11058 2624 11060 2644
rect 11060 2624 11112 2644
rect 11112 2624 11114 2644
rect 11794 2508 11850 2544
rect 12438 3304 12494 3360
rect 12898 7656 12954 7712
rect 13358 9424 13414 9480
rect 13542 8880 13598 8936
rect 13542 8744 13598 8800
rect 13450 7792 13506 7848
rect 12990 6160 13046 6216
rect 12714 4528 12770 4584
rect 12714 3576 12770 3632
rect 11794 2488 11796 2508
rect 11796 2488 11848 2508
rect 11848 2488 11850 2508
rect 14830 14184 14886 14240
rect 14116 14170 14172 14172
rect 14196 14170 14252 14172
rect 14276 14170 14332 14172
rect 14356 14170 14412 14172
rect 14116 14118 14142 14170
rect 14142 14118 14172 14170
rect 14196 14118 14206 14170
rect 14206 14118 14252 14170
rect 14276 14118 14322 14170
rect 14322 14118 14332 14170
rect 14356 14118 14386 14170
rect 14386 14118 14412 14170
rect 14116 14116 14172 14118
rect 14196 14116 14252 14118
rect 14276 14116 14332 14118
rect 14356 14116 14412 14118
rect 14116 13082 14172 13084
rect 14196 13082 14252 13084
rect 14276 13082 14332 13084
rect 14356 13082 14412 13084
rect 14116 13030 14142 13082
rect 14142 13030 14172 13082
rect 14196 13030 14206 13082
rect 14206 13030 14252 13082
rect 14276 13030 14322 13082
rect 14322 13030 14332 13082
rect 14356 13030 14386 13082
rect 14386 13030 14412 13082
rect 14116 13028 14172 13030
rect 14196 13028 14252 13030
rect 14276 13028 14332 13030
rect 14356 13028 14412 13030
rect 13910 12280 13966 12336
rect 14462 12144 14518 12200
rect 13910 11872 13966 11928
rect 14116 11994 14172 11996
rect 14196 11994 14252 11996
rect 14276 11994 14332 11996
rect 14356 11994 14412 11996
rect 14116 11942 14142 11994
rect 14142 11942 14172 11994
rect 14196 11942 14206 11994
rect 14206 11942 14252 11994
rect 14276 11942 14322 11994
rect 14322 11942 14332 11994
rect 14356 11942 14386 11994
rect 14386 11942 14412 11994
rect 14116 11940 14172 11942
rect 14196 11940 14252 11942
rect 14276 11940 14332 11942
rect 14356 11940 14412 11942
rect 14370 11092 14372 11112
rect 14372 11092 14424 11112
rect 14424 11092 14426 11112
rect 14370 11056 14426 11092
rect 13910 10376 13966 10432
rect 14116 10906 14172 10908
rect 14196 10906 14252 10908
rect 14276 10906 14332 10908
rect 14356 10906 14412 10908
rect 14116 10854 14142 10906
rect 14142 10854 14172 10906
rect 14196 10854 14206 10906
rect 14206 10854 14252 10906
rect 14276 10854 14322 10906
rect 14322 10854 14332 10906
rect 14356 10854 14386 10906
rect 14386 10854 14412 10906
rect 14116 10852 14172 10854
rect 14196 10852 14252 10854
rect 14276 10852 14332 10854
rect 14356 10852 14412 10854
rect 14738 12552 14794 12608
rect 14646 10920 14702 10976
rect 15106 15272 15162 15328
rect 15106 14592 15162 14648
rect 14922 12008 14978 12064
rect 14830 10240 14886 10296
rect 16210 16224 16266 16280
rect 16210 15272 16266 15328
rect 15566 11736 15622 11792
rect 15106 11056 15162 11112
rect 15382 10920 15438 10976
rect 15290 10784 15346 10840
rect 14116 9818 14172 9820
rect 14196 9818 14252 9820
rect 14276 9818 14332 9820
rect 14356 9818 14412 9820
rect 14116 9766 14142 9818
rect 14142 9766 14172 9818
rect 14196 9766 14206 9818
rect 14206 9766 14252 9818
rect 14276 9766 14322 9818
rect 14322 9766 14332 9818
rect 14356 9766 14386 9818
rect 14386 9766 14412 9818
rect 14116 9764 14172 9766
rect 14196 9764 14252 9766
rect 14276 9764 14332 9766
rect 14356 9764 14412 9766
rect 14554 9560 14610 9616
rect 13818 8608 13874 8664
rect 13634 8472 13690 8528
rect 14002 9052 14004 9072
rect 14004 9052 14056 9072
rect 14056 9052 14058 9072
rect 14002 9016 14058 9052
rect 14116 8730 14172 8732
rect 14196 8730 14252 8732
rect 14276 8730 14332 8732
rect 14356 8730 14412 8732
rect 14116 8678 14142 8730
rect 14142 8678 14172 8730
rect 14196 8678 14206 8730
rect 14206 8678 14252 8730
rect 14276 8678 14322 8730
rect 14322 8678 14332 8730
rect 14356 8678 14386 8730
rect 14386 8678 14412 8730
rect 14116 8676 14172 8678
rect 14196 8676 14252 8678
rect 14276 8676 14332 8678
rect 14356 8676 14412 8678
rect 14462 8472 14518 8528
rect 13634 8064 13690 8120
rect 13910 8200 13966 8256
rect 13818 7948 13874 7984
rect 13818 7928 13820 7948
rect 13820 7928 13872 7948
rect 13872 7928 13874 7948
rect 13634 7520 13690 7576
rect 13542 3984 13598 4040
rect 14116 7642 14172 7644
rect 14196 7642 14252 7644
rect 14276 7642 14332 7644
rect 14356 7642 14412 7644
rect 14116 7590 14142 7642
rect 14142 7590 14172 7642
rect 14196 7590 14206 7642
rect 14206 7590 14252 7642
rect 14276 7590 14322 7642
rect 14322 7590 14332 7642
rect 14356 7590 14386 7642
rect 14386 7590 14412 7642
rect 14116 7588 14172 7590
rect 14196 7588 14252 7590
rect 14276 7588 14332 7590
rect 14356 7588 14412 7590
rect 13634 3032 13690 3088
rect 14462 7248 14518 7304
rect 14116 6554 14172 6556
rect 14196 6554 14252 6556
rect 14276 6554 14332 6556
rect 14356 6554 14412 6556
rect 14116 6502 14142 6554
rect 14142 6502 14172 6554
rect 14196 6502 14206 6554
rect 14206 6502 14252 6554
rect 14276 6502 14322 6554
rect 14322 6502 14332 6554
rect 14356 6502 14386 6554
rect 14386 6502 14412 6554
rect 14116 6500 14172 6502
rect 14196 6500 14252 6502
rect 14276 6500 14332 6502
rect 14356 6500 14412 6502
rect 14116 5466 14172 5468
rect 14196 5466 14252 5468
rect 14276 5466 14332 5468
rect 14356 5466 14412 5468
rect 14116 5414 14142 5466
rect 14142 5414 14172 5466
rect 14196 5414 14206 5466
rect 14206 5414 14252 5466
rect 14276 5414 14322 5466
rect 14322 5414 14332 5466
rect 14356 5414 14386 5466
rect 14386 5414 14412 5466
rect 14116 5412 14172 5414
rect 14196 5412 14252 5414
rect 14276 5412 14332 5414
rect 14356 5412 14412 5414
rect 14094 4664 14150 4720
rect 14116 4378 14172 4380
rect 14196 4378 14252 4380
rect 14276 4378 14332 4380
rect 14356 4378 14412 4380
rect 14116 4326 14142 4378
rect 14142 4326 14172 4378
rect 14196 4326 14206 4378
rect 14206 4326 14252 4378
rect 14276 4326 14322 4378
rect 14322 4326 14332 4378
rect 14356 4326 14386 4378
rect 14386 4326 14412 4378
rect 14116 4324 14172 4326
rect 14196 4324 14252 4326
rect 14276 4324 14332 4326
rect 14356 4324 14412 4326
rect 14116 3290 14172 3292
rect 14196 3290 14252 3292
rect 14276 3290 14332 3292
rect 14356 3290 14412 3292
rect 14116 3238 14142 3290
rect 14142 3238 14172 3290
rect 14196 3238 14206 3290
rect 14206 3238 14252 3290
rect 14276 3238 14322 3290
rect 14322 3238 14332 3290
rect 14356 3238 14386 3290
rect 14386 3238 14412 3290
rect 14116 3236 14172 3238
rect 14196 3236 14252 3238
rect 14276 3236 14332 3238
rect 14356 3236 14412 3238
rect 14646 8336 14702 8392
rect 14646 7384 14702 7440
rect 14922 8472 14978 8528
rect 15290 10104 15346 10160
rect 14830 6976 14886 7032
rect 14922 6704 14978 6760
rect 10966 992 11022 1048
rect 14002 2352 14058 2408
rect 14116 2202 14172 2204
rect 14196 2202 14252 2204
rect 14276 2202 14332 2204
rect 14356 2202 14412 2204
rect 14116 2150 14142 2202
rect 14142 2150 14172 2202
rect 14196 2150 14206 2202
rect 14206 2150 14252 2202
rect 14276 2150 14322 2202
rect 14322 2150 14332 2202
rect 14356 2150 14386 2202
rect 14386 2150 14412 2202
rect 14116 2148 14172 2150
rect 14196 2148 14252 2150
rect 14276 2148 14332 2150
rect 14356 2148 14412 2150
rect 14738 1808 14794 1864
rect 14922 6024 14978 6080
rect 15106 8064 15162 8120
rect 15290 7792 15346 7848
rect 15014 4392 15070 4448
rect 14830 1400 14886 1456
rect 15106 3576 15162 3632
rect 15014 584 15070 640
rect 3054 176 3110 232
rect 15474 9424 15530 9480
rect 15750 11192 15806 11248
rect 15658 9288 15714 9344
rect 15658 6432 15714 6488
rect 15750 6296 15806 6352
rect 15750 6160 15806 6216
rect 15750 4564 15752 4584
rect 15752 4564 15804 4584
rect 15804 4564 15806 4584
rect 15750 4528 15806 4564
rect 16302 12552 16358 12608
rect 16118 8608 16174 8664
rect 15842 4120 15898 4176
rect 16394 2624 16450 2680
rect 15106 176 15162 232
<< metal3 >>
rect 0 16690 480 16720
rect 7649 16690 7715 16693
rect 0 16688 7715 16690
rect 0 16632 7654 16688
rect 7710 16632 7715 16688
rect 0 16630 7715 16632
rect 0 16600 480 16630
rect 7649 16627 7715 16630
rect 15009 16690 15075 16693
rect 17520 16690 18000 16720
rect 15009 16688 18000 16690
rect 15009 16632 15014 16688
rect 15070 16632 18000 16688
rect 15009 16630 18000 16632
rect 15009 16627 15075 16630
rect 17520 16600 18000 16630
rect 0 16282 480 16312
rect 4061 16282 4127 16285
rect 0 16280 4127 16282
rect 0 16224 4066 16280
rect 4122 16224 4127 16280
rect 0 16222 4127 16224
rect 0 16192 480 16222
rect 4061 16219 4127 16222
rect 16205 16282 16271 16285
rect 17520 16282 18000 16312
rect 16205 16280 18000 16282
rect 16205 16224 16210 16280
rect 16266 16224 18000 16280
rect 16205 16222 18000 16224
rect 16205 16219 16271 16222
rect 17520 16192 18000 16222
rect 0 15874 480 15904
rect 2681 15874 2747 15877
rect 0 15872 2747 15874
rect 0 15816 2686 15872
rect 2742 15816 2747 15872
rect 0 15814 2747 15816
rect 0 15784 480 15814
rect 2681 15811 2747 15814
rect 13353 15874 13419 15877
rect 17520 15874 18000 15904
rect 13353 15872 18000 15874
rect 13353 15816 13358 15872
rect 13414 15816 18000 15872
rect 13353 15814 18000 15816
rect 13353 15811 13419 15814
rect 17520 15784 18000 15814
rect 0 15466 480 15496
rect 3969 15466 4035 15469
rect 0 15464 4035 15466
rect 0 15408 3974 15464
rect 4030 15408 4035 15464
rect 0 15406 4035 15408
rect 0 15376 480 15406
rect 3969 15403 4035 15406
rect 14089 15466 14155 15469
rect 17520 15466 18000 15496
rect 14089 15464 18000 15466
rect 14089 15408 14094 15464
rect 14150 15408 18000 15464
rect 14089 15406 18000 15408
rect 14089 15403 14155 15406
rect 17520 15376 18000 15406
rect 15101 15330 15167 15333
rect 16205 15330 16271 15333
rect 15101 15328 16271 15330
rect 15101 15272 15106 15328
rect 15162 15272 16210 15328
rect 16266 15272 16271 15328
rect 15101 15270 16271 15272
rect 15101 15267 15167 15270
rect 16205 15267 16271 15270
rect 0 15058 480 15088
rect 4061 15058 4127 15061
rect 0 15056 4127 15058
rect 0 15000 4066 15056
rect 4122 15000 4127 15056
rect 0 14998 4127 15000
rect 0 14968 480 14998
rect 4061 14995 4127 14998
rect 13905 15058 13971 15061
rect 17520 15058 18000 15088
rect 13905 15056 18000 15058
rect 13905 15000 13910 15056
rect 13966 15000 18000 15056
rect 13905 14998 18000 15000
rect 13905 14995 13971 14998
rect 17520 14968 18000 14998
rect 6208 14720 6528 14721
rect 0 14650 480 14680
rect 6208 14656 6216 14720
rect 6280 14656 6296 14720
rect 6360 14656 6376 14720
rect 6440 14656 6456 14720
rect 6520 14656 6528 14720
rect 6208 14655 6528 14656
rect 11472 14720 11792 14721
rect 11472 14656 11480 14720
rect 11544 14656 11560 14720
rect 11624 14656 11640 14720
rect 11704 14656 11720 14720
rect 11784 14656 11792 14720
rect 11472 14655 11792 14656
rect 4061 14650 4127 14653
rect 0 14648 4127 14650
rect 0 14592 4066 14648
rect 4122 14592 4127 14648
rect 0 14590 4127 14592
rect 0 14560 480 14590
rect 4061 14587 4127 14590
rect 15101 14650 15167 14653
rect 17520 14650 18000 14680
rect 15101 14648 18000 14650
rect 15101 14592 15106 14648
rect 15162 14592 18000 14648
rect 15101 14590 18000 14592
rect 15101 14587 15167 14590
rect 17520 14560 18000 14590
rect 0 14242 480 14272
rect 14825 14242 14891 14245
rect 17520 14242 18000 14272
rect 0 14182 3434 14242
rect 0 14152 480 14182
rect 3374 13970 3434 14182
rect 14825 14240 18000 14242
rect 14825 14184 14830 14240
rect 14886 14184 18000 14240
rect 14825 14182 18000 14184
rect 14825 14179 14891 14182
rect 3576 14176 3896 14177
rect 3576 14112 3584 14176
rect 3648 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3896 14176
rect 3576 14111 3896 14112
rect 8840 14176 9160 14177
rect 8840 14112 8848 14176
rect 8912 14112 8928 14176
rect 8992 14112 9008 14176
rect 9072 14112 9088 14176
rect 9152 14112 9160 14176
rect 8840 14111 9160 14112
rect 14104 14176 14424 14177
rect 14104 14112 14112 14176
rect 14176 14112 14192 14176
rect 14256 14112 14272 14176
rect 14336 14112 14352 14176
rect 14416 14112 14424 14176
rect 17520 14152 18000 14182
rect 14104 14111 14424 14112
rect 5441 13970 5507 13973
rect 3374 13968 5507 13970
rect 3374 13912 5446 13968
rect 5502 13912 5507 13968
rect 3374 13910 5507 13912
rect 5441 13907 5507 13910
rect 0 13834 480 13864
rect 3509 13834 3575 13837
rect 0 13832 3575 13834
rect 0 13776 3514 13832
rect 3570 13776 3575 13832
rect 0 13774 3575 13776
rect 0 13744 480 13774
rect 3509 13771 3575 13774
rect 10501 13834 10567 13837
rect 12065 13834 12131 13837
rect 17520 13834 18000 13864
rect 10501 13832 18000 13834
rect 10501 13776 10506 13832
rect 10562 13776 12070 13832
rect 12126 13776 18000 13832
rect 10501 13774 18000 13776
rect 10501 13771 10567 13774
rect 12065 13771 12131 13774
rect 17520 13744 18000 13774
rect 6208 13632 6528 13633
rect 6208 13568 6216 13632
rect 6280 13568 6296 13632
rect 6360 13568 6376 13632
rect 6440 13568 6456 13632
rect 6520 13568 6528 13632
rect 6208 13567 6528 13568
rect 11472 13632 11792 13633
rect 11472 13568 11480 13632
rect 11544 13568 11560 13632
rect 11624 13568 11640 13632
rect 11704 13568 11720 13632
rect 11784 13568 11792 13632
rect 11472 13567 11792 13568
rect 0 13290 480 13320
rect 2313 13290 2379 13293
rect 0 13288 2379 13290
rect 0 13232 2318 13288
rect 2374 13232 2379 13288
rect 0 13230 2379 13232
rect 0 13200 480 13230
rect 2313 13227 2379 13230
rect 13813 13290 13879 13293
rect 17520 13290 18000 13320
rect 13813 13288 18000 13290
rect 13813 13232 13818 13288
rect 13874 13232 18000 13288
rect 13813 13230 18000 13232
rect 13813 13227 13879 13230
rect 17520 13200 18000 13230
rect 3576 13088 3896 13089
rect 3576 13024 3584 13088
rect 3648 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3896 13088
rect 3576 13023 3896 13024
rect 8840 13088 9160 13089
rect 8840 13024 8848 13088
rect 8912 13024 8928 13088
rect 8992 13024 9008 13088
rect 9072 13024 9088 13088
rect 9152 13024 9160 13088
rect 8840 13023 9160 13024
rect 14104 13088 14424 13089
rect 14104 13024 14112 13088
rect 14176 13024 14192 13088
rect 14256 13024 14272 13088
rect 14336 13024 14352 13088
rect 14416 13024 14424 13088
rect 14104 13023 14424 13024
rect 12801 13020 12867 13021
rect 12750 13018 12756 13020
rect 12710 12958 12756 13018
rect 12820 13016 12867 13020
rect 12862 12960 12867 13016
rect 12750 12956 12756 12958
rect 12820 12956 12867 12960
rect 12801 12955 12867 12956
rect 0 12882 480 12912
rect 3325 12882 3391 12885
rect 17520 12882 18000 12912
rect 0 12880 3391 12882
rect 0 12824 3330 12880
rect 3386 12824 3391 12880
rect 0 12822 3391 12824
rect 0 12792 480 12822
rect 3325 12819 3391 12822
rect 16438 12822 18000 12882
rect 12893 12610 12959 12613
rect 13670 12610 13676 12612
rect 12893 12608 13676 12610
rect 12893 12552 12898 12608
rect 12954 12552 13676 12608
rect 12893 12550 13676 12552
rect 12893 12547 12959 12550
rect 13670 12548 13676 12550
rect 13740 12548 13746 12612
rect 14733 12610 14799 12613
rect 16297 12610 16363 12613
rect 16438 12610 16498 12822
rect 17520 12792 18000 12822
rect 14733 12608 16498 12610
rect 14733 12552 14738 12608
rect 14794 12552 16302 12608
rect 16358 12552 16498 12608
rect 14733 12550 16498 12552
rect 14733 12547 14799 12550
rect 16297 12547 16363 12550
rect 6208 12544 6528 12545
rect 0 12474 480 12504
rect 6208 12480 6216 12544
rect 6280 12480 6296 12544
rect 6360 12480 6376 12544
rect 6440 12480 6456 12544
rect 6520 12480 6528 12544
rect 6208 12479 6528 12480
rect 11472 12544 11792 12545
rect 11472 12480 11480 12544
rect 11544 12480 11560 12544
rect 11624 12480 11640 12544
rect 11704 12480 11720 12544
rect 11784 12480 11792 12544
rect 11472 12479 11792 12480
rect 4521 12474 4587 12477
rect 17520 12474 18000 12504
rect 0 12472 4587 12474
rect 0 12416 4526 12472
rect 4582 12416 4587 12472
rect 0 12414 4587 12416
rect 0 12384 480 12414
rect 4521 12411 4587 12414
rect 12160 12414 18000 12474
rect 3417 12338 3483 12341
rect 9029 12338 9095 12341
rect 3417 12336 9095 12338
rect 3417 12280 3422 12336
rect 3478 12280 9034 12336
rect 9090 12280 9095 12336
rect 3417 12278 9095 12280
rect 3417 12275 3483 12278
rect 9029 12275 9095 12278
rect 12014 12276 12020 12340
rect 12084 12338 12090 12340
rect 12160 12338 12220 12414
rect 17520 12384 18000 12414
rect 12801 12340 12867 12341
rect 13905 12340 13971 12341
rect 12084 12278 12220 12338
rect 12084 12276 12090 12278
rect 12750 12276 12756 12340
rect 12820 12338 12867 12340
rect 12820 12336 12912 12338
rect 12862 12280 12912 12336
rect 12820 12278 12912 12280
rect 12820 12276 12867 12278
rect 13854 12276 13860 12340
rect 13924 12338 13971 12340
rect 13924 12336 14016 12338
rect 13966 12280 14016 12336
rect 13924 12278 14016 12280
rect 13924 12276 13971 12278
rect 12801 12275 12867 12276
rect 13905 12275 13971 12276
rect 9397 12202 9463 12205
rect 14457 12202 14523 12205
rect 9397 12200 14523 12202
rect 9397 12144 9402 12200
rect 9458 12144 14462 12200
rect 14518 12144 14523 12200
rect 9397 12142 14523 12144
rect 9397 12139 9463 12142
rect 14457 12139 14523 12142
rect 0 12066 480 12096
rect 6637 12066 6703 12069
rect 7925 12066 7991 12069
rect 0 12006 3434 12066
rect 0 11976 480 12006
rect 3374 11794 3434 12006
rect 6637 12064 7991 12066
rect 6637 12008 6642 12064
rect 6698 12008 7930 12064
rect 7986 12008 7991 12064
rect 6637 12006 7991 12008
rect 6637 12003 6703 12006
rect 7925 12003 7991 12006
rect 14917 12066 14983 12069
rect 17520 12066 18000 12096
rect 14917 12064 18000 12066
rect 14917 12008 14922 12064
rect 14978 12008 18000 12064
rect 14917 12006 18000 12008
rect 14917 12003 14983 12006
rect 3576 12000 3896 12001
rect 3576 11936 3584 12000
rect 3648 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3896 12000
rect 3576 11935 3896 11936
rect 8840 12000 9160 12001
rect 8840 11936 8848 12000
rect 8912 11936 8928 12000
rect 8992 11936 9008 12000
rect 9072 11936 9088 12000
rect 9152 11936 9160 12000
rect 8840 11935 9160 11936
rect 14104 12000 14424 12001
rect 14104 11936 14112 12000
rect 14176 11936 14192 12000
rect 14256 11936 14272 12000
rect 14336 11936 14352 12000
rect 14416 11936 14424 12000
rect 17520 11976 18000 12006
rect 14104 11935 14424 11936
rect 13905 11930 13971 11933
rect 11470 11928 13971 11930
rect 11470 11872 13910 11928
rect 13966 11872 13971 11928
rect 11470 11870 13971 11872
rect 4613 11794 4679 11797
rect 10593 11794 10659 11797
rect 11470 11794 11530 11870
rect 13905 11867 13971 11870
rect 3374 11792 11530 11794
rect 3374 11736 4618 11792
rect 4674 11736 10598 11792
rect 10654 11736 11530 11792
rect 3374 11734 11530 11736
rect 12525 11794 12591 11797
rect 15561 11794 15627 11797
rect 12525 11792 15627 11794
rect 12525 11736 12530 11792
rect 12586 11736 15566 11792
rect 15622 11736 15627 11792
rect 12525 11734 15627 11736
rect 4613 11731 4679 11734
rect 10593 11731 10659 11734
rect 12525 11731 12591 11734
rect 15561 11731 15627 11734
rect 0 11658 480 11688
rect 2589 11658 2655 11661
rect 0 11656 2655 11658
rect 0 11600 2594 11656
rect 2650 11600 2655 11656
rect 0 11598 2655 11600
rect 0 11568 480 11598
rect 2589 11595 2655 11598
rect 5901 11658 5967 11661
rect 9581 11658 9647 11661
rect 5901 11656 9647 11658
rect 5901 11600 5906 11656
rect 5962 11600 9586 11656
rect 9642 11600 9647 11656
rect 5901 11598 9647 11600
rect 5901 11595 5967 11598
rect 9581 11595 9647 11598
rect 10961 11658 11027 11661
rect 12249 11658 12315 11661
rect 10961 11656 12315 11658
rect 10961 11600 10966 11656
rect 11022 11600 12254 11656
rect 12310 11600 12315 11656
rect 10961 11598 12315 11600
rect 10961 11595 11027 11598
rect 12249 11595 12315 11598
rect 13302 11596 13308 11660
rect 13372 11658 13378 11660
rect 17520 11658 18000 11688
rect 13372 11598 18000 11658
rect 13372 11596 13378 11598
rect 17520 11568 18000 11598
rect 6208 11456 6528 11457
rect 6208 11392 6216 11456
rect 6280 11392 6296 11456
rect 6360 11392 6376 11456
rect 6440 11392 6456 11456
rect 6520 11392 6528 11456
rect 6208 11391 6528 11392
rect 11472 11456 11792 11457
rect 11472 11392 11480 11456
rect 11544 11392 11560 11456
rect 11624 11392 11640 11456
rect 11704 11392 11720 11456
rect 11784 11392 11792 11456
rect 11472 11391 11792 11392
rect 5022 11324 5028 11388
rect 5092 11386 5098 11388
rect 5165 11386 5231 11389
rect 5092 11384 5231 11386
rect 5092 11328 5170 11384
rect 5226 11328 5231 11384
rect 5092 11326 5231 11328
rect 5092 11324 5098 11326
rect 5165 11323 5231 11326
rect 6913 11386 6979 11389
rect 7741 11386 7807 11389
rect 6913 11384 7807 11386
rect 6913 11328 6918 11384
rect 6974 11328 7746 11384
rect 7802 11328 7807 11384
rect 6913 11326 7807 11328
rect 6913 11323 6979 11326
rect 7741 11323 7807 11326
rect 12617 11386 12683 11389
rect 12893 11386 12959 11389
rect 12617 11384 12959 11386
rect 12617 11328 12622 11384
rect 12678 11328 12898 11384
rect 12954 11328 12959 11384
rect 12617 11326 12959 11328
rect 12617 11323 12683 11326
rect 12893 11323 12959 11326
rect 0 11250 480 11280
rect 3877 11250 3943 11253
rect 0 11248 3943 11250
rect 0 11192 3882 11248
rect 3938 11192 3943 11248
rect 0 11190 3943 11192
rect 0 11160 480 11190
rect 3877 11187 3943 11190
rect 4061 11250 4127 11253
rect 4061 11248 4170 11250
rect 4061 11192 4066 11248
rect 4122 11192 4170 11248
rect 4061 11187 4170 11192
rect 4838 11188 4844 11252
rect 4908 11250 4914 11252
rect 5165 11250 5231 11253
rect 12014 11250 12020 11252
rect 4908 11248 12020 11250
rect 4908 11192 5170 11248
rect 5226 11192 12020 11248
rect 4908 11190 12020 11192
rect 4908 11188 4914 11190
rect 5165 11187 5231 11190
rect 12014 11188 12020 11190
rect 12084 11188 12090 11252
rect 15745 11250 15811 11253
rect 17520 11250 18000 11280
rect 15745 11248 18000 11250
rect 15745 11192 15750 11248
rect 15806 11192 18000 11248
rect 15745 11190 18000 11192
rect 15745 11187 15811 11190
rect 4110 11114 4170 11187
rect 17520 11160 18000 11190
rect 8293 11114 8359 11117
rect 4110 11112 8359 11114
rect 4110 11056 8298 11112
rect 8354 11056 8359 11112
rect 4110 11054 8359 11056
rect 8293 11051 8359 11054
rect 12249 11114 12315 11117
rect 13261 11114 13327 11117
rect 12249 11112 13327 11114
rect 12249 11056 12254 11112
rect 12310 11056 13266 11112
rect 13322 11056 13327 11112
rect 12249 11054 13327 11056
rect 12249 11051 12315 11054
rect 13261 11051 13327 11054
rect 14365 11114 14431 11117
rect 14365 11112 14704 11114
rect 14365 11056 14370 11112
rect 14426 11056 14704 11112
rect 14365 11054 14704 11056
rect 14365 11051 14431 11054
rect 14644 10981 14704 11054
rect 14958 11052 14964 11116
rect 15028 11114 15034 11116
rect 15101 11114 15167 11117
rect 15028 11112 15167 11114
rect 15028 11056 15106 11112
rect 15162 11056 15167 11112
rect 15028 11054 15167 11056
rect 15028 11052 15034 11054
rect 15101 11051 15167 11054
rect 4337 10978 4403 10981
rect 7925 10978 7991 10981
rect 4337 10976 7991 10978
rect 4337 10920 4342 10976
rect 4398 10920 7930 10976
rect 7986 10920 7991 10976
rect 4337 10918 7991 10920
rect 4337 10915 4403 10918
rect 7925 10915 7991 10918
rect 13077 10978 13143 10981
rect 13261 10978 13327 10981
rect 13077 10976 13327 10978
rect 13077 10920 13082 10976
rect 13138 10920 13266 10976
rect 13322 10920 13327 10976
rect 13077 10918 13327 10920
rect 13077 10915 13143 10918
rect 13261 10915 13327 10918
rect 14641 10976 14707 10981
rect 15377 10978 15443 10981
rect 14641 10920 14646 10976
rect 14702 10920 14707 10976
rect 14641 10915 14707 10920
rect 14782 10976 15443 10978
rect 14782 10920 15382 10976
rect 15438 10920 15443 10976
rect 14782 10918 15443 10920
rect 3576 10912 3896 10913
rect 0 10842 480 10872
rect 3576 10848 3584 10912
rect 3648 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3896 10912
rect 3576 10847 3896 10848
rect 8840 10912 9160 10913
rect 8840 10848 8848 10912
rect 8912 10848 8928 10912
rect 8992 10848 9008 10912
rect 9072 10848 9088 10912
rect 9152 10848 9160 10912
rect 8840 10847 9160 10848
rect 14104 10912 14424 10913
rect 14104 10848 14112 10912
rect 14176 10848 14192 10912
rect 14256 10848 14272 10912
rect 14336 10848 14352 10912
rect 14416 10848 14424 10912
rect 14104 10847 14424 10848
rect 3325 10842 3391 10845
rect 4337 10842 4403 10845
rect 5165 10842 5231 10845
rect 0 10840 3434 10842
rect 0 10784 3330 10840
rect 3386 10784 3434 10840
rect 0 10782 3434 10784
rect 0 10752 480 10782
rect 3325 10779 3434 10782
rect 4337 10840 5231 10842
rect 4337 10784 4342 10840
rect 4398 10784 5170 10840
rect 5226 10784 5231 10840
rect 4337 10782 5231 10784
rect 4337 10779 4403 10782
rect 5165 10779 5231 10782
rect 10358 10780 10364 10844
rect 10428 10842 10434 10844
rect 10685 10842 10751 10845
rect 10428 10840 10751 10842
rect 10428 10784 10690 10840
rect 10746 10784 10751 10840
rect 10428 10782 10751 10784
rect 10428 10780 10434 10782
rect 10685 10779 10751 10782
rect 11973 10842 12039 10845
rect 12525 10842 12591 10845
rect 13537 10842 13603 10845
rect 11973 10840 12591 10842
rect 11973 10784 11978 10840
rect 12034 10784 12530 10840
rect 12586 10784 12591 10840
rect 11973 10782 12591 10784
rect 11973 10779 12039 10782
rect 12525 10779 12591 10782
rect 13310 10840 13603 10842
rect 13310 10784 13542 10840
rect 13598 10784 13603 10840
rect 13310 10782 13603 10784
rect 3374 10706 3434 10779
rect 6177 10706 6243 10709
rect 11789 10706 11855 10709
rect 3374 10704 6243 10706
rect 3374 10648 6182 10704
rect 6238 10648 6243 10704
rect 3374 10646 6243 10648
rect 6177 10643 6243 10646
rect 7606 10704 11855 10706
rect 7606 10648 11794 10704
rect 11850 10648 11855 10704
rect 7606 10646 11855 10648
rect 5165 10570 5231 10573
rect 7606 10570 7666 10646
rect 11789 10643 11855 10646
rect 11973 10706 12039 10709
rect 12893 10706 12959 10709
rect 11973 10704 12959 10706
rect 11973 10648 11978 10704
rect 12034 10648 12898 10704
rect 12954 10648 12959 10704
rect 11973 10646 12959 10648
rect 11973 10643 12039 10646
rect 12893 10643 12959 10646
rect 5165 10568 7666 10570
rect 5165 10512 5170 10568
rect 5226 10512 7666 10568
rect 5165 10510 7666 10512
rect 8201 10570 8267 10573
rect 12617 10570 12683 10573
rect 8201 10568 12683 10570
rect 8201 10512 8206 10568
rect 8262 10512 12622 10568
rect 12678 10512 12683 10568
rect 8201 10510 12683 10512
rect 5165 10507 5231 10510
rect 8201 10507 8267 10510
rect 12617 10507 12683 10510
rect 0 10434 480 10464
rect 3693 10434 3759 10437
rect 0 10432 3759 10434
rect 0 10376 3698 10432
rect 3754 10376 3759 10432
rect 0 10374 3759 10376
rect 0 10344 480 10374
rect 3693 10371 3759 10374
rect 12433 10434 12499 10437
rect 13310 10434 13370 10782
rect 13537 10779 13603 10782
rect 13629 10706 13695 10709
rect 14782 10706 14842 10918
rect 15377 10915 15443 10918
rect 15285 10842 15351 10845
rect 17520 10842 18000 10872
rect 15285 10840 18000 10842
rect 15285 10784 15290 10840
rect 15346 10784 18000 10840
rect 15285 10782 18000 10784
rect 15285 10779 15351 10782
rect 17520 10752 18000 10782
rect 13629 10704 14842 10706
rect 13629 10648 13634 10704
rect 13690 10648 14842 10704
rect 13629 10646 14842 10648
rect 13629 10643 13695 10646
rect 12433 10432 13370 10434
rect 12433 10376 12438 10432
rect 12494 10376 13370 10432
rect 12433 10374 13370 10376
rect 13905 10434 13971 10437
rect 17520 10434 18000 10464
rect 13905 10432 18000 10434
rect 13905 10376 13910 10432
rect 13966 10376 18000 10432
rect 13905 10374 18000 10376
rect 12433 10371 12499 10374
rect 13905 10371 13971 10374
rect 6208 10368 6528 10369
rect 6208 10304 6216 10368
rect 6280 10304 6296 10368
rect 6360 10304 6376 10368
rect 6440 10304 6456 10368
rect 6520 10304 6528 10368
rect 6208 10303 6528 10304
rect 11472 10368 11792 10369
rect 11472 10304 11480 10368
rect 11544 10304 11560 10368
rect 11624 10304 11640 10368
rect 11704 10304 11720 10368
rect 11784 10304 11792 10368
rect 17520 10344 18000 10374
rect 11472 10303 11792 10304
rect 3417 10300 3483 10301
rect 3366 10236 3372 10300
rect 3436 10298 3483 10300
rect 5901 10298 5967 10301
rect 3436 10296 5967 10298
rect 3478 10240 5906 10296
rect 5962 10240 5967 10296
rect 3436 10238 5967 10240
rect 3436 10236 3483 10238
rect 3417 10235 3483 10236
rect 5901 10235 5967 10238
rect 9857 10298 9923 10301
rect 9990 10298 9996 10300
rect 9857 10296 9996 10298
rect 9857 10240 9862 10296
rect 9918 10240 9996 10296
rect 9857 10238 9996 10240
rect 9857 10235 9923 10238
rect 9990 10236 9996 10238
rect 10060 10236 10066 10300
rect 10777 10298 10843 10301
rect 11278 10298 11284 10300
rect 10777 10296 11284 10298
rect 10777 10240 10782 10296
rect 10838 10240 11284 10296
rect 10777 10238 11284 10240
rect 10777 10235 10843 10238
rect 11278 10236 11284 10238
rect 11348 10236 11354 10300
rect 12893 10298 12959 10301
rect 14825 10298 14891 10301
rect 12893 10296 14891 10298
rect 12893 10240 12898 10296
rect 12954 10240 14830 10296
rect 14886 10240 14891 10296
rect 12893 10238 14891 10240
rect 12893 10235 12959 10238
rect 14825 10235 14891 10238
rect 5717 10162 5783 10165
rect 6821 10162 6887 10165
rect 5717 10160 6887 10162
rect 5717 10104 5722 10160
rect 5778 10104 6826 10160
rect 6882 10104 6887 10160
rect 5717 10102 6887 10104
rect 5717 10099 5783 10102
rect 6821 10099 6887 10102
rect 9213 10162 9279 10165
rect 15285 10162 15351 10165
rect 9213 10160 15351 10162
rect 9213 10104 9218 10160
rect 9274 10104 15290 10160
rect 15346 10104 15351 10160
rect 9213 10102 15351 10104
rect 9213 10099 9279 10102
rect 15285 10099 15351 10102
rect 1853 10026 1919 10029
rect 9857 10026 9923 10029
rect 12893 10026 12959 10029
rect 1853 10024 9322 10026
rect 1853 9968 1858 10024
rect 1914 9968 9322 10024
rect 1853 9966 9322 9968
rect 1853 9963 1919 9966
rect 0 9890 480 9920
rect 2497 9890 2563 9893
rect 0 9888 2563 9890
rect 0 9832 2502 9888
rect 2558 9832 2563 9888
rect 0 9830 2563 9832
rect 0 9800 480 9830
rect 2497 9827 2563 9830
rect 4153 9890 4219 9893
rect 4286 9890 4292 9892
rect 4153 9888 4292 9890
rect 4153 9832 4158 9888
rect 4214 9832 4292 9888
rect 4153 9830 4292 9832
rect 4153 9827 4219 9830
rect 4286 9828 4292 9830
rect 4356 9828 4362 9892
rect 4705 9890 4771 9893
rect 5022 9890 5028 9892
rect 4705 9888 5028 9890
rect 4705 9832 4710 9888
rect 4766 9832 5028 9888
rect 4705 9830 5028 9832
rect 4705 9827 4771 9830
rect 5022 9828 5028 9830
rect 5092 9828 5098 9892
rect 5901 9890 5967 9893
rect 8385 9890 8451 9893
rect 5901 9888 8451 9890
rect 5901 9832 5906 9888
rect 5962 9832 8390 9888
rect 8446 9832 8451 9888
rect 5901 9830 8451 9832
rect 9262 9890 9322 9966
rect 9857 10024 12959 10026
rect 9857 9968 9862 10024
rect 9918 9968 12898 10024
rect 12954 9968 12959 10024
rect 9857 9966 12959 9968
rect 9857 9963 9923 9966
rect 12893 9963 12959 9966
rect 13118 9964 13124 10028
rect 13188 10026 13194 10028
rect 13188 9966 14658 10026
rect 13188 9964 13194 9966
rect 12433 9890 12499 9893
rect 13854 9890 13860 9892
rect 9262 9888 13860 9890
rect 9262 9832 12438 9888
rect 12494 9832 13860 9888
rect 9262 9830 13860 9832
rect 5901 9827 5967 9830
rect 8385 9827 8451 9830
rect 12433 9827 12499 9830
rect 13854 9828 13860 9830
rect 13924 9828 13930 9892
rect 14598 9890 14658 9966
rect 17520 9890 18000 9920
rect 14598 9830 18000 9890
rect 3576 9824 3896 9825
rect 3576 9760 3584 9824
rect 3648 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3896 9824
rect 3576 9759 3896 9760
rect 8840 9824 9160 9825
rect 8840 9760 8848 9824
rect 8912 9760 8928 9824
rect 8992 9760 9008 9824
rect 9072 9760 9088 9824
rect 9152 9760 9160 9824
rect 8840 9759 9160 9760
rect 14104 9824 14424 9825
rect 14104 9760 14112 9824
rect 14176 9760 14192 9824
rect 14256 9760 14272 9824
rect 14336 9760 14352 9824
rect 14416 9760 14424 9824
rect 17520 9800 18000 9830
rect 14104 9759 14424 9760
rect 6545 9754 6611 9757
rect 7005 9754 7071 9757
rect 6545 9752 7071 9754
rect 6545 9696 6550 9752
rect 6606 9696 7010 9752
rect 7066 9696 7071 9752
rect 6545 9694 7071 9696
rect 6545 9691 6611 9694
rect 7005 9691 7071 9694
rect 10869 9754 10935 9757
rect 12382 9754 12388 9756
rect 10869 9752 12388 9754
rect 10869 9696 10874 9752
rect 10930 9696 12388 9752
rect 10869 9694 12388 9696
rect 10869 9691 10935 9694
rect 12382 9692 12388 9694
rect 12452 9692 12458 9756
rect 12525 9754 12591 9757
rect 13169 9754 13235 9757
rect 13302 9754 13308 9756
rect 12525 9752 13308 9754
rect 12525 9696 12530 9752
rect 12586 9696 13174 9752
rect 13230 9696 13308 9752
rect 12525 9694 13308 9696
rect 12525 9691 12591 9694
rect 13169 9691 13235 9694
rect 13302 9692 13308 9694
rect 13372 9692 13378 9756
rect 2681 9618 2747 9621
rect 4245 9618 4311 9621
rect 2681 9616 4311 9618
rect 2681 9560 2686 9616
rect 2742 9560 4250 9616
rect 4306 9560 4311 9616
rect 2681 9558 4311 9560
rect 2681 9555 2747 9558
rect 4245 9555 4311 9558
rect 6269 9618 6335 9621
rect 10041 9618 10107 9621
rect 6269 9616 10107 9618
rect 6269 9560 6274 9616
rect 6330 9560 10046 9616
rect 10102 9560 10107 9616
rect 6269 9558 10107 9560
rect 6269 9555 6335 9558
rect 10041 9555 10107 9558
rect 13670 9556 13676 9620
rect 13740 9618 13746 9620
rect 14549 9618 14615 9621
rect 13740 9616 14615 9618
rect 13740 9560 14554 9616
rect 14610 9560 14615 9616
rect 13740 9558 14615 9560
rect 13740 9556 13746 9558
rect 14549 9555 14615 9558
rect 0 9482 480 9512
rect 4705 9482 4771 9485
rect 9254 9482 9260 9484
rect 0 9422 3296 9482
rect 0 9392 480 9422
rect 3236 9349 3296 9422
rect 4705 9480 9260 9482
rect 4705 9424 4710 9480
rect 4766 9424 9260 9480
rect 4705 9422 9260 9424
rect 4705 9419 4771 9422
rect 9254 9420 9260 9422
rect 9324 9420 9330 9484
rect 9765 9482 9831 9485
rect 10685 9482 10751 9485
rect 13353 9482 13419 9485
rect 15469 9482 15535 9485
rect 17520 9482 18000 9512
rect 9765 9480 10751 9482
rect 9765 9424 9770 9480
rect 9826 9424 10690 9480
rect 10746 9424 10751 9480
rect 9765 9422 10751 9424
rect 9765 9419 9831 9422
rect 10685 9419 10751 9422
rect 11286 9422 13232 9482
rect 3233 9346 3299 9349
rect 5574 9346 5580 9348
rect 3233 9344 5580 9346
rect 3233 9288 3238 9344
rect 3294 9288 5580 9344
rect 3233 9286 5580 9288
rect 3233 9283 3299 9286
rect 5574 9284 5580 9286
rect 5644 9284 5650 9348
rect 10777 9346 10843 9349
rect 11286 9346 11346 9422
rect 10777 9344 11346 9346
rect 10777 9288 10782 9344
rect 10838 9288 11346 9344
rect 10777 9286 11346 9288
rect 12341 9346 12407 9349
rect 12985 9346 13051 9349
rect 12341 9344 13051 9346
rect 12341 9288 12346 9344
rect 12402 9288 12990 9344
rect 13046 9288 13051 9344
rect 12341 9286 13051 9288
rect 13172 9346 13232 9422
rect 13353 9480 18000 9482
rect 13353 9424 13358 9480
rect 13414 9424 15474 9480
rect 15530 9424 18000 9480
rect 13353 9422 18000 9424
rect 13353 9419 13419 9422
rect 15469 9419 15535 9422
rect 17520 9392 18000 9422
rect 15653 9346 15719 9349
rect 13172 9344 15762 9346
rect 13172 9288 15658 9344
rect 15714 9288 15762 9344
rect 13172 9286 15762 9288
rect 10777 9283 10843 9286
rect 12341 9283 12407 9286
rect 12985 9283 13051 9286
rect 15653 9283 15762 9286
rect 6208 9280 6528 9281
rect 6208 9216 6216 9280
rect 6280 9216 6296 9280
rect 6360 9216 6376 9280
rect 6440 9216 6456 9280
rect 6520 9216 6528 9280
rect 6208 9215 6528 9216
rect 11472 9280 11792 9281
rect 11472 9216 11480 9280
rect 11544 9216 11560 9280
rect 11624 9216 11640 9280
rect 11704 9216 11720 9280
rect 11784 9216 11792 9280
rect 11472 9215 11792 9216
rect 2773 9210 2839 9213
rect 4102 9210 4108 9212
rect 2773 9208 4108 9210
rect 2773 9152 2778 9208
rect 2834 9152 4108 9208
rect 2773 9150 4108 9152
rect 2773 9147 2839 9150
rect 4102 9148 4108 9150
rect 4172 9210 4178 9212
rect 4245 9210 4311 9213
rect 4172 9208 4311 9210
rect 4172 9152 4250 9208
rect 4306 9152 4311 9208
rect 4172 9150 4311 9152
rect 4172 9148 4178 9150
rect 4245 9147 4311 9150
rect 8201 9210 8267 9213
rect 8702 9210 8708 9212
rect 8201 9208 8708 9210
rect 8201 9152 8206 9208
rect 8262 9152 8708 9208
rect 8201 9150 8708 9152
rect 8201 9147 8267 9150
rect 8702 9148 8708 9150
rect 8772 9148 8778 9212
rect 12249 9210 12315 9213
rect 13077 9210 13143 9213
rect 12249 9208 13143 9210
rect 12249 9152 12254 9208
rect 12310 9152 13082 9208
rect 13138 9152 13143 9208
rect 12249 9150 13143 9152
rect 12249 9147 12315 9150
rect 13077 9147 13143 9150
rect 0 9074 480 9104
rect 1945 9074 2011 9077
rect 8569 9074 8635 9077
rect 0 9072 2011 9074
rect 0 9016 1950 9072
rect 2006 9016 2011 9072
rect 0 9014 2011 9016
rect 0 8984 480 9014
rect 1945 9011 2011 9014
rect 2500 9072 8635 9074
rect 2500 9016 8574 9072
rect 8630 9016 8635 9072
rect 2500 9014 8635 9016
rect 2500 8941 2560 9014
rect 8569 9011 8635 9014
rect 9121 9074 9187 9077
rect 13997 9074 14063 9077
rect 9121 9072 14063 9074
rect 9121 9016 9126 9072
rect 9182 9016 14002 9072
rect 14058 9016 14063 9072
rect 9121 9014 14063 9016
rect 15702 9074 15762 9283
rect 17520 9074 18000 9104
rect 15702 9014 18000 9074
rect 9121 9011 9187 9014
rect 13997 9011 14063 9014
rect 17520 8984 18000 9014
rect 2497 8936 2563 8941
rect 8017 8938 8083 8941
rect 2497 8880 2502 8936
rect 2558 8880 2563 8936
rect 2497 8875 2563 8880
rect 3420 8936 8083 8938
rect 3420 8880 8022 8936
rect 8078 8880 8083 8936
rect 3420 8878 8083 8880
rect 1393 8802 1459 8805
rect 3420 8802 3480 8878
rect 8017 8875 8083 8878
rect 8753 8938 8819 8941
rect 12709 8938 12775 8941
rect 13537 8938 13603 8941
rect 8753 8936 12634 8938
rect 8753 8880 8758 8936
rect 8814 8880 12634 8936
rect 8753 8878 12634 8880
rect 8753 8875 8819 8878
rect 9489 8804 9555 8805
rect 1393 8800 3480 8802
rect 1393 8744 1398 8800
rect 1454 8744 3480 8800
rect 1393 8742 3480 8744
rect 1393 8739 1459 8742
rect 9438 8740 9444 8804
rect 9508 8802 9555 8804
rect 9508 8800 9600 8802
rect 9550 8744 9600 8800
rect 9508 8742 9600 8744
rect 9508 8740 9555 8742
rect 9806 8740 9812 8804
rect 9876 8802 9882 8804
rect 9949 8802 10015 8805
rect 11329 8804 11395 8805
rect 9876 8800 10015 8802
rect 9876 8744 9954 8800
rect 10010 8744 10015 8800
rect 9876 8742 10015 8744
rect 9876 8740 9882 8742
rect 9489 8739 9555 8740
rect 9949 8739 10015 8742
rect 11278 8740 11284 8804
rect 11348 8802 11395 8804
rect 11881 8802 11947 8805
rect 12198 8802 12204 8804
rect 11348 8800 11440 8802
rect 11390 8744 11440 8800
rect 11348 8742 11440 8744
rect 11881 8800 12204 8802
rect 11881 8744 11886 8800
rect 11942 8744 12204 8800
rect 11881 8742 12204 8744
rect 11348 8740 11395 8742
rect 11329 8739 11395 8740
rect 11881 8739 11947 8742
rect 12198 8740 12204 8742
rect 12268 8740 12274 8804
rect 12574 8802 12634 8878
rect 12709 8936 13603 8938
rect 12709 8880 12714 8936
rect 12770 8880 13542 8936
rect 13598 8880 13603 8936
rect 12709 8878 13603 8880
rect 12709 8875 12775 8878
rect 13537 8875 13603 8878
rect 13537 8802 13603 8805
rect 12574 8800 13603 8802
rect 12574 8744 13542 8800
rect 13598 8744 13603 8800
rect 12574 8742 13603 8744
rect 13537 8739 13603 8742
rect 3576 8736 3896 8737
rect 0 8666 480 8696
rect 3576 8672 3584 8736
rect 3648 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3896 8736
rect 3576 8671 3896 8672
rect 8840 8736 9160 8737
rect 8840 8672 8848 8736
rect 8912 8672 8928 8736
rect 8992 8672 9008 8736
rect 9072 8672 9088 8736
rect 9152 8672 9160 8736
rect 8840 8671 9160 8672
rect 14104 8736 14424 8737
rect 14104 8672 14112 8736
rect 14176 8672 14192 8736
rect 14256 8672 14272 8736
rect 14336 8672 14352 8736
rect 14416 8672 14424 8736
rect 14104 8671 14424 8672
rect 2681 8666 2747 8669
rect 3182 8666 3188 8668
rect 0 8664 3188 8666
rect 0 8608 2686 8664
rect 2742 8608 3188 8664
rect 0 8606 3188 8608
rect 0 8576 480 8606
rect 2681 8603 2747 8606
rect 3182 8604 3188 8606
rect 3252 8604 3258 8668
rect 10041 8666 10107 8669
rect 13813 8666 13879 8669
rect 10041 8664 13879 8666
rect 10041 8608 10046 8664
rect 10102 8608 13818 8664
rect 13874 8608 13879 8664
rect 10041 8606 13879 8608
rect 10041 8603 10107 8606
rect 13813 8603 13879 8606
rect 16113 8666 16179 8669
rect 17520 8666 18000 8696
rect 16113 8664 18000 8666
rect 16113 8608 16118 8664
rect 16174 8608 18000 8664
rect 16113 8606 18000 8608
rect 16113 8603 16179 8606
rect 17520 8576 18000 8606
rect 9397 8530 9463 8533
rect 12065 8530 12131 8533
rect 9397 8528 12131 8530
rect 9397 8472 9402 8528
rect 9458 8472 12070 8528
rect 12126 8472 12131 8528
rect 9397 8470 12131 8472
rect 9397 8467 9463 8470
rect 12065 8467 12131 8470
rect 13629 8530 13695 8533
rect 14457 8530 14523 8533
rect 14917 8530 14983 8533
rect 13629 8528 14983 8530
rect 13629 8472 13634 8528
rect 13690 8472 14462 8528
rect 14518 8472 14922 8528
rect 14978 8472 14983 8528
rect 13629 8470 14983 8472
rect 13629 8467 13695 8470
rect 14457 8467 14523 8470
rect 14917 8467 14983 8470
rect 3049 8396 3115 8397
rect 2998 8332 3004 8396
rect 3068 8394 3115 8396
rect 8201 8394 8267 8397
rect 3068 8392 8267 8394
rect 3110 8336 8206 8392
rect 8262 8336 8267 8392
rect 3068 8334 8267 8336
rect 3068 8332 3115 8334
rect 3049 8331 3115 8332
rect 8201 8331 8267 8334
rect 9857 8394 9923 8397
rect 10041 8394 10107 8397
rect 9857 8392 10107 8394
rect 9857 8336 9862 8392
rect 9918 8336 10046 8392
rect 10102 8336 10107 8392
rect 9857 8334 10107 8336
rect 9857 8331 9923 8334
rect 10041 8331 10107 8334
rect 11237 8394 11303 8397
rect 14641 8394 14707 8397
rect 11237 8392 14707 8394
rect 11237 8336 11242 8392
rect 11298 8336 14646 8392
rect 14702 8336 14707 8392
rect 11237 8334 14707 8336
rect 11237 8331 11303 8334
rect 14641 8331 14707 8334
rect 0 8258 480 8288
rect 4061 8258 4127 8261
rect 0 8256 4127 8258
rect 0 8200 4066 8256
rect 4122 8200 4127 8256
rect 0 8198 4127 8200
rect 0 8168 480 8198
rect 4061 8195 4127 8198
rect 7833 8258 7899 8261
rect 9489 8258 9555 8261
rect 7833 8256 9555 8258
rect 7833 8200 7838 8256
rect 7894 8200 9494 8256
rect 9550 8200 9555 8256
rect 7833 8198 9555 8200
rect 7833 8195 7899 8198
rect 9489 8195 9555 8198
rect 9673 8258 9739 8261
rect 10542 8258 10548 8260
rect 9673 8256 10548 8258
rect 9673 8200 9678 8256
rect 9734 8200 10548 8256
rect 9673 8198 10548 8200
rect 9673 8195 9739 8198
rect 10542 8196 10548 8198
rect 10612 8196 10618 8260
rect 13905 8258 13971 8261
rect 17520 8258 18000 8288
rect 13905 8256 18000 8258
rect 13905 8200 13910 8256
rect 13966 8200 18000 8256
rect 13905 8198 18000 8200
rect 13905 8195 13971 8198
rect 6208 8192 6528 8193
rect 6208 8128 6216 8192
rect 6280 8128 6296 8192
rect 6360 8128 6376 8192
rect 6440 8128 6456 8192
rect 6520 8128 6528 8192
rect 6208 8127 6528 8128
rect 11472 8192 11792 8193
rect 11472 8128 11480 8192
rect 11544 8128 11560 8192
rect 11624 8128 11640 8192
rect 11704 8128 11720 8192
rect 11784 8128 11792 8192
rect 17520 8168 18000 8198
rect 11472 8127 11792 8128
rect 8477 8122 8543 8125
rect 10777 8122 10843 8125
rect 8477 8120 10843 8122
rect 8477 8064 8482 8120
rect 8538 8064 10782 8120
rect 10838 8064 10843 8120
rect 8477 8062 10843 8064
rect 8477 8059 8543 8062
rect 10777 8059 10843 8062
rect 13629 8122 13695 8125
rect 15101 8122 15167 8125
rect 13629 8120 15167 8122
rect 13629 8064 13634 8120
rect 13690 8064 15106 8120
rect 15162 8064 15167 8120
rect 13629 8062 15167 8064
rect 13629 8059 13695 8062
rect 15101 8059 15167 8062
rect 9438 7924 9444 7988
rect 9508 7986 9514 7988
rect 13813 7986 13879 7989
rect 9508 7984 13879 7986
rect 9508 7928 13818 7984
rect 13874 7928 13879 7984
rect 9508 7926 13879 7928
rect 9508 7924 9514 7926
rect 13813 7923 13879 7926
rect 0 7850 480 7880
rect 4153 7850 4219 7853
rect 4429 7850 4495 7853
rect 0 7848 4219 7850
rect 0 7792 4158 7848
rect 4214 7792 4219 7848
rect 0 7790 4219 7792
rect 0 7760 480 7790
rect 4153 7787 4219 7790
rect 4294 7848 4495 7850
rect 4294 7792 4434 7848
rect 4490 7792 4495 7848
rect 4294 7790 4495 7792
rect 3576 7648 3896 7649
rect 3576 7584 3584 7648
rect 3648 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3896 7648
rect 3576 7583 3896 7584
rect 4294 7581 4354 7790
rect 4429 7787 4495 7790
rect 5717 7850 5783 7853
rect 5717 7848 9322 7850
rect 5717 7792 5722 7848
rect 5778 7792 9322 7848
rect 5717 7790 9322 7792
rect 5717 7787 5783 7790
rect 9262 7714 9322 7790
rect 9438 7788 9444 7852
rect 9508 7850 9514 7852
rect 11697 7850 11763 7853
rect 9508 7848 11763 7850
rect 9508 7792 11702 7848
rect 11758 7792 11763 7848
rect 9508 7790 11763 7792
rect 9508 7788 9514 7790
rect 11697 7787 11763 7790
rect 13445 7850 13511 7853
rect 15285 7850 15351 7853
rect 17520 7850 18000 7880
rect 13445 7848 14842 7850
rect 13445 7792 13450 7848
rect 13506 7792 14842 7848
rect 13445 7790 14842 7792
rect 13445 7787 13511 7790
rect 12341 7714 12407 7717
rect 12893 7714 12959 7717
rect 9262 7712 12959 7714
rect 9262 7656 12346 7712
rect 12402 7656 12898 7712
rect 12954 7656 12959 7712
rect 9262 7654 12959 7656
rect 12341 7651 12407 7654
rect 12893 7651 12959 7654
rect 8840 7648 9160 7649
rect 8840 7584 8848 7648
rect 8912 7584 8928 7648
rect 8992 7584 9008 7648
rect 9072 7584 9088 7648
rect 9152 7584 9160 7648
rect 8840 7583 9160 7584
rect 14104 7648 14424 7649
rect 14104 7584 14112 7648
rect 14176 7584 14192 7648
rect 14256 7584 14272 7648
rect 14336 7584 14352 7648
rect 14416 7584 14424 7648
rect 14104 7583 14424 7584
rect 4245 7576 4354 7581
rect 4245 7520 4250 7576
rect 4306 7520 4354 7576
rect 4245 7518 4354 7520
rect 4245 7515 4311 7518
rect 9254 7516 9260 7580
rect 9324 7578 9330 7580
rect 13629 7578 13695 7581
rect 9324 7576 13695 7578
rect 9324 7520 13634 7576
rect 13690 7520 13695 7576
rect 9324 7518 13695 7520
rect 9324 7516 9330 7518
rect 13629 7515 13695 7518
rect 0 7442 480 7472
rect 1577 7442 1643 7445
rect 0 7440 1643 7442
rect 0 7384 1582 7440
rect 1638 7384 1643 7440
rect 0 7382 1643 7384
rect 0 7352 480 7382
rect 1577 7379 1643 7382
rect 8293 7442 8359 7445
rect 9438 7442 9444 7444
rect 8293 7440 9444 7442
rect 8293 7384 8298 7440
rect 8354 7384 9444 7440
rect 8293 7382 9444 7384
rect 8293 7379 8359 7382
rect 9438 7380 9444 7382
rect 9508 7380 9514 7444
rect 14641 7442 14707 7445
rect 9814 7440 14707 7442
rect 9814 7384 14646 7440
rect 14702 7384 14707 7440
rect 9814 7382 14707 7384
rect 14782 7442 14842 7790
rect 15285 7848 18000 7850
rect 15285 7792 15290 7848
rect 15346 7792 18000 7848
rect 15285 7790 18000 7792
rect 15285 7787 15351 7790
rect 17520 7760 18000 7790
rect 17520 7442 18000 7472
rect 14782 7382 18000 7442
rect 2589 7306 2655 7309
rect 9489 7306 9555 7309
rect 9814 7308 9874 7382
rect 14641 7379 14707 7382
rect 17520 7352 18000 7382
rect 2589 7304 9555 7306
rect 2589 7248 2594 7304
rect 2650 7248 9494 7304
rect 9550 7248 9555 7304
rect 2589 7246 9555 7248
rect 2589 7243 2655 7246
rect 9489 7243 9555 7246
rect 9806 7244 9812 7308
rect 9876 7244 9882 7308
rect 11053 7306 11119 7309
rect 14457 7306 14523 7309
rect 11053 7304 14523 7306
rect 11053 7248 11058 7304
rect 11114 7248 14462 7304
rect 14518 7248 14523 7304
rect 11053 7246 14523 7248
rect 11053 7243 11119 7246
rect 14457 7243 14523 7246
rect 8477 7170 8543 7173
rect 10685 7170 10751 7173
rect 8477 7168 10751 7170
rect 8477 7112 8482 7168
rect 8538 7112 10690 7168
rect 10746 7112 10751 7168
rect 8477 7110 10751 7112
rect 8477 7107 8543 7110
rect 10685 7107 10751 7110
rect 6208 7104 6528 7105
rect 0 7034 480 7064
rect 6208 7040 6216 7104
rect 6280 7040 6296 7104
rect 6360 7040 6376 7104
rect 6440 7040 6456 7104
rect 6520 7040 6528 7104
rect 6208 7039 6528 7040
rect 11472 7104 11792 7105
rect 11472 7040 11480 7104
rect 11544 7040 11560 7104
rect 11624 7040 11640 7104
rect 11704 7040 11720 7104
rect 11784 7040 11792 7104
rect 11472 7039 11792 7040
rect 3417 7034 3483 7037
rect 0 7032 3483 7034
rect 0 6976 3422 7032
rect 3478 6976 3483 7032
rect 0 6974 3483 6976
rect 0 6944 480 6974
rect 3417 6971 3483 6974
rect 8518 6972 8524 7036
rect 8588 7034 8594 7036
rect 8753 7034 8819 7037
rect 11237 7034 11303 7037
rect 8588 7032 11303 7034
rect 8588 6976 8758 7032
rect 8814 6976 11242 7032
rect 11298 6976 11303 7032
rect 8588 6974 11303 6976
rect 8588 6972 8594 6974
rect 8753 6971 8819 6974
rect 11237 6971 11303 6974
rect 14825 7034 14891 7037
rect 17520 7034 18000 7064
rect 14825 7032 18000 7034
rect 14825 6976 14830 7032
rect 14886 6976 18000 7032
rect 14825 6974 18000 6976
rect 14825 6971 14891 6974
rect 17520 6944 18000 6974
rect 1301 6898 1367 6901
rect 2773 6898 2839 6901
rect 3417 6900 3483 6901
rect 3366 6898 3372 6900
rect 1301 6896 2839 6898
rect 1301 6840 1306 6896
rect 1362 6840 2778 6896
rect 2834 6840 2839 6896
rect 1301 6838 2839 6840
rect 3326 6838 3372 6898
rect 3436 6896 3483 6900
rect 3478 6840 3483 6896
rect 1301 6835 1367 6838
rect 2773 6835 2839 6838
rect 3366 6836 3372 6838
rect 3436 6836 3483 6840
rect 7598 6836 7604 6900
rect 7668 6898 7674 6900
rect 8109 6898 8175 6901
rect 7668 6896 8175 6898
rect 7668 6840 8114 6896
rect 8170 6840 8175 6896
rect 7668 6838 8175 6840
rect 7668 6836 7674 6838
rect 3417 6835 3483 6836
rect 8109 6835 8175 6838
rect 7281 6762 7347 6765
rect 8845 6762 8911 6765
rect 7281 6760 8911 6762
rect 7281 6704 7286 6760
rect 7342 6704 8850 6760
rect 8906 6704 8911 6760
rect 7281 6702 8911 6704
rect 7281 6699 7347 6702
rect 8845 6699 8911 6702
rect 9121 6762 9187 6765
rect 9949 6762 10015 6765
rect 9121 6760 10015 6762
rect 9121 6704 9126 6760
rect 9182 6704 9954 6760
rect 10010 6704 10015 6760
rect 9121 6702 10015 6704
rect 9121 6699 9187 6702
rect 9949 6699 10015 6702
rect 11789 6762 11855 6765
rect 14917 6762 14983 6765
rect 11789 6760 14983 6762
rect 11789 6704 11794 6760
rect 11850 6704 14922 6760
rect 14978 6704 14983 6760
rect 11789 6702 14983 6704
rect 11789 6699 11855 6702
rect 14917 6699 14983 6702
rect 4102 6564 4108 6628
rect 4172 6626 4178 6628
rect 4337 6626 4403 6629
rect 4172 6624 4403 6626
rect 4172 6568 4342 6624
rect 4398 6568 4403 6624
rect 4172 6566 4403 6568
rect 4172 6564 4178 6566
rect 4337 6563 4403 6566
rect 3576 6560 3896 6561
rect 0 6490 480 6520
rect 3576 6496 3584 6560
rect 3648 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3896 6560
rect 3576 6495 3896 6496
rect 8840 6560 9160 6561
rect 8840 6496 8848 6560
rect 8912 6496 8928 6560
rect 8992 6496 9008 6560
rect 9072 6496 9088 6560
rect 9152 6496 9160 6560
rect 8840 6495 9160 6496
rect 14104 6560 14424 6561
rect 14104 6496 14112 6560
rect 14176 6496 14192 6560
rect 14256 6496 14272 6560
rect 14336 6496 14352 6560
rect 14416 6496 14424 6560
rect 14104 6495 14424 6496
rect 2865 6490 2931 6493
rect 0 6488 2931 6490
rect 0 6432 2870 6488
rect 2926 6432 2931 6488
rect 0 6430 2931 6432
rect 0 6400 480 6430
rect 2865 6427 2931 6430
rect 15653 6490 15719 6493
rect 17520 6490 18000 6520
rect 15653 6488 18000 6490
rect 15653 6432 15658 6488
rect 15714 6432 18000 6488
rect 15653 6430 18000 6432
rect 15653 6427 15719 6430
rect 17520 6400 18000 6430
rect 12198 6292 12204 6356
rect 12268 6354 12274 6356
rect 15745 6354 15811 6357
rect 12268 6352 15811 6354
rect 12268 6296 15750 6352
rect 15806 6296 15811 6352
rect 12268 6294 15811 6296
rect 12268 6292 12274 6294
rect 15745 6291 15811 6294
rect 4797 6218 4863 6221
rect 5441 6218 5507 6221
rect 8293 6218 8359 6221
rect 4797 6216 8359 6218
rect 4797 6160 4802 6216
rect 4858 6160 5446 6216
rect 5502 6160 8298 6216
rect 8354 6160 8359 6216
rect 4797 6158 8359 6160
rect 4797 6155 4863 6158
rect 5441 6155 5507 6158
rect 8293 6155 8359 6158
rect 9121 6218 9187 6221
rect 12985 6218 13051 6221
rect 15745 6218 15811 6221
rect 9121 6216 15811 6218
rect 9121 6160 9126 6216
rect 9182 6160 12990 6216
rect 13046 6160 15750 6216
rect 15806 6160 15811 6216
rect 9121 6158 15811 6160
rect 9121 6155 9187 6158
rect 12985 6155 13051 6158
rect 15745 6155 15811 6158
rect 0 6082 480 6112
rect 3509 6082 3575 6085
rect 0 6080 3575 6082
rect 0 6024 3514 6080
rect 3570 6024 3575 6080
rect 0 6022 3575 6024
rect 0 5992 480 6022
rect 3509 6019 3575 6022
rect 4429 6082 4495 6085
rect 4838 6082 4844 6084
rect 4429 6080 4844 6082
rect 4429 6024 4434 6080
rect 4490 6024 4844 6080
rect 4429 6022 4844 6024
rect 4429 6019 4495 6022
rect 4838 6020 4844 6022
rect 4908 6020 4914 6084
rect 6821 6082 6887 6085
rect 7557 6082 7623 6085
rect 8201 6082 8267 6085
rect 6821 6080 8267 6082
rect 6821 6024 6826 6080
rect 6882 6024 7562 6080
rect 7618 6024 8206 6080
rect 8262 6024 8267 6080
rect 6821 6022 8267 6024
rect 6821 6019 6887 6022
rect 7557 6019 7623 6022
rect 8201 6019 8267 6022
rect 14917 6082 14983 6085
rect 17520 6082 18000 6112
rect 14917 6080 18000 6082
rect 14917 6024 14922 6080
rect 14978 6024 18000 6080
rect 14917 6022 18000 6024
rect 14917 6019 14983 6022
rect 6208 6016 6528 6017
rect 6208 5952 6216 6016
rect 6280 5952 6296 6016
rect 6360 5952 6376 6016
rect 6440 5952 6456 6016
rect 6520 5952 6528 6016
rect 6208 5951 6528 5952
rect 11472 6016 11792 6017
rect 11472 5952 11480 6016
rect 11544 5952 11560 6016
rect 11624 5952 11640 6016
rect 11704 5952 11720 6016
rect 11784 5952 11792 6016
rect 17520 5992 18000 6022
rect 11472 5951 11792 5952
rect 8702 5884 8708 5948
rect 8772 5946 8778 5948
rect 8937 5946 9003 5949
rect 8772 5944 9003 5946
rect 8772 5888 8942 5944
rect 8998 5888 9003 5944
rect 8772 5886 9003 5888
rect 8772 5884 8778 5886
rect 8937 5883 9003 5886
rect 10133 5946 10199 5949
rect 10358 5946 10364 5948
rect 10133 5944 10364 5946
rect 10133 5888 10138 5944
rect 10194 5888 10364 5944
rect 10133 5886 10364 5888
rect 10133 5883 10199 5886
rect 10358 5884 10364 5886
rect 10428 5884 10434 5948
rect 2405 5810 2471 5813
rect 2957 5810 3023 5813
rect 6729 5810 6795 5813
rect 9673 5810 9739 5813
rect 2405 5808 9739 5810
rect 2405 5752 2410 5808
rect 2466 5752 2962 5808
rect 3018 5752 6734 5808
rect 6790 5752 9678 5808
rect 9734 5752 9739 5808
rect 2405 5750 9739 5752
rect 2405 5747 2471 5750
rect 2957 5747 3023 5750
rect 6729 5747 6795 5750
rect 9673 5747 9739 5750
rect 10041 5810 10107 5813
rect 12157 5810 12223 5813
rect 10041 5808 12223 5810
rect 10041 5752 10046 5808
rect 10102 5752 12162 5808
rect 12218 5752 12223 5808
rect 10041 5750 12223 5752
rect 10041 5747 10107 5750
rect 12157 5747 12223 5750
rect 0 5674 480 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 480 5614
rect 1301 5611 1367 5614
rect 6821 5674 6887 5677
rect 9990 5674 9996 5676
rect 6821 5672 9996 5674
rect 6821 5616 6826 5672
rect 6882 5616 9996 5672
rect 6821 5614 9996 5616
rect 6821 5611 6887 5614
rect 9990 5612 9996 5614
rect 10060 5674 10066 5676
rect 11973 5674 12039 5677
rect 10060 5672 12039 5674
rect 10060 5616 11978 5672
rect 12034 5616 12039 5672
rect 10060 5614 12039 5616
rect 10060 5612 10066 5614
rect 11973 5611 12039 5614
rect 12341 5674 12407 5677
rect 17520 5674 18000 5704
rect 12341 5672 18000 5674
rect 12341 5616 12346 5672
rect 12402 5616 18000 5672
rect 12341 5614 18000 5616
rect 12341 5611 12407 5614
rect 17520 5584 18000 5614
rect 10317 5538 10383 5541
rect 11145 5538 11211 5541
rect 10317 5536 11211 5538
rect 10317 5480 10322 5536
rect 10378 5480 11150 5536
rect 11206 5480 11211 5536
rect 10317 5478 11211 5480
rect 10317 5475 10383 5478
rect 11145 5475 11211 5478
rect 3576 5472 3896 5473
rect 3576 5408 3584 5472
rect 3648 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3896 5472
rect 3576 5407 3896 5408
rect 8840 5472 9160 5473
rect 8840 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 9008 5472
rect 9072 5408 9088 5472
rect 9152 5408 9160 5472
rect 8840 5407 9160 5408
rect 14104 5472 14424 5473
rect 14104 5408 14112 5472
rect 14176 5408 14192 5472
rect 14256 5408 14272 5472
rect 14336 5408 14352 5472
rect 14416 5408 14424 5472
rect 14104 5407 14424 5408
rect 3049 5402 3115 5405
rect 614 5400 3115 5402
rect 614 5344 3054 5400
rect 3110 5344 3115 5400
rect 614 5342 3115 5344
rect 0 5266 480 5296
rect 614 5266 674 5342
rect 3049 5339 3115 5342
rect 4337 5402 4403 5405
rect 7925 5402 7991 5405
rect 4337 5400 7991 5402
rect 4337 5344 4342 5400
rect 4398 5344 7930 5400
rect 7986 5344 7991 5400
rect 4337 5342 7991 5344
rect 4337 5339 4403 5342
rect 7925 5339 7991 5342
rect 10409 5402 10475 5405
rect 10409 5400 10978 5402
rect 10409 5344 10414 5400
rect 10470 5344 10978 5400
rect 10409 5342 10978 5344
rect 10409 5339 10475 5342
rect 0 5206 674 5266
rect 4613 5266 4679 5269
rect 5625 5266 5691 5269
rect 8109 5266 8175 5269
rect 9857 5268 9923 5269
rect 9806 5266 9812 5268
rect 4613 5264 8175 5266
rect 4613 5208 4618 5264
rect 4674 5208 5630 5264
rect 5686 5208 8114 5264
rect 8170 5208 8175 5264
rect 4613 5206 8175 5208
rect 9766 5206 9812 5266
rect 9876 5264 9923 5268
rect 9918 5208 9923 5264
rect 0 5176 480 5206
rect 4613 5203 4679 5206
rect 5625 5203 5691 5206
rect 8109 5203 8175 5206
rect 9806 5204 9812 5206
rect 9876 5204 9923 5208
rect 9857 5203 9923 5204
rect 10409 5266 10475 5269
rect 10777 5266 10843 5269
rect 10409 5264 10843 5266
rect 10409 5208 10414 5264
rect 10470 5208 10782 5264
rect 10838 5208 10843 5264
rect 10409 5206 10843 5208
rect 10918 5266 10978 5342
rect 17520 5266 18000 5296
rect 10918 5206 18000 5266
rect 10409 5203 10475 5206
rect 10777 5203 10843 5206
rect 17520 5176 18000 5206
rect 3601 5130 3667 5133
rect 4286 5130 4292 5132
rect 3601 5128 4292 5130
rect 3601 5072 3606 5128
rect 3662 5072 4292 5128
rect 3601 5070 4292 5072
rect 3601 5067 3667 5070
rect 4286 5068 4292 5070
rect 4356 5068 4362 5132
rect 4705 5130 4771 5133
rect 6269 5130 6335 5133
rect 4705 5128 6335 5130
rect 4705 5072 4710 5128
rect 4766 5072 6274 5128
rect 6330 5072 6335 5128
rect 4705 5070 6335 5072
rect 4705 5067 4771 5070
rect 6269 5067 6335 5070
rect 9397 5130 9463 5133
rect 9397 5128 13600 5130
rect 9397 5072 9402 5128
rect 9458 5072 13600 5128
rect 9397 5070 13600 5072
rect 9397 5067 9463 5070
rect 6208 4928 6528 4929
rect 0 4858 480 4888
rect 6208 4864 6216 4928
rect 6280 4864 6296 4928
rect 6360 4864 6376 4928
rect 6440 4864 6456 4928
rect 6520 4864 6528 4928
rect 6208 4863 6528 4864
rect 11472 4928 11792 4929
rect 11472 4864 11480 4928
rect 11544 4864 11560 4928
rect 11624 4864 11640 4928
rect 11704 4864 11720 4928
rect 11784 4864 11792 4928
rect 11472 4863 11792 4864
rect 2865 4858 2931 4861
rect 0 4856 2931 4858
rect 0 4800 2870 4856
rect 2926 4800 2931 4856
rect 0 4798 2931 4800
rect 0 4768 480 4798
rect 2865 4795 2931 4798
rect 11973 4858 12039 4861
rect 12198 4858 12204 4860
rect 11973 4856 12204 4858
rect 11973 4800 11978 4856
rect 12034 4800 12204 4856
rect 11973 4798 12204 4800
rect 11973 4795 12039 4798
rect 12198 4796 12204 4798
rect 12268 4796 12274 4860
rect 13540 4858 13600 5070
rect 17520 4858 18000 4888
rect 13540 4798 18000 4858
rect 17520 4768 18000 4798
rect 12341 4722 12407 4725
rect 14089 4722 14155 4725
rect 12341 4720 14155 4722
rect 12341 4664 12346 4720
rect 12402 4664 14094 4720
rect 14150 4664 14155 4720
rect 12341 4662 14155 4664
rect 12341 4659 12407 4662
rect 14089 4659 14155 4662
rect 12709 4586 12775 4589
rect 15745 4586 15811 4589
rect 12709 4584 15811 4586
rect 12709 4528 12714 4584
rect 12770 4528 15750 4584
rect 15806 4528 15811 4584
rect 12709 4526 15811 4528
rect 12709 4523 12775 4526
rect 15745 4523 15811 4526
rect 0 4450 480 4480
rect 1393 4450 1459 4453
rect 0 4448 1459 4450
rect 0 4392 1398 4448
rect 1454 4392 1459 4448
rect 0 4390 1459 4392
rect 0 4360 480 4390
rect 1393 4387 1459 4390
rect 15009 4450 15075 4453
rect 17520 4450 18000 4480
rect 15009 4448 18000 4450
rect 15009 4392 15014 4448
rect 15070 4392 18000 4448
rect 15009 4390 18000 4392
rect 15009 4387 15075 4390
rect 3576 4384 3896 4385
rect 3576 4320 3584 4384
rect 3648 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3896 4384
rect 3576 4319 3896 4320
rect 8840 4384 9160 4385
rect 8840 4320 8848 4384
rect 8912 4320 8928 4384
rect 8992 4320 9008 4384
rect 9072 4320 9088 4384
rect 9152 4320 9160 4384
rect 8840 4319 9160 4320
rect 14104 4384 14424 4385
rect 14104 4320 14112 4384
rect 14176 4320 14192 4384
rect 14256 4320 14272 4384
rect 14336 4320 14352 4384
rect 14416 4320 14424 4384
rect 17520 4360 18000 4390
rect 14104 4319 14424 4320
rect 8109 4178 8175 4181
rect 8937 4178 9003 4181
rect 8109 4176 9003 4178
rect 8109 4120 8114 4176
rect 8170 4120 8942 4176
rect 8998 4120 9003 4176
rect 8109 4118 9003 4120
rect 8109 4115 8175 4118
rect 8937 4115 9003 4118
rect 9949 4178 10015 4181
rect 11789 4178 11855 4181
rect 15837 4178 15903 4181
rect 9949 4176 15903 4178
rect 9949 4120 9954 4176
rect 10010 4120 11794 4176
rect 11850 4120 15842 4176
rect 15898 4120 15903 4176
rect 9949 4118 15903 4120
rect 9949 4115 10015 4118
rect 11789 4115 11855 4118
rect 15837 4115 15903 4118
rect 0 4042 480 4072
rect 1669 4042 1735 4045
rect 7833 4042 7899 4045
rect 0 4040 1735 4042
rect 0 3984 1674 4040
rect 1730 3984 1735 4040
rect 0 3982 1735 3984
rect 0 3952 480 3982
rect 1669 3979 1735 3982
rect 3742 4040 7899 4042
rect 3742 3984 7838 4040
rect 7894 3984 7899 4040
rect 3742 3982 7899 3984
rect 3601 3770 3667 3773
rect 3742 3770 3802 3982
rect 7833 3979 7899 3982
rect 8293 4042 8359 4045
rect 8937 4042 9003 4045
rect 8293 4040 9003 4042
rect 8293 3984 8298 4040
rect 8354 3984 8942 4040
rect 8998 3984 9003 4040
rect 8293 3982 9003 3984
rect 8293 3979 8359 3982
rect 8937 3979 9003 3982
rect 13537 4042 13603 4045
rect 17520 4042 18000 4072
rect 13537 4040 18000 4042
rect 13537 3984 13542 4040
rect 13598 3984 18000 4040
rect 13537 3982 18000 3984
rect 13537 3979 13603 3982
rect 17520 3952 18000 3982
rect 8845 3906 8911 3909
rect 10409 3906 10475 3909
rect 8845 3904 10475 3906
rect 8845 3848 8850 3904
rect 8906 3848 10414 3904
rect 10470 3848 10475 3904
rect 8845 3846 10475 3848
rect 8845 3843 8911 3846
rect 10409 3843 10475 3846
rect 6208 3840 6528 3841
rect 6208 3776 6216 3840
rect 6280 3776 6296 3840
rect 6360 3776 6376 3840
rect 6440 3776 6456 3840
rect 6520 3776 6528 3840
rect 6208 3775 6528 3776
rect 11472 3840 11792 3841
rect 11472 3776 11480 3840
rect 11544 3776 11560 3840
rect 11624 3776 11640 3840
rect 11704 3776 11720 3840
rect 11784 3776 11792 3840
rect 11472 3775 11792 3776
rect 3601 3768 3802 3770
rect 3601 3712 3606 3768
rect 3662 3712 3802 3768
rect 3601 3710 3802 3712
rect 3601 3707 3667 3710
rect 8518 3708 8524 3772
rect 8588 3770 8594 3772
rect 8845 3770 8911 3773
rect 8588 3768 8911 3770
rect 8588 3712 8850 3768
rect 8906 3712 8911 3768
rect 8588 3710 8911 3712
rect 8588 3708 8594 3710
rect 8845 3707 8911 3710
rect 0 3634 480 3664
rect 3877 3634 3943 3637
rect 0 3632 3943 3634
rect 0 3576 3882 3632
rect 3938 3576 3943 3632
rect 0 3574 3943 3576
rect 0 3544 480 3574
rect 3877 3571 3943 3574
rect 8753 3634 8819 3637
rect 9254 3634 9260 3636
rect 8753 3632 9260 3634
rect 8753 3576 8758 3632
rect 8814 3576 9260 3632
rect 8753 3574 9260 3576
rect 8753 3571 8819 3574
rect 9254 3572 9260 3574
rect 9324 3572 9330 3636
rect 9765 3634 9831 3637
rect 10358 3634 10364 3636
rect 9765 3632 10364 3634
rect 9765 3576 9770 3632
rect 9826 3576 10364 3632
rect 9765 3574 10364 3576
rect 9765 3571 9831 3574
rect 10358 3572 10364 3574
rect 10428 3634 10434 3636
rect 10685 3634 10751 3637
rect 10428 3632 10751 3634
rect 10428 3576 10690 3632
rect 10746 3576 10751 3632
rect 10428 3574 10751 3576
rect 10428 3572 10434 3574
rect 10685 3571 10751 3574
rect 11053 3634 11119 3637
rect 12709 3634 12775 3637
rect 11053 3632 12775 3634
rect 11053 3576 11058 3632
rect 11114 3576 12714 3632
rect 12770 3576 12775 3632
rect 11053 3574 12775 3576
rect 11053 3571 11119 3574
rect 12709 3571 12775 3574
rect 15101 3634 15167 3637
rect 17520 3634 18000 3664
rect 15101 3632 18000 3634
rect 15101 3576 15106 3632
rect 15162 3576 18000 3632
rect 15101 3574 18000 3576
rect 15101 3571 15167 3574
rect 17520 3544 18000 3574
rect 2681 3498 2747 3501
rect 3601 3498 3667 3501
rect 2681 3496 3667 3498
rect 2681 3440 2686 3496
rect 2742 3440 3606 3496
rect 3662 3440 3667 3496
rect 2681 3438 3667 3440
rect 2681 3435 2747 3438
rect 3601 3435 3667 3438
rect 3877 3498 3943 3501
rect 9121 3498 9187 3501
rect 3877 3496 9187 3498
rect 3877 3440 3882 3496
rect 3938 3440 9126 3496
rect 9182 3440 9187 3496
rect 3877 3438 9187 3440
rect 3877 3435 3943 3438
rect 5352 3365 5412 3438
rect 9121 3435 9187 3438
rect 10777 3498 10843 3501
rect 11789 3498 11855 3501
rect 14958 3498 14964 3500
rect 10777 3496 14964 3498
rect 10777 3440 10782 3496
rect 10838 3440 11794 3496
rect 11850 3440 14964 3496
rect 10777 3438 14964 3440
rect 10777 3435 10843 3438
rect 11789 3435 11855 3438
rect 14958 3436 14964 3438
rect 15028 3436 15034 3500
rect 5349 3360 5415 3365
rect 5349 3304 5354 3360
rect 5410 3304 5415 3360
rect 5349 3299 5415 3304
rect 10542 3300 10548 3364
rect 10612 3362 10618 3364
rect 12433 3362 12499 3365
rect 10612 3360 12499 3362
rect 10612 3304 12438 3360
rect 12494 3304 12499 3360
rect 10612 3302 12499 3304
rect 10612 3300 10618 3302
rect 12433 3299 12499 3302
rect 3576 3296 3896 3297
rect 3576 3232 3584 3296
rect 3648 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3896 3296
rect 3576 3231 3896 3232
rect 8840 3296 9160 3297
rect 8840 3232 8848 3296
rect 8912 3232 8928 3296
rect 8992 3232 9008 3296
rect 9072 3232 9088 3296
rect 9152 3232 9160 3296
rect 8840 3231 9160 3232
rect 14104 3296 14424 3297
rect 14104 3232 14112 3296
rect 14176 3232 14192 3296
rect 14256 3232 14272 3296
rect 14336 3232 14352 3296
rect 14416 3232 14424 3296
rect 14104 3231 14424 3232
rect 4889 3226 4955 3229
rect 5993 3226 6059 3229
rect 4889 3224 6059 3226
rect 4889 3168 4894 3224
rect 4950 3168 5998 3224
rect 6054 3168 6059 3224
rect 4889 3166 6059 3168
rect 4889 3163 4955 3166
rect 5993 3163 6059 3166
rect 0 3090 480 3120
rect 4061 3090 4127 3093
rect 0 3088 4127 3090
rect 0 3032 4066 3088
rect 4122 3032 4127 3088
rect 0 3030 4127 3032
rect 0 3000 480 3030
rect 4061 3027 4127 3030
rect 4337 3090 4403 3093
rect 9305 3090 9371 3093
rect 4337 3088 9371 3090
rect 4337 3032 4342 3088
rect 4398 3032 9310 3088
rect 9366 3032 9371 3088
rect 4337 3030 9371 3032
rect 4337 3027 4403 3030
rect 9305 3027 9371 3030
rect 10593 3090 10659 3093
rect 11513 3090 11579 3093
rect 10593 3088 11579 3090
rect 10593 3032 10598 3088
rect 10654 3032 11518 3088
rect 11574 3032 11579 3088
rect 10593 3030 11579 3032
rect 10593 3027 10659 3030
rect 11513 3027 11579 3030
rect 13629 3090 13695 3093
rect 17520 3090 18000 3120
rect 13629 3088 18000 3090
rect 13629 3032 13634 3088
rect 13690 3032 18000 3088
rect 13629 3030 18000 3032
rect 13629 3027 13695 3030
rect 17520 3000 18000 3030
rect 2957 2956 3023 2957
rect 2957 2952 3004 2956
rect 3068 2954 3074 2956
rect 3325 2954 3391 2957
rect 4797 2954 4863 2957
rect 6821 2954 6887 2957
rect 2957 2896 2962 2952
rect 2957 2892 3004 2896
rect 3068 2894 3114 2954
rect 3325 2952 6887 2954
rect 3325 2896 3330 2952
rect 3386 2896 4802 2952
rect 4858 2896 6826 2952
rect 6882 2896 6887 2952
rect 3325 2894 6887 2896
rect 3068 2892 3074 2894
rect 2957 2891 3023 2892
rect 3325 2891 3391 2894
rect 4797 2891 4863 2894
rect 6821 2891 6887 2894
rect 8293 2954 8359 2957
rect 10317 2954 10383 2957
rect 8293 2952 10383 2954
rect 8293 2896 8298 2952
rect 8354 2896 10322 2952
rect 10378 2896 10383 2952
rect 8293 2894 10383 2896
rect 8293 2891 8359 2894
rect 10317 2891 10383 2894
rect 10593 2954 10659 2957
rect 11329 2954 11395 2957
rect 11973 2956 12039 2957
rect 11973 2954 12020 2956
rect 10593 2952 11395 2954
rect 10593 2896 10598 2952
rect 10654 2896 11334 2952
rect 11390 2896 11395 2952
rect 10593 2894 11395 2896
rect 11928 2952 12020 2954
rect 11928 2896 11978 2952
rect 11928 2894 12020 2896
rect 10593 2891 10659 2894
rect 11329 2891 11395 2894
rect 11973 2892 12020 2894
rect 12084 2892 12090 2956
rect 11973 2891 12039 2892
rect 3182 2756 3188 2820
rect 3252 2818 3258 2820
rect 5441 2818 5507 2821
rect 5625 2820 5691 2821
rect 3252 2816 5507 2818
rect 3252 2760 5446 2816
rect 5502 2760 5507 2816
rect 3252 2758 5507 2760
rect 3252 2756 3258 2758
rect 5441 2755 5507 2758
rect 5574 2756 5580 2820
rect 5644 2818 5691 2820
rect 5644 2816 5736 2818
rect 5686 2760 5736 2816
rect 5644 2758 5736 2760
rect 5644 2756 5691 2758
rect 5625 2755 5691 2756
rect 6208 2752 6528 2753
rect 0 2682 480 2712
rect 6208 2688 6216 2752
rect 6280 2688 6296 2752
rect 6360 2688 6376 2752
rect 6440 2688 6456 2752
rect 6520 2688 6528 2752
rect 6208 2687 6528 2688
rect 11472 2752 11792 2753
rect 11472 2688 11480 2752
rect 11544 2688 11560 2752
rect 11624 2688 11640 2752
rect 11704 2688 11720 2752
rect 11784 2688 11792 2752
rect 11472 2687 11792 2688
rect 841 2682 907 2685
rect 0 2680 907 2682
rect 0 2624 846 2680
rect 902 2624 907 2680
rect 0 2622 907 2624
rect 0 2592 480 2622
rect 841 2619 907 2622
rect 7465 2682 7531 2685
rect 7598 2682 7604 2684
rect 7465 2680 7604 2682
rect 7465 2624 7470 2680
rect 7526 2624 7604 2680
rect 7465 2622 7604 2624
rect 7465 2619 7531 2622
rect 7598 2620 7604 2622
rect 7668 2620 7674 2684
rect 9990 2620 9996 2684
rect 10060 2682 10066 2684
rect 11053 2682 11119 2685
rect 10060 2680 11119 2682
rect 10060 2624 11058 2680
rect 11114 2624 11119 2680
rect 10060 2622 11119 2624
rect 10060 2620 10066 2622
rect 11053 2619 11119 2622
rect 16389 2682 16455 2685
rect 17520 2682 18000 2712
rect 16389 2680 18000 2682
rect 16389 2624 16394 2680
rect 16450 2624 18000 2680
rect 16389 2622 18000 2624
rect 16389 2619 16455 2622
rect 17520 2592 18000 2622
rect 2681 2546 2747 2549
rect 6913 2546 6979 2549
rect 2681 2544 6979 2546
rect 2681 2488 2686 2544
rect 2742 2488 6918 2544
rect 6974 2488 6979 2544
rect 2681 2486 6979 2488
rect 2681 2483 2747 2486
rect 6913 2483 6979 2486
rect 10317 2546 10383 2549
rect 11789 2546 11855 2549
rect 10317 2544 11855 2546
rect 10317 2488 10322 2544
rect 10378 2488 11794 2544
rect 11850 2488 11855 2544
rect 10317 2486 11855 2488
rect 10317 2483 10383 2486
rect 11789 2483 11855 2486
rect 13997 2410 14063 2413
rect 13997 2408 14658 2410
rect 13997 2352 14002 2408
rect 14058 2352 14658 2408
rect 13997 2350 14658 2352
rect 13997 2347 14063 2350
rect 0 2274 480 2304
rect 3417 2274 3483 2277
rect 0 2272 3483 2274
rect 0 2216 3422 2272
rect 3478 2216 3483 2272
rect 0 2214 3483 2216
rect 14598 2274 14658 2350
rect 17520 2274 18000 2304
rect 14598 2214 18000 2274
rect 0 2184 480 2214
rect 3417 2211 3483 2214
rect 3576 2208 3896 2209
rect 3576 2144 3584 2208
rect 3648 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3896 2208
rect 3576 2143 3896 2144
rect 8840 2208 9160 2209
rect 8840 2144 8848 2208
rect 8912 2144 8928 2208
rect 8992 2144 9008 2208
rect 9072 2144 9088 2208
rect 9152 2144 9160 2208
rect 8840 2143 9160 2144
rect 14104 2208 14424 2209
rect 14104 2144 14112 2208
rect 14176 2144 14192 2208
rect 14256 2144 14272 2208
rect 14336 2144 14352 2208
rect 14416 2144 14424 2208
rect 17520 2184 18000 2214
rect 14104 2143 14424 2144
rect 0 1866 480 1896
rect 1945 1866 2011 1869
rect 0 1864 2011 1866
rect 0 1808 1950 1864
rect 2006 1808 2011 1864
rect 0 1806 2011 1808
rect 0 1776 480 1806
rect 1945 1803 2011 1806
rect 14733 1866 14799 1869
rect 17520 1866 18000 1896
rect 14733 1864 18000 1866
rect 14733 1808 14738 1864
rect 14794 1808 18000 1864
rect 14733 1806 18000 1808
rect 14733 1803 14799 1806
rect 17520 1776 18000 1806
rect 0 1458 480 1488
rect 3233 1458 3299 1461
rect 0 1456 3299 1458
rect 0 1400 3238 1456
rect 3294 1400 3299 1456
rect 0 1398 3299 1400
rect 0 1368 480 1398
rect 3233 1395 3299 1398
rect 14825 1458 14891 1461
rect 17520 1458 18000 1488
rect 14825 1456 18000 1458
rect 14825 1400 14830 1456
rect 14886 1400 18000 1456
rect 14825 1398 18000 1400
rect 14825 1395 14891 1398
rect 17520 1368 18000 1398
rect 0 1050 480 1080
rect 2497 1050 2563 1053
rect 0 1048 2563 1050
rect 0 992 2502 1048
rect 2558 992 2563 1048
rect 0 990 2563 992
rect 0 960 480 990
rect 2497 987 2563 990
rect 10961 1050 11027 1053
rect 17520 1050 18000 1080
rect 10961 1048 18000 1050
rect 10961 992 10966 1048
rect 11022 992 18000 1048
rect 10961 990 18000 992
rect 10961 987 11027 990
rect 17520 960 18000 990
rect 0 642 480 672
rect 3417 642 3483 645
rect 0 640 3483 642
rect 0 584 3422 640
rect 3478 584 3483 640
rect 0 582 3483 584
rect 0 552 480 582
rect 3417 579 3483 582
rect 15009 642 15075 645
rect 17520 642 18000 672
rect 15009 640 18000 642
rect 15009 584 15014 640
rect 15070 584 18000 640
rect 15009 582 18000 584
rect 15009 579 15075 582
rect 17520 552 18000 582
rect 0 234 480 264
rect 3049 234 3115 237
rect 0 232 3115 234
rect 0 176 3054 232
rect 3110 176 3115 232
rect 0 174 3115 176
rect 0 144 480 174
rect 3049 171 3115 174
rect 15101 234 15167 237
rect 17520 234 18000 264
rect 15101 232 18000 234
rect 15101 176 15106 232
rect 15162 176 18000 232
rect 15101 174 18000 176
rect 15101 171 15167 174
rect 17520 144 18000 174
<< via3 >>
rect 6216 14716 6280 14720
rect 6216 14660 6220 14716
rect 6220 14660 6276 14716
rect 6276 14660 6280 14716
rect 6216 14656 6280 14660
rect 6296 14716 6360 14720
rect 6296 14660 6300 14716
rect 6300 14660 6356 14716
rect 6356 14660 6360 14716
rect 6296 14656 6360 14660
rect 6376 14716 6440 14720
rect 6376 14660 6380 14716
rect 6380 14660 6436 14716
rect 6436 14660 6440 14716
rect 6376 14656 6440 14660
rect 6456 14716 6520 14720
rect 6456 14660 6460 14716
rect 6460 14660 6516 14716
rect 6516 14660 6520 14716
rect 6456 14656 6520 14660
rect 11480 14716 11544 14720
rect 11480 14660 11484 14716
rect 11484 14660 11540 14716
rect 11540 14660 11544 14716
rect 11480 14656 11544 14660
rect 11560 14716 11624 14720
rect 11560 14660 11564 14716
rect 11564 14660 11620 14716
rect 11620 14660 11624 14716
rect 11560 14656 11624 14660
rect 11640 14716 11704 14720
rect 11640 14660 11644 14716
rect 11644 14660 11700 14716
rect 11700 14660 11704 14716
rect 11640 14656 11704 14660
rect 11720 14716 11784 14720
rect 11720 14660 11724 14716
rect 11724 14660 11780 14716
rect 11780 14660 11784 14716
rect 11720 14656 11784 14660
rect 3584 14172 3648 14176
rect 3584 14116 3588 14172
rect 3588 14116 3644 14172
rect 3644 14116 3648 14172
rect 3584 14112 3648 14116
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 8848 14172 8912 14176
rect 8848 14116 8852 14172
rect 8852 14116 8908 14172
rect 8908 14116 8912 14172
rect 8848 14112 8912 14116
rect 8928 14172 8992 14176
rect 8928 14116 8932 14172
rect 8932 14116 8988 14172
rect 8988 14116 8992 14172
rect 8928 14112 8992 14116
rect 9008 14172 9072 14176
rect 9008 14116 9012 14172
rect 9012 14116 9068 14172
rect 9068 14116 9072 14172
rect 9008 14112 9072 14116
rect 9088 14172 9152 14176
rect 9088 14116 9092 14172
rect 9092 14116 9148 14172
rect 9148 14116 9152 14172
rect 9088 14112 9152 14116
rect 14112 14172 14176 14176
rect 14112 14116 14116 14172
rect 14116 14116 14172 14172
rect 14172 14116 14176 14172
rect 14112 14112 14176 14116
rect 14192 14172 14256 14176
rect 14192 14116 14196 14172
rect 14196 14116 14252 14172
rect 14252 14116 14256 14172
rect 14192 14112 14256 14116
rect 14272 14172 14336 14176
rect 14272 14116 14276 14172
rect 14276 14116 14332 14172
rect 14332 14116 14336 14172
rect 14272 14112 14336 14116
rect 14352 14172 14416 14176
rect 14352 14116 14356 14172
rect 14356 14116 14412 14172
rect 14412 14116 14416 14172
rect 14352 14112 14416 14116
rect 6216 13628 6280 13632
rect 6216 13572 6220 13628
rect 6220 13572 6276 13628
rect 6276 13572 6280 13628
rect 6216 13568 6280 13572
rect 6296 13628 6360 13632
rect 6296 13572 6300 13628
rect 6300 13572 6356 13628
rect 6356 13572 6360 13628
rect 6296 13568 6360 13572
rect 6376 13628 6440 13632
rect 6376 13572 6380 13628
rect 6380 13572 6436 13628
rect 6436 13572 6440 13628
rect 6376 13568 6440 13572
rect 6456 13628 6520 13632
rect 6456 13572 6460 13628
rect 6460 13572 6516 13628
rect 6516 13572 6520 13628
rect 6456 13568 6520 13572
rect 11480 13628 11544 13632
rect 11480 13572 11484 13628
rect 11484 13572 11540 13628
rect 11540 13572 11544 13628
rect 11480 13568 11544 13572
rect 11560 13628 11624 13632
rect 11560 13572 11564 13628
rect 11564 13572 11620 13628
rect 11620 13572 11624 13628
rect 11560 13568 11624 13572
rect 11640 13628 11704 13632
rect 11640 13572 11644 13628
rect 11644 13572 11700 13628
rect 11700 13572 11704 13628
rect 11640 13568 11704 13572
rect 11720 13628 11784 13632
rect 11720 13572 11724 13628
rect 11724 13572 11780 13628
rect 11780 13572 11784 13628
rect 11720 13568 11784 13572
rect 3584 13084 3648 13088
rect 3584 13028 3588 13084
rect 3588 13028 3644 13084
rect 3644 13028 3648 13084
rect 3584 13024 3648 13028
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 8848 13084 8912 13088
rect 8848 13028 8852 13084
rect 8852 13028 8908 13084
rect 8908 13028 8912 13084
rect 8848 13024 8912 13028
rect 8928 13084 8992 13088
rect 8928 13028 8932 13084
rect 8932 13028 8988 13084
rect 8988 13028 8992 13084
rect 8928 13024 8992 13028
rect 9008 13084 9072 13088
rect 9008 13028 9012 13084
rect 9012 13028 9068 13084
rect 9068 13028 9072 13084
rect 9008 13024 9072 13028
rect 9088 13084 9152 13088
rect 9088 13028 9092 13084
rect 9092 13028 9148 13084
rect 9148 13028 9152 13084
rect 9088 13024 9152 13028
rect 14112 13084 14176 13088
rect 14112 13028 14116 13084
rect 14116 13028 14172 13084
rect 14172 13028 14176 13084
rect 14112 13024 14176 13028
rect 14192 13084 14256 13088
rect 14192 13028 14196 13084
rect 14196 13028 14252 13084
rect 14252 13028 14256 13084
rect 14192 13024 14256 13028
rect 14272 13084 14336 13088
rect 14272 13028 14276 13084
rect 14276 13028 14332 13084
rect 14332 13028 14336 13084
rect 14272 13024 14336 13028
rect 14352 13084 14416 13088
rect 14352 13028 14356 13084
rect 14356 13028 14412 13084
rect 14412 13028 14416 13084
rect 14352 13024 14416 13028
rect 12756 13016 12820 13020
rect 12756 12960 12806 13016
rect 12806 12960 12820 13016
rect 12756 12956 12820 12960
rect 13676 12548 13740 12612
rect 6216 12540 6280 12544
rect 6216 12484 6220 12540
rect 6220 12484 6276 12540
rect 6276 12484 6280 12540
rect 6216 12480 6280 12484
rect 6296 12540 6360 12544
rect 6296 12484 6300 12540
rect 6300 12484 6356 12540
rect 6356 12484 6360 12540
rect 6296 12480 6360 12484
rect 6376 12540 6440 12544
rect 6376 12484 6380 12540
rect 6380 12484 6436 12540
rect 6436 12484 6440 12540
rect 6376 12480 6440 12484
rect 6456 12540 6520 12544
rect 6456 12484 6460 12540
rect 6460 12484 6516 12540
rect 6516 12484 6520 12540
rect 6456 12480 6520 12484
rect 11480 12540 11544 12544
rect 11480 12484 11484 12540
rect 11484 12484 11540 12540
rect 11540 12484 11544 12540
rect 11480 12480 11544 12484
rect 11560 12540 11624 12544
rect 11560 12484 11564 12540
rect 11564 12484 11620 12540
rect 11620 12484 11624 12540
rect 11560 12480 11624 12484
rect 11640 12540 11704 12544
rect 11640 12484 11644 12540
rect 11644 12484 11700 12540
rect 11700 12484 11704 12540
rect 11640 12480 11704 12484
rect 11720 12540 11784 12544
rect 11720 12484 11724 12540
rect 11724 12484 11780 12540
rect 11780 12484 11784 12540
rect 11720 12480 11784 12484
rect 12020 12276 12084 12340
rect 12756 12336 12820 12340
rect 12756 12280 12806 12336
rect 12806 12280 12820 12336
rect 12756 12276 12820 12280
rect 13860 12336 13924 12340
rect 13860 12280 13910 12336
rect 13910 12280 13924 12336
rect 13860 12276 13924 12280
rect 3584 11996 3648 12000
rect 3584 11940 3588 11996
rect 3588 11940 3644 11996
rect 3644 11940 3648 11996
rect 3584 11936 3648 11940
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 8848 11996 8912 12000
rect 8848 11940 8852 11996
rect 8852 11940 8908 11996
rect 8908 11940 8912 11996
rect 8848 11936 8912 11940
rect 8928 11996 8992 12000
rect 8928 11940 8932 11996
rect 8932 11940 8988 11996
rect 8988 11940 8992 11996
rect 8928 11936 8992 11940
rect 9008 11996 9072 12000
rect 9008 11940 9012 11996
rect 9012 11940 9068 11996
rect 9068 11940 9072 11996
rect 9008 11936 9072 11940
rect 9088 11996 9152 12000
rect 9088 11940 9092 11996
rect 9092 11940 9148 11996
rect 9148 11940 9152 11996
rect 9088 11936 9152 11940
rect 14112 11996 14176 12000
rect 14112 11940 14116 11996
rect 14116 11940 14172 11996
rect 14172 11940 14176 11996
rect 14112 11936 14176 11940
rect 14192 11996 14256 12000
rect 14192 11940 14196 11996
rect 14196 11940 14252 11996
rect 14252 11940 14256 11996
rect 14192 11936 14256 11940
rect 14272 11996 14336 12000
rect 14272 11940 14276 11996
rect 14276 11940 14332 11996
rect 14332 11940 14336 11996
rect 14272 11936 14336 11940
rect 14352 11996 14416 12000
rect 14352 11940 14356 11996
rect 14356 11940 14412 11996
rect 14412 11940 14416 11996
rect 14352 11936 14416 11940
rect 13308 11596 13372 11660
rect 6216 11452 6280 11456
rect 6216 11396 6220 11452
rect 6220 11396 6276 11452
rect 6276 11396 6280 11452
rect 6216 11392 6280 11396
rect 6296 11452 6360 11456
rect 6296 11396 6300 11452
rect 6300 11396 6356 11452
rect 6356 11396 6360 11452
rect 6296 11392 6360 11396
rect 6376 11452 6440 11456
rect 6376 11396 6380 11452
rect 6380 11396 6436 11452
rect 6436 11396 6440 11452
rect 6376 11392 6440 11396
rect 6456 11452 6520 11456
rect 6456 11396 6460 11452
rect 6460 11396 6516 11452
rect 6516 11396 6520 11452
rect 6456 11392 6520 11396
rect 11480 11452 11544 11456
rect 11480 11396 11484 11452
rect 11484 11396 11540 11452
rect 11540 11396 11544 11452
rect 11480 11392 11544 11396
rect 11560 11452 11624 11456
rect 11560 11396 11564 11452
rect 11564 11396 11620 11452
rect 11620 11396 11624 11452
rect 11560 11392 11624 11396
rect 11640 11452 11704 11456
rect 11640 11396 11644 11452
rect 11644 11396 11700 11452
rect 11700 11396 11704 11452
rect 11640 11392 11704 11396
rect 11720 11452 11784 11456
rect 11720 11396 11724 11452
rect 11724 11396 11780 11452
rect 11780 11396 11784 11452
rect 11720 11392 11784 11396
rect 5028 11324 5092 11388
rect 4844 11188 4908 11252
rect 12020 11188 12084 11252
rect 14964 11052 15028 11116
rect 3584 10908 3648 10912
rect 3584 10852 3588 10908
rect 3588 10852 3644 10908
rect 3644 10852 3648 10908
rect 3584 10848 3648 10852
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 8848 10908 8912 10912
rect 8848 10852 8852 10908
rect 8852 10852 8908 10908
rect 8908 10852 8912 10908
rect 8848 10848 8912 10852
rect 8928 10908 8992 10912
rect 8928 10852 8932 10908
rect 8932 10852 8988 10908
rect 8988 10852 8992 10908
rect 8928 10848 8992 10852
rect 9008 10908 9072 10912
rect 9008 10852 9012 10908
rect 9012 10852 9068 10908
rect 9068 10852 9072 10908
rect 9008 10848 9072 10852
rect 9088 10908 9152 10912
rect 9088 10852 9092 10908
rect 9092 10852 9148 10908
rect 9148 10852 9152 10908
rect 9088 10848 9152 10852
rect 14112 10908 14176 10912
rect 14112 10852 14116 10908
rect 14116 10852 14172 10908
rect 14172 10852 14176 10908
rect 14112 10848 14176 10852
rect 14192 10908 14256 10912
rect 14192 10852 14196 10908
rect 14196 10852 14252 10908
rect 14252 10852 14256 10908
rect 14192 10848 14256 10852
rect 14272 10908 14336 10912
rect 14272 10852 14276 10908
rect 14276 10852 14332 10908
rect 14332 10852 14336 10908
rect 14272 10848 14336 10852
rect 14352 10908 14416 10912
rect 14352 10852 14356 10908
rect 14356 10852 14412 10908
rect 14412 10852 14416 10908
rect 14352 10848 14416 10852
rect 10364 10780 10428 10844
rect 6216 10364 6280 10368
rect 6216 10308 6220 10364
rect 6220 10308 6276 10364
rect 6276 10308 6280 10364
rect 6216 10304 6280 10308
rect 6296 10364 6360 10368
rect 6296 10308 6300 10364
rect 6300 10308 6356 10364
rect 6356 10308 6360 10364
rect 6296 10304 6360 10308
rect 6376 10364 6440 10368
rect 6376 10308 6380 10364
rect 6380 10308 6436 10364
rect 6436 10308 6440 10364
rect 6376 10304 6440 10308
rect 6456 10364 6520 10368
rect 6456 10308 6460 10364
rect 6460 10308 6516 10364
rect 6516 10308 6520 10364
rect 6456 10304 6520 10308
rect 11480 10364 11544 10368
rect 11480 10308 11484 10364
rect 11484 10308 11540 10364
rect 11540 10308 11544 10364
rect 11480 10304 11544 10308
rect 11560 10364 11624 10368
rect 11560 10308 11564 10364
rect 11564 10308 11620 10364
rect 11620 10308 11624 10364
rect 11560 10304 11624 10308
rect 11640 10364 11704 10368
rect 11640 10308 11644 10364
rect 11644 10308 11700 10364
rect 11700 10308 11704 10364
rect 11640 10304 11704 10308
rect 11720 10364 11784 10368
rect 11720 10308 11724 10364
rect 11724 10308 11780 10364
rect 11780 10308 11784 10364
rect 11720 10304 11784 10308
rect 3372 10296 3436 10300
rect 3372 10240 3422 10296
rect 3422 10240 3436 10296
rect 3372 10236 3436 10240
rect 9996 10236 10060 10300
rect 11284 10236 11348 10300
rect 4292 9828 4356 9892
rect 5028 9828 5092 9892
rect 13124 9964 13188 10028
rect 13860 9828 13924 9892
rect 3584 9820 3648 9824
rect 3584 9764 3588 9820
rect 3588 9764 3644 9820
rect 3644 9764 3648 9820
rect 3584 9760 3648 9764
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 8848 9820 8912 9824
rect 8848 9764 8852 9820
rect 8852 9764 8908 9820
rect 8908 9764 8912 9820
rect 8848 9760 8912 9764
rect 8928 9820 8992 9824
rect 8928 9764 8932 9820
rect 8932 9764 8988 9820
rect 8988 9764 8992 9820
rect 8928 9760 8992 9764
rect 9008 9820 9072 9824
rect 9008 9764 9012 9820
rect 9012 9764 9068 9820
rect 9068 9764 9072 9820
rect 9008 9760 9072 9764
rect 9088 9820 9152 9824
rect 9088 9764 9092 9820
rect 9092 9764 9148 9820
rect 9148 9764 9152 9820
rect 9088 9760 9152 9764
rect 14112 9820 14176 9824
rect 14112 9764 14116 9820
rect 14116 9764 14172 9820
rect 14172 9764 14176 9820
rect 14112 9760 14176 9764
rect 14192 9820 14256 9824
rect 14192 9764 14196 9820
rect 14196 9764 14252 9820
rect 14252 9764 14256 9820
rect 14192 9760 14256 9764
rect 14272 9820 14336 9824
rect 14272 9764 14276 9820
rect 14276 9764 14332 9820
rect 14332 9764 14336 9820
rect 14272 9760 14336 9764
rect 14352 9820 14416 9824
rect 14352 9764 14356 9820
rect 14356 9764 14412 9820
rect 14412 9764 14416 9820
rect 14352 9760 14416 9764
rect 12388 9692 12452 9756
rect 13308 9692 13372 9756
rect 13676 9556 13740 9620
rect 9260 9420 9324 9484
rect 5580 9284 5644 9348
rect 6216 9276 6280 9280
rect 6216 9220 6220 9276
rect 6220 9220 6276 9276
rect 6276 9220 6280 9276
rect 6216 9216 6280 9220
rect 6296 9276 6360 9280
rect 6296 9220 6300 9276
rect 6300 9220 6356 9276
rect 6356 9220 6360 9276
rect 6296 9216 6360 9220
rect 6376 9276 6440 9280
rect 6376 9220 6380 9276
rect 6380 9220 6436 9276
rect 6436 9220 6440 9276
rect 6376 9216 6440 9220
rect 6456 9276 6520 9280
rect 6456 9220 6460 9276
rect 6460 9220 6516 9276
rect 6516 9220 6520 9276
rect 6456 9216 6520 9220
rect 11480 9276 11544 9280
rect 11480 9220 11484 9276
rect 11484 9220 11540 9276
rect 11540 9220 11544 9276
rect 11480 9216 11544 9220
rect 11560 9276 11624 9280
rect 11560 9220 11564 9276
rect 11564 9220 11620 9276
rect 11620 9220 11624 9276
rect 11560 9216 11624 9220
rect 11640 9276 11704 9280
rect 11640 9220 11644 9276
rect 11644 9220 11700 9276
rect 11700 9220 11704 9276
rect 11640 9216 11704 9220
rect 11720 9276 11784 9280
rect 11720 9220 11724 9276
rect 11724 9220 11780 9276
rect 11780 9220 11784 9276
rect 11720 9216 11784 9220
rect 4108 9148 4172 9212
rect 8708 9148 8772 9212
rect 9444 8800 9508 8804
rect 9444 8744 9494 8800
rect 9494 8744 9508 8800
rect 9444 8740 9508 8744
rect 9812 8740 9876 8804
rect 11284 8800 11348 8804
rect 11284 8744 11334 8800
rect 11334 8744 11348 8800
rect 11284 8740 11348 8744
rect 12204 8740 12268 8804
rect 3584 8732 3648 8736
rect 3584 8676 3588 8732
rect 3588 8676 3644 8732
rect 3644 8676 3648 8732
rect 3584 8672 3648 8676
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 8848 8732 8912 8736
rect 8848 8676 8852 8732
rect 8852 8676 8908 8732
rect 8908 8676 8912 8732
rect 8848 8672 8912 8676
rect 8928 8732 8992 8736
rect 8928 8676 8932 8732
rect 8932 8676 8988 8732
rect 8988 8676 8992 8732
rect 8928 8672 8992 8676
rect 9008 8732 9072 8736
rect 9008 8676 9012 8732
rect 9012 8676 9068 8732
rect 9068 8676 9072 8732
rect 9008 8672 9072 8676
rect 9088 8732 9152 8736
rect 9088 8676 9092 8732
rect 9092 8676 9148 8732
rect 9148 8676 9152 8732
rect 9088 8672 9152 8676
rect 14112 8732 14176 8736
rect 14112 8676 14116 8732
rect 14116 8676 14172 8732
rect 14172 8676 14176 8732
rect 14112 8672 14176 8676
rect 14192 8732 14256 8736
rect 14192 8676 14196 8732
rect 14196 8676 14252 8732
rect 14252 8676 14256 8732
rect 14192 8672 14256 8676
rect 14272 8732 14336 8736
rect 14272 8676 14276 8732
rect 14276 8676 14332 8732
rect 14332 8676 14336 8732
rect 14272 8672 14336 8676
rect 14352 8732 14416 8736
rect 14352 8676 14356 8732
rect 14356 8676 14412 8732
rect 14412 8676 14416 8732
rect 14352 8672 14416 8676
rect 3188 8604 3252 8668
rect 3004 8392 3068 8396
rect 3004 8336 3054 8392
rect 3054 8336 3068 8392
rect 3004 8332 3068 8336
rect 10548 8196 10612 8260
rect 6216 8188 6280 8192
rect 6216 8132 6220 8188
rect 6220 8132 6276 8188
rect 6276 8132 6280 8188
rect 6216 8128 6280 8132
rect 6296 8188 6360 8192
rect 6296 8132 6300 8188
rect 6300 8132 6356 8188
rect 6356 8132 6360 8188
rect 6296 8128 6360 8132
rect 6376 8188 6440 8192
rect 6376 8132 6380 8188
rect 6380 8132 6436 8188
rect 6436 8132 6440 8188
rect 6376 8128 6440 8132
rect 6456 8188 6520 8192
rect 6456 8132 6460 8188
rect 6460 8132 6516 8188
rect 6516 8132 6520 8188
rect 6456 8128 6520 8132
rect 11480 8188 11544 8192
rect 11480 8132 11484 8188
rect 11484 8132 11540 8188
rect 11540 8132 11544 8188
rect 11480 8128 11544 8132
rect 11560 8188 11624 8192
rect 11560 8132 11564 8188
rect 11564 8132 11620 8188
rect 11620 8132 11624 8188
rect 11560 8128 11624 8132
rect 11640 8188 11704 8192
rect 11640 8132 11644 8188
rect 11644 8132 11700 8188
rect 11700 8132 11704 8188
rect 11640 8128 11704 8132
rect 11720 8188 11784 8192
rect 11720 8132 11724 8188
rect 11724 8132 11780 8188
rect 11780 8132 11784 8188
rect 11720 8128 11784 8132
rect 9444 7924 9508 7988
rect 3584 7644 3648 7648
rect 3584 7588 3588 7644
rect 3588 7588 3644 7644
rect 3644 7588 3648 7644
rect 3584 7584 3648 7588
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 9444 7788 9508 7852
rect 8848 7644 8912 7648
rect 8848 7588 8852 7644
rect 8852 7588 8908 7644
rect 8908 7588 8912 7644
rect 8848 7584 8912 7588
rect 8928 7644 8992 7648
rect 8928 7588 8932 7644
rect 8932 7588 8988 7644
rect 8988 7588 8992 7644
rect 8928 7584 8992 7588
rect 9008 7644 9072 7648
rect 9008 7588 9012 7644
rect 9012 7588 9068 7644
rect 9068 7588 9072 7644
rect 9008 7584 9072 7588
rect 9088 7644 9152 7648
rect 9088 7588 9092 7644
rect 9092 7588 9148 7644
rect 9148 7588 9152 7644
rect 9088 7584 9152 7588
rect 14112 7644 14176 7648
rect 14112 7588 14116 7644
rect 14116 7588 14172 7644
rect 14172 7588 14176 7644
rect 14112 7584 14176 7588
rect 14192 7644 14256 7648
rect 14192 7588 14196 7644
rect 14196 7588 14252 7644
rect 14252 7588 14256 7644
rect 14192 7584 14256 7588
rect 14272 7644 14336 7648
rect 14272 7588 14276 7644
rect 14276 7588 14332 7644
rect 14332 7588 14336 7644
rect 14272 7584 14336 7588
rect 14352 7644 14416 7648
rect 14352 7588 14356 7644
rect 14356 7588 14412 7644
rect 14412 7588 14416 7644
rect 14352 7584 14416 7588
rect 9260 7516 9324 7580
rect 9444 7380 9508 7444
rect 9812 7244 9876 7308
rect 6216 7100 6280 7104
rect 6216 7044 6220 7100
rect 6220 7044 6276 7100
rect 6276 7044 6280 7100
rect 6216 7040 6280 7044
rect 6296 7100 6360 7104
rect 6296 7044 6300 7100
rect 6300 7044 6356 7100
rect 6356 7044 6360 7100
rect 6296 7040 6360 7044
rect 6376 7100 6440 7104
rect 6376 7044 6380 7100
rect 6380 7044 6436 7100
rect 6436 7044 6440 7100
rect 6376 7040 6440 7044
rect 6456 7100 6520 7104
rect 6456 7044 6460 7100
rect 6460 7044 6516 7100
rect 6516 7044 6520 7100
rect 6456 7040 6520 7044
rect 11480 7100 11544 7104
rect 11480 7044 11484 7100
rect 11484 7044 11540 7100
rect 11540 7044 11544 7100
rect 11480 7040 11544 7044
rect 11560 7100 11624 7104
rect 11560 7044 11564 7100
rect 11564 7044 11620 7100
rect 11620 7044 11624 7100
rect 11560 7040 11624 7044
rect 11640 7100 11704 7104
rect 11640 7044 11644 7100
rect 11644 7044 11700 7100
rect 11700 7044 11704 7100
rect 11640 7040 11704 7044
rect 11720 7100 11784 7104
rect 11720 7044 11724 7100
rect 11724 7044 11780 7100
rect 11780 7044 11784 7100
rect 11720 7040 11784 7044
rect 8524 6972 8588 7036
rect 3372 6896 3436 6900
rect 3372 6840 3422 6896
rect 3422 6840 3436 6896
rect 3372 6836 3436 6840
rect 7604 6836 7668 6900
rect 4108 6564 4172 6628
rect 3584 6556 3648 6560
rect 3584 6500 3588 6556
rect 3588 6500 3644 6556
rect 3644 6500 3648 6556
rect 3584 6496 3648 6500
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 8848 6556 8912 6560
rect 8848 6500 8852 6556
rect 8852 6500 8908 6556
rect 8908 6500 8912 6556
rect 8848 6496 8912 6500
rect 8928 6556 8992 6560
rect 8928 6500 8932 6556
rect 8932 6500 8988 6556
rect 8988 6500 8992 6556
rect 8928 6496 8992 6500
rect 9008 6556 9072 6560
rect 9008 6500 9012 6556
rect 9012 6500 9068 6556
rect 9068 6500 9072 6556
rect 9008 6496 9072 6500
rect 9088 6556 9152 6560
rect 9088 6500 9092 6556
rect 9092 6500 9148 6556
rect 9148 6500 9152 6556
rect 9088 6496 9152 6500
rect 14112 6556 14176 6560
rect 14112 6500 14116 6556
rect 14116 6500 14172 6556
rect 14172 6500 14176 6556
rect 14112 6496 14176 6500
rect 14192 6556 14256 6560
rect 14192 6500 14196 6556
rect 14196 6500 14252 6556
rect 14252 6500 14256 6556
rect 14192 6496 14256 6500
rect 14272 6556 14336 6560
rect 14272 6500 14276 6556
rect 14276 6500 14332 6556
rect 14332 6500 14336 6556
rect 14272 6496 14336 6500
rect 14352 6556 14416 6560
rect 14352 6500 14356 6556
rect 14356 6500 14412 6556
rect 14412 6500 14416 6556
rect 14352 6496 14416 6500
rect 12204 6292 12268 6356
rect 4844 6020 4908 6084
rect 6216 6012 6280 6016
rect 6216 5956 6220 6012
rect 6220 5956 6276 6012
rect 6276 5956 6280 6012
rect 6216 5952 6280 5956
rect 6296 6012 6360 6016
rect 6296 5956 6300 6012
rect 6300 5956 6356 6012
rect 6356 5956 6360 6012
rect 6296 5952 6360 5956
rect 6376 6012 6440 6016
rect 6376 5956 6380 6012
rect 6380 5956 6436 6012
rect 6436 5956 6440 6012
rect 6376 5952 6440 5956
rect 6456 6012 6520 6016
rect 6456 5956 6460 6012
rect 6460 5956 6516 6012
rect 6516 5956 6520 6012
rect 6456 5952 6520 5956
rect 11480 6012 11544 6016
rect 11480 5956 11484 6012
rect 11484 5956 11540 6012
rect 11540 5956 11544 6012
rect 11480 5952 11544 5956
rect 11560 6012 11624 6016
rect 11560 5956 11564 6012
rect 11564 5956 11620 6012
rect 11620 5956 11624 6012
rect 11560 5952 11624 5956
rect 11640 6012 11704 6016
rect 11640 5956 11644 6012
rect 11644 5956 11700 6012
rect 11700 5956 11704 6012
rect 11640 5952 11704 5956
rect 11720 6012 11784 6016
rect 11720 5956 11724 6012
rect 11724 5956 11780 6012
rect 11780 5956 11784 6012
rect 11720 5952 11784 5956
rect 8708 5884 8772 5948
rect 10364 5884 10428 5948
rect 9996 5612 10060 5676
rect 3584 5468 3648 5472
rect 3584 5412 3588 5468
rect 3588 5412 3644 5468
rect 3644 5412 3648 5468
rect 3584 5408 3648 5412
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 8848 5468 8912 5472
rect 8848 5412 8852 5468
rect 8852 5412 8908 5468
rect 8908 5412 8912 5468
rect 8848 5408 8912 5412
rect 8928 5468 8992 5472
rect 8928 5412 8932 5468
rect 8932 5412 8988 5468
rect 8988 5412 8992 5468
rect 8928 5408 8992 5412
rect 9008 5468 9072 5472
rect 9008 5412 9012 5468
rect 9012 5412 9068 5468
rect 9068 5412 9072 5468
rect 9008 5408 9072 5412
rect 9088 5468 9152 5472
rect 9088 5412 9092 5468
rect 9092 5412 9148 5468
rect 9148 5412 9152 5468
rect 9088 5408 9152 5412
rect 14112 5468 14176 5472
rect 14112 5412 14116 5468
rect 14116 5412 14172 5468
rect 14172 5412 14176 5468
rect 14112 5408 14176 5412
rect 14192 5468 14256 5472
rect 14192 5412 14196 5468
rect 14196 5412 14252 5468
rect 14252 5412 14256 5468
rect 14192 5408 14256 5412
rect 14272 5468 14336 5472
rect 14272 5412 14276 5468
rect 14276 5412 14332 5468
rect 14332 5412 14336 5468
rect 14272 5408 14336 5412
rect 14352 5468 14416 5472
rect 14352 5412 14356 5468
rect 14356 5412 14412 5468
rect 14412 5412 14416 5468
rect 14352 5408 14416 5412
rect 9812 5264 9876 5268
rect 9812 5208 9862 5264
rect 9862 5208 9876 5264
rect 9812 5204 9876 5208
rect 4292 5068 4356 5132
rect 6216 4924 6280 4928
rect 6216 4868 6220 4924
rect 6220 4868 6276 4924
rect 6276 4868 6280 4924
rect 6216 4864 6280 4868
rect 6296 4924 6360 4928
rect 6296 4868 6300 4924
rect 6300 4868 6356 4924
rect 6356 4868 6360 4924
rect 6296 4864 6360 4868
rect 6376 4924 6440 4928
rect 6376 4868 6380 4924
rect 6380 4868 6436 4924
rect 6436 4868 6440 4924
rect 6376 4864 6440 4868
rect 6456 4924 6520 4928
rect 6456 4868 6460 4924
rect 6460 4868 6516 4924
rect 6516 4868 6520 4924
rect 6456 4864 6520 4868
rect 11480 4924 11544 4928
rect 11480 4868 11484 4924
rect 11484 4868 11540 4924
rect 11540 4868 11544 4924
rect 11480 4864 11544 4868
rect 11560 4924 11624 4928
rect 11560 4868 11564 4924
rect 11564 4868 11620 4924
rect 11620 4868 11624 4924
rect 11560 4864 11624 4868
rect 11640 4924 11704 4928
rect 11640 4868 11644 4924
rect 11644 4868 11700 4924
rect 11700 4868 11704 4924
rect 11640 4864 11704 4868
rect 11720 4924 11784 4928
rect 11720 4868 11724 4924
rect 11724 4868 11780 4924
rect 11780 4868 11784 4924
rect 11720 4864 11784 4868
rect 12204 4796 12268 4860
rect 3584 4380 3648 4384
rect 3584 4324 3588 4380
rect 3588 4324 3644 4380
rect 3644 4324 3648 4380
rect 3584 4320 3648 4324
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 8848 4380 8912 4384
rect 8848 4324 8852 4380
rect 8852 4324 8908 4380
rect 8908 4324 8912 4380
rect 8848 4320 8912 4324
rect 8928 4380 8992 4384
rect 8928 4324 8932 4380
rect 8932 4324 8988 4380
rect 8988 4324 8992 4380
rect 8928 4320 8992 4324
rect 9008 4380 9072 4384
rect 9008 4324 9012 4380
rect 9012 4324 9068 4380
rect 9068 4324 9072 4380
rect 9008 4320 9072 4324
rect 9088 4380 9152 4384
rect 9088 4324 9092 4380
rect 9092 4324 9148 4380
rect 9148 4324 9152 4380
rect 9088 4320 9152 4324
rect 14112 4380 14176 4384
rect 14112 4324 14116 4380
rect 14116 4324 14172 4380
rect 14172 4324 14176 4380
rect 14112 4320 14176 4324
rect 14192 4380 14256 4384
rect 14192 4324 14196 4380
rect 14196 4324 14252 4380
rect 14252 4324 14256 4380
rect 14192 4320 14256 4324
rect 14272 4380 14336 4384
rect 14272 4324 14276 4380
rect 14276 4324 14332 4380
rect 14332 4324 14336 4380
rect 14272 4320 14336 4324
rect 14352 4380 14416 4384
rect 14352 4324 14356 4380
rect 14356 4324 14412 4380
rect 14412 4324 14416 4380
rect 14352 4320 14416 4324
rect 6216 3836 6280 3840
rect 6216 3780 6220 3836
rect 6220 3780 6276 3836
rect 6276 3780 6280 3836
rect 6216 3776 6280 3780
rect 6296 3836 6360 3840
rect 6296 3780 6300 3836
rect 6300 3780 6356 3836
rect 6356 3780 6360 3836
rect 6296 3776 6360 3780
rect 6376 3836 6440 3840
rect 6376 3780 6380 3836
rect 6380 3780 6436 3836
rect 6436 3780 6440 3836
rect 6376 3776 6440 3780
rect 6456 3836 6520 3840
rect 6456 3780 6460 3836
rect 6460 3780 6516 3836
rect 6516 3780 6520 3836
rect 6456 3776 6520 3780
rect 11480 3836 11544 3840
rect 11480 3780 11484 3836
rect 11484 3780 11540 3836
rect 11540 3780 11544 3836
rect 11480 3776 11544 3780
rect 11560 3836 11624 3840
rect 11560 3780 11564 3836
rect 11564 3780 11620 3836
rect 11620 3780 11624 3836
rect 11560 3776 11624 3780
rect 11640 3836 11704 3840
rect 11640 3780 11644 3836
rect 11644 3780 11700 3836
rect 11700 3780 11704 3836
rect 11640 3776 11704 3780
rect 11720 3836 11784 3840
rect 11720 3780 11724 3836
rect 11724 3780 11780 3836
rect 11780 3780 11784 3836
rect 11720 3776 11784 3780
rect 8524 3708 8588 3772
rect 9260 3572 9324 3636
rect 10364 3572 10428 3636
rect 14964 3436 15028 3500
rect 10548 3300 10612 3364
rect 3584 3292 3648 3296
rect 3584 3236 3588 3292
rect 3588 3236 3644 3292
rect 3644 3236 3648 3292
rect 3584 3232 3648 3236
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 8848 3292 8912 3296
rect 8848 3236 8852 3292
rect 8852 3236 8908 3292
rect 8908 3236 8912 3292
rect 8848 3232 8912 3236
rect 8928 3292 8992 3296
rect 8928 3236 8932 3292
rect 8932 3236 8988 3292
rect 8988 3236 8992 3292
rect 8928 3232 8992 3236
rect 9008 3292 9072 3296
rect 9008 3236 9012 3292
rect 9012 3236 9068 3292
rect 9068 3236 9072 3292
rect 9008 3232 9072 3236
rect 9088 3292 9152 3296
rect 9088 3236 9092 3292
rect 9092 3236 9148 3292
rect 9148 3236 9152 3292
rect 9088 3232 9152 3236
rect 14112 3292 14176 3296
rect 14112 3236 14116 3292
rect 14116 3236 14172 3292
rect 14172 3236 14176 3292
rect 14112 3232 14176 3236
rect 14192 3292 14256 3296
rect 14192 3236 14196 3292
rect 14196 3236 14252 3292
rect 14252 3236 14256 3292
rect 14192 3232 14256 3236
rect 14272 3292 14336 3296
rect 14272 3236 14276 3292
rect 14276 3236 14332 3292
rect 14332 3236 14336 3292
rect 14272 3232 14336 3236
rect 14352 3292 14416 3296
rect 14352 3236 14356 3292
rect 14356 3236 14412 3292
rect 14412 3236 14416 3292
rect 14352 3232 14416 3236
rect 3004 2952 3068 2956
rect 3004 2896 3018 2952
rect 3018 2896 3068 2952
rect 3004 2892 3068 2896
rect 12020 2952 12084 2956
rect 12020 2896 12034 2952
rect 12034 2896 12084 2952
rect 12020 2892 12084 2896
rect 3188 2756 3252 2820
rect 5580 2816 5644 2820
rect 5580 2760 5630 2816
rect 5630 2760 5644 2816
rect 5580 2756 5644 2760
rect 6216 2748 6280 2752
rect 6216 2692 6220 2748
rect 6220 2692 6276 2748
rect 6276 2692 6280 2748
rect 6216 2688 6280 2692
rect 6296 2748 6360 2752
rect 6296 2692 6300 2748
rect 6300 2692 6356 2748
rect 6356 2692 6360 2748
rect 6296 2688 6360 2692
rect 6376 2748 6440 2752
rect 6376 2692 6380 2748
rect 6380 2692 6436 2748
rect 6436 2692 6440 2748
rect 6376 2688 6440 2692
rect 6456 2748 6520 2752
rect 6456 2692 6460 2748
rect 6460 2692 6516 2748
rect 6516 2692 6520 2748
rect 6456 2688 6520 2692
rect 11480 2748 11544 2752
rect 11480 2692 11484 2748
rect 11484 2692 11540 2748
rect 11540 2692 11544 2748
rect 11480 2688 11544 2692
rect 11560 2748 11624 2752
rect 11560 2692 11564 2748
rect 11564 2692 11620 2748
rect 11620 2692 11624 2748
rect 11560 2688 11624 2692
rect 11640 2748 11704 2752
rect 11640 2692 11644 2748
rect 11644 2692 11700 2748
rect 11700 2692 11704 2748
rect 11640 2688 11704 2692
rect 11720 2748 11784 2752
rect 11720 2692 11724 2748
rect 11724 2692 11780 2748
rect 11780 2692 11784 2748
rect 11720 2688 11784 2692
rect 7604 2620 7668 2684
rect 9996 2620 10060 2684
rect 3584 2204 3648 2208
rect 3584 2148 3588 2204
rect 3588 2148 3644 2204
rect 3644 2148 3648 2204
rect 3584 2144 3648 2148
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 8848 2204 8912 2208
rect 8848 2148 8852 2204
rect 8852 2148 8908 2204
rect 8908 2148 8912 2204
rect 8848 2144 8912 2148
rect 8928 2204 8992 2208
rect 8928 2148 8932 2204
rect 8932 2148 8988 2204
rect 8988 2148 8992 2204
rect 8928 2144 8992 2148
rect 9008 2204 9072 2208
rect 9008 2148 9012 2204
rect 9012 2148 9068 2204
rect 9068 2148 9072 2204
rect 9008 2144 9072 2148
rect 9088 2204 9152 2208
rect 9088 2148 9092 2204
rect 9092 2148 9148 2204
rect 9148 2148 9152 2204
rect 9088 2144 9152 2148
rect 14112 2204 14176 2208
rect 14112 2148 14116 2204
rect 14116 2148 14172 2204
rect 14172 2148 14176 2204
rect 14112 2144 14176 2148
rect 14192 2204 14256 2208
rect 14192 2148 14196 2204
rect 14196 2148 14252 2204
rect 14252 2148 14256 2204
rect 14192 2144 14256 2148
rect 14272 2204 14336 2208
rect 14272 2148 14276 2204
rect 14276 2148 14332 2204
rect 14332 2148 14336 2204
rect 14272 2144 14336 2148
rect 14352 2204 14416 2208
rect 14352 2148 14356 2204
rect 14356 2148 14412 2204
rect 14412 2148 14416 2204
rect 14352 2144 14416 2148
<< metal4 >>
rect 3576 14176 3896 14736
rect 3576 14112 3584 14176
rect 3648 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3896 14176
rect 3576 13088 3896 14112
rect 3576 13024 3584 13088
rect 3648 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3896 13088
rect 3576 12000 3896 13024
rect 3576 11936 3584 12000
rect 3648 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3896 12000
rect 3576 10912 3896 11936
rect 6208 14720 6528 14736
rect 6208 14656 6216 14720
rect 6280 14656 6296 14720
rect 6360 14656 6376 14720
rect 6440 14656 6456 14720
rect 6520 14656 6528 14720
rect 6208 13632 6528 14656
rect 6208 13568 6216 13632
rect 6280 13568 6296 13632
rect 6360 13568 6376 13632
rect 6440 13568 6456 13632
rect 6520 13568 6528 13632
rect 6208 12544 6528 13568
rect 6208 12480 6216 12544
rect 6280 12480 6296 12544
rect 6360 12480 6376 12544
rect 6440 12480 6456 12544
rect 6520 12480 6528 12544
rect 6208 11456 6528 12480
rect 6208 11392 6216 11456
rect 6280 11392 6296 11456
rect 6360 11392 6376 11456
rect 6440 11392 6456 11456
rect 6520 11392 6528 11456
rect 5027 11388 5093 11389
rect 5027 11324 5028 11388
rect 5092 11324 5093 11388
rect 5027 11323 5093 11324
rect 4843 11252 4909 11253
rect 4843 11188 4844 11252
rect 4908 11188 4909 11252
rect 4843 11187 4909 11188
rect 3576 10848 3584 10912
rect 3648 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3896 10912
rect 3371 10300 3437 10301
rect 3371 10236 3372 10300
rect 3436 10236 3437 10300
rect 3371 10235 3437 10236
rect 3187 8668 3253 8669
rect 3187 8604 3188 8668
rect 3252 8604 3253 8668
rect 3187 8603 3253 8604
rect 3003 8396 3069 8397
rect 3003 8332 3004 8396
rect 3068 8332 3069 8396
rect 3003 8331 3069 8332
rect 3006 2957 3066 8331
rect 3003 2956 3069 2957
rect 3003 2892 3004 2956
rect 3068 2892 3069 2956
rect 3003 2891 3069 2892
rect 3190 2821 3250 8603
rect 3374 6901 3434 10235
rect 3576 9824 3896 10848
rect 4291 9892 4357 9893
rect 4291 9828 4292 9892
rect 4356 9828 4357 9892
rect 4291 9827 4357 9828
rect 3576 9760 3584 9824
rect 3648 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3896 9824
rect 3576 8736 3896 9760
rect 4107 9212 4173 9213
rect 4107 9148 4108 9212
rect 4172 9148 4173 9212
rect 4107 9147 4173 9148
rect 3576 8672 3584 8736
rect 3648 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3896 8736
rect 3576 7648 3896 8672
rect 3576 7584 3584 7648
rect 3648 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3896 7648
rect 3371 6900 3437 6901
rect 3371 6836 3372 6900
rect 3436 6836 3437 6900
rect 3371 6835 3437 6836
rect 3576 6560 3896 7584
rect 4110 6629 4170 9147
rect 4107 6628 4173 6629
rect 4107 6564 4108 6628
rect 4172 6564 4173 6628
rect 4107 6563 4173 6564
rect 3576 6496 3584 6560
rect 3648 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3896 6560
rect 3576 5472 3896 6496
rect 3576 5408 3584 5472
rect 3648 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3896 5472
rect 3576 4384 3896 5408
rect 4294 5133 4354 9827
rect 4846 6085 4906 11187
rect 5030 9893 5090 11323
rect 6208 10368 6528 11392
rect 6208 10304 6216 10368
rect 6280 10304 6296 10368
rect 6360 10304 6376 10368
rect 6440 10304 6456 10368
rect 6520 10304 6528 10368
rect 5027 9892 5093 9893
rect 5027 9828 5028 9892
rect 5092 9828 5093 9892
rect 5027 9827 5093 9828
rect 5579 9348 5645 9349
rect 5579 9284 5580 9348
rect 5644 9284 5645 9348
rect 5579 9283 5645 9284
rect 4843 6084 4909 6085
rect 4843 6020 4844 6084
rect 4908 6020 4909 6084
rect 4843 6019 4909 6020
rect 4291 5132 4357 5133
rect 4291 5068 4292 5132
rect 4356 5068 4357 5132
rect 4291 5067 4357 5068
rect 3576 4320 3584 4384
rect 3648 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3896 4384
rect 3576 3296 3896 4320
rect 3576 3232 3584 3296
rect 3648 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3896 3296
rect 3187 2820 3253 2821
rect 3187 2756 3188 2820
rect 3252 2756 3253 2820
rect 3187 2755 3253 2756
rect 3576 2208 3896 3232
rect 5582 2821 5642 9283
rect 6208 9280 6528 10304
rect 6208 9216 6216 9280
rect 6280 9216 6296 9280
rect 6360 9216 6376 9280
rect 6440 9216 6456 9280
rect 6520 9216 6528 9280
rect 6208 8192 6528 9216
rect 8840 14176 9160 14736
rect 8840 14112 8848 14176
rect 8912 14112 8928 14176
rect 8992 14112 9008 14176
rect 9072 14112 9088 14176
rect 9152 14112 9160 14176
rect 8840 13088 9160 14112
rect 8840 13024 8848 13088
rect 8912 13024 8928 13088
rect 8992 13024 9008 13088
rect 9072 13024 9088 13088
rect 9152 13024 9160 13088
rect 8840 12000 9160 13024
rect 8840 11936 8848 12000
rect 8912 11936 8928 12000
rect 8992 11936 9008 12000
rect 9072 11936 9088 12000
rect 9152 11936 9160 12000
rect 8840 10912 9160 11936
rect 8840 10848 8848 10912
rect 8912 10848 8928 10912
rect 8992 10848 9008 10912
rect 9072 10848 9088 10912
rect 9152 10848 9160 10912
rect 8840 9824 9160 10848
rect 11472 14720 11792 14736
rect 11472 14656 11480 14720
rect 11544 14656 11560 14720
rect 11624 14656 11640 14720
rect 11704 14656 11720 14720
rect 11784 14656 11792 14720
rect 11472 13632 11792 14656
rect 11472 13568 11480 13632
rect 11544 13568 11560 13632
rect 11624 13568 11640 13632
rect 11704 13568 11720 13632
rect 11784 13568 11792 13632
rect 11472 12544 11792 13568
rect 14104 14176 14424 14736
rect 14104 14112 14112 14176
rect 14176 14112 14192 14176
rect 14256 14112 14272 14176
rect 14336 14112 14352 14176
rect 14416 14112 14424 14176
rect 14104 13088 14424 14112
rect 14104 13024 14112 13088
rect 14176 13024 14192 13088
rect 14256 13024 14272 13088
rect 14336 13024 14352 13088
rect 14416 13024 14424 13088
rect 12755 13020 12821 13021
rect 12755 12956 12756 13020
rect 12820 12956 12821 13020
rect 12755 12955 12821 12956
rect 11472 12480 11480 12544
rect 11544 12480 11560 12544
rect 11624 12480 11640 12544
rect 11704 12480 11720 12544
rect 11784 12480 11792 12544
rect 11472 11456 11792 12480
rect 12758 12341 12818 12955
rect 13675 12612 13741 12613
rect 13675 12548 13676 12612
rect 13740 12548 13741 12612
rect 13675 12547 13741 12548
rect 12019 12340 12085 12341
rect 12019 12276 12020 12340
rect 12084 12276 12085 12340
rect 12019 12275 12085 12276
rect 12755 12340 12821 12341
rect 12755 12276 12756 12340
rect 12820 12276 12821 12340
rect 12755 12275 12821 12276
rect 11472 11392 11480 11456
rect 11544 11392 11560 11456
rect 11624 11392 11640 11456
rect 11704 11392 11720 11456
rect 11784 11392 11792 11456
rect 10363 10844 10429 10845
rect 10363 10780 10364 10844
rect 10428 10780 10429 10844
rect 10363 10779 10429 10780
rect 9995 10300 10061 10301
rect 9995 10236 9996 10300
rect 10060 10236 10061 10300
rect 9995 10235 10061 10236
rect 8840 9760 8848 9824
rect 8912 9760 8928 9824
rect 8992 9760 9008 9824
rect 9072 9760 9088 9824
rect 9152 9760 9160 9824
rect 8707 9212 8773 9213
rect 8707 9148 8708 9212
rect 8772 9148 8773 9212
rect 8707 9147 8773 9148
rect 6208 8128 6216 8192
rect 6280 8128 6296 8192
rect 6360 8128 6376 8192
rect 6440 8128 6456 8192
rect 6520 8128 6528 8192
rect 6208 7104 6528 8128
rect 6208 7040 6216 7104
rect 6280 7040 6296 7104
rect 6360 7040 6376 7104
rect 6440 7040 6456 7104
rect 6520 7040 6528 7104
rect 6208 6016 6528 7040
rect 8523 7036 8589 7037
rect 8523 6972 8524 7036
rect 8588 6972 8589 7036
rect 8523 6971 8589 6972
rect 7603 6900 7669 6901
rect 7603 6836 7604 6900
rect 7668 6836 7669 6900
rect 7603 6835 7669 6836
rect 6208 5952 6216 6016
rect 6280 5952 6296 6016
rect 6360 5952 6376 6016
rect 6440 5952 6456 6016
rect 6520 5952 6528 6016
rect 6208 4928 6528 5952
rect 6208 4864 6216 4928
rect 6280 4864 6296 4928
rect 6360 4864 6376 4928
rect 6440 4864 6456 4928
rect 6520 4864 6528 4928
rect 6208 3840 6528 4864
rect 6208 3776 6216 3840
rect 6280 3776 6296 3840
rect 6360 3776 6376 3840
rect 6440 3776 6456 3840
rect 6520 3776 6528 3840
rect 5579 2820 5645 2821
rect 5579 2756 5580 2820
rect 5644 2756 5645 2820
rect 5579 2755 5645 2756
rect 3576 2144 3584 2208
rect 3648 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3896 2208
rect 3576 2128 3896 2144
rect 6208 2752 6528 3776
rect 6208 2688 6216 2752
rect 6280 2688 6296 2752
rect 6360 2688 6376 2752
rect 6440 2688 6456 2752
rect 6520 2688 6528 2752
rect 6208 2128 6528 2688
rect 7606 2685 7666 6835
rect 8526 3773 8586 6971
rect 8710 5949 8770 9147
rect 8840 8736 9160 9760
rect 9259 9484 9325 9485
rect 9259 9420 9260 9484
rect 9324 9420 9325 9484
rect 9259 9419 9325 9420
rect 8840 8672 8848 8736
rect 8912 8672 8928 8736
rect 8992 8672 9008 8736
rect 9072 8672 9088 8736
rect 9152 8672 9160 8736
rect 8840 7648 9160 8672
rect 8840 7584 8848 7648
rect 8912 7584 8928 7648
rect 8992 7584 9008 7648
rect 9072 7584 9088 7648
rect 9152 7584 9160 7648
rect 8840 6560 9160 7584
rect 9262 7581 9322 9419
rect 9443 8804 9509 8805
rect 9443 8740 9444 8804
rect 9508 8740 9509 8804
rect 9443 8739 9509 8740
rect 9811 8804 9877 8805
rect 9811 8740 9812 8804
rect 9876 8740 9877 8804
rect 9811 8739 9877 8740
rect 9446 7989 9506 8739
rect 9443 7988 9509 7989
rect 9443 7924 9444 7988
rect 9508 7924 9509 7988
rect 9443 7923 9509 7924
rect 9443 7852 9509 7853
rect 9443 7788 9444 7852
rect 9508 7788 9509 7852
rect 9443 7787 9509 7788
rect 9259 7580 9325 7581
rect 9259 7516 9260 7580
rect 9324 7516 9325 7580
rect 9259 7515 9325 7516
rect 8840 6496 8848 6560
rect 8912 6496 8928 6560
rect 8992 6496 9008 6560
rect 9072 6496 9088 6560
rect 9152 6496 9160 6560
rect 8707 5948 8773 5949
rect 8707 5884 8708 5948
rect 8772 5884 8773 5948
rect 8707 5883 8773 5884
rect 8840 5472 9160 6496
rect 8840 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 9008 5472
rect 9072 5408 9088 5472
rect 9152 5408 9160 5472
rect 8840 4384 9160 5408
rect 8840 4320 8848 4384
rect 8912 4320 8928 4384
rect 8992 4320 9008 4384
rect 9072 4320 9088 4384
rect 9152 4320 9160 4384
rect 8523 3772 8589 3773
rect 8523 3708 8524 3772
rect 8588 3708 8589 3772
rect 8523 3707 8589 3708
rect 8840 3296 9160 4320
rect 9262 3637 9322 7515
rect 9446 7445 9506 7787
rect 9443 7444 9509 7445
rect 9443 7380 9444 7444
rect 9508 7380 9509 7444
rect 9443 7379 9509 7380
rect 9814 7309 9874 8739
rect 9811 7308 9877 7309
rect 9811 7244 9812 7308
rect 9876 7244 9877 7308
rect 9811 7243 9877 7244
rect 9814 5269 9874 7243
rect 9998 5677 10058 10235
rect 10366 5949 10426 10779
rect 11472 10368 11792 11392
rect 12022 11253 12082 12275
rect 13307 11660 13373 11661
rect 13307 11596 13308 11660
rect 13372 11596 13373 11660
rect 13307 11595 13373 11596
rect 12019 11252 12085 11253
rect 12019 11188 12020 11252
rect 12084 11188 12085 11252
rect 12019 11187 12085 11188
rect 11472 10304 11480 10368
rect 11544 10304 11560 10368
rect 11624 10304 11640 10368
rect 11704 10304 11720 10368
rect 11784 10304 11792 10368
rect 11283 10300 11349 10301
rect 11283 10236 11284 10300
rect 11348 10236 11349 10300
rect 11283 10235 11349 10236
rect 11286 8805 11346 10235
rect 11472 9280 11792 10304
rect 11472 9216 11480 9280
rect 11544 9216 11560 9280
rect 11624 9216 11640 9280
rect 11704 9216 11720 9280
rect 11784 9216 11792 9280
rect 11283 8804 11349 8805
rect 11283 8740 11284 8804
rect 11348 8740 11349 8804
rect 11283 8739 11349 8740
rect 10547 8260 10613 8261
rect 10547 8196 10548 8260
rect 10612 8196 10613 8260
rect 10547 8195 10613 8196
rect 10363 5948 10429 5949
rect 10363 5884 10364 5948
rect 10428 5884 10429 5948
rect 10363 5883 10429 5884
rect 9995 5676 10061 5677
rect 9995 5612 9996 5676
rect 10060 5612 10061 5676
rect 9995 5611 10061 5612
rect 9811 5268 9877 5269
rect 9811 5204 9812 5268
rect 9876 5204 9877 5268
rect 9811 5203 9877 5204
rect 9259 3636 9325 3637
rect 9259 3572 9260 3636
rect 9324 3572 9325 3636
rect 9259 3571 9325 3572
rect 8840 3232 8848 3296
rect 8912 3232 8928 3296
rect 8992 3232 9008 3296
rect 9072 3232 9088 3296
rect 9152 3232 9160 3296
rect 7603 2684 7669 2685
rect 7603 2620 7604 2684
rect 7668 2620 7669 2684
rect 7603 2619 7669 2620
rect 8840 2208 9160 3232
rect 9998 2685 10058 5611
rect 10366 3637 10426 5883
rect 10363 3636 10429 3637
rect 10363 3572 10364 3636
rect 10428 3572 10429 3636
rect 10363 3571 10429 3572
rect 10550 3365 10610 8195
rect 11472 8192 11792 9216
rect 11472 8128 11480 8192
rect 11544 8128 11560 8192
rect 11624 8128 11640 8192
rect 11704 8128 11720 8192
rect 11784 8128 11792 8192
rect 11472 7104 11792 8128
rect 11472 7040 11480 7104
rect 11544 7040 11560 7104
rect 11624 7040 11640 7104
rect 11704 7040 11720 7104
rect 11784 7040 11792 7104
rect 11472 6016 11792 7040
rect 11472 5952 11480 6016
rect 11544 5952 11560 6016
rect 11624 5952 11640 6016
rect 11704 5952 11720 6016
rect 11784 5952 11792 6016
rect 11472 4928 11792 5952
rect 11472 4864 11480 4928
rect 11544 4864 11560 4928
rect 11624 4864 11640 4928
rect 11704 4864 11720 4928
rect 11784 4864 11792 4928
rect 11472 3840 11792 4864
rect 11472 3776 11480 3840
rect 11544 3776 11560 3840
rect 11624 3776 11640 3840
rect 11704 3776 11720 3840
rect 11784 3776 11792 3840
rect 10547 3364 10613 3365
rect 10547 3300 10548 3364
rect 10612 3300 10613 3364
rect 10547 3299 10613 3300
rect 11472 2752 11792 3776
rect 12022 2957 12082 11187
rect 13123 10028 13189 10029
rect 13123 9964 13124 10028
rect 13188 9964 13189 10028
rect 13123 9963 13189 9964
rect 12387 9756 12453 9757
rect 12387 9692 12388 9756
rect 12452 9754 12453 9756
rect 13126 9754 13186 9963
rect 13310 9757 13370 11595
rect 12452 9694 13186 9754
rect 13307 9756 13373 9757
rect 12452 9692 12453 9694
rect 12387 9691 12453 9692
rect 13307 9692 13308 9756
rect 13372 9692 13373 9756
rect 13307 9691 13373 9692
rect 13678 9621 13738 12547
rect 13859 12340 13925 12341
rect 13859 12276 13860 12340
rect 13924 12276 13925 12340
rect 13859 12275 13925 12276
rect 13862 9893 13922 12275
rect 14104 12000 14424 13024
rect 14104 11936 14112 12000
rect 14176 11936 14192 12000
rect 14256 11936 14272 12000
rect 14336 11936 14352 12000
rect 14416 11936 14424 12000
rect 14104 10912 14424 11936
rect 14963 11116 15029 11117
rect 14963 11052 14964 11116
rect 15028 11052 15029 11116
rect 14963 11051 15029 11052
rect 14104 10848 14112 10912
rect 14176 10848 14192 10912
rect 14256 10848 14272 10912
rect 14336 10848 14352 10912
rect 14416 10848 14424 10912
rect 13859 9892 13925 9893
rect 13859 9828 13860 9892
rect 13924 9828 13925 9892
rect 13859 9827 13925 9828
rect 14104 9824 14424 10848
rect 14104 9760 14112 9824
rect 14176 9760 14192 9824
rect 14256 9760 14272 9824
rect 14336 9760 14352 9824
rect 14416 9760 14424 9824
rect 13675 9620 13741 9621
rect 13675 9556 13676 9620
rect 13740 9556 13741 9620
rect 13675 9555 13741 9556
rect 12203 8804 12269 8805
rect 12203 8740 12204 8804
rect 12268 8740 12269 8804
rect 12203 8739 12269 8740
rect 12206 6357 12266 8739
rect 14104 8736 14424 9760
rect 14104 8672 14112 8736
rect 14176 8672 14192 8736
rect 14256 8672 14272 8736
rect 14336 8672 14352 8736
rect 14416 8672 14424 8736
rect 14104 7648 14424 8672
rect 14104 7584 14112 7648
rect 14176 7584 14192 7648
rect 14256 7584 14272 7648
rect 14336 7584 14352 7648
rect 14416 7584 14424 7648
rect 14104 6560 14424 7584
rect 14104 6496 14112 6560
rect 14176 6496 14192 6560
rect 14256 6496 14272 6560
rect 14336 6496 14352 6560
rect 14416 6496 14424 6560
rect 12203 6356 12269 6357
rect 12203 6292 12204 6356
rect 12268 6292 12269 6356
rect 12203 6291 12269 6292
rect 12206 4861 12266 6291
rect 14104 5472 14424 6496
rect 14104 5408 14112 5472
rect 14176 5408 14192 5472
rect 14256 5408 14272 5472
rect 14336 5408 14352 5472
rect 14416 5408 14424 5472
rect 12203 4860 12269 4861
rect 12203 4796 12204 4860
rect 12268 4796 12269 4860
rect 12203 4795 12269 4796
rect 14104 4384 14424 5408
rect 14104 4320 14112 4384
rect 14176 4320 14192 4384
rect 14256 4320 14272 4384
rect 14336 4320 14352 4384
rect 14416 4320 14424 4384
rect 14104 3296 14424 4320
rect 14966 3501 15026 11051
rect 14963 3500 15029 3501
rect 14963 3436 14964 3500
rect 15028 3436 15029 3500
rect 14963 3435 15029 3436
rect 14104 3232 14112 3296
rect 14176 3232 14192 3296
rect 14256 3232 14272 3296
rect 14336 3232 14352 3296
rect 14416 3232 14424 3296
rect 12019 2956 12085 2957
rect 12019 2892 12020 2956
rect 12084 2892 12085 2956
rect 12019 2891 12085 2892
rect 11472 2688 11480 2752
rect 11544 2688 11560 2752
rect 11624 2688 11640 2752
rect 11704 2688 11720 2752
rect 11784 2688 11792 2752
rect 9995 2684 10061 2685
rect 9995 2620 9996 2684
rect 10060 2620 10061 2684
rect 9995 2619 10061 2620
rect 8840 2144 8848 2208
rect 8912 2144 8928 2208
rect 8992 2144 9008 2208
rect 9072 2144 9088 2208
rect 9152 2144 9160 2208
rect 8840 2128 9160 2144
rect 11472 2128 11792 2688
rect 14104 2208 14424 3232
rect 14104 2144 14112 2208
rect 14176 2144 14192 2208
rect 14256 2144 14272 2208
rect 14336 2144 14352 2208
rect 14416 2144 14424 2208
rect 14104 2128 14424 2144
use sky130_fd_sc_hd__fill_1  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1472 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1472 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_10 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1605641404
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10
timestamp 1605641404
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2208 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2208 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4416 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4232 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 3220 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1605641404
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_21
timestamp 1605641404
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_32
timestamp 1605641404
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_43
timestamp 1605641404
transform 1 0 5060 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45
timestamp 1605641404
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 5428 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5428 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1605641404
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56
timestamp 1605641404
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _31_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 7268 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1605641404
transform 1 0 8280 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1605641404
transform 1 0 7084 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74
timestamp 1605641404
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_65
timestamp 1605641404
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1605641404
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_87
timestamp 1605641404
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1605641404
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1605641404
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1605641404
transform 1 0 9292 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _52_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 9108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_98
timestamp 1605641404
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1605641404
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1605641404
transform 1 0 10304 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_109
timestamp 1605641404
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1605641404
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1605641404
transform 1 0 11316 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1605641404
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1605641404
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13708 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14352 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13616 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1605641404
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_142
timestamp 1605641404
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1605641404
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_136
timestamp 1605641404
transform 1 0 13616 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1605641404
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1605641404
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14720 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1605641404
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1605641404
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15456 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1605641404
transform 1 0 16008 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1605641404
transform 1 0 16008 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 16836 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 16836 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1472 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2300 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_10
timestamp 1605641404
transform 1 0 2024 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1605641404
transform 1 0 3312 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1605641404
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1605641404
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1605641404
transform 1 0 6716 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5704 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_48
timestamp 1605641404
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59
timestamp 1605641404
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1605641404
transform 1 0 7728 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 8372 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_70
timestamp 1605641404
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_76
timestamp 1605641404
transform 1 0 8096 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1605641404
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_102
timestamp 1605641404
transform 1 0 10488 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1605641404
transform 1 0 10764 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12328 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1605641404
transform 1 0 11132 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 12144 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_118
timestamp 1605641404
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13800 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_2_131
timestamp 1605641404
transform 1 0 13156 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_137
timestamp 1605641404
transform 1 0 13708 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1605641404
transform 1 0 16008 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_147
timestamp 1605641404
transform 1 0 14628 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_160
timestamp 1605641404
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1605641404
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 16836 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2392 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_12
timestamp 1605641404
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4048 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_30
timestamp 1605641404
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_41
timestamp 1605641404
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1605641404
transform 1 0 6072 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5060 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_52
timestamp 1605641404
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1605641404
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8464 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1605641404
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 10580 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 9476 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1605641404
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_100
timestamp 1605641404
transform 1 0 10304 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1605641404
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14076 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_139
timestamp 1605641404
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15732 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1605641404
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1605641404
transform 1 0 16284 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 16836 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1472 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_20
timestamp 1605641404
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3220 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1605641404
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5704 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_48
timestamp 1605641404
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7360 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1605641404
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 8832 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 10028 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1605641404
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1605641404
transform 1 0 12144 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11040 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_106
timestamp 1605641404
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_117
timestamp 1605641404
transform 1 0 11868 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1605641404
transform 1 0 14168 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1605641404
transform 1 0 13156 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_129
timestamp 1605641404
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_140
timestamp 1605641404
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1605641404
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_163
timestamp 1605641404
transform 1 0 16100 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 16836 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_167
timestamp 1605641404
transform 1 0 16468 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 2116 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_9
timestamp 1605641404
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_20
timestamp 1605641404
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 3128 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1605641404
transform 1 0 4140 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_31
timestamp 1605641404
transform 1 0 3956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1605641404
transform 1 0 6164 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1605641404
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_42
timestamp 1605641404
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1605641404
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1605641404
transform 1 0 8556 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_77
timestamp 1605641404
transform 1 0 8188 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9568 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_90
timestamp 1605641404
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1605641404
transform 1 0 11224 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_108
timestamp 1605641404
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp 1605641404
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1605641404
transform 1 0 14260 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1605641404
transform 1 0 13892 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 14812 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_147
timestamp 1605641404
transform 1 0 14628 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1605641404
transform 1 0 16284 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 16836 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1605641404
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_8
timestamp 1605641404
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1605641404
transform 1 0 1840 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1605641404
transform 1 0 1472 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_17
timestamp 1605641404
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 2024 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2852 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4508 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4140 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1605641404
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp 1605641404
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1605641404
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_42
timestamp 1605641404
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1605641404
transform 1 0 5704 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1605641404
transform 1 0 5152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1605641404
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_53
timestamp 1605641404
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1605641404
transform 1 0 6164 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5980 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8096 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1605641404
transform 1 0 7084 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1605641404
transform 1 0 7728 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_6_69
timestamp 1605641404
transform 1 0 7452 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp 1605641404
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1605641404
transform 1 0 9752 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10212 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10028 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1605641404
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1605641404
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_97
timestamp 1605641404
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_106
timestamp 1605641404
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11040 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1605641404
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_115
timestamp 1605641404
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_117
timestamp 1605641404
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12052 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1605641404
transform 1 0 11868 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12512 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13064 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1605641404
transform 1 0 13616 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1605641404
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_133
timestamp 1605641404
transform 1 0 13340 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1605641404
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1605641404
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14812 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1605641404
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1605641404
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1605641404
transform 1 0 16100 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1605641404
transform 1 0 16284 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 16836 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 16836 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_167
timestamp 1605641404
transform 1 0 16468 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1605641404
transform 1 0 1472 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1605641404
transform 1 0 2024 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_8
timestamp 1605641404
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_19
timestamp 1605641404
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1605641404
transform 1 0 3036 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1605641404
transform 1 0 3404 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1605641404
transform 1 0 4876 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5244 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_61
timestamp 1605641404
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6900 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1605641404
transform 1 0 8372 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1605641404
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 11592 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 11316 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1605641404
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1605641404
transform 1 0 13616 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1605641404
transform 1 0 13248 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_130
timestamp 1605641404
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_135
timestamp 1605641404
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_140
timestamp 1605641404
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1605641404
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1605641404
transform 1 0 16100 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 16836 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_167
timestamp 1605641404
transform 1 0 16468 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1564 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1605641404
transform 1 0 4232 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1605641404
transform 1 0 3220 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_21
timestamp 1605641404
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_32
timestamp 1605641404
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1605641404
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1605641404
transform 1 0 5244 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_43
timestamp 1605641404
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1605641404
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1605641404
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1605641404
transform 1 0 7820 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 8280 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1605641404
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_76
timestamp 1605641404
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1605641404
transform 1 0 9936 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 10304 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_94
timestamp 1605641404
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_116
timestamp 1605641404
transform 1 0 11776 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1605641404
transform 1 0 12788 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14352 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13340 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_131
timestamp 1605641404
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_142
timestamp 1605641404
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1605641404
transform 1 0 15364 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_153
timestamp 1605641404
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1605641404
transform 1 0 16192 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 16836 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1605641404
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1605641404
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4876 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1605641404
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_36
timestamp 1605641404
transform 1 0 4416 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_40
timestamp 1605641404
transform 1 0 4784 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1605641404
transform 1 0 6532 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_57
timestamp 1605641404
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1605641404
transform 1 0 8280 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7360 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_77
timestamp 1605641404
transform 1 0 8188 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10488 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1605641404
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_87
timestamp 1605641404
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12420 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_118
timestamp 1605641404
transform 1 0 11960 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_122
timestamp 1605641404
transform 1 0 12328 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13432 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_132
timestamp 1605641404
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_143
timestamp 1605641404
transform 1 0 14260 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1605641404
transform 1 0 14628 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1605641404
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1605641404
transform 1 0 16100 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 16836 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_167
timestamp 1605641404
transform 1 0 16468 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_19
timestamp 1605641404
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1605641404
transform 1 0 4048 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 4416 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 3036 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1605641404
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1605641404
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1605641404
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_52
timestamp 1605641404
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1605641404
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1605641404
transform 1 0 7268 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7544 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_66
timestamp 1605641404
transform 1 0 7176 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10304 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9292 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_86
timestamp 1605641404
transform 1 0 9016 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_98
timestamp 1605641404
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1605641404
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1605641404
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12696 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14352 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_142
timestamp 1605641404
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15364 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_153
timestamp 1605641404
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1605641404
transform 1 0 16192 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 16836 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 1932 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1605641404
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_18
timestamp 1605641404
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1605641404
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1605641404
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5336 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 5060 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_62
timestamp 1605641404
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1605641404
transform 1 0 6992 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7728 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_12_68
timestamp 1605641404
transform 1 0 7360 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1605641404
transform 1 0 9936 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10488 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_93
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_100
timestamp 1605641404
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 11500 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_111
timestamp 1605641404
transform 1 0 11316 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 13524 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 13156 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_129
timestamp 1605641404
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1605641404
transform 1 0 13432 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1605641404
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_163
timestamp 1605641404
transform 1 0 16100 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 16836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1605641404
transform 1 0 16468 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_7
timestamp 1605641404
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1605641404
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1605641404
transform 1 0 1564 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_20
timestamp 1605641404
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2116 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 1932 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1605641404
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_25
timestamp 1605641404
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 3588 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_36
timestamp 1605641404
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_38
timestamp 1605641404
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1605641404
transform 1 0 4508 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1605641404
transform 1 0 4784 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 3128 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1605641404
transform 1 0 6624 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1605641404
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5520 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_44
timestamp 1605641404
transform 1 0 5152 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1605641404
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_46
timestamp 1605641404
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_57
timestamp 1605641404
transform 1 0 6348 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1605641404
transform 1 0 8556 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1605641404
transform 1 0 8188 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1605641404
transform 1 0 7176 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_78
timestamp 1605641404
transform 1 0 8280 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_64
timestamp 1605641404
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 1605641404
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_86
timestamp 1605641404
transform 1 0 9016 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_85
timestamp 1605641404
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1605641404
transform 1 0 9108 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_96
timestamp 1605641404
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_96
timestamp 1605641404
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1605641404
transform 1 0 10120 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10120 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11132 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1605641404
transform 1 0 11132 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12328 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_107
timestamp 1605641404
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1605641404
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_107
timestamp 1605641404
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_118
timestamp 1605641404
transform 1 0 11960 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13524 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1605641404
transform 1 0 13432 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1605641404
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_143
timestamp 1605641404
transform 1 0 14260 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_131
timestamp 1605641404
transform 1 0 13156 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14812 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1605641404
transform 1 0 16284 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1605641404
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_163
timestamp 1605641404
transform 1 0 16100 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 16836 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 16836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_167
timestamp 1605641404
transform 1 0 16468 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1605641404
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 3036 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1605641404
transform 1 0 4048 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1605641404
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_41
timestamp 1605641404
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5060 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1605641404
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1605641404
transform 1 0 8096 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8648 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_71
timestamp 1605641404
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_75
timestamp 1605641404
transform 1 0 8004 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_80
timestamp 1605641404
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 10304 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1605641404
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 11960 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_116
timestamp 1605641404
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1605641404
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_123
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1605641404
transform 1 0 13708 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1605641404
transform 1 0 12696 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_135
timestamp 1605641404
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14904 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_146
timestamp 1605641404
transform 1 0 14536 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1605641404
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 16836 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 1932 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1605641404
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1605641404
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 4692 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1605641404
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_36
timestamp 1605641404
transform 1 0 4416 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5980 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4968 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_51
timestamp 1605641404
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7912 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1605641404
transform 1 0 7636 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1605641404
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10120 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1605641404
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_96
timestamp 1605641404
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 11132 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_107
timestamp 1605641404
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1605641404
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12788 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_143
timestamp 1605641404
transform 1 0 14260 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1605641404
transform 1 0 14628 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1605641404
transform 1 0 16284 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1605641404
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1605641404
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 16836 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1748 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 3496 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_23
timestamp 1605641404
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_42 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4968 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1605641404
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1605641404
transform 1 0 6900 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7360 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_66
timestamp 1605641404
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10304 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9200 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_84
timestamp 1605641404
transform 1 0 8832 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_97
timestamp 1605641404
transform 1 0 10028 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1605641404
transform 1 0 11316 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1605641404
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1605641404
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_123
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12696 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 14352 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1605641404
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1605641404
transform 1 0 16008 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_160
timestamp 1605641404
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1605641404
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 16836 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1605641404
transform 1 0 1472 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 2944 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 1932 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_7
timestamp 1605641404
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_18
timestamp 1605641404
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1605641404
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6164 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_48
timestamp 1605641404
transform 1 0 5520 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_54
timestamp 1605641404
transform 1 0 6072 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 7176 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_64
timestamp 1605641404
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_82
timestamp 1605641404
transform 1 0 8648 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1605641404
transform 1 0 9844 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1605641404
transform 1 0 9016 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10396 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1605641404
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_99
timestamp 1605641404
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1605641404
transform 1 0 12144 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_117
timestamp 1605641404
transform 1 0 11868 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_124
timestamp 1605641404
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1605641404
transform 1 0 13708 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12696 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_135
timestamp 1605641404
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_140
timestamp 1605641404
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1605641404
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1605641404
transform 1 0 16100 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 16836 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_167
timestamp 1605641404
transform 1 0 16468 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 2300 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2944 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 1932 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_18
timestamp 1605641404
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1605641404
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 4692 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4692 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_36
timestamp 1605641404
transform 1 0 4416 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1605641404
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_32
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_38
timestamp 1605641404
transform 1 0 4600 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5704 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_48
timestamp 1605641404
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_62
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1605641404
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7360 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1605641404
transform 1 0 7544 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_66
timestamp 1605641404
transform 1 0 7176 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_79
timestamp 1605641404
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1605641404
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1605641404
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1605641404
transform 1 0 8832 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9660 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1605641404
transform 1 0 9200 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1605641404
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_102
timestamp 1605641404
transform 1 0 10488 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1605641404
transform 1 0 10672 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1605641404
transform 1 0 10764 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 11224 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_109
timestamp 1605641404
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1605641404
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_108
timestamp 1605641404
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12972 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13892 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1605641404
transform 1 0 12880 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1605641404
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1605641404
transform 1 0 14444 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_126
timestamp 1605641404
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_137
timestamp 1605641404
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14904 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1605641404
transform 1 0 15548 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_149
timestamp 1605641404
transform 1 0 14812 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1605641404
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1605641404
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1605641404
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_166
timestamp 1605641404
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 16836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 16836 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 2024 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp 1605641404
transform 1 0 1932 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_19
timestamp 1605641404
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 4140 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 3036 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_30
timestamp 1605641404
transform 1 0 3864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1605641404
transform 1 0 6164 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_42
timestamp 1605641404
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1605641404
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_58
timestamp 1605641404
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1605641404
transform 1 0 8648 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_78
timestamp 1605641404
transform 1 0 8280 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1605641404
transform 1 0 9660 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_91
timestamp 1605641404
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_102
timestamp 1605641404
transform 1 0 10488 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1605641404
transform 1 0 10856 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_109
timestamp 1605641404
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1605641404
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1605641404
transform 1 0 14076 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1605641404
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15364 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_150
timestamp 1605641404
transform 1 0 14904 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_154
timestamp 1605641404
transform 1 0 15272 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1605641404
transform 1 0 16192 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 16836 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 2024 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_9
timestamp 1605641404
transform 1 0 1932 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_19 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2852 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4140 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 5152 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_42
timestamp 1605641404
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_53
timestamp 1605641404
transform 1 0 5980 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 1605641404
transform 1 0 6716 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6900 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1605641404
transform 1 0 8648 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_72
timestamp 1605641404
transform 1 0 7728 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1605641404
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10212 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_91
timestamp 1605641404
transform 1 0 9476 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_94
timestamp 1605641404
transform 1 0 9752 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_98
timestamp 1605641404
transform 1 0 10120 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12604 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_108
timestamp 1605641404
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1605641404
transform 1 0 12052 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_123
timestamp 1605641404
transform 1 0 12420 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_134
timestamp 1605641404
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1605641404
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14628 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15456 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_153
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1605641404
transform 1 0 16284 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 16836 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 570 0 626 480 6 bottom_grid_pin_0_
port 0 nsew default tristate
rlabel metal2 s 11794 0 11850 480 6 bottom_grid_pin_10_
port 1 nsew default tristate
rlabel metal2 s 12898 0 12954 480 6 bottom_grid_pin_11_
port 2 nsew default tristate
rlabel metal2 s 14094 0 14150 480 6 bottom_grid_pin_12_
port 3 nsew default tristate
rlabel metal2 s 15198 0 15254 480 6 bottom_grid_pin_13_
port 4 nsew default tristate
rlabel metal2 s 16302 0 16358 480 6 bottom_grid_pin_14_
port 5 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 bottom_grid_pin_15_
port 6 nsew default tristate
rlabel metal2 s 1674 0 1730 480 6 bottom_grid_pin_1_
port 7 nsew default tristate
rlabel metal2 s 2778 0 2834 480 6 bottom_grid_pin_2_
port 8 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 bottom_grid_pin_3_
port 9 nsew default tristate
rlabel metal2 s 5078 0 5134 480 6 bottom_grid_pin_4_
port 10 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 bottom_grid_pin_5_
port 11 nsew default tristate
rlabel metal2 s 7286 0 7342 480 6 bottom_grid_pin_6_
port 12 nsew default tristate
rlabel metal2 s 8390 0 8446 480 6 bottom_grid_pin_7_
port 13 nsew default tristate
rlabel metal2 s 9586 0 9642 480 6 bottom_grid_pin_8_
port 14 nsew default tristate
rlabel metal2 s 10690 0 10746 480 6 bottom_grid_pin_9_
port 15 nsew default tristate
rlabel metal2 s 6734 16520 6790 17000 6 ccff_head
port 16 nsew default input
rlabel metal2 s 11242 16520 11298 17000 6 ccff_tail
port 17 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_in[0]
port 18 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[10]
port 19 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[11]
port 20 nsew default input
rlabel metal3 s 0 13744 480 13864 6 chanx_left_in[12]
port 21 nsew default input
rlabel metal3 s 0 14152 480 14272 6 chanx_left_in[13]
port 22 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[14]
port 23 nsew default input
rlabel metal3 s 0 14968 480 15088 6 chanx_left_in[15]
port 24 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[16]
port 25 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[17]
port 26 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chanx_left_in[18]
port 27 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_in[19]
port 28 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[1]
port 29 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[2]
port 30 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_left_in[3]
port 31 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[4]
port 32 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[5]
port 33 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[6]
port 34 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[7]
port 35 nsew default input
rlabel metal3 s 0 11976 480 12096 6 chanx_left_in[8]
port 36 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_in[9]
port 37 nsew default input
rlabel metal3 s 0 144 480 264 6 chanx_left_out[0]
port 38 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[10]
port 39 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 chanx_left_out[11]
port 40 nsew default tristate
rlabel metal3 s 0 5176 480 5296 6 chanx_left_out[12]
port 41 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[13]
port 42 nsew default tristate
rlabel metal3 s 0 5992 480 6112 6 chanx_left_out[14]
port 43 nsew default tristate
rlabel metal3 s 0 6400 480 6520 6 chanx_left_out[15]
port 44 nsew default tristate
rlabel metal3 s 0 6944 480 7064 6 chanx_left_out[16]
port 45 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[17]
port 46 nsew default tristate
rlabel metal3 s 0 7760 480 7880 6 chanx_left_out[18]
port 47 nsew default tristate
rlabel metal3 s 0 8168 480 8288 6 chanx_left_out[19]
port 48 nsew default tristate
rlabel metal3 s 0 552 480 672 6 chanx_left_out[1]
port 49 nsew default tristate
rlabel metal3 s 0 960 480 1080 6 chanx_left_out[2]
port 50 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[3]
port 51 nsew default tristate
rlabel metal3 s 0 1776 480 1896 6 chanx_left_out[4]
port 52 nsew default tristate
rlabel metal3 s 0 2184 480 2304 6 chanx_left_out[5]
port 53 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[6]
port 54 nsew default tristate
rlabel metal3 s 0 3000 480 3120 6 chanx_left_out[7]
port 55 nsew default tristate
rlabel metal3 s 0 3544 480 3664 6 chanx_left_out[8]
port 56 nsew default tristate
rlabel metal3 s 0 3952 480 4072 6 chanx_left_out[9]
port 57 nsew default tristate
rlabel metal3 s 17520 8576 18000 8696 6 chanx_right_in[0]
port 58 nsew default input
rlabel metal3 s 17520 12792 18000 12912 6 chanx_right_in[10]
port 59 nsew default input
rlabel metal3 s 17520 13200 18000 13320 6 chanx_right_in[11]
port 60 nsew default input
rlabel metal3 s 17520 13744 18000 13864 6 chanx_right_in[12]
port 61 nsew default input
rlabel metal3 s 17520 14152 18000 14272 6 chanx_right_in[13]
port 62 nsew default input
rlabel metal3 s 17520 14560 18000 14680 6 chanx_right_in[14]
port 63 nsew default input
rlabel metal3 s 17520 14968 18000 15088 6 chanx_right_in[15]
port 64 nsew default input
rlabel metal3 s 17520 15376 18000 15496 6 chanx_right_in[16]
port 65 nsew default input
rlabel metal3 s 17520 15784 18000 15904 6 chanx_right_in[17]
port 66 nsew default input
rlabel metal3 s 17520 16192 18000 16312 6 chanx_right_in[18]
port 67 nsew default input
rlabel metal3 s 17520 16600 18000 16720 6 chanx_right_in[19]
port 68 nsew default input
rlabel metal3 s 17520 8984 18000 9104 6 chanx_right_in[1]
port 69 nsew default input
rlabel metal3 s 17520 9392 18000 9512 6 chanx_right_in[2]
port 70 nsew default input
rlabel metal3 s 17520 9800 18000 9920 6 chanx_right_in[3]
port 71 nsew default input
rlabel metal3 s 17520 10344 18000 10464 6 chanx_right_in[4]
port 72 nsew default input
rlabel metal3 s 17520 10752 18000 10872 6 chanx_right_in[5]
port 73 nsew default input
rlabel metal3 s 17520 11160 18000 11280 6 chanx_right_in[6]
port 74 nsew default input
rlabel metal3 s 17520 11568 18000 11688 6 chanx_right_in[7]
port 75 nsew default input
rlabel metal3 s 17520 11976 18000 12096 6 chanx_right_in[8]
port 76 nsew default input
rlabel metal3 s 17520 12384 18000 12504 6 chanx_right_in[9]
port 77 nsew default input
rlabel metal3 s 17520 144 18000 264 6 chanx_right_out[0]
port 78 nsew default tristate
rlabel metal3 s 17520 4360 18000 4480 6 chanx_right_out[10]
port 79 nsew default tristate
rlabel metal3 s 17520 4768 18000 4888 6 chanx_right_out[11]
port 80 nsew default tristate
rlabel metal3 s 17520 5176 18000 5296 6 chanx_right_out[12]
port 81 nsew default tristate
rlabel metal3 s 17520 5584 18000 5704 6 chanx_right_out[13]
port 82 nsew default tristate
rlabel metal3 s 17520 5992 18000 6112 6 chanx_right_out[14]
port 83 nsew default tristate
rlabel metal3 s 17520 6400 18000 6520 6 chanx_right_out[15]
port 84 nsew default tristate
rlabel metal3 s 17520 6944 18000 7064 6 chanx_right_out[16]
port 85 nsew default tristate
rlabel metal3 s 17520 7352 18000 7472 6 chanx_right_out[17]
port 86 nsew default tristate
rlabel metal3 s 17520 7760 18000 7880 6 chanx_right_out[18]
port 87 nsew default tristate
rlabel metal3 s 17520 8168 18000 8288 6 chanx_right_out[19]
port 88 nsew default tristate
rlabel metal3 s 17520 552 18000 672 6 chanx_right_out[1]
port 89 nsew default tristate
rlabel metal3 s 17520 960 18000 1080 6 chanx_right_out[2]
port 90 nsew default tristate
rlabel metal3 s 17520 1368 18000 1488 6 chanx_right_out[3]
port 91 nsew default tristate
rlabel metal3 s 17520 1776 18000 1896 6 chanx_right_out[4]
port 92 nsew default tristate
rlabel metal3 s 17520 2184 18000 2304 6 chanx_right_out[5]
port 93 nsew default tristate
rlabel metal3 s 17520 2592 18000 2712 6 chanx_right_out[6]
port 94 nsew default tristate
rlabel metal3 s 17520 3000 18000 3120 6 chanx_right_out[7]
port 95 nsew default tristate
rlabel metal3 s 17520 3544 18000 3664 6 chanx_right_out[8]
port 96 nsew default tristate
rlabel metal3 s 17520 3952 18000 4072 6 chanx_right_out[9]
port 97 nsew default tristate
rlabel metal2 s 2226 16520 2282 17000 6 prog_clk
port 98 nsew default input
rlabel metal2 s 15750 16520 15806 17000 6 top_grid_pin_0_
port 99 nsew default tristate
rlabel metal4 s 3576 2128 3896 14736 6 VPWR
port 100 nsew default input
rlabel metal4 s 6208 2128 6528 14736 6 VGND
port 101 nsew default input
<< properties >>
string FIXED_BBOX 0 0 18000 17000
<< end >>
