VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 2.400 18.320 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 2.400 53.680 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 2.400 89.720 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 2.400 125.080 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 2.400 161.120 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 2.400 ;
    END
  END address[6]
  PIN address[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 2.400 ;
    END
  END address[7]
  PIN address[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 2.400 196.480 ;
    END
  END address[8]
  PIN address[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 2.400 ;
    END
  END address[9]
  PIN bottom_width_0_height_0__pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 2.400 ;
    END
  END bottom_width_0_height_0__pin_10_
  PIN bottom_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.490 247.600 41.770 250.000 ;
    END
  END bottom_width_0_height_0__pin_14_
  PIN bottom_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 124.480 250.000 125.080 ;
    END
  END bottom_width_0_height_0__pin_2_
  PIN bottom_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 247.600 14.170 250.000 ;
    END
  END bottom_width_0_height_0__pin_6_
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 2.400 ;
    END
  END clk
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 74.160 250.000 74.760 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 24.520 250.000 25.120 ;
    END
  END enable
  PIN left_width_0_height_0__pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.750 247.600 125.030 250.000 ;
    END
  END left_width_0_height_0__pin_11_
  PIN left_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 247.600 69.370 250.000 ;
    END
  END left_width_0_height_0__pin_3_
  PIN left_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.150 247.600 97.430 250.000 ;
    END
  END left_width_0_height_0__pin_7_
  PIN reset
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 2.400 ;
    END
  END reset
  PIN right_width_0_height_0__pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 2.400 232.520 ;
    END
  END right_width_0_height_0__pin_13_
  PIN right_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 152.350 247.600 152.630 250.000 ;
    END
  END right_width_0_height_0__pin_1_
  PIN right_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.410 247.600 180.690 250.000 ;
    END
  END right_width_0_height_0__pin_5_
  PIN right_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.010 247.600 208.290 250.000 ;
    END
  END right_width_0_height_0__pin_9_
  PIN set
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 2.400 ;
    END
  END set
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 174.120 250.000 174.720 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 2.400 ;
    END
  END top_width_0_height_0__pin_12_
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 235.610 247.600 235.890 250.000 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 224.440 250.000 225.040 ;
    END
  END top_width_0_height_0__pin_8_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 236.880 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 236.725 ;
      LAYER met1 ;
        RECT 0.530 0.380 244.260 236.880 ;
      LAYER met2 ;
        RECT 0.550 247.320 13.610 247.930 ;
        RECT 14.450 247.320 41.210 247.930 ;
        RECT 42.050 247.320 68.810 247.930 ;
        RECT 69.650 247.320 96.870 247.930 ;
        RECT 97.710 247.320 124.470 247.930 ;
        RECT 125.310 247.320 152.070 247.930 ;
        RECT 152.910 247.320 180.130 247.930 ;
        RECT 180.970 247.320 207.730 247.930 ;
        RECT 208.570 247.320 235.330 247.930 ;
        RECT 236.170 247.320 247.850 247.930 ;
        RECT 0.550 2.680 247.850 247.320 ;
        RECT 0.550 0.270 13.610 2.680 ;
        RECT 14.450 0.270 41.210 2.680 ;
        RECT 42.050 0.270 68.810 2.680 ;
        RECT 69.650 0.270 96.870 2.680 ;
        RECT 97.710 0.270 124.470 2.680 ;
        RECT 125.310 0.270 152.070 2.680 ;
        RECT 152.910 0.270 180.130 2.680 ;
        RECT 180.970 0.270 207.730 2.680 ;
        RECT 208.570 0.270 235.330 2.680 ;
        RECT 236.170 0.270 247.850 2.680 ;
      LAYER met3 ;
        RECT 0.310 232.920 248.130 236.805 ;
        RECT 2.800 231.520 248.130 232.920 ;
        RECT 0.310 225.440 248.130 231.520 ;
        RECT 0.310 224.040 247.200 225.440 ;
        RECT 0.310 196.880 248.130 224.040 ;
        RECT 2.800 195.480 248.130 196.880 ;
        RECT 0.310 175.120 248.130 195.480 ;
        RECT 0.310 173.720 247.200 175.120 ;
        RECT 0.310 161.520 248.130 173.720 ;
        RECT 2.800 160.120 248.130 161.520 ;
        RECT 0.310 125.480 248.130 160.120 ;
        RECT 2.800 124.080 247.200 125.480 ;
        RECT 0.310 90.120 248.130 124.080 ;
        RECT 2.800 88.720 248.130 90.120 ;
        RECT 0.310 75.160 248.130 88.720 ;
        RECT 0.310 73.760 247.200 75.160 ;
        RECT 0.310 54.080 248.130 73.760 ;
        RECT 2.800 52.680 248.130 54.080 ;
        RECT 0.310 25.520 248.130 52.680 ;
        RECT 0.310 24.120 247.200 25.520 ;
        RECT 0.310 18.720 248.130 24.120 ;
        RECT 2.800 17.320 248.130 18.720 ;
        RECT 0.310 10.715 248.130 17.320 ;
      LAYER met4 ;
        RECT 96.895 10.640 97.440 236.880 ;
        RECT 99.840 10.640 248.105 236.880 ;
  END
END grid_clb
END LIBRARY

